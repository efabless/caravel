magic
tech sky130A
magscale 1 2
timestamp 1675851710
<< viali >>
rect 2881 18377 2915 18411
rect 18429 18377 18463 18411
rect 2421 18309 2455 18343
rect 6009 18309 6043 18343
rect 5457 18241 5491 18275
rect 8217 18241 8251 18275
rect 10517 18241 10551 18275
rect 857 18173 891 18207
rect 1593 18173 1627 18207
rect 3617 18173 3651 18207
rect 3985 18173 4019 18207
rect 4169 18173 4203 18207
rect 4537 18173 4571 18207
rect 6745 18173 6779 18207
rect 7941 18173 7975 18207
rect 8769 18173 8803 18207
rect 11713 18173 11747 18207
rect 12725 18173 12759 18207
rect 12909 18173 12943 18207
rect 14197 18173 14231 18207
rect 14933 18173 14967 18207
rect 16589 18173 16623 18207
rect 17969 18173 18003 18207
rect 1225 18105 1259 18139
rect 3341 18105 3375 18139
rect 6377 18105 6411 18139
rect 7021 18105 7055 18139
rect 10425 18105 10459 18139
rect 13921 18105 13955 18139
rect 14841 18105 14875 18139
rect 1777 18037 1811 18071
rect 4445 18037 4479 18071
rect 5549 18037 5583 18071
rect 5641 18037 5675 18071
rect 7573 18037 7607 18071
rect 8033 18037 8067 18071
rect 9413 18037 9447 18071
rect 9965 18037 9999 18071
rect 10333 18037 10367 18071
rect 11161 18037 11195 18071
rect 15485 18037 15519 18071
rect 15945 18037 15979 18071
rect 17785 18037 17819 18071
rect 3433 17833 3467 17867
rect 4546 17765 4580 17799
rect 7849 17765 7883 17799
rect 9965 17765 9999 17799
rect 16543 17765 16577 17799
rect 17417 17765 17451 17799
rect 2881 17697 2915 17731
rect 5181 17697 5215 17731
rect 12633 17697 12667 17731
rect 12909 17697 12943 17731
rect 14749 17697 14783 17731
rect 17141 17697 17175 17731
rect 581 17629 615 17663
rect 857 17629 891 17663
rect 4813 17629 4847 17663
rect 12357 17629 12391 17663
rect 12541 17629 12575 17663
rect 13369 17629 13403 17663
rect 15117 17629 15151 17663
rect 3065 17561 3099 17595
rect 17233 17561 17267 17595
rect 2329 17493 2363 17527
rect 6469 17493 6503 17527
rect 9137 17493 9171 17527
rect 11437 17493 11471 17527
rect 12449 17493 12483 17527
rect 17141 17493 17175 17527
rect 2513 17289 2547 17323
rect 2697 17289 2731 17323
rect 5549 17289 5583 17323
rect 8263 17289 8297 17323
rect 15577 17289 15611 17323
rect 857 17221 891 17255
rect 12081 17221 12115 17255
rect 3065 17153 3099 17187
rect 6837 17153 6871 17187
rect 8815 17153 8849 17187
rect 10241 17153 10275 17187
rect 11529 17153 11563 17187
rect 13829 17153 13863 17187
rect 16497 17153 16531 17187
rect 1132 17085 1166 17119
rect 1225 17085 1259 17119
rect 2145 17085 2179 17119
rect 4261 17085 4295 17119
rect 6469 17085 6503 17119
rect 10609 17085 10643 17119
rect 12449 17085 12483 17119
rect 12725 17085 12759 17119
rect 13185 17085 13219 17119
rect 16129 17085 16163 17119
rect 14105 17017 14139 17051
rect 2513 16949 2547 16983
rect 3617 16949 3651 16983
rect 11621 16949 11655 16983
rect 11713 16949 11747 16983
rect 12633 16949 12667 16983
rect 17923 16949 17957 16983
rect 2145 16745 2179 16779
rect 4261 16745 4295 16779
rect 7803 16745 7837 16779
rect 18245 16745 18279 16779
rect 1409 16677 1443 16711
rect 4169 16677 4203 16711
rect 7021 16677 7055 16711
rect 1317 16609 1351 16643
rect 1777 16609 1811 16643
rect 2053 16609 2087 16643
rect 2881 16609 2915 16643
rect 3249 16609 3283 16643
rect 3525 16609 3559 16643
rect 4077 16609 4111 16643
rect 4813 16609 4847 16643
rect 9229 16609 9263 16643
rect 9597 16609 9631 16643
rect 9965 16609 9999 16643
rect 12817 16609 12851 16643
rect 13277 16609 13311 16643
rect 14197 16609 14231 16643
rect 14933 16609 14967 16643
rect 17785 16609 17819 16643
rect 18429 16609 18463 16643
rect 2421 16541 2455 16575
rect 4629 16541 4663 16575
rect 14289 16541 14323 16575
rect 15209 16541 15243 16575
rect 1639 16473 1673 16507
rect 2329 16473 2363 16507
rect 5733 16473 5767 16507
rect 11253 16473 11287 16507
rect 13461 16473 13495 16507
rect 1501 16405 1535 16439
rect 2237 16405 2271 16439
rect 12725 16405 12759 16439
rect 13921 16405 13955 16439
rect 16681 16405 16715 16439
rect 17141 16405 17175 16439
rect 5917 16201 5951 16235
rect 12449 16201 12483 16235
rect 13829 16201 13863 16235
rect 18429 16133 18463 16167
rect 4169 16065 4203 16099
rect 16497 16065 16531 16099
rect 2421 15997 2455 16031
rect 2605 15997 2639 16031
rect 6653 15997 6687 16031
rect 8401 15997 8435 16031
rect 16129 15997 16163 16031
rect 4445 15929 4479 15963
rect 8769 15929 8803 15963
rect 11161 15929 11195 15963
rect 15301 15929 15335 15963
rect 2513 15861 2547 15895
rect 10057 15861 10091 15895
rect 17923 15861 17957 15895
rect 3249 15657 3283 15691
rect 5733 15657 5767 15691
rect 11989 15657 12023 15691
rect 12725 15657 12759 15691
rect 14013 15657 14047 15691
rect 18245 15657 18279 15691
rect 4537 15589 4571 15623
rect 7021 15589 7055 15623
rect 13921 15589 13955 15623
rect 7757 15521 7791 15555
rect 12817 15521 12851 15555
rect 16497 15521 16531 15555
rect 17969 15521 18003 15555
rect 18429 15521 18463 15555
rect 8033 15453 8067 15487
rect 10241 15453 10275 15487
rect 10517 15453 10551 15487
rect 12909 15453 12943 15487
rect 13829 15453 13863 15487
rect 9505 15317 9539 15351
rect 12357 15317 12391 15351
rect 14381 15317 14415 15351
rect 15209 15317 15243 15351
rect 5917 15113 5951 15147
rect 8125 15113 8159 15147
rect 11253 15113 11287 15147
rect 14013 15113 14047 15147
rect 14749 15045 14783 15079
rect 2145 14977 2179 15011
rect 2789 14977 2823 15011
rect 6377 14977 6411 15011
rect 13093 14977 13127 15011
rect 15301 14977 15335 15011
rect 2053 14909 2087 14943
rect 2867 14909 2901 14943
rect 3433 14909 3467 14943
rect 3617 14909 3651 14943
rect 4077 14909 4111 14943
rect 4169 14909 4203 14943
rect 4261 14909 4295 14943
rect 5181 14909 5215 14943
rect 5825 14909 5859 14943
rect 11345 14909 11379 14943
rect 11989 14909 12023 14943
rect 12449 14909 12483 14943
rect 12541 14909 12575 14943
rect 12633 14909 12667 14943
rect 13001 14909 13035 14943
rect 13185 14909 13219 14943
rect 13829 14909 13863 14943
rect 13921 14909 13955 14943
rect 14381 14909 14415 14943
rect 15117 14909 15151 14943
rect 16221 14909 16255 14943
rect 1961 14841 1995 14875
rect 4629 14841 4663 14875
rect 4997 14841 5031 14875
rect 6653 14841 6687 14875
rect 8769 14841 8803 14875
rect 16497 14841 16531 14875
rect 1593 14773 1627 14807
rect 3157 14773 3191 14807
rect 3525 14773 3559 14807
rect 4445 14773 4479 14807
rect 10057 14773 10091 14807
rect 11897 14773 11931 14807
rect 12265 14773 12299 14807
rect 14289 14773 14323 14807
rect 15209 14773 15243 14807
rect 17969 14773 18003 14807
rect 2329 14569 2363 14603
rect 2789 14569 2823 14603
rect 3249 14569 3283 14603
rect 7665 14569 7699 14603
rect 11069 14569 11103 14603
rect 11621 14569 11655 14603
rect 12633 14569 12667 14603
rect 13277 14569 13311 14603
rect 15025 14569 15059 14603
rect 17141 14569 17175 14603
rect 857 14501 891 14535
rect 4077 14501 4111 14535
rect 9137 14501 9171 14535
rect 14013 14501 14047 14535
rect 15117 14501 15151 14535
rect 18245 14501 18279 14535
rect 581 14433 615 14467
rect 3157 14433 3191 14467
rect 3801 14433 3835 14467
rect 4629 14433 4663 14467
rect 4813 14433 4847 14467
rect 5181 14433 5215 14467
rect 11345 14433 11379 14467
rect 11896 14433 11930 14467
rect 11989 14433 12023 14467
rect 12909 14433 12943 14467
rect 13002 14433 13036 14467
rect 13921 14433 13955 14467
rect 15485 14433 15519 14467
rect 15639 14433 15673 14467
rect 16405 14433 16439 14467
rect 16681 14433 16715 14467
rect 3433 14365 3467 14399
rect 3893 14365 3927 14399
rect 4077 14365 4111 14399
rect 4721 14365 4755 14399
rect 5549 14365 5583 14399
rect 9413 14365 9447 14399
rect 11069 14365 11103 14399
rect 14105 14365 14139 14399
rect 16129 14365 16163 14399
rect 16313 14365 16347 14399
rect 17785 14365 17819 14399
rect 18061 14297 18095 14331
rect 6975 14229 7009 14263
rect 10057 14229 10091 14263
rect 11253 14229 11287 14263
rect 13553 14229 13587 14263
rect 15669 14229 15703 14263
rect 16221 14229 16255 14263
rect 5089 14025 5123 14059
rect 7021 14025 7055 14059
rect 10517 14025 10551 14059
rect 14289 14025 14323 14059
rect 15209 14025 15243 14059
rect 17969 14025 18003 14059
rect 6377 13889 6411 13923
rect 8769 13889 8803 13923
rect 13737 13889 13771 13923
rect 13829 13889 13863 13923
rect 16497 13889 16531 13923
rect 2881 13821 2915 13855
rect 7389 13821 7423 13855
rect 7757 13821 7791 13855
rect 8309 13821 8343 13855
rect 11345 13821 11379 13855
rect 14749 13821 14783 13855
rect 15485 13821 15519 13855
rect 16221 13821 16255 13855
rect 9045 13753 9079 13787
rect 13921 13753 13955 13787
rect 14565 13753 14599 13787
rect 3065 13685 3099 13719
rect 11253 13685 11287 13719
rect 3249 13481 3283 13515
rect 5273 13481 5307 13515
rect 7573 13481 7607 13515
rect 13093 13481 13127 13515
rect 16313 13481 16347 13515
rect 15025 13413 15059 13447
rect 17785 13413 17819 13447
rect 581 13345 615 13379
rect 2421 13345 2455 13379
rect 4537 13345 4571 13379
rect 10241 13345 10275 13379
rect 14381 13345 14415 13379
rect 17693 13345 17727 13379
rect 949 13277 983 13311
rect 6745 13277 6779 13311
rect 7021 13277 7055 13311
rect 9045 13277 9079 13311
rect 9321 13277 9355 13311
rect 10517 13277 10551 13311
rect 17877 13277 17911 13311
rect 11989 13141 12023 13175
rect 17325 13141 17359 13175
rect 1593 12937 1627 12971
rect 11253 12937 11287 12971
rect 16773 12937 16807 12971
rect 17969 12937 18003 12971
rect 2145 12801 2179 12835
rect 3249 12801 3283 12835
rect 3433 12801 3467 12835
rect 7573 12801 7607 12835
rect 7757 12801 7791 12835
rect 11437 12801 11471 12835
rect 12357 12801 12391 12835
rect 13921 12801 13955 12835
rect 17233 12801 17267 12835
rect 2053 12733 2087 12767
rect 4445 12733 4479 12767
rect 7849 12733 7883 12767
rect 11161 12733 11195 12767
rect 12541 12733 12575 12767
rect 12633 12733 12667 12767
rect 12725 12733 12759 12767
rect 14197 12733 14231 12767
rect 14657 12733 14691 12767
rect 14841 12733 14875 12767
rect 15301 12733 15335 12767
rect 16037 12733 16071 12767
rect 16221 12733 16255 12767
rect 16405 12733 16439 12767
rect 17509 12733 17543 12767
rect 1961 12665 1995 12699
rect 3157 12665 3191 12699
rect 4712 12665 4746 12699
rect 7205 12665 7239 12699
rect 11437 12665 11471 12699
rect 16773 12665 16807 12699
rect 17325 12665 17359 12699
rect 2789 12597 2823 12631
rect 5825 12597 5859 12631
rect 8217 12597 8251 12631
rect 14289 12393 14323 12427
rect 15669 12393 15703 12427
rect 5917 12325 5951 12359
rect 11161 12325 11195 12359
rect 11345 12325 11379 12359
rect 13921 12325 13955 12359
rect 16313 12325 16347 12359
rect 16681 12325 16715 12359
rect 17141 12325 17175 12359
rect 17601 12325 17635 12359
rect 2053 12257 2087 12291
rect 3341 12257 3375 12291
rect 3608 12257 3642 12291
rect 5273 12257 5307 12291
rect 5366 12257 5400 12291
rect 5641 12257 5675 12291
rect 6101 12257 6135 12291
rect 6193 12257 6227 12291
rect 9229 12257 9263 12291
rect 9597 12257 9631 12291
rect 11437 12257 11471 12291
rect 12541 12257 12575 12291
rect 13737 12257 13771 12291
rect 15117 12257 15151 12291
rect 16129 12257 16163 12291
rect 16589 12257 16623 12291
rect 16773 12257 16807 12291
rect 17509 12257 17543 12291
rect 17693 12257 17727 12291
rect 18429 12257 18463 12291
rect 7205 12189 7239 12223
rect 14013 12189 14047 12223
rect 14102 12189 14136 12223
rect 14196 12189 14230 12223
rect 14933 12189 14967 12223
rect 15025 12189 15059 12223
rect 15209 12189 15243 12223
rect 15945 12189 15979 12223
rect 4721 12121 4755 12155
rect 11161 12121 11195 12155
rect 18245 12121 18279 12155
rect 1961 12053 1995 12087
rect 6193 12053 6227 12087
rect 7803 12053 7837 12087
rect 12633 12053 12667 12087
rect 14749 12053 14783 12087
rect 7757 11849 7791 11883
rect 8033 11781 8067 11815
rect 1593 11713 1627 11747
rect 6469 11713 6503 11747
rect 12909 11713 12943 11747
rect 16589 11713 16623 11747
rect 1961 11645 1995 11679
rect 6009 11645 6043 11679
rect 7113 11645 7147 11679
rect 7205 11645 7239 11679
rect 7389 11645 7423 11679
rect 8033 11645 8067 11679
rect 8217 11645 8251 11679
rect 8769 11645 8803 11679
rect 9137 11645 9171 11679
rect 12817 11645 12851 11679
rect 15577 11645 15611 11679
rect 16313 11645 16347 11679
rect 7757 11577 7791 11611
rect 16856 11577 16890 11611
rect 3387 11509 3421 11543
rect 4537 11509 4571 11543
rect 10563 11509 10597 11543
rect 12357 11509 12391 11543
rect 12725 11509 12759 11543
rect 14289 11509 14323 11543
rect 16037 11509 16071 11543
rect 17969 11509 18003 11543
rect 18429 11509 18463 11543
rect 1685 11305 1719 11339
rect 2053 11305 2087 11339
rect 5549 11305 5583 11339
rect 8309 11305 8343 11339
rect 9597 11237 9631 11271
rect 3801 11169 3835 11203
rect 3985 11169 4019 11203
rect 5181 11169 5215 11203
rect 5274 11169 5308 11203
rect 9965 11169 9999 11203
rect 14013 11169 14047 11203
rect 14197 11169 14231 11203
rect 14749 11169 14783 11203
rect 17141 11169 17175 11203
rect 17295 11169 17329 11203
rect 17785 11169 17819 11203
rect 17878 11169 17912 11203
rect 1501 11101 1535 11135
rect 1593 11101 1627 11135
rect 10241 11101 10275 11135
rect 14105 11101 14139 11135
rect 15117 11101 15151 11135
rect 18153 11033 18187 11067
rect 3985 10965 4019 10999
rect 11713 10965 11747 10999
rect 16543 10965 16577 10999
rect 17325 10965 17359 10999
rect 2697 10761 2731 10795
rect 6469 10761 6503 10795
rect 7757 10761 7791 10795
rect 11161 10761 11195 10795
rect 15485 10761 15519 10795
rect 16957 10761 16991 10795
rect 17601 10761 17635 10795
rect 2145 10625 2179 10659
rect 3157 10625 3191 10659
rect 3341 10625 3375 10659
rect 4445 10625 4479 10659
rect 4537 10625 4571 10659
rect 11805 10625 11839 10659
rect 12817 10625 12851 10659
rect 2053 10557 2087 10591
rect 4261 10557 4295 10591
rect 6377 10557 6411 10591
rect 6653 10557 6687 10591
rect 6745 10557 6779 10591
rect 7665 10557 7699 10591
rect 8125 10557 8159 10591
rect 11529 10557 11563 10591
rect 15577 10557 15611 10591
rect 3065 10489 3099 10523
rect 12541 10489 12575 10523
rect 2421 10421 2455 10455
rect 4077 10421 4111 10455
rect 6929 10421 6963 10455
rect 11621 10421 11655 10455
rect 12173 10421 12207 10455
rect 12633 10421 12667 10455
rect 765 10217 799 10251
rect 3801 10217 3835 10251
rect 6561 10217 6595 10251
rect 7205 10217 7239 10251
rect 11897 10217 11931 10251
rect 12817 10217 12851 10251
rect 5273 10149 5307 10183
rect 8125 10149 8159 10183
rect 11345 10149 11379 10183
rect 17509 10149 17543 10183
rect 581 10081 615 10115
rect 1041 10081 1075 10115
rect 3801 10081 3835 10115
rect 5181 10081 5215 10115
rect 5365 10081 5399 10115
rect 5825 10081 5859 10115
rect 6285 10081 6319 10115
rect 7021 10081 7055 10115
rect 11161 10081 11195 10115
rect 11713 10081 11747 10115
rect 11897 10081 11931 10115
rect 12357 10081 12391 10115
rect 12449 10081 12483 10115
rect 12633 10081 12667 10115
rect 13277 10081 13311 10115
rect 13553 10081 13587 10115
rect 17417 10081 17451 10115
rect 17693 10081 17727 10115
rect 3893 10013 3927 10047
rect 4077 10013 4111 10047
rect 5641 10013 5675 10047
rect 6561 10013 6595 10047
rect 6837 10013 6871 10047
rect 7849 10013 7883 10047
rect 10885 10013 10919 10047
rect 13461 10013 13495 10047
rect 6009 9877 6043 9911
rect 6377 9877 6411 9911
rect 9597 9877 9631 9911
rect 10977 9877 11011 9911
rect 13093 9877 13127 9911
rect 17417 9877 17451 9911
rect 13001 9673 13035 9707
rect 8769 9605 8803 9639
rect 15945 9605 15979 9639
rect 17969 9605 18003 9639
rect 2145 9537 2179 9571
rect 4445 9537 4479 9571
rect 4537 9537 4571 9571
rect 7113 9537 7147 9571
rect 11897 9537 11931 9571
rect 15025 9537 15059 9571
rect 1961 9469 1995 9503
rect 2881 9469 2915 9503
rect 3065 9469 3099 9503
rect 7021 9469 7055 9503
rect 7205 9469 7239 9503
rect 9045 9469 9079 9503
rect 10149 9469 10183 9503
rect 11989 9469 12023 9503
rect 15209 9469 15243 9503
rect 15301 9469 15335 9503
rect 16221 9469 16255 9503
rect 16589 9469 16623 9503
rect 16856 9469 16890 9503
rect 2053 9401 2087 9435
rect 8769 9401 8803 9435
rect 15945 9401 15979 9435
rect 1593 9333 1627 9367
rect 2973 9333 3007 9367
rect 3985 9333 4019 9367
rect 4353 9333 4387 9367
rect 7757 9333 7791 9367
rect 8953 9333 8987 9367
rect 10149 9333 10183 9367
rect 12357 9333 12391 9367
rect 15025 9333 15059 9367
rect 16129 9333 16163 9367
rect 2329 9129 2363 9163
rect 3617 9129 3651 9163
rect 5181 9129 5215 9163
rect 7205 9129 7239 9163
rect 9367 9129 9401 9163
rect 11759 9129 11793 9163
rect 13001 9129 13035 9163
rect 18245 9129 18279 9163
rect 857 9061 891 9095
rect 13921 9061 13955 9095
rect 14197 9061 14231 9095
rect 3157 8993 3191 9027
rect 3249 8993 3283 9027
rect 3433 8993 3467 9027
rect 6305 8993 6339 9027
rect 9965 8993 9999 9027
rect 13645 8993 13679 9027
rect 14749 8993 14783 9027
rect 15117 8993 15151 9027
rect 17969 8993 18003 9027
rect 18429 8993 18463 9027
rect 581 8925 615 8959
rect 6561 8925 6595 8959
rect 7573 8925 7607 8959
rect 7941 8925 7975 8959
rect 10333 8925 10367 8959
rect 13093 8925 13127 8959
rect 13277 8925 13311 8959
rect 16543 8925 16577 8959
rect 13737 8857 13771 8891
rect 2881 8789 2915 8823
rect 12633 8789 12667 8823
rect 13645 8789 13679 8823
rect 2605 8585 2639 8619
rect 2973 8585 3007 8619
rect 6929 8585 6963 8619
rect 8125 8585 8159 8619
rect 8861 8585 8895 8619
rect 11161 8585 11195 8619
rect 13553 8585 13587 8619
rect 14013 8585 14047 8619
rect 17923 8585 17957 8619
rect 8033 8517 8067 8551
rect 8217 8449 8251 8483
rect 11621 8449 11655 8483
rect 11805 8449 11839 8483
rect 16129 8449 16163 8483
rect 2513 8381 2547 8415
rect 2789 8381 2823 8415
rect 3249 8381 3283 8415
rect 5549 8381 5583 8415
rect 6745 8381 6779 8415
rect 7021 8381 7055 8415
rect 7941 8381 7975 8415
rect 9137 8381 9171 8415
rect 11529 8381 11563 8415
rect 13553 8381 13587 8415
rect 13737 8381 13771 8415
rect 16497 8381 16531 8415
rect 3341 8313 3375 8347
rect 5273 8313 5307 8347
rect 6561 8313 6595 8347
rect 10793 8245 10827 8279
rect 2421 8041 2455 8075
rect 3249 8041 3283 8075
rect 15945 8041 15979 8075
rect 16589 8041 16623 8075
rect 17785 8041 17819 8075
rect 4537 7973 4571 8007
rect 10333 7973 10367 8007
rect 11161 7973 11195 8007
rect 14381 7973 14415 8007
rect 15669 7973 15703 8007
rect 5181 7905 5215 7939
rect 7941 7905 7975 7939
rect 8309 7905 8343 7939
rect 9045 7905 9079 7939
rect 10885 7905 10919 7939
rect 14933 7905 14967 7939
rect 15025 7905 15059 7939
rect 15301 7905 15335 7939
rect 16589 7905 16623 7939
rect 16773 7905 16807 7939
rect 17141 7905 17175 7939
rect 673 7837 707 7871
rect 949 7837 983 7871
rect 5549 7837 5583 7871
rect 8125 7837 8159 7871
rect 8861 7837 8895 7871
rect 17325 7837 17359 7871
rect 17417 7837 17451 7871
rect 7941 7769 7975 7803
rect 10057 7769 10091 7803
rect 15209 7769 15243 7803
rect 6975 7701 7009 7735
rect 13093 7701 13127 7735
rect 14749 7701 14783 7735
rect 1593 7497 1627 7531
rect 9873 7497 9907 7531
rect 15577 7497 15611 7531
rect 17233 7497 17267 7531
rect 3617 7429 3651 7463
rect 8953 7429 8987 7463
rect 9229 7429 9263 7463
rect 2145 7361 2179 7395
rect 3157 7361 3191 7395
rect 4445 7361 4479 7395
rect 4537 7361 4571 7395
rect 9045 7361 9079 7395
rect 9321 7361 9355 7395
rect 11805 7361 11839 7395
rect 12817 7361 12851 7395
rect 14105 7361 14139 7395
rect 1961 7293 1995 7327
rect 3249 7293 3283 7327
rect 4353 7293 4387 7327
rect 6837 7293 6871 7327
rect 8861 7293 8895 7327
rect 9965 7293 9999 7327
rect 10793 7293 10827 7327
rect 11529 7293 11563 7327
rect 12541 7293 12575 7327
rect 13829 7293 13863 7327
rect 15945 7293 15979 7327
rect 16129 7293 16163 7327
rect 16405 7293 16439 7327
rect 17417 7293 17451 7327
rect 17509 7293 17543 7327
rect 17601 7293 17635 7327
rect 2053 7225 2087 7259
rect 6377 7225 6411 7259
rect 8953 7225 8987 7259
rect 10701 7225 10735 7259
rect 2697 7157 2731 7191
rect 3985 7157 4019 7191
rect 5089 7157 5123 7191
rect 11161 7157 11195 7191
rect 11621 7157 11655 7191
rect 12173 7157 12207 7191
rect 12633 7157 12667 7191
rect 16037 7157 16071 7191
rect 11897 6953 11931 6987
rect 15393 6953 15427 6987
rect 2053 6817 2087 6851
rect 5181 6817 5215 6851
rect 5273 6817 5307 6851
rect 5733 6817 5767 6851
rect 10149 6817 10183 6851
rect 12541 6817 12575 6851
rect 12808 6817 12842 6851
rect 14933 6817 14967 6851
rect 15669 6817 15703 6851
rect 17969 6817 18003 6851
rect 18429 6817 18463 6851
rect 14749 6749 14783 6783
rect 15393 6749 15427 6783
rect 5549 6681 5583 6715
rect 13921 6681 13955 6715
rect 15117 6681 15151 6715
rect 15577 6681 15611 6715
rect 1961 6613 1995 6647
rect 5641 6613 5675 6647
rect 10412 6613 10446 6647
rect 14197 6613 14231 6647
rect 18245 6613 18279 6647
rect 12633 6409 12667 6443
rect 13645 6409 13679 6443
rect 14565 6409 14599 6443
rect 1593 6273 1627 6307
rect 1961 6273 1995 6307
rect 4261 6273 4295 6307
rect 6377 6273 6411 6307
rect 13001 6273 13035 6307
rect 15945 6273 15979 6307
rect 6745 6205 6779 6239
rect 8769 6205 8803 6239
rect 12909 6205 12943 6239
rect 16313 6205 16347 6239
rect 3433 6137 3467 6171
rect 4537 6137 4571 6171
rect 8217 6137 8251 6171
rect 9045 6137 9079 6171
rect 10793 6137 10827 6171
rect 17785 6137 17819 6171
rect 6009 6069 6043 6103
rect 2329 5865 2363 5899
rect 5181 5865 5215 5899
rect 6285 5865 6319 5899
rect 8585 5865 8619 5899
rect 8953 5865 8987 5899
rect 17693 5865 17727 5899
rect 581 5729 615 5763
rect 4629 5729 4663 5763
rect 4813 5729 4847 5763
rect 5365 5729 5399 5763
rect 5457 5729 5491 5763
rect 8125 5729 8159 5763
rect 8309 5729 8343 5763
rect 15025 5729 15059 5763
rect 17417 5729 17451 5763
rect 17693 5729 17727 5763
rect 857 5661 891 5695
rect 5549 5661 5583 5695
rect 5641 5661 5675 5695
rect 15301 5661 15335 5695
rect 4813 5593 4847 5627
rect 8309 5593 8343 5627
rect 16773 5593 16807 5627
rect 17601 5593 17635 5627
rect 2881 5525 2915 5559
rect 3617 5525 3651 5559
rect 4169 5525 4203 5559
rect 1685 5321 1719 5355
rect 6561 5321 6595 5355
rect 7665 5253 7699 5287
rect 2237 5185 2271 5219
rect 8125 5185 8159 5219
rect 8769 5185 8803 5219
rect 13093 5185 13127 5219
rect 13553 5185 13587 5219
rect 15577 5185 15611 5219
rect 15945 5185 15979 5219
rect 6745 5117 6779 5151
rect 6837 5117 6871 5151
rect 7205 5117 7239 5151
rect 7481 5117 7515 5151
rect 8033 5117 8067 5151
rect 8217 5117 8251 5151
rect 12725 5117 12759 5151
rect 2053 5049 2087 5083
rect 7113 5049 7147 5083
rect 9045 5049 9079 5083
rect 13829 5049 13863 5083
rect 16221 5049 16255 5083
rect 2145 4981 2179 5015
rect 10517 4981 10551 5015
rect 11299 4981 11333 5015
rect 17693 4981 17727 5015
rect 1961 4777 1995 4811
rect 3065 4777 3099 4811
rect 3617 4777 3651 4811
rect 4537 4777 4571 4811
rect 7941 4777 7975 4811
rect 12357 4777 12391 4811
rect 14013 4777 14047 4811
rect 14749 4777 14783 4811
rect 15209 4777 15243 4811
rect 2881 4709 2915 4743
rect 8401 4709 8435 4743
rect 9413 4709 9447 4743
rect 1869 4641 1903 4675
rect 2789 4641 2823 4675
rect 3341 4641 3375 4675
rect 3892 4641 3926 4675
rect 3985 4641 4019 4675
rect 4813 4641 4847 4675
rect 7573 4641 7607 4675
rect 7727 4641 7761 4675
rect 8309 4641 8343 4675
rect 8493 4641 8527 4675
rect 8953 4641 8987 4675
rect 9045 4641 9079 4675
rect 9321 4641 9355 4675
rect 10241 4641 10275 4675
rect 12541 4641 12575 4675
rect 12817 4641 12851 4675
rect 13737 4641 13771 4675
rect 13829 4641 13863 4675
rect 4537 4573 4571 4607
rect 10517 4573 10551 4607
rect 12633 4573 12667 4607
rect 14013 4573 14047 4607
rect 11989 4505 12023 4539
rect 12725 4505 12759 4539
rect 3249 4437 3283 4471
rect 4721 4437 4755 4471
rect 8769 4437 8803 4471
rect 857 4233 891 4267
rect 3433 4233 3467 4267
rect 5733 4233 5767 4267
rect 8953 4233 8987 4267
rect 14289 4233 14323 4267
rect 17785 4233 17819 4267
rect 6929 4165 6963 4199
rect 11437 4165 11471 4199
rect 12541 4165 12575 4199
rect 14197 4165 14231 4199
rect 15025 4165 15059 4199
rect 15393 4165 15427 4199
rect 17049 4165 17083 4199
rect 1041 4097 1075 4131
rect 1593 4097 1627 4131
rect 3985 4097 4019 4131
rect 4537 4097 4571 4131
rect 7113 4097 7147 4131
rect 8769 4097 8803 4131
rect 11161 4097 11195 4131
rect 11529 4097 11563 4131
rect 14381 4097 14415 4131
rect 15209 4097 15243 4131
rect 16957 4097 16991 4131
rect 17141 4097 17175 4131
rect 765 4029 799 4063
rect 1777 4029 1811 4063
rect 1869 4029 1903 4063
rect 1961 4029 1995 4063
rect 3341 4029 3375 4063
rect 3525 4029 3559 4063
rect 4353 4029 4387 4063
rect 5089 4029 5123 4063
rect 5273 4029 5307 4063
rect 5733 4029 5767 4063
rect 6009 4029 6043 4063
rect 6837 4029 6871 4063
rect 9045 4029 9079 4063
rect 11345 4029 11379 4063
rect 11621 4029 11655 4063
rect 12817 4029 12851 4063
rect 13001 4029 13035 4063
rect 14105 4029 14139 4063
rect 15485 4029 15519 4063
rect 17601 4029 17635 4063
rect 17694 4029 17728 4063
rect 1041 3961 1075 3995
rect 5917 3961 5951 3995
rect 7113 3961 7147 3995
rect 17325 3961 17359 3995
rect 8769 3893 8803 3927
rect 12725 3893 12759 3927
rect 17233 3893 17267 3927
rect 857 3689 891 3723
rect 4537 3689 4571 3723
rect 5457 3689 5491 3723
rect 5917 3689 5951 3723
rect 7573 3689 7607 3723
rect 9965 3689 9999 3723
rect 11161 3689 11195 3723
rect 14749 3689 14783 3723
rect 15209 3689 15243 3723
rect 16037 3689 16071 3723
rect 17601 3689 17635 3723
rect 18245 3689 18279 3723
rect 14381 3621 14415 3655
rect 16497 3621 16531 3655
rect 949 3553 983 3587
rect 4151 3553 4185 3587
rect 4261 3553 4295 3587
rect 4353 3575 4387 3609
rect 5549 3553 5583 3587
rect 5641 3553 5675 3587
rect 7941 3553 7975 3587
rect 10333 3553 10367 3587
rect 11253 3553 11287 3587
rect 11437 3553 11471 3587
rect 15117 3553 15151 3587
rect 16405 3553 16439 3587
rect 17141 3553 17175 3587
rect 17601 3553 17635 3587
rect 17969 3553 18003 3587
rect 18429 3553 18463 3587
rect 5181 3485 5215 3519
rect 8033 3485 8067 3519
rect 8125 3485 8159 3519
rect 10425 3485 10459 3519
rect 10517 3485 10551 3519
rect 15301 3485 15335 3519
rect 16681 3485 16715 3519
rect 17279 3485 17313 3519
rect 10977 3417 11011 3451
rect 5273 3349 5307 3383
rect 17417 3349 17451 3383
rect 5181 3145 5215 3179
rect 7021 3145 7055 3179
rect 10241 3145 10275 3179
rect 11253 3145 11287 3179
rect 12449 3145 12483 3179
rect 14105 3145 14139 3179
rect 15209 3077 15243 3111
rect 2421 3009 2455 3043
rect 7573 3009 7607 3043
rect 9689 3009 9723 3043
rect 9781 3009 9815 3043
rect 11897 3009 11931 3043
rect 13001 3009 13035 3043
rect 13645 3009 13679 3043
rect 2237 2941 2271 2975
rect 5273 2941 5307 2975
rect 12909 2941 12943 2975
rect 13553 2941 13587 2975
rect 13737 2941 13771 2975
rect 14473 2941 14507 2975
rect 14749 2941 14783 2975
rect 14933 2941 14967 2975
rect 15117 2941 15151 2975
rect 15393 2941 15427 2975
rect 7481 2873 7515 2907
rect 1777 2805 1811 2839
rect 2145 2805 2179 2839
rect 7389 2805 7423 2839
rect 9873 2805 9907 2839
rect 11621 2805 11655 2839
rect 11713 2805 11747 2839
rect 12817 2805 12851 2839
rect 1041 2601 1075 2635
rect 1409 2601 1443 2635
rect 2145 2601 2179 2635
rect 2881 2601 2915 2635
rect 3341 2601 3375 2635
rect 5365 2601 5399 2635
rect 8217 2601 8251 2635
rect 8585 2601 8619 2635
rect 15117 2601 15151 2635
rect 15485 2601 15519 2635
rect 1501 2533 1535 2567
rect 8677 2533 8711 2567
rect 12449 2533 12483 2567
rect 14197 2533 14231 2567
rect 17141 2533 17175 2567
rect 18429 2533 18463 2567
rect 2329 2465 2363 2499
rect 3249 2465 3283 2499
rect 5733 2465 5767 2499
rect 17325 2465 17359 2499
rect 17417 2465 17451 2499
rect 17969 2465 18003 2499
rect 1685 2397 1719 2431
rect 3433 2397 3467 2431
rect 5825 2397 5859 2431
rect 6009 2397 6043 2431
rect 8861 2397 8895 2431
rect 14841 2397 14875 2431
rect 15025 2397 15059 2431
rect 17417 2261 17451 2295
rect 3617 2057 3651 2091
rect 6377 2057 6411 2091
rect 7665 2057 7699 2091
rect 9873 2057 9907 2091
rect 10425 2057 10459 2091
rect 11529 2057 11563 2091
rect 13737 2057 13771 2091
rect 14841 2057 14875 2091
rect 15945 2057 15979 2091
rect 5365 1989 5399 2023
rect 3065 1921 3099 1955
rect 6929 1921 6963 1955
rect 8125 1921 8159 1955
rect 8309 1921 8343 1955
rect 8953 1921 8987 1955
rect 10609 1921 10643 1955
rect 12173 1921 12207 1955
rect 13185 1921 13219 1955
rect 14381 1921 14415 1955
rect 16497 1921 16531 1955
rect 17509 1921 17543 1955
rect 3157 1853 3191 1887
rect 3985 1853 4019 1887
rect 4353 1853 4387 1887
rect 4721 1853 4755 1887
rect 5181 1853 5215 1887
rect 5457 1853 5491 1887
rect 6837 1853 6871 1887
rect 9137 1853 9171 1887
rect 9321 1853 9355 1887
rect 9964 1853 9998 1887
rect 10057 1853 10091 1887
rect 10333 1853 10367 1887
rect 11989 1853 12023 1887
rect 12633 1853 12667 1887
rect 12817 1853 12851 1887
rect 13001 1853 13035 1887
rect 14197 1853 14231 1887
rect 10609 1785 10643 1819
rect 16313 1785 16347 1819
rect 17417 1785 17451 1819
rect 18337 1785 18371 1819
rect 3249 1717 3283 1751
rect 4721 1717 4755 1751
rect 5457 1717 5491 1751
rect 6745 1717 6779 1751
rect 8033 1717 8067 1751
rect 9321 1717 9355 1751
rect 11897 1717 11931 1751
rect 14105 1717 14139 1751
rect 16405 1717 16439 1751
rect 16957 1717 16991 1751
rect 17325 1717 17359 1751
rect 3433 1513 3467 1547
rect 5917 1513 5951 1547
rect 7205 1513 7239 1547
rect 9965 1513 9999 1547
rect 11713 1513 11747 1547
rect 12357 1513 12391 1547
rect 17141 1513 17175 1547
rect 17509 1513 17543 1547
rect 18245 1513 18279 1547
rect 8861 1445 8895 1479
rect 10241 1445 10275 1479
rect 11069 1445 11103 1479
rect 14749 1445 14783 1479
rect 17601 1445 17635 1479
rect 3065 1377 3099 1411
rect 5549 1377 5583 1411
rect 5642 1377 5676 1411
rect 6837 1377 6871 1411
rect 8769 1377 8803 1411
rect 9965 1377 9999 1411
rect 10057 1377 10091 1411
rect 10793 1377 10827 1411
rect 11345 1377 11379 1411
rect 11438 1377 11472 1411
rect 13369 1377 13403 1411
rect 14841 1377 14875 1411
rect 16129 1377 16163 1411
rect 18153 1377 18187 1411
rect 3157 1309 3191 1343
rect 6745 1309 6779 1343
rect 11069 1309 11103 1343
rect 13461 1309 13495 1343
rect 16221 1309 16255 1343
rect 17693 1309 17727 1343
rect 13737 1241 13771 1275
rect 16497 1241 16531 1275
rect 10885 1173 10919 1207
rect 5365 969 5399 1003
rect 5457 969 5491 1003
rect 11345 969 11379 1003
rect 17233 969 17267 1003
rect 17969 969 18003 1003
rect 18429 969 18463 1003
rect 11437 901 11471 935
rect 5549 833 5583 867
rect 11621 833 11655 867
rect 5273 765 5307 799
rect 11345 765 11379 799
rect 17785 765 17819 799
<< metal1 >>
rect 184 18522 18860 18544
rect 184 18470 1556 18522
rect 1608 18470 1620 18522
rect 1672 18470 1684 18522
rect 1736 18470 1748 18522
rect 1800 18470 1812 18522
rect 1864 18470 4656 18522
rect 4708 18470 4720 18522
rect 4772 18470 4784 18522
rect 4836 18470 4848 18522
rect 4900 18470 4912 18522
rect 4964 18470 7756 18522
rect 7808 18470 7820 18522
rect 7872 18470 7884 18522
rect 7936 18470 7948 18522
rect 8000 18470 8012 18522
rect 8064 18470 10856 18522
rect 10908 18470 10920 18522
rect 10972 18470 10984 18522
rect 11036 18470 11048 18522
rect 11100 18470 11112 18522
rect 11164 18470 13956 18522
rect 14008 18470 14020 18522
rect 14072 18470 14084 18522
rect 14136 18470 14148 18522
rect 14200 18470 14212 18522
rect 14264 18470 17056 18522
rect 17108 18470 17120 18522
rect 17172 18470 17184 18522
rect 17236 18470 17248 18522
rect 17300 18470 17312 18522
rect 17364 18470 18860 18522
rect 184 18448 18860 18470
rect 2869 18411 2927 18417
rect 2869 18377 2881 18411
rect 2915 18408 2927 18411
rect 4246 18408 4252 18420
rect 2915 18380 4252 18408
rect 2915 18377 2927 18380
rect 2869 18371 2927 18377
rect 4246 18368 4252 18380
rect 4304 18368 4310 18420
rect 18414 18408 18420 18420
rect 18375 18380 18420 18408
rect 18414 18368 18420 18380
rect 18472 18368 18478 18420
rect 2409 18343 2467 18349
rect 2409 18309 2421 18343
rect 2455 18340 2467 18343
rect 5810 18340 5816 18352
rect 2455 18312 5816 18340
rect 2455 18309 2467 18312
rect 2409 18303 2467 18309
rect 5810 18300 5816 18312
rect 5868 18300 5874 18352
rect 5997 18343 6055 18349
rect 5997 18309 6009 18343
rect 6043 18340 6055 18343
rect 9858 18340 9864 18352
rect 6043 18312 9864 18340
rect 6043 18309 6055 18312
rect 5997 18303 6055 18309
rect 9858 18300 9864 18312
rect 9916 18300 9922 18352
rect 5445 18275 5503 18281
rect 5445 18241 5457 18275
rect 5491 18272 5503 18275
rect 5718 18272 5724 18284
rect 5491 18244 5724 18272
rect 5491 18241 5503 18244
rect 5445 18235 5503 18241
rect 5718 18232 5724 18244
rect 5776 18232 5782 18284
rect 8202 18272 8208 18284
rect 8163 18244 8208 18272
rect 8202 18232 8208 18244
rect 8260 18272 8266 18284
rect 10505 18275 10563 18281
rect 10505 18272 10517 18275
rect 8260 18244 10517 18272
rect 8260 18232 8266 18244
rect 10505 18241 10517 18244
rect 10551 18241 10563 18275
rect 12986 18272 12992 18284
rect 10505 18235 10563 18241
rect 12728 18244 12992 18272
rect 845 18207 903 18213
rect 845 18173 857 18207
rect 891 18204 903 18207
rect 1394 18204 1400 18216
rect 891 18176 1400 18204
rect 891 18173 903 18176
rect 845 18167 903 18173
rect 1394 18164 1400 18176
rect 1452 18204 1458 18216
rect 1581 18207 1639 18213
rect 1581 18204 1593 18207
rect 1452 18176 1593 18204
rect 1452 18164 1458 18176
rect 1581 18173 1593 18176
rect 1627 18173 1639 18207
rect 3605 18207 3663 18213
rect 3605 18204 3617 18207
rect 1581 18167 1639 18173
rect 2792 18176 3617 18204
rect 2792 18148 2820 18176
rect 3605 18173 3617 18176
rect 3651 18173 3663 18207
rect 3970 18204 3976 18216
rect 3931 18176 3976 18204
rect 3605 18167 3663 18173
rect 1213 18139 1271 18145
rect 1213 18105 1225 18139
rect 1259 18136 1271 18139
rect 2774 18136 2780 18148
rect 1259 18108 2780 18136
rect 1259 18105 1271 18108
rect 1213 18099 1271 18105
rect 2774 18096 2780 18108
rect 2832 18096 2838 18148
rect 2866 18096 2872 18148
rect 2924 18136 2930 18148
rect 3329 18139 3387 18145
rect 3329 18136 3341 18139
rect 2924 18108 3341 18136
rect 2924 18096 2930 18108
rect 3329 18105 3341 18108
rect 3375 18105 3387 18139
rect 3620 18136 3648 18167
rect 3970 18164 3976 18176
rect 4028 18164 4034 18216
rect 4154 18204 4160 18216
rect 4115 18176 4160 18204
rect 4154 18164 4160 18176
rect 4212 18164 4218 18216
rect 4522 18204 4528 18216
rect 4483 18176 4528 18204
rect 4522 18164 4528 18176
rect 4580 18164 4586 18216
rect 6733 18207 6791 18213
rect 6733 18173 6745 18207
rect 6779 18173 6791 18207
rect 6733 18167 6791 18173
rect 3878 18136 3884 18148
rect 3620 18108 3884 18136
rect 3329 18099 3387 18105
rect 3878 18096 3884 18108
rect 3936 18136 3942 18148
rect 6365 18139 6423 18145
rect 6365 18136 6377 18139
rect 3936 18108 6377 18136
rect 3936 18096 3942 18108
rect 6365 18105 6377 18108
rect 6411 18136 6423 18139
rect 6748 18136 6776 18167
rect 6822 18164 6828 18216
rect 6880 18204 6886 18216
rect 7929 18207 7987 18213
rect 7929 18204 7941 18207
rect 6880 18176 7941 18204
rect 6880 18164 6886 18176
rect 7929 18173 7941 18176
rect 7975 18173 7987 18207
rect 8754 18204 8760 18216
rect 8715 18176 8760 18204
rect 7929 18167 7987 18173
rect 8754 18164 8760 18176
rect 8812 18164 8818 18216
rect 11330 18164 11336 18216
rect 11388 18204 11394 18216
rect 12728 18213 12756 18244
rect 12986 18232 12992 18244
rect 13044 18232 13050 18284
rect 11701 18207 11759 18213
rect 11701 18204 11713 18207
rect 11388 18176 11713 18204
rect 11388 18164 11394 18176
rect 11701 18173 11713 18176
rect 11747 18173 11759 18207
rect 11701 18167 11759 18173
rect 12713 18207 12771 18213
rect 12713 18173 12725 18207
rect 12759 18173 12771 18207
rect 12894 18204 12900 18216
rect 12855 18176 12900 18204
rect 12713 18167 12771 18173
rect 12894 18164 12900 18176
rect 12952 18164 12958 18216
rect 14185 18207 14243 18213
rect 14185 18173 14197 18207
rect 14231 18204 14243 18207
rect 14366 18204 14372 18216
rect 14231 18176 14372 18204
rect 14231 18173 14243 18176
rect 14185 18167 14243 18173
rect 14366 18164 14372 18176
rect 14424 18164 14430 18216
rect 14918 18204 14924 18216
rect 14879 18176 14924 18204
rect 14918 18164 14924 18176
rect 14976 18164 14982 18216
rect 16577 18207 16635 18213
rect 16577 18173 16589 18207
rect 16623 18204 16635 18207
rect 16666 18204 16672 18216
rect 16623 18176 16672 18204
rect 16623 18173 16635 18176
rect 16577 18167 16635 18173
rect 16666 18164 16672 18176
rect 16724 18164 16730 18216
rect 17957 18207 18015 18213
rect 17957 18173 17969 18207
rect 18003 18204 18015 18207
rect 18414 18204 18420 18216
rect 18003 18176 18420 18204
rect 18003 18173 18015 18176
rect 17957 18167 18015 18173
rect 18414 18164 18420 18176
rect 18472 18164 18478 18216
rect 6411 18108 6776 18136
rect 7009 18139 7067 18145
rect 6411 18105 6423 18108
rect 6365 18099 6423 18105
rect 7009 18105 7021 18139
rect 7055 18136 7067 18139
rect 9214 18136 9220 18148
rect 7055 18108 9220 18136
rect 7055 18105 7067 18108
rect 7009 18099 7067 18105
rect 9214 18096 9220 18108
rect 9272 18096 9278 18148
rect 10413 18139 10471 18145
rect 10413 18105 10425 18139
rect 10459 18136 10471 18139
rect 13814 18136 13820 18148
rect 10459 18108 13820 18136
rect 10459 18105 10471 18108
rect 10413 18099 10471 18105
rect 13814 18096 13820 18108
rect 13872 18096 13878 18148
rect 13909 18139 13967 18145
rect 13909 18105 13921 18139
rect 13955 18136 13967 18139
rect 14642 18136 14648 18148
rect 13955 18108 14648 18136
rect 13955 18105 13967 18108
rect 13909 18099 13967 18105
rect 14642 18096 14648 18108
rect 14700 18096 14706 18148
rect 14826 18136 14832 18148
rect 14787 18108 14832 18136
rect 14826 18096 14832 18108
rect 14884 18096 14890 18148
rect 1765 18071 1823 18077
rect 1765 18037 1777 18071
rect 1811 18068 1823 18071
rect 2498 18068 2504 18080
rect 1811 18040 2504 18068
rect 1811 18037 1823 18040
rect 1765 18031 1823 18037
rect 2498 18028 2504 18040
rect 2556 18028 2562 18080
rect 4430 18068 4436 18080
rect 4391 18040 4436 18068
rect 4430 18028 4436 18040
rect 4488 18028 4494 18080
rect 5534 18068 5540 18080
rect 5495 18040 5540 18068
rect 5534 18028 5540 18040
rect 5592 18028 5598 18080
rect 5626 18028 5632 18080
rect 5684 18068 5690 18080
rect 7558 18068 7564 18080
rect 5684 18040 5729 18068
rect 7519 18040 7564 18068
rect 5684 18028 5690 18040
rect 7558 18028 7564 18040
rect 7616 18028 7622 18080
rect 8021 18071 8079 18077
rect 8021 18037 8033 18071
rect 8067 18068 8079 18071
rect 8110 18068 8116 18080
rect 8067 18040 8116 18068
rect 8067 18037 8079 18040
rect 8021 18031 8079 18037
rect 8110 18028 8116 18040
rect 8168 18028 8174 18080
rect 9122 18028 9128 18080
rect 9180 18068 9186 18080
rect 9401 18071 9459 18077
rect 9401 18068 9413 18071
rect 9180 18040 9413 18068
rect 9180 18028 9186 18040
rect 9401 18037 9413 18040
rect 9447 18037 9459 18071
rect 9950 18068 9956 18080
rect 9911 18040 9956 18068
rect 9401 18031 9459 18037
rect 9950 18028 9956 18040
rect 10008 18028 10014 18080
rect 10318 18068 10324 18080
rect 10279 18040 10324 18068
rect 10318 18028 10324 18040
rect 10376 18028 10382 18080
rect 11149 18071 11207 18077
rect 11149 18037 11161 18071
rect 11195 18068 11207 18071
rect 11238 18068 11244 18080
rect 11195 18040 11244 18068
rect 11195 18037 11207 18040
rect 11149 18031 11207 18037
rect 11238 18028 11244 18040
rect 11296 18028 11302 18080
rect 13262 18028 13268 18080
rect 13320 18068 13326 18080
rect 15473 18071 15531 18077
rect 15473 18068 15485 18071
rect 13320 18040 15485 18068
rect 13320 18028 13326 18040
rect 15473 18037 15485 18040
rect 15519 18037 15531 18071
rect 15930 18068 15936 18080
rect 15891 18040 15936 18068
rect 15473 18031 15531 18037
rect 15930 18028 15936 18040
rect 15988 18028 15994 18080
rect 16574 18028 16580 18080
rect 16632 18068 16638 18080
rect 17773 18071 17831 18077
rect 17773 18068 17785 18071
rect 16632 18040 17785 18068
rect 16632 18028 16638 18040
rect 17773 18037 17785 18040
rect 17819 18037 17831 18071
rect 17773 18031 17831 18037
rect 184 17978 18920 18000
rect 184 17926 3106 17978
rect 3158 17926 3170 17978
rect 3222 17926 3234 17978
rect 3286 17926 3298 17978
rect 3350 17926 3362 17978
rect 3414 17926 6206 17978
rect 6258 17926 6270 17978
rect 6322 17926 6334 17978
rect 6386 17926 6398 17978
rect 6450 17926 6462 17978
rect 6514 17926 9306 17978
rect 9358 17926 9370 17978
rect 9422 17926 9434 17978
rect 9486 17926 9498 17978
rect 9550 17926 9562 17978
rect 9614 17926 12406 17978
rect 12458 17926 12470 17978
rect 12522 17926 12534 17978
rect 12586 17926 12598 17978
rect 12650 17926 12662 17978
rect 12714 17926 15506 17978
rect 15558 17926 15570 17978
rect 15622 17926 15634 17978
rect 15686 17926 15698 17978
rect 15750 17926 15762 17978
rect 15814 17926 18606 17978
rect 18658 17926 18670 17978
rect 18722 17926 18734 17978
rect 18786 17926 18798 17978
rect 18850 17926 18862 17978
rect 18914 17926 18920 17978
rect 184 17904 18920 17926
rect 3050 17824 3056 17876
rect 3108 17864 3114 17876
rect 3421 17867 3479 17873
rect 3421 17864 3433 17867
rect 3108 17836 3433 17864
rect 3108 17824 3114 17836
rect 3421 17833 3433 17836
rect 3467 17864 3479 17867
rect 3970 17864 3976 17876
rect 3467 17836 3976 17864
rect 3467 17833 3479 17836
rect 3421 17827 3479 17833
rect 3970 17824 3976 17836
rect 4028 17824 4034 17876
rect 13630 17824 13636 17876
rect 13688 17864 13694 17876
rect 13688 17836 16252 17864
rect 13688 17824 13694 17836
rect 2406 17796 2412 17808
rect 2070 17768 2412 17796
rect 2406 17756 2412 17768
rect 2464 17796 2470 17808
rect 4154 17796 4160 17808
rect 2464 17768 4160 17796
rect 2464 17756 2470 17768
rect 4154 17756 4160 17768
rect 4212 17756 4218 17808
rect 4430 17756 4436 17808
rect 4488 17796 4494 17808
rect 4534 17799 4592 17805
rect 4534 17796 4546 17799
rect 4488 17768 4546 17796
rect 4488 17756 4494 17768
rect 4534 17765 4546 17768
rect 4580 17765 4592 17799
rect 4534 17759 4592 17765
rect 7558 17756 7564 17808
rect 7616 17796 7622 17808
rect 7837 17799 7895 17805
rect 7837 17796 7849 17799
rect 7616 17768 7849 17796
rect 7616 17756 7622 17768
rect 7837 17765 7849 17768
rect 7883 17765 7895 17799
rect 7837 17759 7895 17765
rect 9858 17756 9864 17808
rect 9916 17796 9922 17808
rect 9953 17799 10011 17805
rect 9953 17796 9965 17799
rect 9916 17768 9965 17796
rect 9916 17756 9922 17768
rect 9953 17765 9965 17768
rect 9999 17765 10011 17799
rect 13648 17796 13676 17824
rect 9953 17759 10011 17765
rect 12636 17768 13676 17796
rect 2682 17688 2688 17740
rect 2740 17728 2746 17740
rect 2869 17731 2927 17737
rect 2869 17728 2881 17731
rect 2740 17700 2881 17728
rect 2740 17688 2746 17700
rect 2869 17697 2881 17700
rect 2915 17697 2927 17731
rect 2869 17691 2927 17697
rect 4246 17688 4252 17740
rect 4304 17728 4310 17740
rect 5169 17731 5227 17737
rect 5169 17728 5181 17731
rect 4304 17700 5181 17728
rect 4304 17688 4310 17700
rect 5169 17697 5181 17700
rect 5215 17697 5227 17731
rect 5169 17691 5227 17697
rect 12434 17688 12440 17740
rect 12492 17728 12498 17740
rect 12636 17737 12664 17768
rect 16114 17756 16120 17808
rect 16172 17756 16178 17808
rect 16224 17796 16252 17836
rect 16531 17799 16589 17805
rect 16531 17796 16543 17799
rect 16224 17768 16543 17796
rect 16531 17765 16543 17768
rect 16577 17796 16589 17799
rect 17405 17799 17463 17805
rect 17405 17796 17417 17799
rect 16577 17768 17417 17796
rect 16577 17765 16589 17768
rect 16531 17759 16589 17765
rect 17405 17765 17417 17768
rect 17451 17765 17463 17799
rect 17405 17759 17463 17765
rect 12621 17731 12679 17737
rect 12621 17728 12633 17731
rect 12492 17700 12633 17728
rect 12492 17688 12498 17700
rect 12621 17697 12633 17700
rect 12667 17697 12679 17731
rect 12894 17728 12900 17740
rect 12855 17700 12900 17728
rect 12621 17691 12679 17697
rect 12894 17688 12900 17700
rect 12952 17688 12958 17740
rect 14737 17731 14795 17737
rect 14737 17697 14749 17731
rect 14783 17728 14795 17731
rect 14826 17728 14832 17740
rect 14783 17700 14832 17728
rect 14783 17697 14795 17700
rect 14737 17691 14795 17697
rect 14826 17688 14832 17700
rect 14884 17688 14890 17740
rect 16132 17728 16160 17756
rect 16758 17728 16764 17740
rect 16132 17700 16764 17728
rect 16758 17688 16764 17700
rect 16816 17688 16822 17740
rect 17129 17731 17187 17737
rect 17129 17697 17141 17731
rect 17175 17697 17187 17731
rect 17129 17691 17187 17697
rect 566 17660 572 17672
rect 527 17632 572 17660
rect 566 17620 572 17632
rect 624 17620 630 17672
rect 842 17660 848 17672
rect 803 17632 848 17660
rect 842 17620 848 17632
rect 900 17620 906 17672
rect 4801 17663 4859 17669
rect 4801 17629 4813 17663
rect 4847 17629 4859 17663
rect 4801 17623 4859 17629
rect 12345 17663 12403 17669
rect 12345 17629 12357 17663
rect 12391 17629 12403 17663
rect 12345 17623 12403 17629
rect 12529 17663 12587 17669
rect 12529 17629 12541 17663
rect 12575 17660 12587 17663
rect 12575 17632 12756 17660
rect 12575 17629 12587 17632
rect 12529 17623 12587 17629
rect 2774 17552 2780 17604
rect 2832 17592 2838 17604
rect 3053 17595 3111 17601
rect 3053 17592 3065 17595
rect 2832 17564 3065 17592
rect 2832 17552 2838 17564
rect 3053 17561 3065 17564
rect 3099 17561 3111 17595
rect 4816 17592 4844 17623
rect 5166 17592 5172 17604
rect 4816 17564 5172 17592
rect 3053 17555 3111 17561
rect 5166 17552 5172 17564
rect 5224 17552 5230 17604
rect 9214 17552 9220 17604
rect 9272 17592 9278 17604
rect 11514 17592 11520 17604
rect 9272 17564 11520 17592
rect 9272 17552 9278 17564
rect 11514 17552 11520 17564
rect 11572 17552 11578 17604
rect 11974 17552 11980 17604
rect 12032 17592 12038 17604
rect 12360 17592 12388 17623
rect 12728 17592 12756 17632
rect 12802 17620 12808 17672
rect 12860 17660 12866 17672
rect 13357 17663 13415 17669
rect 13357 17660 13369 17663
rect 12860 17632 13369 17660
rect 12860 17620 12866 17632
rect 13357 17629 13369 17632
rect 13403 17629 13415 17663
rect 15102 17660 15108 17672
rect 15063 17632 15108 17660
rect 13357 17623 13415 17629
rect 15102 17620 15108 17632
rect 15160 17620 15166 17672
rect 17144 17660 17172 17691
rect 15856 17632 17172 17660
rect 13078 17592 13084 17604
rect 12032 17564 12572 17592
rect 12728 17564 13084 17592
rect 12032 17552 12038 17564
rect 2038 17484 2044 17536
rect 2096 17524 2102 17536
rect 2317 17527 2375 17533
rect 2317 17524 2329 17527
rect 2096 17496 2329 17524
rect 2096 17484 2102 17496
rect 2317 17493 2329 17496
rect 2363 17493 2375 17527
rect 2317 17487 2375 17493
rect 4430 17484 4436 17536
rect 4488 17524 4494 17536
rect 6457 17527 6515 17533
rect 6457 17524 6469 17527
rect 4488 17496 6469 17524
rect 4488 17484 4494 17496
rect 6457 17493 6469 17496
rect 6503 17493 6515 17527
rect 6457 17487 6515 17493
rect 7006 17484 7012 17536
rect 7064 17524 7070 17536
rect 9125 17527 9183 17533
rect 9125 17524 9137 17527
rect 7064 17496 9137 17524
rect 7064 17484 7070 17496
rect 9125 17493 9137 17496
rect 9171 17493 9183 17527
rect 11422 17524 11428 17536
rect 11383 17496 11428 17524
rect 9125 17487 9183 17493
rect 11422 17484 11428 17496
rect 11480 17484 11486 17536
rect 11882 17484 11888 17536
rect 11940 17524 11946 17536
rect 12437 17527 12495 17533
rect 12437 17524 12449 17527
rect 11940 17496 12449 17524
rect 11940 17484 11946 17496
rect 12437 17493 12449 17496
rect 12483 17493 12495 17527
rect 12544 17524 12572 17564
rect 13078 17552 13084 17564
rect 13136 17552 13142 17604
rect 12710 17524 12716 17536
rect 12544 17496 12716 17524
rect 12437 17487 12495 17493
rect 12710 17484 12716 17496
rect 12768 17524 12774 17536
rect 15856 17524 15884 17632
rect 16298 17552 16304 17604
rect 16356 17592 16362 17604
rect 17221 17595 17279 17601
rect 17221 17592 17233 17595
rect 16356 17564 17233 17592
rect 16356 17552 16362 17564
rect 17221 17561 17233 17564
rect 17267 17561 17279 17595
rect 17221 17555 17279 17561
rect 12768 17496 15884 17524
rect 12768 17484 12774 17496
rect 16850 17484 16856 17536
rect 16908 17524 16914 17536
rect 17129 17527 17187 17533
rect 17129 17524 17141 17527
rect 16908 17496 17141 17524
rect 16908 17484 16914 17496
rect 17129 17493 17141 17496
rect 17175 17493 17187 17527
rect 17129 17487 17187 17493
rect 184 17434 18860 17456
rect 184 17382 1556 17434
rect 1608 17382 1620 17434
rect 1672 17382 1684 17434
rect 1736 17382 1748 17434
rect 1800 17382 1812 17434
rect 1864 17382 4656 17434
rect 4708 17382 4720 17434
rect 4772 17382 4784 17434
rect 4836 17382 4848 17434
rect 4900 17382 4912 17434
rect 4964 17382 7756 17434
rect 7808 17382 7820 17434
rect 7872 17382 7884 17434
rect 7936 17382 7948 17434
rect 8000 17382 8012 17434
rect 8064 17382 10856 17434
rect 10908 17382 10920 17434
rect 10972 17382 10984 17434
rect 11036 17382 11048 17434
rect 11100 17382 11112 17434
rect 11164 17382 13956 17434
rect 14008 17382 14020 17434
rect 14072 17382 14084 17434
rect 14136 17382 14148 17434
rect 14200 17382 14212 17434
rect 14264 17382 17056 17434
rect 17108 17382 17120 17434
rect 17172 17382 17184 17434
rect 17236 17382 17248 17434
rect 17300 17382 17312 17434
rect 17364 17382 18860 17434
rect 184 17360 18860 17382
rect 1394 17280 1400 17332
rect 1452 17320 1458 17332
rect 2501 17323 2559 17329
rect 2501 17320 2513 17323
rect 1452 17292 2513 17320
rect 1452 17280 1458 17292
rect 2501 17289 2513 17292
rect 2547 17289 2559 17323
rect 2682 17320 2688 17332
rect 2643 17292 2688 17320
rect 2501 17283 2559 17289
rect 842 17252 848 17264
rect 803 17224 848 17252
rect 842 17212 848 17224
rect 900 17212 906 17264
rect 2516 17252 2544 17283
rect 2682 17280 2688 17292
rect 2740 17280 2746 17332
rect 5537 17323 5595 17329
rect 5537 17289 5549 17323
rect 5583 17320 5595 17323
rect 5626 17320 5632 17332
rect 5583 17292 5632 17320
rect 5583 17289 5595 17292
rect 5537 17283 5595 17289
rect 5626 17280 5632 17292
rect 5684 17280 5690 17332
rect 8251 17323 8309 17329
rect 8251 17289 8263 17323
rect 8297 17320 8309 17323
rect 8754 17320 8760 17332
rect 8297 17292 8760 17320
rect 8297 17289 8309 17292
rect 8251 17283 8309 17289
rect 8754 17280 8760 17292
rect 8812 17280 8818 17332
rect 12986 17320 12992 17332
rect 9508 17292 12992 17320
rect 2590 17252 2596 17264
rect 2516 17224 2596 17252
rect 2590 17212 2596 17224
rect 2648 17212 2654 17264
rect 3050 17184 3056 17196
rect 3011 17156 3056 17184
rect 3050 17144 3056 17156
rect 3108 17144 3114 17196
rect 5810 17144 5816 17196
rect 5868 17184 5874 17196
rect 6825 17187 6883 17193
rect 6825 17184 6837 17187
rect 5868 17156 6837 17184
rect 5868 17144 5874 17156
rect 6825 17153 6837 17156
rect 6871 17153 6883 17187
rect 6825 17147 6883 17153
rect 8803 17187 8861 17193
rect 8803 17153 8815 17187
rect 8849 17184 8861 17187
rect 9508 17184 9536 17292
rect 12986 17280 12992 17292
rect 13044 17280 13050 17332
rect 13170 17280 13176 17332
rect 13228 17320 13234 17332
rect 15565 17323 15623 17329
rect 13228 17292 15240 17320
rect 13228 17280 13234 17292
rect 12069 17255 12127 17261
rect 12069 17221 12081 17255
rect 12115 17252 12127 17255
rect 12802 17252 12808 17264
rect 12115 17224 12808 17252
rect 12115 17221 12127 17224
rect 12069 17215 12127 17221
rect 12802 17212 12808 17224
rect 12860 17212 12866 17264
rect 12894 17212 12900 17264
rect 12952 17252 12958 17264
rect 13446 17252 13452 17264
rect 12952 17224 13452 17252
rect 12952 17212 12958 17224
rect 13446 17212 13452 17224
rect 13504 17212 13510 17264
rect 8849 17156 9536 17184
rect 10229 17187 10287 17193
rect 8849 17153 8861 17156
rect 8803 17147 8861 17153
rect 10229 17153 10241 17187
rect 10275 17184 10287 17187
rect 11238 17184 11244 17196
rect 10275 17156 11244 17184
rect 10275 17153 10287 17156
rect 10229 17147 10287 17153
rect 11238 17144 11244 17156
rect 11296 17144 11302 17196
rect 11517 17187 11575 17193
rect 11517 17153 11529 17187
rect 11563 17184 11575 17187
rect 13814 17184 13820 17196
rect 11563 17156 13032 17184
rect 13775 17156 13820 17184
rect 11563 17153 11575 17156
rect 11517 17147 11575 17153
rect 1118 17116 1124 17128
rect 1079 17088 1124 17116
rect 1118 17076 1124 17088
rect 1176 17076 1182 17128
rect 1210 17076 1216 17128
rect 1268 17116 1274 17128
rect 2133 17119 2191 17125
rect 1268 17088 1313 17116
rect 1268 17076 1274 17088
rect 2133 17085 2145 17119
rect 2179 17085 2191 17119
rect 2133 17079 2191 17085
rect 2148 17048 2176 17079
rect 2406 17076 2412 17128
rect 2464 17116 2470 17128
rect 2682 17116 2688 17128
rect 2464 17088 2688 17116
rect 2464 17076 2470 17088
rect 2682 17076 2688 17088
rect 2740 17076 2746 17128
rect 4249 17119 4307 17125
rect 4249 17085 4261 17119
rect 4295 17116 4307 17119
rect 4430 17116 4436 17128
rect 4295 17088 4436 17116
rect 4295 17085 4307 17088
rect 4249 17079 4307 17085
rect 4430 17076 4436 17088
rect 4488 17076 4494 17128
rect 5902 17076 5908 17128
rect 5960 17116 5966 17128
rect 6457 17119 6515 17125
rect 6457 17116 6469 17119
rect 5960 17088 6469 17116
rect 5960 17076 5966 17088
rect 6457 17085 6469 17088
rect 6503 17085 6515 17119
rect 6457 17079 6515 17085
rect 10597 17119 10655 17125
rect 10597 17085 10609 17119
rect 10643 17085 10655 17119
rect 10597 17079 10655 17085
rect 4798 17048 4804 17060
rect 2148 17020 4804 17048
rect 4798 17008 4804 17020
rect 4856 17008 4862 17060
rect 7374 17008 7380 17060
rect 7432 17008 7438 17060
rect 9214 17008 9220 17060
rect 9272 17008 9278 17060
rect 10612 17048 10640 17079
rect 12434 17076 12440 17128
rect 12492 17116 12498 17128
rect 12710 17116 12716 17128
rect 12492 17088 12537 17116
rect 12671 17088 12716 17116
rect 12492 17076 12498 17088
rect 12710 17076 12716 17088
rect 12768 17076 12774 17128
rect 12894 17048 12900 17060
rect 10612 17020 12900 17048
rect 12894 17008 12900 17020
rect 12952 17008 12958 17060
rect 2498 16980 2504 16992
rect 2459 16952 2504 16980
rect 2498 16940 2504 16952
rect 2556 16940 2562 16992
rect 3605 16983 3663 16989
rect 3605 16949 3617 16983
rect 3651 16980 3663 16983
rect 4338 16980 4344 16992
rect 3651 16952 4344 16980
rect 3651 16949 3663 16952
rect 3605 16943 3663 16949
rect 4338 16940 4344 16952
rect 4396 16940 4402 16992
rect 11606 16980 11612 16992
rect 11567 16952 11612 16980
rect 11606 16940 11612 16952
rect 11664 16940 11670 16992
rect 11698 16940 11704 16992
rect 11756 16980 11762 16992
rect 12621 16983 12679 16989
rect 11756 16952 11801 16980
rect 11756 16940 11762 16952
rect 12621 16949 12633 16983
rect 12667 16980 12679 16983
rect 13004 16980 13032 17156
rect 13814 17144 13820 17156
rect 13872 17144 13878 17196
rect 13078 17076 13084 17128
rect 13136 17116 13142 17128
rect 13173 17119 13231 17125
rect 13173 17116 13185 17119
rect 13136 17088 13185 17116
rect 13136 17076 13142 17088
rect 13173 17085 13185 17088
rect 13219 17116 13231 17119
rect 13354 17116 13360 17128
rect 13219 17088 13360 17116
rect 13219 17085 13231 17088
rect 13173 17079 13231 17085
rect 13354 17076 13360 17088
rect 13412 17076 13418 17128
rect 15212 17116 15240 17292
rect 15565 17289 15577 17323
rect 15611 17320 15623 17323
rect 16666 17320 16672 17332
rect 15611 17292 16672 17320
rect 15611 17289 15623 17292
rect 15565 17283 15623 17289
rect 16666 17280 16672 17292
rect 16724 17280 16730 17332
rect 16485 17187 16543 17193
rect 16485 17153 16497 17187
rect 16531 17184 16543 17187
rect 18230 17184 18236 17196
rect 16531 17156 18236 17184
rect 16531 17153 16543 17156
rect 16485 17147 16543 17153
rect 18230 17144 18236 17156
rect 18288 17144 18294 17196
rect 16022 17116 16028 17128
rect 15212 17102 16028 17116
rect 15226 17088 16028 17102
rect 16022 17076 16028 17088
rect 16080 17076 16086 17128
rect 16117 17119 16175 17125
rect 16117 17085 16129 17119
rect 16163 17116 16175 17119
rect 16206 17116 16212 17128
rect 16163 17088 16212 17116
rect 16163 17085 16175 17088
rect 16117 17079 16175 17085
rect 16206 17076 16212 17088
rect 16264 17076 16270 17128
rect 14090 17048 14096 17060
rect 14051 17020 14096 17048
rect 14090 17008 14096 17020
rect 14148 17008 14154 17060
rect 17494 17008 17500 17060
rect 17552 17008 17558 17060
rect 13722 16980 13728 16992
rect 12667 16952 13728 16980
rect 12667 16949 12679 16952
rect 12621 16943 12679 16949
rect 13722 16940 13728 16952
rect 13780 16940 13786 16992
rect 13998 16940 14004 16992
rect 14056 16980 14062 16992
rect 16574 16980 16580 16992
rect 14056 16952 16580 16980
rect 14056 16940 14062 16952
rect 16574 16940 16580 16952
rect 16632 16940 16638 16992
rect 17770 16940 17776 16992
rect 17828 16980 17834 16992
rect 17911 16983 17969 16989
rect 17911 16980 17923 16983
rect 17828 16952 17923 16980
rect 17828 16940 17834 16952
rect 17911 16949 17923 16952
rect 17957 16949 17969 16983
rect 17911 16943 17969 16949
rect 184 16890 18920 16912
rect 184 16838 3106 16890
rect 3158 16838 3170 16890
rect 3222 16838 3234 16890
rect 3286 16838 3298 16890
rect 3350 16838 3362 16890
rect 3414 16838 6206 16890
rect 6258 16838 6270 16890
rect 6322 16838 6334 16890
rect 6386 16838 6398 16890
rect 6450 16838 6462 16890
rect 6514 16838 9306 16890
rect 9358 16838 9370 16890
rect 9422 16838 9434 16890
rect 9486 16838 9498 16890
rect 9550 16838 9562 16890
rect 9614 16838 12406 16890
rect 12458 16838 12470 16890
rect 12522 16838 12534 16890
rect 12586 16838 12598 16890
rect 12650 16838 12662 16890
rect 12714 16838 15506 16890
rect 15558 16838 15570 16890
rect 15622 16838 15634 16890
rect 15686 16838 15698 16890
rect 15750 16838 15762 16890
rect 15814 16838 18606 16890
rect 18658 16838 18670 16890
rect 18722 16838 18734 16890
rect 18786 16838 18798 16890
rect 18850 16838 18862 16890
rect 18914 16838 18920 16890
rect 184 16816 18920 16838
rect 1210 16736 1216 16788
rect 1268 16776 1274 16788
rect 2133 16779 2191 16785
rect 2133 16776 2145 16779
rect 1268 16748 2145 16776
rect 1268 16736 1274 16748
rect 2133 16745 2145 16748
rect 2179 16745 2191 16779
rect 2133 16739 2191 16745
rect 2498 16736 2504 16788
rect 2556 16776 2562 16788
rect 4249 16779 4307 16785
rect 4249 16776 4261 16779
rect 2556 16748 4261 16776
rect 2556 16736 2562 16748
rect 4249 16745 4261 16748
rect 4295 16745 4307 16779
rect 4249 16739 4307 16745
rect 7791 16779 7849 16785
rect 7791 16745 7803 16779
rect 7837 16776 7849 16779
rect 11330 16776 11336 16788
rect 7837 16748 11336 16776
rect 7837 16745 7849 16748
rect 7791 16739 7849 16745
rect 11330 16736 11336 16748
rect 11388 16736 11394 16788
rect 11606 16736 11612 16788
rect 11664 16776 11670 16788
rect 12710 16776 12716 16788
rect 11664 16748 12716 16776
rect 11664 16736 11670 16748
rect 12710 16736 12716 16748
rect 12768 16736 12774 16788
rect 13998 16776 14004 16788
rect 12820 16748 14004 16776
rect 1118 16668 1124 16720
rect 1176 16708 1182 16720
rect 1397 16711 1455 16717
rect 1397 16708 1409 16711
rect 1176 16680 1409 16708
rect 1176 16668 1182 16680
rect 1397 16677 1409 16680
rect 1443 16677 1455 16711
rect 1397 16671 1455 16677
rect 1780 16680 2452 16708
rect 1780 16649 1808 16680
rect 2148 16652 2176 16680
rect 1305 16643 1363 16649
rect 1305 16609 1317 16643
rect 1351 16640 1363 16643
rect 1765 16643 1823 16649
rect 1351 16612 1716 16640
rect 1351 16609 1363 16612
rect 1305 16603 1363 16609
rect 1688 16572 1716 16612
rect 1765 16609 1777 16643
rect 1811 16609 1823 16643
rect 2038 16640 2044 16652
rect 1765 16603 1823 16609
rect 1872 16612 2044 16640
rect 1872 16572 1900 16612
rect 2038 16600 2044 16612
rect 2096 16600 2102 16652
rect 2130 16600 2136 16652
rect 2188 16600 2194 16652
rect 2424 16581 2452 16680
rect 2590 16668 2596 16720
rect 2648 16708 2654 16720
rect 4157 16711 4215 16717
rect 4157 16708 4169 16711
rect 2648 16680 4169 16708
rect 2648 16668 2654 16680
rect 4157 16677 4169 16680
rect 4203 16677 4215 16711
rect 5626 16708 5632 16720
rect 4157 16671 4215 16677
rect 4632 16680 5632 16708
rect 2682 16600 2688 16652
rect 2740 16640 2746 16652
rect 2740 16612 2820 16640
rect 2740 16600 2746 16612
rect 1688 16544 1900 16572
rect 2409 16575 2467 16581
rect 2409 16541 2421 16575
rect 2455 16541 2467 16575
rect 2792 16572 2820 16612
rect 2866 16600 2872 16652
rect 2924 16640 2930 16652
rect 3237 16643 3295 16649
rect 3237 16640 3249 16643
rect 2924 16612 3249 16640
rect 2924 16600 2930 16612
rect 3237 16609 3249 16612
rect 3283 16609 3295 16643
rect 3513 16643 3571 16649
rect 3513 16640 3525 16643
rect 3237 16603 3295 16609
rect 3344 16612 3525 16640
rect 3344 16572 3372 16612
rect 3513 16609 3525 16612
rect 3559 16640 3571 16643
rect 4062 16640 4068 16652
rect 3559 16612 3924 16640
rect 4023 16612 4068 16640
rect 3559 16609 3571 16612
rect 3513 16603 3571 16609
rect 2792 16544 3372 16572
rect 3896 16572 3924 16612
rect 4062 16600 4068 16612
rect 4120 16600 4126 16652
rect 4632 16640 4660 16680
rect 5626 16668 5632 16680
rect 5684 16668 5690 16720
rect 7006 16708 7012 16720
rect 6967 16680 7012 16708
rect 7006 16668 7012 16680
rect 7064 16668 7070 16720
rect 7466 16668 7472 16720
rect 7524 16708 7530 16720
rect 12820 16708 12848 16748
rect 13998 16736 14004 16748
rect 14056 16736 14062 16788
rect 14090 16736 14096 16788
rect 14148 16776 14154 16788
rect 18233 16779 18291 16785
rect 18233 16776 18245 16779
rect 14148 16748 18245 16776
rect 14148 16736 14154 16748
rect 18233 16745 18245 16748
rect 18279 16745 18291 16779
rect 18233 16739 18291 16745
rect 7524 16680 8234 16708
rect 9508 16680 12848 16708
rect 13188 16680 13584 16708
rect 7524 16668 7530 16680
rect 4798 16640 4804 16652
rect 4172 16612 4660 16640
rect 4711 16612 4804 16640
rect 4172 16572 4200 16612
rect 4798 16600 4804 16612
rect 4856 16640 4862 16652
rect 4856 16612 8524 16640
rect 4856 16600 4862 16612
rect 3896 16544 4200 16572
rect 2409 16535 2467 16541
rect 4522 16532 4528 16584
rect 4580 16572 4586 16584
rect 4617 16575 4675 16581
rect 4617 16572 4629 16575
rect 4580 16544 4629 16572
rect 4580 16532 4586 16544
rect 4617 16541 4629 16544
rect 4663 16541 4675 16575
rect 8496 16572 8524 16612
rect 9122 16600 9128 16652
rect 9180 16640 9186 16652
rect 9217 16643 9275 16649
rect 9217 16640 9229 16643
rect 9180 16612 9229 16640
rect 9180 16600 9186 16612
rect 9217 16609 9229 16612
rect 9263 16609 9275 16643
rect 9508 16640 9536 16680
rect 9217 16603 9275 16609
rect 9324 16612 9536 16640
rect 9585 16643 9643 16649
rect 9324 16572 9352 16612
rect 9585 16609 9597 16643
rect 9631 16640 9643 16643
rect 9858 16640 9864 16652
rect 9631 16612 9864 16640
rect 9631 16609 9643 16612
rect 9585 16603 9643 16609
rect 9858 16600 9864 16612
rect 9916 16600 9922 16652
rect 9950 16600 9956 16652
rect 10008 16640 10014 16652
rect 12805 16643 12863 16649
rect 10008 16612 10053 16640
rect 10008 16600 10014 16612
rect 12805 16609 12817 16643
rect 12851 16640 12863 16643
rect 13188 16640 13216 16680
rect 12851 16612 13216 16640
rect 13265 16643 13323 16649
rect 12851 16609 12863 16612
rect 12805 16603 12863 16609
rect 13265 16609 13277 16643
rect 13311 16609 13323 16643
rect 13265 16603 13323 16609
rect 8496 16544 9352 16572
rect 4617 16535 4675 16541
rect 11330 16532 11336 16584
rect 11388 16572 11394 16584
rect 13280 16572 13308 16603
rect 11388 16544 13308 16572
rect 11388 16532 11394 16544
rect 1627 16507 1685 16513
rect 1627 16473 1639 16507
rect 1673 16504 1685 16507
rect 2317 16507 2375 16513
rect 2317 16504 2329 16507
rect 1673 16476 2329 16504
rect 1673 16473 1685 16476
rect 1627 16467 1685 16473
rect 2317 16473 2329 16476
rect 2363 16504 2375 16507
rect 2590 16504 2596 16516
rect 2363 16476 2596 16504
rect 2363 16473 2375 16476
rect 2317 16467 2375 16473
rect 2590 16464 2596 16476
rect 2648 16464 2654 16516
rect 5721 16507 5779 16513
rect 5721 16473 5733 16507
rect 5767 16504 5779 16507
rect 5810 16504 5816 16516
rect 5767 16476 5816 16504
rect 5767 16473 5779 16476
rect 5721 16467 5779 16473
rect 5810 16464 5816 16476
rect 5868 16504 5874 16516
rect 7098 16504 7104 16516
rect 5868 16476 7104 16504
rect 5868 16464 5874 16476
rect 7098 16464 7104 16476
rect 7156 16464 7162 16516
rect 10042 16464 10048 16516
rect 10100 16504 10106 16516
rect 11241 16507 11299 16513
rect 11241 16504 11253 16507
rect 10100 16476 11253 16504
rect 10100 16464 10106 16476
rect 11241 16473 11253 16476
rect 11287 16473 11299 16507
rect 11241 16467 11299 16473
rect 11514 16464 11520 16516
rect 11572 16504 11578 16516
rect 13170 16504 13176 16516
rect 11572 16476 13176 16504
rect 11572 16464 11578 16476
rect 13170 16464 13176 16476
rect 13228 16464 13234 16516
rect 13446 16504 13452 16516
rect 13407 16476 13452 16504
rect 13446 16464 13452 16476
rect 13504 16464 13510 16516
rect 13556 16504 13584 16680
rect 13814 16668 13820 16720
rect 13872 16708 13878 16720
rect 16758 16708 16764 16720
rect 13872 16680 14964 16708
rect 16422 16680 16764 16708
rect 13872 16668 13878 16680
rect 13630 16600 13636 16652
rect 13688 16640 13694 16652
rect 14936 16649 14964 16680
rect 16758 16668 16764 16680
rect 16816 16708 16822 16720
rect 17494 16708 17500 16720
rect 16816 16680 17500 16708
rect 16816 16668 16822 16680
rect 17494 16668 17500 16680
rect 17552 16668 17558 16720
rect 14185 16643 14243 16649
rect 14185 16640 14197 16643
rect 13688 16612 14197 16640
rect 13688 16600 13694 16612
rect 14185 16609 14197 16612
rect 14231 16609 14243 16643
rect 14185 16603 14243 16609
rect 14921 16643 14979 16649
rect 14921 16609 14933 16643
rect 14967 16609 14979 16643
rect 17770 16640 17776 16652
rect 17731 16612 17776 16640
rect 14921 16603 14979 16609
rect 17770 16600 17776 16612
rect 17828 16600 17834 16652
rect 18414 16640 18420 16652
rect 18375 16612 18420 16640
rect 18414 16600 18420 16612
rect 18472 16600 18478 16652
rect 14274 16572 14280 16584
rect 14235 16544 14280 16572
rect 14274 16532 14280 16544
rect 14332 16532 14338 16584
rect 15197 16575 15255 16581
rect 15197 16541 15209 16575
rect 15243 16572 15255 16575
rect 15930 16572 15936 16584
rect 15243 16544 15936 16572
rect 15243 16541 15255 16544
rect 15197 16535 15255 16541
rect 15930 16532 15936 16544
rect 15988 16532 15994 16584
rect 13556 16476 14872 16504
rect 1489 16439 1547 16445
rect 1489 16405 1501 16439
rect 1535 16436 1547 16439
rect 2222 16436 2228 16448
rect 1535 16408 2228 16436
rect 1535 16405 1547 16408
rect 1489 16399 1547 16405
rect 2222 16396 2228 16408
rect 2280 16396 2286 16448
rect 12710 16436 12716 16448
rect 12623 16408 12716 16436
rect 12710 16396 12716 16408
rect 12768 16436 12774 16448
rect 13262 16436 13268 16448
rect 12768 16408 13268 16436
rect 12768 16396 12774 16408
rect 13262 16396 13268 16408
rect 13320 16396 13326 16448
rect 13909 16439 13967 16445
rect 13909 16405 13921 16439
rect 13955 16436 13967 16439
rect 14274 16436 14280 16448
rect 13955 16408 14280 16436
rect 13955 16405 13967 16408
rect 13909 16399 13967 16405
rect 14274 16396 14280 16408
rect 14332 16396 14338 16448
rect 14844 16436 14872 16476
rect 16390 16436 16396 16448
rect 14844 16408 16396 16436
rect 16390 16396 16396 16408
rect 16448 16436 16454 16448
rect 16669 16439 16727 16445
rect 16669 16436 16681 16439
rect 16448 16408 16681 16436
rect 16448 16396 16454 16408
rect 16669 16405 16681 16408
rect 16715 16405 16727 16439
rect 16669 16399 16727 16405
rect 16758 16396 16764 16448
rect 16816 16436 16822 16448
rect 17129 16439 17187 16445
rect 17129 16436 17141 16439
rect 16816 16408 17141 16436
rect 16816 16396 16822 16408
rect 17129 16405 17141 16408
rect 17175 16405 17187 16439
rect 17129 16399 17187 16405
rect 184 16346 18860 16368
rect 184 16294 1556 16346
rect 1608 16294 1620 16346
rect 1672 16294 1684 16346
rect 1736 16294 1748 16346
rect 1800 16294 1812 16346
rect 1864 16294 4656 16346
rect 4708 16294 4720 16346
rect 4772 16294 4784 16346
rect 4836 16294 4848 16346
rect 4900 16294 4912 16346
rect 4964 16294 7756 16346
rect 7808 16294 7820 16346
rect 7872 16294 7884 16346
rect 7936 16294 7948 16346
rect 8000 16294 8012 16346
rect 8064 16294 10856 16346
rect 10908 16294 10920 16346
rect 10972 16294 10984 16346
rect 11036 16294 11048 16346
rect 11100 16294 11112 16346
rect 11164 16294 13956 16346
rect 14008 16294 14020 16346
rect 14072 16294 14084 16346
rect 14136 16294 14148 16346
rect 14200 16294 14212 16346
rect 14264 16294 17056 16346
rect 17108 16294 17120 16346
rect 17172 16294 17184 16346
rect 17236 16294 17248 16346
rect 17300 16294 17312 16346
rect 17364 16294 18860 16346
rect 184 16272 18860 16294
rect 5534 16192 5540 16244
rect 5592 16232 5598 16244
rect 5905 16235 5963 16241
rect 5905 16232 5917 16235
rect 5592 16204 5917 16232
rect 5592 16192 5598 16204
rect 5905 16201 5917 16204
rect 5951 16201 5963 16235
rect 5905 16195 5963 16201
rect 10318 16192 10324 16244
rect 10376 16232 10382 16244
rect 12437 16235 12495 16241
rect 12437 16232 12449 16235
rect 10376 16204 12449 16232
rect 10376 16192 10382 16204
rect 12437 16201 12449 16204
rect 12483 16201 12495 16235
rect 13814 16232 13820 16244
rect 13775 16204 13820 16232
rect 12437 16195 12495 16201
rect 13814 16192 13820 16204
rect 13872 16192 13878 16244
rect 18414 16164 18420 16176
rect 18375 16136 18420 16164
rect 18414 16124 18420 16136
rect 18472 16124 18478 16176
rect 4157 16099 4215 16105
rect 4157 16065 4169 16099
rect 4203 16096 4215 16099
rect 5166 16096 5172 16108
rect 4203 16068 5172 16096
rect 4203 16065 4215 16068
rect 4157 16059 4215 16065
rect 5166 16056 5172 16068
rect 5224 16056 5230 16108
rect 5626 16056 5632 16108
rect 5684 16056 5690 16108
rect 16485 16099 16543 16105
rect 16485 16065 16497 16099
rect 16531 16096 16543 16099
rect 16758 16096 16764 16108
rect 16531 16068 16764 16096
rect 16531 16065 16543 16068
rect 16485 16059 16543 16065
rect 16758 16056 16764 16068
rect 16816 16056 16822 16108
rect 2314 15988 2320 16040
rect 2372 16028 2378 16040
rect 2409 16031 2467 16037
rect 2409 16028 2421 16031
rect 2372 16000 2421 16028
rect 2372 15988 2378 16000
rect 2409 15997 2421 16000
rect 2455 15997 2467 16031
rect 2590 16028 2596 16040
rect 2551 16000 2596 16028
rect 2409 15991 2467 15997
rect 2590 15988 2596 16000
rect 2648 15988 2654 16040
rect 4338 15920 4344 15972
rect 4396 15960 4402 15972
rect 4433 15963 4491 15969
rect 4433 15960 4445 15963
rect 4396 15932 4445 15960
rect 4396 15920 4402 15932
rect 4433 15929 4445 15932
rect 4479 15929 4491 15963
rect 5644 15960 5672 16056
rect 6641 16031 6699 16037
rect 6641 15997 6653 16031
rect 6687 16028 6699 16031
rect 7006 16028 7012 16040
rect 6687 16000 7012 16028
rect 6687 15997 6699 16000
rect 6641 15991 6699 15997
rect 7006 15988 7012 16000
rect 7064 15988 7070 16040
rect 8389 16031 8447 16037
rect 8389 15997 8401 16031
rect 8435 16028 8447 16031
rect 11330 16028 11336 16040
rect 8435 16000 11336 16028
rect 8435 15997 8447 16000
rect 8389 15991 8447 15997
rect 11330 15988 11336 16000
rect 11388 15988 11394 16040
rect 16117 16031 16175 16037
rect 16117 15997 16129 16031
rect 16163 16028 16175 16031
rect 16206 16028 16212 16040
rect 16163 16000 16212 16028
rect 16163 15997 16175 16000
rect 16117 15991 16175 15997
rect 16206 15988 16212 16000
rect 16264 15988 16270 16040
rect 6546 15960 6552 15972
rect 5644 15946 6552 15960
rect 5658 15932 6552 15946
rect 4433 15923 4491 15929
rect 6546 15920 6552 15932
rect 6604 15920 6610 15972
rect 8757 15963 8815 15969
rect 8757 15929 8769 15963
rect 8803 15960 8815 15963
rect 9030 15960 9036 15972
rect 8803 15932 9036 15960
rect 8803 15929 8815 15932
rect 8757 15923 8815 15929
rect 9030 15920 9036 15932
rect 9088 15920 9094 15972
rect 11146 15960 11152 15972
rect 11107 15932 11152 15960
rect 11146 15920 11152 15932
rect 11204 15960 11210 15972
rect 11422 15960 11428 15972
rect 11204 15932 11428 15960
rect 11204 15920 11210 15932
rect 11422 15920 11428 15932
rect 11480 15920 11486 15972
rect 15010 15920 15016 15972
rect 15068 15960 15074 15972
rect 15289 15963 15347 15969
rect 15289 15960 15301 15963
rect 15068 15932 15301 15960
rect 15068 15920 15074 15932
rect 15289 15929 15301 15932
rect 15335 15929 15347 15963
rect 15289 15923 15347 15929
rect 17494 15920 17500 15972
rect 17552 15920 17558 15972
rect 2501 15895 2559 15901
rect 2501 15861 2513 15895
rect 2547 15892 2559 15895
rect 3602 15892 3608 15904
rect 2547 15864 3608 15892
rect 2547 15861 2559 15864
rect 2501 15855 2559 15861
rect 3602 15852 3608 15864
rect 3660 15852 3666 15904
rect 8018 15852 8024 15904
rect 8076 15892 8082 15904
rect 10045 15895 10103 15901
rect 10045 15892 10057 15895
rect 8076 15864 10057 15892
rect 8076 15852 8082 15864
rect 10045 15861 10057 15864
rect 10091 15861 10103 15895
rect 10045 15855 10103 15861
rect 17862 15852 17868 15904
rect 17920 15901 17926 15904
rect 17920 15895 17969 15901
rect 17920 15861 17923 15895
rect 17957 15861 17969 15895
rect 17920 15855 17969 15861
rect 17920 15852 17926 15855
rect 184 15802 18920 15824
rect 184 15750 3106 15802
rect 3158 15750 3170 15802
rect 3222 15750 3234 15802
rect 3286 15750 3298 15802
rect 3350 15750 3362 15802
rect 3414 15750 6206 15802
rect 6258 15750 6270 15802
rect 6322 15750 6334 15802
rect 6386 15750 6398 15802
rect 6450 15750 6462 15802
rect 6514 15750 9306 15802
rect 9358 15750 9370 15802
rect 9422 15750 9434 15802
rect 9486 15750 9498 15802
rect 9550 15750 9562 15802
rect 9614 15750 12406 15802
rect 12458 15750 12470 15802
rect 12522 15750 12534 15802
rect 12586 15750 12598 15802
rect 12650 15750 12662 15802
rect 12714 15750 15506 15802
rect 15558 15750 15570 15802
rect 15622 15750 15634 15802
rect 15686 15750 15698 15802
rect 15750 15750 15762 15802
rect 15814 15750 18606 15802
rect 18658 15750 18670 15802
rect 18722 15750 18734 15802
rect 18786 15750 18798 15802
rect 18850 15750 18862 15802
rect 18914 15750 18920 15802
rect 184 15728 18920 15750
rect 3237 15691 3295 15697
rect 3237 15657 3249 15691
rect 3283 15688 3295 15691
rect 4062 15688 4068 15700
rect 3283 15660 4068 15688
rect 3283 15657 3295 15660
rect 3237 15651 3295 15657
rect 4062 15648 4068 15660
rect 4120 15648 4126 15700
rect 5721 15691 5779 15697
rect 5721 15657 5733 15691
rect 5767 15688 5779 15691
rect 6822 15688 6828 15700
rect 5767 15660 6828 15688
rect 5767 15657 5779 15660
rect 5721 15651 5779 15657
rect 6822 15648 6828 15660
rect 6880 15648 6886 15700
rect 11146 15688 11152 15700
rect 7024 15660 11152 15688
rect 4430 15580 4436 15632
rect 4488 15620 4494 15632
rect 7024 15629 7052 15660
rect 11146 15648 11152 15660
rect 11204 15648 11210 15700
rect 11974 15688 11980 15700
rect 11935 15660 11980 15688
rect 11974 15648 11980 15660
rect 12032 15648 12038 15700
rect 12713 15691 12771 15697
rect 12713 15657 12725 15691
rect 12759 15688 12771 15691
rect 12802 15688 12808 15700
rect 12759 15660 12808 15688
rect 12759 15657 12771 15660
rect 12713 15651 12771 15657
rect 12802 15648 12808 15660
rect 12860 15648 12866 15700
rect 14001 15691 14059 15697
rect 14001 15657 14013 15691
rect 14047 15688 14059 15691
rect 14274 15688 14280 15700
rect 14047 15660 14280 15688
rect 14047 15657 14059 15660
rect 14001 15651 14059 15657
rect 14274 15648 14280 15660
rect 14332 15648 14338 15700
rect 18230 15688 18236 15700
rect 18191 15660 18236 15688
rect 18230 15648 18236 15660
rect 18288 15648 18294 15700
rect 4525 15623 4583 15629
rect 4525 15620 4537 15623
rect 4488 15592 4537 15620
rect 4488 15580 4494 15592
rect 4525 15589 4537 15592
rect 4571 15589 4583 15623
rect 4525 15583 4583 15589
rect 7009 15623 7067 15629
rect 7009 15589 7021 15623
rect 7055 15589 7067 15623
rect 8018 15620 8024 15632
rect 7009 15583 7067 15589
rect 7760 15592 8024 15620
rect 7760 15561 7788 15592
rect 8018 15580 8024 15592
rect 8076 15580 8082 15632
rect 8294 15580 8300 15632
rect 8352 15620 8358 15632
rect 8352 15592 8510 15620
rect 8352 15580 8358 15592
rect 11514 15580 11520 15632
rect 11572 15580 11578 15632
rect 13446 15580 13452 15632
rect 13504 15620 13510 15632
rect 13909 15623 13967 15629
rect 13909 15620 13921 15623
rect 13504 15592 13921 15620
rect 13504 15580 13510 15592
rect 13909 15589 13921 15592
rect 13955 15620 13967 15623
rect 14366 15620 14372 15632
rect 13955 15592 14372 15620
rect 13955 15589 13967 15592
rect 13909 15583 13967 15589
rect 14366 15580 14372 15592
rect 14424 15620 14430 15632
rect 16298 15620 16304 15632
rect 14424 15592 16304 15620
rect 14424 15580 14430 15592
rect 16298 15580 16304 15592
rect 16356 15620 16362 15632
rect 17862 15620 17868 15632
rect 16356 15592 17868 15620
rect 16356 15580 16362 15592
rect 17862 15580 17868 15592
rect 17920 15580 17926 15632
rect 7745 15555 7803 15561
rect 7745 15521 7757 15555
rect 7791 15521 7803 15555
rect 12802 15552 12808 15564
rect 12715 15524 12808 15552
rect 7745 15515 7803 15521
rect 12802 15512 12808 15524
rect 12860 15552 12866 15564
rect 13262 15552 13268 15564
rect 12860 15524 13268 15552
rect 12860 15512 12866 15524
rect 13262 15512 13268 15524
rect 13320 15512 13326 15564
rect 16482 15552 16488 15564
rect 16443 15524 16488 15552
rect 16482 15512 16488 15524
rect 16540 15512 16546 15564
rect 17957 15555 18015 15561
rect 17957 15521 17969 15555
rect 18003 15552 18015 15555
rect 18417 15555 18475 15561
rect 18417 15552 18429 15555
rect 18003 15524 18429 15552
rect 18003 15521 18015 15524
rect 17957 15515 18015 15521
rect 18417 15521 18429 15524
rect 18463 15552 18475 15555
rect 19058 15552 19064 15564
rect 18463 15524 19064 15552
rect 18463 15521 18475 15524
rect 18417 15515 18475 15521
rect 19058 15512 19064 15524
rect 19116 15512 19122 15564
rect 7650 15444 7656 15496
rect 7708 15484 7714 15496
rect 8021 15487 8079 15493
rect 8021 15484 8033 15487
rect 7708 15456 8033 15484
rect 7708 15444 7714 15456
rect 8021 15453 8033 15456
rect 8067 15453 8079 15487
rect 10226 15484 10232 15496
rect 10187 15456 10232 15484
rect 8021 15447 8079 15453
rect 10226 15444 10232 15456
rect 10284 15444 10290 15496
rect 10505 15487 10563 15493
rect 10505 15453 10517 15487
rect 10551 15484 10563 15487
rect 11514 15484 11520 15496
rect 10551 15456 11520 15484
rect 10551 15453 10563 15456
rect 10505 15447 10563 15453
rect 11514 15444 11520 15456
rect 11572 15444 11578 15496
rect 12894 15484 12900 15496
rect 12855 15456 12900 15484
rect 12894 15444 12900 15456
rect 12952 15444 12958 15496
rect 13814 15484 13820 15496
rect 13775 15456 13820 15484
rect 13814 15444 13820 15456
rect 13872 15444 13878 15496
rect 9490 15348 9496 15360
rect 9451 15320 9496 15348
rect 9490 15308 9496 15320
rect 9548 15308 9554 15360
rect 12342 15348 12348 15360
rect 12303 15320 12348 15348
rect 12342 15308 12348 15320
rect 12400 15308 12406 15360
rect 14369 15351 14427 15357
rect 14369 15317 14381 15351
rect 14415 15348 14427 15351
rect 14826 15348 14832 15360
rect 14415 15320 14832 15348
rect 14415 15317 14427 15320
rect 14369 15311 14427 15317
rect 14826 15308 14832 15320
rect 14884 15308 14890 15360
rect 15010 15308 15016 15360
rect 15068 15348 15074 15360
rect 15197 15351 15255 15357
rect 15197 15348 15209 15351
rect 15068 15320 15209 15348
rect 15068 15308 15074 15320
rect 15197 15317 15209 15320
rect 15243 15317 15255 15351
rect 15197 15311 15255 15317
rect 184 15258 18860 15280
rect 184 15206 1556 15258
rect 1608 15206 1620 15258
rect 1672 15206 1684 15258
rect 1736 15206 1748 15258
rect 1800 15206 1812 15258
rect 1864 15206 4656 15258
rect 4708 15206 4720 15258
rect 4772 15206 4784 15258
rect 4836 15206 4848 15258
rect 4900 15206 4912 15258
rect 4964 15206 7756 15258
rect 7808 15206 7820 15258
rect 7872 15206 7884 15258
rect 7936 15206 7948 15258
rect 8000 15206 8012 15258
rect 8064 15206 10856 15258
rect 10908 15206 10920 15258
rect 10972 15206 10984 15258
rect 11036 15206 11048 15258
rect 11100 15206 11112 15258
rect 11164 15206 13956 15258
rect 14008 15206 14020 15258
rect 14072 15206 14084 15258
rect 14136 15206 14148 15258
rect 14200 15206 14212 15258
rect 14264 15206 17056 15258
rect 17108 15206 17120 15258
rect 17172 15206 17184 15258
rect 17236 15206 17248 15258
rect 17300 15206 17312 15258
rect 17364 15206 18860 15258
rect 184 15184 18860 15206
rect 5902 15144 5908 15156
rect 5863 15116 5908 15144
rect 5902 15104 5908 15116
rect 5960 15104 5966 15156
rect 8113 15147 8171 15153
rect 6472 15116 8064 15144
rect 6472 15076 6500 15116
rect 5184 15048 6500 15076
rect 8036 15076 8064 15116
rect 8113 15113 8125 15147
rect 8159 15144 8171 15147
rect 8202 15144 8208 15156
rect 8159 15116 8208 15144
rect 8159 15113 8171 15116
rect 8113 15107 8171 15113
rect 8202 15104 8208 15116
rect 8260 15104 8266 15156
rect 9858 15104 9864 15156
rect 9916 15144 9922 15156
rect 11241 15147 11299 15153
rect 11241 15144 11253 15147
rect 9916 15116 11253 15144
rect 9916 15104 9922 15116
rect 11241 15113 11253 15116
rect 11287 15113 11299 15147
rect 11241 15107 11299 15113
rect 12986 15104 12992 15156
rect 13044 15144 13050 15156
rect 13630 15144 13636 15156
rect 13044 15116 13636 15144
rect 13044 15104 13050 15116
rect 13630 15104 13636 15116
rect 13688 15104 13694 15156
rect 14001 15147 14059 15153
rect 14001 15113 14013 15147
rect 14047 15144 14059 15147
rect 15102 15144 15108 15156
rect 14047 15116 15108 15144
rect 14047 15113 14059 15116
rect 14001 15107 14059 15113
rect 15102 15104 15108 15116
rect 15160 15104 15166 15156
rect 8754 15076 8760 15088
rect 8036 15048 8760 15076
rect 2130 15008 2136 15020
rect 2091 14980 2136 15008
rect 2130 14968 2136 14980
rect 2188 14968 2194 15020
rect 2222 14968 2228 15020
rect 2280 15008 2286 15020
rect 2777 15011 2835 15017
rect 2777 15008 2789 15011
rect 2280 14980 2789 15008
rect 2280 14968 2286 14980
rect 2777 14977 2789 14980
rect 2823 15008 2835 15011
rect 2823 14980 3464 15008
rect 2823 14977 2835 14980
rect 2777 14971 2835 14977
rect 2041 14943 2099 14949
rect 2041 14909 2053 14943
rect 2087 14940 2099 14943
rect 2590 14940 2596 14952
rect 2087 14912 2596 14940
rect 2087 14909 2099 14912
rect 2041 14903 2099 14909
rect 2590 14900 2596 14912
rect 2648 14940 2654 14952
rect 3436 14949 3464 14980
rect 3620 14980 4292 15008
rect 3620 14952 3648 14980
rect 2855 14943 2913 14949
rect 2855 14940 2867 14943
rect 2648 14912 2867 14940
rect 2648 14900 2654 14912
rect 2855 14909 2867 14912
rect 2901 14909 2913 14943
rect 2855 14903 2913 14909
rect 3421 14943 3479 14949
rect 3421 14909 3433 14943
rect 3467 14909 3479 14943
rect 3602 14940 3608 14952
rect 3563 14912 3608 14940
rect 3421 14903 3479 14909
rect 1949 14875 2007 14881
rect 1949 14841 1961 14875
rect 1995 14872 2007 14875
rect 2682 14872 2688 14884
rect 1995 14844 2688 14872
rect 1995 14841 2007 14844
rect 1949 14835 2007 14841
rect 2682 14832 2688 14844
rect 2740 14832 2746 14884
rect 3436 14872 3464 14903
rect 3602 14900 3608 14912
rect 3660 14900 3666 14952
rect 4062 14940 4068 14952
rect 4023 14912 4068 14940
rect 4062 14900 4068 14912
rect 4120 14900 4126 14952
rect 4264 14949 4292 14980
rect 5184 14949 5212 15048
rect 8754 15036 8760 15048
rect 8812 15076 8818 15088
rect 9490 15076 9496 15088
rect 8812 15048 9496 15076
rect 8812 15036 8818 15048
rect 9490 15036 9496 15048
rect 9548 15036 9554 15088
rect 11974 15036 11980 15088
rect 12032 15036 12038 15088
rect 14737 15079 14795 15085
rect 14737 15045 14749 15079
rect 14783 15045 14795 15079
rect 14737 15039 14795 15045
rect 6365 15011 6423 15017
rect 6365 14977 6377 15011
rect 6411 15008 6423 15011
rect 6638 15008 6644 15020
rect 6411 14980 6644 15008
rect 6411 14977 6423 14980
rect 6365 14971 6423 14977
rect 6638 14968 6644 14980
rect 6696 14968 6702 15020
rect 11992 15008 12020 15036
rect 13081 15011 13139 15017
rect 11992 14980 12572 15008
rect 4157 14943 4215 14949
rect 4157 14909 4169 14943
rect 4203 14909 4215 14943
rect 4157 14903 4215 14909
rect 4249 14943 4307 14949
rect 4249 14909 4261 14943
rect 4295 14909 4307 14943
rect 4249 14903 4307 14909
rect 5169 14943 5227 14949
rect 5169 14909 5181 14943
rect 5215 14909 5227 14943
rect 5810 14940 5816 14952
rect 5771 14912 5816 14940
rect 5169 14903 5227 14909
rect 4172 14872 4200 14903
rect 5810 14900 5816 14912
rect 5868 14900 5874 14952
rect 8110 14940 8116 14952
rect 7774 14912 8116 14940
rect 8110 14900 8116 14912
rect 8168 14900 8174 14952
rect 11330 14940 11336 14952
rect 11291 14912 11336 14940
rect 11330 14900 11336 14912
rect 11388 14900 11394 14952
rect 11977 14943 12035 14949
rect 11977 14909 11989 14943
rect 12023 14940 12035 14943
rect 12342 14940 12348 14952
rect 12023 14912 12348 14940
rect 12023 14909 12035 14912
rect 11977 14903 12035 14909
rect 12342 14900 12348 14912
rect 12400 14900 12406 14952
rect 12544 14949 12572 14980
rect 13081 14977 13093 15011
rect 13127 15008 13139 15011
rect 13127 14980 13860 15008
rect 13127 14977 13139 14980
rect 13081 14971 13139 14977
rect 12437 14943 12495 14949
rect 12437 14909 12449 14943
rect 12483 14909 12495 14943
rect 12437 14903 12495 14909
rect 12529 14943 12587 14949
rect 12529 14909 12541 14943
rect 12575 14909 12587 14943
rect 12529 14903 12587 14909
rect 12621 14943 12679 14949
rect 12621 14909 12633 14943
rect 12667 14940 12679 14943
rect 12894 14940 12900 14952
rect 12667 14912 12900 14940
rect 12667 14909 12679 14912
rect 12621 14903 12679 14909
rect 3436 14844 4200 14872
rect 4617 14875 4675 14881
rect 4617 14841 4629 14875
rect 4663 14872 4675 14875
rect 4982 14872 4988 14884
rect 4663 14844 4988 14872
rect 4663 14841 4675 14844
rect 4617 14835 4675 14841
rect 4982 14832 4988 14844
rect 5040 14832 5046 14884
rect 6641 14875 6699 14881
rect 6641 14841 6653 14875
rect 6687 14872 6699 14875
rect 6914 14872 6920 14884
rect 6687 14844 6920 14872
rect 6687 14841 6699 14844
rect 6641 14835 6699 14841
rect 6914 14832 6920 14844
rect 6972 14832 6978 14884
rect 8757 14875 8815 14881
rect 8757 14872 8769 14875
rect 7944 14844 8769 14872
rect 842 14764 848 14816
rect 900 14804 906 14816
rect 1581 14807 1639 14813
rect 1581 14804 1593 14807
rect 900 14776 1593 14804
rect 900 14764 906 14776
rect 1581 14773 1593 14776
rect 1627 14773 1639 14807
rect 1581 14767 1639 14773
rect 2958 14764 2964 14816
rect 3016 14804 3022 14816
rect 3145 14807 3203 14813
rect 3145 14804 3157 14807
rect 3016 14776 3157 14804
rect 3016 14764 3022 14776
rect 3145 14773 3157 14776
rect 3191 14773 3203 14807
rect 3510 14804 3516 14816
rect 3471 14776 3516 14804
rect 3145 14767 3203 14773
rect 3510 14764 3516 14776
rect 3568 14764 3574 14816
rect 4433 14807 4491 14813
rect 4433 14773 4445 14807
rect 4479 14804 4491 14807
rect 4798 14804 4804 14816
rect 4479 14776 4804 14804
rect 4479 14773 4491 14776
rect 4433 14767 4491 14773
rect 4798 14764 4804 14776
rect 4856 14764 4862 14816
rect 7558 14764 7564 14816
rect 7616 14804 7622 14816
rect 7944 14804 7972 14844
rect 8757 14841 8769 14844
rect 8803 14841 8815 14875
rect 12452 14872 12480 14903
rect 12894 14900 12900 14912
rect 12952 14900 12958 14952
rect 12986 14900 12992 14952
rect 13044 14940 13050 14952
rect 13832 14949 13860 14980
rect 13173 14943 13231 14949
rect 13044 14912 13089 14940
rect 13044 14900 13050 14912
rect 13173 14909 13185 14943
rect 13219 14909 13231 14943
rect 13173 14903 13231 14909
rect 13817 14943 13875 14949
rect 13817 14909 13829 14943
rect 13863 14909 13875 14943
rect 13817 14903 13875 14909
rect 13188 14872 13216 14903
rect 13906 14900 13912 14952
rect 13964 14940 13970 14952
rect 14369 14943 14427 14949
rect 13964 14912 14009 14940
rect 13964 14900 13970 14912
rect 14369 14909 14381 14943
rect 14415 14940 14427 14943
rect 14752 14940 14780 15039
rect 15194 14968 15200 15020
rect 15252 15008 15258 15020
rect 15289 15011 15347 15017
rect 15289 15008 15301 15011
rect 15252 14980 15301 15008
rect 15252 14968 15258 14980
rect 15289 14977 15301 14980
rect 15335 14977 15347 15011
rect 16850 15008 16856 15020
rect 15289 14971 15347 14977
rect 15396 14980 16856 15008
rect 14415 14912 14780 14940
rect 14415 14909 14427 14912
rect 14369 14903 14427 14909
rect 14826 14900 14832 14952
rect 14884 14940 14890 14952
rect 15105 14943 15163 14949
rect 15105 14940 15117 14943
rect 14884 14912 15117 14940
rect 14884 14900 14890 14912
rect 15105 14909 15117 14912
rect 15151 14909 15163 14943
rect 15105 14903 15163 14909
rect 12452 14844 13216 14872
rect 8757 14835 8815 14841
rect 13004 14816 13032 14844
rect 13722 14832 13728 14884
rect 13780 14872 13786 14884
rect 15396 14872 15424 14980
rect 16850 14968 16856 14980
rect 16908 14968 16914 15020
rect 16206 14940 16212 14952
rect 16167 14912 16212 14940
rect 16206 14900 16212 14912
rect 16264 14900 16270 14952
rect 17586 14900 17592 14952
rect 17644 14900 17650 14952
rect 13780 14844 15424 14872
rect 16485 14875 16543 14881
rect 13780 14832 13786 14844
rect 16485 14841 16497 14875
rect 16531 14872 16543 14875
rect 16758 14872 16764 14884
rect 16531 14844 16764 14872
rect 16531 14841 16543 14844
rect 16485 14835 16543 14841
rect 16758 14832 16764 14844
rect 16816 14832 16822 14884
rect 7616 14776 7972 14804
rect 7616 14764 7622 14776
rect 9030 14764 9036 14816
rect 9088 14804 9094 14816
rect 10045 14807 10103 14813
rect 10045 14804 10057 14807
rect 9088 14776 10057 14804
rect 9088 14764 9094 14776
rect 10045 14773 10057 14776
rect 10091 14773 10103 14807
rect 10045 14767 10103 14773
rect 11330 14764 11336 14816
rect 11388 14804 11394 14816
rect 11885 14807 11943 14813
rect 11885 14804 11897 14807
rect 11388 14776 11897 14804
rect 11388 14764 11394 14776
rect 11885 14773 11897 14776
rect 11931 14773 11943 14807
rect 12250 14804 12256 14816
rect 12211 14776 12256 14804
rect 11885 14767 11943 14773
rect 12250 14764 12256 14776
rect 12308 14764 12314 14816
rect 12986 14764 12992 14816
rect 13044 14764 13050 14816
rect 14274 14804 14280 14816
rect 14235 14776 14280 14804
rect 14274 14764 14280 14776
rect 14332 14764 14338 14816
rect 14642 14764 14648 14816
rect 14700 14804 14706 14816
rect 14826 14804 14832 14816
rect 14700 14776 14832 14804
rect 14700 14764 14706 14776
rect 14826 14764 14832 14776
rect 14884 14804 14890 14816
rect 15197 14807 15255 14813
rect 15197 14804 15209 14807
rect 14884 14776 15209 14804
rect 14884 14764 14890 14776
rect 15197 14773 15209 14776
rect 15243 14804 15255 14807
rect 16574 14804 16580 14816
rect 15243 14776 16580 14804
rect 15243 14773 15255 14776
rect 15197 14767 15255 14773
rect 16574 14764 16580 14776
rect 16632 14764 16638 14816
rect 17954 14804 17960 14816
rect 17915 14776 17960 14804
rect 17954 14764 17960 14776
rect 18012 14764 18018 14816
rect 184 14714 18920 14736
rect 184 14662 3106 14714
rect 3158 14662 3170 14714
rect 3222 14662 3234 14714
rect 3286 14662 3298 14714
rect 3350 14662 3362 14714
rect 3414 14662 6206 14714
rect 6258 14662 6270 14714
rect 6322 14662 6334 14714
rect 6386 14662 6398 14714
rect 6450 14662 6462 14714
rect 6514 14662 9306 14714
rect 9358 14662 9370 14714
rect 9422 14662 9434 14714
rect 9486 14662 9498 14714
rect 9550 14662 9562 14714
rect 9614 14662 12406 14714
rect 12458 14662 12470 14714
rect 12522 14662 12534 14714
rect 12586 14662 12598 14714
rect 12650 14662 12662 14714
rect 12714 14662 15506 14714
rect 15558 14662 15570 14714
rect 15622 14662 15634 14714
rect 15686 14662 15698 14714
rect 15750 14662 15762 14714
rect 15814 14662 18606 14714
rect 18658 14662 18670 14714
rect 18722 14662 18734 14714
rect 18786 14662 18798 14714
rect 18850 14662 18862 14714
rect 18914 14662 18920 14714
rect 184 14640 18920 14662
rect 2317 14603 2375 14609
rect 2317 14569 2329 14603
rect 2363 14600 2375 14603
rect 2590 14600 2596 14612
rect 2363 14572 2596 14600
rect 2363 14569 2375 14572
rect 2317 14563 2375 14569
rect 2590 14560 2596 14572
rect 2648 14560 2654 14612
rect 2682 14560 2688 14612
rect 2740 14600 2746 14612
rect 2777 14603 2835 14609
rect 2777 14600 2789 14603
rect 2740 14572 2789 14600
rect 2740 14560 2746 14572
rect 2777 14569 2789 14572
rect 2823 14569 2835 14603
rect 2777 14563 2835 14569
rect 2958 14560 2964 14612
rect 3016 14600 3022 14612
rect 3237 14603 3295 14609
rect 3237 14600 3249 14603
rect 3016 14572 3249 14600
rect 3016 14560 3022 14572
rect 3237 14569 3249 14572
rect 3283 14569 3295 14603
rect 4982 14600 4988 14612
rect 3237 14563 3295 14569
rect 3804 14572 4988 14600
rect 842 14532 848 14544
rect 803 14504 848 14532
rect 842 14492 848 14504
rect 900 14492 906 14544
rect 2130 14492 2136 14544
rect 2188 14532 2194 14544
rect 3804 14532 3832 14572
rect 4982 14560 4988 14572
rect 5040 14560 5046 14612
rect 7650 14600 7656 14612
rect 7611 14572 7656 14600
rect 7650 14560 7656 14572
rect 7708 14560 7714 14612
rect 11057 14603 11115 14609
rect 11057 14569 11069 14603
rect 11103 14600 11115 14603
rect 11514 14600 11520 14612
rect 11103 14572 11520 14600
rect 11103 14569 11115 14572
rect 11057 14563 11115 14569
rect 11514 14560 11520 14572
rect 11572 14560 11578 14612
rect 11609 14603 11667 14609
rect 11609 14569 11621 14603
rect 11655 14600 11667 14603
rect 11698 14600 11704 14612
rect 11655 14572 11704 14600
rect 11655 14569 11667 14572
rect 11609 14563 11667 14569
rect 11698 14560 11704 14572
rect 11756 14560 11762 14612
rect 12621 14603 12679 14609
rect 12621 14569 12633 14603
rect 12667 14600 12679 14603
rect 12802 14600 12808 14612
rect 12667 14572 12808 14600
rect 12667 14569 12679 14572
rect 12621 14563 12679 14569
rect 12802 14560 12808 14572
rect 12860 14560 12866 14612
rect 13265 14603 13323 14609
rect 13265 14569 13277 14603
rect 13311 14600 13323 14603
rect 14274 14600 14280 14612
rect 13311 14572 14280 14600
rect 13311 14569 13323 14572
rect 13265 14563 13323 14569
rect 14274 14560 14280 14572
rect 14332 14560 14338 14612
rect 14366 14560 14372 14612
rect 14424 14600 14430 14612
rect 15013 14603 15071 14609
rect 15013 14600 15025 14603
rect 14424 14572 15025 14600
rect 14424 14560 14430 14572
rect 15013 14569 15025 14572
rect 15059 14600 15071 14603
rect 16666 14600 16672 14612
rect 15059 14572 16672 14600
rect 15059 14569 15071 14572
rect 15013 14563 15071 14569
rect 16666 14560 16672 14572
rect 16724 14560 16730 14612
rect 16758 14560 16764 14612
rect 16816 14600 16822 14612
rect 17129 14603 17187 14609
rect 17129 14600 17141 14603
rect 16816 14572 17141 14600
rect 16816 14560 16822 14572
rect 17129 14569 17141 14572
rect 17175 14569 17187 14603
rect 17129 14563 17187 14569
rect 2188 14504 3832 14532
rect 2188 14492 2194 14504
rect 566 14464 572 14476
rect 527 14436 572 14464
rect 566 14424 572 14436
rect 624 14424 630 14476
rect 2314 14464 2320 14476
rect 1978 14436 2320 14464
rect 2314 14424 2320 14436
rect 2372 14464 2378 14476
rect 2498 14464 2504 14476
rect 2372 14436 2504 14464
rect 2372 14424 2378 14436
rect 2498 14424 2504 14436
rect 2556 14424 2562 14476
rect 3142 14464 3148 14476
rect 3103 14436 3148 14464
rect 3142 14424 3148 14436
rect 3200 14424 3206 14476
rect 3804 14473 3832 14504
rect 4065 14535 4123 14541
rect 4065 14501 4077 14535
rect 4111 14532 4123 14535
rect 4111 14504 4660 14532
rect 4111 14501 4123 14504
rect 4065 14495 4123 14501
rect 4632 14473 4660 14504
rect 6546 14492 6552 14544
rect 6604 14492 6610 14544
rect 9125 14535 9183 14541
rect 9125 14501 9137 14535
rect 9171 14532 9183 14535
rect 13722 14532 13728 14544
rect 9171 14504 10088 14532
rect 9171 14501 9183 14504
rect 9125 14495 9183 14501
rect 3789 14467 3847 14473
rect 3789 14433 3801 14467
rect 3835 14433 3847 14467
rect 3789 14427 3847 14433
rect 4617 14467 4675 14473
rect 4617 14433 4629 14467
rect 4663 14433 4675 14467
rect 4798 14464 4804 14476
rect 4759 14436 4804 14464
rect 4617 14427 4675 14433
rect 4798 14424 4804 14436
rect 4856 14424 4862 14476
rect 5166 14464 5172 14476
rect 5079 14436 5172 14464
rect 5166 14424 5172 14436
rect 5224 14464 5230 14476
rect 6564 14464 6592 14492
rect 7466 14464 7472 14476
rect 5224 14436 5672 14464
rect 6564 14436 7472 14464
rect 5224 14424 5230 14436
rect 3421 14399 3479 14405
rect 3421 14365 3433 14399
rect 3467 14396 3479 14399
rect 3510 14396 3516 14408
rect 3467 14368 3516 14396
rect 3467 14365 3479 14368
rect 3421 14359 3479 14365
rect 3510 14356 3516 14368
rect 3568 14396 3574 14408
rect 3881 14399 3939 14405
rect 3881 14396 3893 14399
rect 3568 14368 3893 14396
rect 3568 14356 3574 14368
rect 3881 14365 3893 14368
rect 3927 14365 3939 14399
rect 3881 14359 3939 14365
rect 4062 14356 4068 14408
rect 4120 14396 4126 14408
rect 4709 14399 4767 14405
rect 4120 14368 4213 14396
rect 4120 14356 4126 14368
rect 4709 14365 4721 14399
rect 4755 14396 4767 14399
rect 5537 14399 5595 14405
rect 5537 14396 5549 14399
rect 4755 14368 5549 14396
rect 4755 14365 4767 14368
rect 4709 14359 4767 14365
rect 5537 14365 5549 14368
rect 5583 14365 5595 14399
rect 5644 14396 5672 14436
rect 7466 14424 7472 14436
rect 7524 14464 7530 14476
rect 7524 14450 8050 14464
rect 7524 14436 8064 14450
rect 7524 14424 7530 14436
rect 6638 14396 6644 14408
rect 5644 14368 6644 14396
rect 5537 14359 5595 14365
rect 6638 14356 6644 14368
rect 6696 14356 6702 14408
rect 8036 14396 8064 14436
rect 8110 14396 8116 14408
rect 8036 14368 8116 14396
rect 8110 14356 8116 14368
rect 8168 14356 8174 14408
rect 9401 14399 9459 14405
rect 9401 14365 9413 14399
rect 9447 14365 9459 14399
rect 9401 14359 9459 14365
rect 4080 14260 4108 14356
rect 7006 14269 7012 14272
rect 6963 14263 7012 14269
rect 6963 14260 6975 14263
rect 4080 14232 6975 14260
rect 6963 14229 6975 14232
rect 7009 14229 7012 14263
rect 6963 14223 7012 14229
rect 7006 14220 7012 14223
rect 7064 14220 7070 14272
rect 9122 14220 9128 14272
rect 9180 14260 9186 14272
rect 9416 14260 9444 14359
rect 10060 14272 10088 14504
rect 12406 14504 13728 14532
rect 11330 14464 11336 14476
rect 11291 14436 11336 14464
rect 11330 14424 11336 14436
rect 11388 14424 11394 14476
rect 11882 14464 11888 14476
rect 11843 14436 11888 14464
rect 11882 14424 11888 14436
rect 11940 14424 11946 14476
rect 11977 14467 12035 14473
rect 11977 14433 11989 14467
rect 12023 14464 12035 14467
rect 12406 14464 12434 14504
rect 13722 14492 13728 14504
rect 13780 14492 13786 14544
rect 14001 14535 14059 14541
rect 14001 14501 14013 14535
rect 14047 14532 14059 14535
rect 14642 14532 14648 14544
rect 14047 14504 14648 14532
rect 14047 14501 14059 14504
rect 14001 14495 14059 14501
rect 14642 14492 14648 14504
rect 14700 14492 14706 14544
rect 15105 14535 15163 14541
rect 15105 14501 15117 14535
rect 15151 14532 15163 14535
rect 17954 14532 17960 14544
rect 15151 14504 17960 14532
rect 15151 14501 15163 14504
rect 15105 14495 15163 14501
rect 17954 14492 17960 14504
rect 18012 14532 18018 14544
rect 18233 14535 18291 14541
rect 18233 14532 18245 14535
rect 18012 14504 18245 14532
rect 18012 14492 18018 14504
rect 18233 14501 18245 14504
rect 18279 14501 18291 14535
rect 18233 14495 18291 14501
rect 12894 14464 12900 14476
rect 12023 14436 12434 14464
rect 12855 14436 12900 14464
rect 12023 14433 12035 14436
rect 11977 14427 12035 14433
rect 12894 14424 12900 14436
rect 12952 14424 12958 14476
rect 12986 14424 12992 14476
rect 13044 14464 13050 14476
rect 13909 14467 13967 14473
rect 13044 14436 13089 14464
rect 13044 14424 13050 14436
rect 13909 14433 13921 14467
rect 13955 14464 13967 14467
rect 14274 14464 14280 14476
rect 13955 14436 14280 14464
rect 13955 14433 13967 14436
rect 13909 14427 13967 14433
rect 14274 14424 14280 14436
rect 14332 14424 14338 14476
rect 15473 14467 15531 14473
rect 15473 14433 15485 14467
rect 15519 14433 15531 14467
rect 15473 14427 15531 14433
rect 15627 14467 15685 14473
rect 15627 14433 15639 14467
rect 15673 14464 15685 14467
rect 15746 14464 15752 14476
rect 15673 14436 15752 14464
rect 15673 14433 15685 14436
rect 15627 14427 15685 14433
rect 11057 14399 11115 14405
rect 11057 14365 11069 14399
rect 11103 14396 11115 14399
rect 12250 14396 12256 14408
rect 11103 14368 12256 14396
rect 11103 14365 11115 14368
rect 11057 14359 11115 14365
rect 12250 14356 12256 14368
rect 12308 14356 12314 14408
rect 14093 14399 14151 14405
rect 14093 14365 14105 14399
rect 14139 14396 14151 14399
rect 15194 14396 15200 14408
rect 14139 14368 15200 14396
rect 14139 14365 14151 14368
rect 14093 14359 14151 14365
rect 12894 14288 12900 14340
rect 12952 14328 12958 14340
rect 13906 14328 13912 14340
rect 12952 14300 13912 14328
rect 12952 14288 12958 14300
rect 13906 14288 13912 14300
rect 13964 14328 13970 14340
rect 14108 14328 14136 14359
rect 15194 14356 15200 14368
rect 15252 14396 15258 14408
rect 15488 14396 15516 14427
rect 15746 14424 15752 14436
rect 15804 14424 15810 14476
rect 15930 14424 15936 14476
rect 15988 14464 15994 14476
rect 16390 14464 16396 14476
rect 15988 14436 16396 14464
rect 15988 14424 15994 14436
rect 16390 14424 16396 14436
rect 16448 14424 16454 14476
rect 16574 14424 16580 14476
rect 16632 14464 16638 14476
rect 16669 14467 16727 14473
rect 16669 14464 16681 14467
rect 16632 14436 16681 14464
rect 16632 14424 16638 14436
rect 16669 14433 16681 14436
rect 16715 14464 16727 14467
rect 16942 14464 16948 14476
rect 16715 14436 16948 14464
rect 16715 14433 16727 14436
rect 16669 14427 16727 14433
rect 16942 14424 16948 14436
rect 17000 14424 17006 14476
rect 15252 14368 15516 14396
rect 16117 14399 16175 14405
rect 15252 14356 15258 14368
rect 16117 14365 16129 14399
rect 16163 14365 16175 14399
rect 16117 14359 16175 14365
rect 13964 14300 14136 14328
rect 13964 14288 13970 14300
rect 14642 14288 14648 14340
rect 14700 14328 14706 14340
rect 16132 14328 16160 14359
rect 16298 14356 16304 14408
rect 16356 14396 16362 14408
rect 17773 14399 17831 14405
rect 16356 14368 16401 14396
rect 16356 14356 16362 14368
rect 17773 14365 17785 14399
rect 17819 14396 17831 14399
rect 17954 14396 17960 14408
rect 17819 14368 17960 14396
rect 17819 14365 17831 14368
rect 17773 14359 17831 14365
rect 17954 14356 17960 14368
rect 18012 14356 18018 14408
rect 17494 14328 17500 14340
rect 14700 14300 17500 14328
rect 14700 14288 14706 14300
rect 17494 14288 17500 14300
rect 17552 14328 17558 14340
rect 18049 14331 18107 14337
rect 18049 14328 18061 14331
rect 17552 14300 18061 14328
rect 17552 14288 17558 14300
rect 18049 14297 18061 14300
rect 18095 14297 18107 14331
rect 18049 14291 18107 14297
rect 10042 14260 10048 14272
rect 9180 14232 9444 14260
rect 10003 14232 10048 14260
rect 9180 14220 9186 14232
rect 10042 14220 10048 14232
rect 10100 14220 10106 14272
rect 11241 14263 11299 14269
rect 11241 14229 11253 14263
rect 11287 14260 11299 14263
rect 11330 14260 11336 14272
rect 11287 14232 11336 14260
rect 11287 14229 11299 14232
rect 11241 14223 11299 14229
rect 11330 14220 11336 14232
rect 11388 14220 11394 14272
rect 13538 14260 13544 14272
rect 13499 14232 13544 14260
rect 13538 14220 13544 14232
rect 13596 14220 13602 14272
rect 15286 14220 15292 14272
rect 15344 14260 15350 14272
rect 15657 14263 15715 14269
rect 15657 14260 15669 14263
rect 15344 14232 15669 14260
rect 15344 14220 15350 14232
rect 15657 14229 15669 14232
rect 15703 14229 15715 14263
rect 15657 14223 15715 14229
rect 15746 14220 15752 14272
rect 15804 14260 15810 14272
rect 16114 14260 16120 14272
rect 15804 14232 16120 14260
rect 15804 14220 15810 14232
rect 16114 14220 16120 14232
rect 16172 14260 16178 14272
rect 16209 14263 16267 14269
rect 16209 14260 16221 14263
rect 16172 14232 16221 14260
rect 16172 14220 16178 14232
rect 16209 14229 16221 14232
rect 16255 14229 16267 14263
rect 16209 14223 16267 14229
rect 184 14170 18860 14192
rect 184 14118 1556 14170
rect 1608 14118 1620 14170
rect 1672 14118 1684 14170
rect 1736 14118 1748 14170
rect 1800 14118 1812 14170
rect 1864 14118 4656 14170
rect 4708 14118 4720 14170
rect 4772 14118 4784 14170
rect 4836 14118 4848 14170
rect 4900 14118 4912 14170
rect 4964 14118 7756 14170
rect 7808 14118 7820 14170
rect 7872 14118 7884 14170
rect 7936 14118 7948 14170
rect 8000 14118 8012 14170
rect 8064 14118 10856 14170
rect 10908 14118 10920 14170
rect 10972 14118 10984 14170
rect 11036 14118 11048 14170
rect 11100 14118 11112 14170
rect 11164 14118 13956 14170
rect 14008 14118 14020 14170
rect 14072 14118 14084 14170
rect 14136 14118 14148 14170
rect 14200 14118 14212 14170
rect 14264 14118 17056 14170
rect 17108 14118 17120 14170
rect 17172 14118 17184 14170
rect 17236 14118 17248 14170
rect 17300 14118 17312 14170
rect 17364 14118 18860 14170
rect 184 14096 18860 14118
rect 3878 14016 3884 14068
rect 3936 14056 3942 14068
rect 5077 14059 5135 14065
rect 5077 14056 5089 14059
rect 3936 14028 5089 14056
rect 3936 14016 3942 14028
rect 5077 14025 5089 14028
rect 5123 14056 5135 14059
rect 5626 14056 5632 14068
rect 5123 14028 5632 14056
rect 5123 14025 5135 14028
rect 5077 14019 5135 14025
rect 5626 14016 5632 14028
rect 5684 14016 5690 14068
rect 6914 14016 6920 14068
rect 6972 14056 6978 14068
rect 7009 14059 7067 14065
rect 7009 14056 7021 14059
rect 6972 14028 7021 14056
rect 6972 14016 6978 14028
rect 7009 14025 7021 14028
rect 7055 14025 7067 14059
rect 8202 14056 8208 14068
rect 7009 14019 7067 14025
rect 7300 14028 8208 14056
rect 3142 13948 3148 14000
rect 3200 13988 3206 14000
rect 7300 13988 7328 14028
rect 8202 14016 8208 14028
rect 8260 14056 8266 14068
rect 10505 14059 10563 14065
rect 10505 14056 10517 14059
rect 8260 14028 10517 14056
rect 8260 14016 8266 14028
rect 10505 14025 10517 14028
rect 10551 14025 10563 14059
rect 13814 14056 13820 14068
rect 10505 14019 10563 14025
rect 13740 14028 13820 14056
rect 3200 13960 7328 13988
rect 3200 13948 3206 13960
rect 5718 13880 5724 13932
rect 5776 13920 5782 13932
rect 6365 13923 6423 13929
rect 6365 13920 6377 13923
rect 5776 13892 6377 13920
rect 5776 13880 5782 13892
rect 6365 13889 6377 13892
rect 6411 13889 6423 13923
rect 6365 13883 6423 13889
rect 8757 13923 8815 13929
rect 8757 13889 8769 13923
rect 8803 13920 8815 13923
rect 9122 13920 9128 13932
rect 8803 13892 9128 13920
rect 8803 13889 8815 13892
rect 8757 13883 8815 13889
rect 9122 13880 9128 13892
rect 9180 13880 9186 13932
rect 10042 13880 10048 13932
rect 10100 13920 10106 13932
rect 13740 13929 13768 14028
rect 13814 14016 13820 14028
rect 13872 14016 13878 14068
rect 14274 14056 14280 14068
rect 14235 14028 14280 14056
rect 14274 14016 14280 14028
rect 14332 14016 14338 14068
rect 15194 14056 15200 14068
rect 15155 14028 15200 14056
rect 15194 14016 15200 14028
rect 15252 14016 15258 14068
rect 17954 14056 17960 14068
rect 15304 14028 17540 14056
rect 17915 14028 17960 14056
rect 13725 13923 13783 13929
rect 10100 13892 13676 13920
rect 10100 13880 10106 13892
rect 2222 13812 2228 13864
rect 2280 13852 2286 13864
rect 2869 13855 2927 13861
rect 2869 13852 2881 13855
rect 2280 13824 2881 13852
rect 2280 13812 2286 13824
rect 2869 13821 2881 13824
rect 2915 13821 2927 13855
rect 2869 13815 2927 13821
rect 5626 13812 5632 13864
rect 5684 13852 5690 13864
rect 7377 13855 7435 13861
rect 7377 13852 7389 13855
rect 5684 13824 7389 13852
rect 5684 13812 5690 13824
rect 7377 13821 7389 13824
rect 7423 13852 7435 13855
rect 7742 13852 7748 13864
rect 7423 13824 7748 13852
rect 7423 13821 7435 13824
rect 7377 13815 7435 13821
rect 7742 13812 7748 13824
rect 7800 13852 7806 13864
rect 8294 13852 8300 13864
rect 7800 13824 8300 13852
rect 7800 13812 7806 13824
rect 8294 13812 8300 13824
rect 8352 13812 8358 13864
rect 11333 13855 11391 13861
rect 11333 13821 11345 13855
rect 11379 13852 11391 13855
rect 13538 13852 13544 13864
rect 11379 13824 13544 13852
rect 11379 13821 11391 13824
rect 11333 13815 11391 13821
rect 13538 13812 13544 13824
rect 13596 13812 13602 13864
rect 13648 13852 13676 13892
rect 13725 13889 13737 13923
rect 13771 13889 13783 13923
rect 13725 13883 13783 13889
rect 13817 13923 13875 13929
rect 13817 13889 13829 13923
rect 13863 13920 13875 13923
rect 14366 13920 14372 13932
rect 13863 13892 14372 13920
rect 13863 13889 13875 13892
rect 13817 13883 13875 13889
rect 14366 13880 14372 13892
rect 14424 13880 14430 13932
rect 15304 13920 15332 14028
rect 17512 13988 17540 14028
rect 17954 14016 17960 14028
rect 18012 14016 18018 14068
rect 18046 13988 18052 14000
rect 17512 13960 18052 13988
rect 18046 13948 18052 13960
rect 18104 13948 18110 14000
rect 14476 13892 15332 13920
rect 16485 13923 16543 13929
rect 14476 13852 14504 13892
rect 16485 13889 16497 13923
rect 16531 13920 16543 13923
rect 18230 13920 18236 13932
rect 16531 13892 18236 13920
rect 16531 13889 16543 13892
rect 16485 13883 16543 13889
rect 18230 13880 18236 13892
rect 18288 13880 18294 13932
rect 14734 13852 14740 13864
rect 13648 13824 14504 13852
rect 14695 13824 14740 13852
rect 14734 13812 14740 13824
rect 14792 13812 14798 13864
rect 15473 13855 15531 13861
rect 15473 13821 15485 13855
rect 15519 13852 15531 13855
rect 15838 13852 15844 13864
rect 15519 13824 15844 13852
rect 15519 13821 15531 13824
rect 15473 13815 15531 13821
rect 15838 13812 15844 13824
rect 15896 13812 15902 13864
rect 16206 13852 16212 13864
rect 16167 13824 16212 13852
rect 16206 13812 16212 13824
rect 16264 13812 16270 13864
rect 17586 13812 17592 13864
rect 17644 13812 17650 13864
rect 2958 13676 2964 13728
rect 3016 13716 3022 13728
rect 3053 13719 3111 13725
rect 3053 13716 3065 13719
rect 3016 13688 3065 13716
rect 3016 13676 3022 13688
rect 3053 13685 3065 13688
rect 3099 13685 3111 13719
rect 8312 13716 8340 13812
rect 8386 13744 8392 13796
rect 8444 13784 8450 13796
rect 9033 13787 9091 13793
rect 9033 13784 9045 13787
rect 8444 13756 9045 13784
rect 8444 13744 8450 13756
rect 9033 13753 9045 13756
rect 9079 13753 9091 13787
rect 13909 13787 13967 13793
rect 9033 13747 9091 13753
rect 9140 13756 9522 13784
rect 9140 13716 9168 13756
rect 8312 13688 9168 13716
rect 9416 13716 9444 13756
rect 13909 13753 13921 13787
rect 13955 13784 13967 13787
rect 14553 13787 14611 13793
rect 14553 13784 14565 13787
rect 13955 13756 14565 13784
rect 13955 13753 13967 13756
rect 13909 13747 13967 13753
rect 14553 13753 14565 13756
rect 14599 13753 14611 13787
rect 14553 13747 14611 13753
rect 9674 13716 9680 13728
rect 9416 13688 9680 13716
rect 3053 13679 3111 13685
rect 9674 13676 9680 13688
rect 9732 13676 9738 13728
rect 11238 13716 11244 13728
rect 11199 13688 11244 13716
rect 11238 13676 11244 13688
rect 11296 13676 11302 13728
rect 184 13626 18920 13648
rect 184 13574 3106 13626
rect 3158 13574 3170 13626
rect 3222 13574 3234 13626
rect 3286 13574 3298 13626
rect 3350 13574 3362 13626
rect 3414 13574 6206 13626
rect 6258 13574 6270 13626
rect 6322 13574 6334 13626
rect 6386 13574 6398 13626
rect 6450 13574 6462 13626
rect 6514 13574 9306 13626
rect 9358 13574 9370 13626
rect 9422 13574 9434 13626
rect 9486 13574 9498 13626
rect 9550 13574 9562 13626
rect 9614 13574 12406 13626
rect 12458 13574 12470 13626
rect 12522 13574 12534 13626
rect 12586 13574 12598 13626
rect 12650 13574 12662 13626
rect 12714 13574 15506 13626
rect 15558 13574 15570 13626
rect 15622 13574 15634 13626
rect 15686 13574 15698 13626
rect 15750 13574 15762 13626
rect 15814 13574 18606 13626
rect 18658 13574 18670 13626
rect 18722 13574 18734 13626
rect 18786 13574 18798 13626
rect 18850 13574 18862 13626
rect 18914 13574 18920 13626
rect 184 13552 18920 13574
rect 3237 13515 3295 13521
rect 3237 13512 3249 13515
rect 2746 13484 3249 13512
rect 2314 13444 2320 13456
rect 1978 13416 2320 13444
rect 2314 13404 2320 13416
rect 2372 13404 2378 13456
rect 566 13376 572 13388
rect 527 13348 572 13376
rect 566 13336 572 13348
rect 624 13376 630 13388
rect 624 13348 1072 13376
rect 624 13336 630 13348
rect 934 13308 940 13320
rect 895 13280 940 13308
rect 934 13268 940 13280
rect 992 13268 998 13320
rect 1044 13308 1072 13348
rect 2222 13336 2228 13388
rect 2280 13376 2286 13388
rect 2409 13379 2467 13385
rect 2409 13376 2421 13379
rect 2280 13348 2421 13376
rect 2280 13336 2286 13348
rect 2409 13345 2421 13348
rect 2455 13345 2467 13379
rect 2409 13339 2467 13345
rect 2746 13320 2774 13484
rect 3237 13481 3249 13484
rect 3283 13512 3295 13515
rect 5166 13512 5172 13524
rect 3283 13484 5172 13512
rect 3283 13481 3295 13484
rect 3237 13475 3295 13481
rect 5166 13472 5172 13484
rect 5224 13472 5230 13524
rect 5261 13515 5319 13521
rect 5261 13481 5273 13515
rect 5307 13512 5319 13515
rect 5718 13512 5724 13524
rect 5307 13484 5724 13512
rect 5307 13481 5319 13484
rect 5261 13475 5319 13481
rect 5718 13472 5724 13484
rect 5776 13472 5782 13524
rect 7561 13515 7619 13521
rect 7561 13481 7573 13515
rect 7607 13512 7619 13515
rect 8386 13512 8392 13524
rect 7607 13484 8392 13512
rect 7607 13481 7619 13484
rect 7561 13475 7619 13481
rect 8386 13472 8392 13484
rect 8444 13472 8450 13524
rect 13081 13515 13139 13521
rect 13081 13481 13093 13515
rect 13127 13512 13139 13515
rect 13814 13512 13820 13524
rect 13127 13484 13820 13512
rect 13127 13481 13139 13484
rect 13081 13475 13139 13481
rect 6638 13404 6644 13456
rect 6696 13444 6702 13456
rect 6696 13416 7052 13444
rect 6696 13404 6702 13416
rect 4522 13376 4528 13388
rect 4483 13348 4528 13376
rect 4522 13336 4528 13348
rect 4580 13336 4586 13388
rect 5626 13336 5632 13388
rect 5684 13336 5690 13388
rect 2746 13308 2780 13320
rect 1044 13280 2780 13308
rect 2774 13268 2780 13280
rect 2832 13268 2838 13320
rect 6730 13308 6736 13320
rect 6691 13280 6736 13308
rect 6730 13268 6736 13280
rect 6788 13268 6794 13320
rect 7024 13317 7052 13416
rect 7742 13404 7748 13456
rect 7800 13444 7806 13456
rect 7800 13416 7866 13444
rect 7800 13404 7806 13416
rect 9950 13336 9956 13388
rect 10008 13376 10014 13388
rect 10226 13376 10232 13388
rect 10008 13348 10232 13376
rect 10008 13336 10014 13348
rect 10226 13336 10232 13348
rect 10284 13336 10290 13388
rect 11606 13336 11612 13388
rect 11664 13336 11670 13388
rect 7009 13311 7067 13317
rect 7009 13277 7021 13311
rect 7055 13308 7067 13311
rect 7650 13308 7656 13320
rect 7055 13280 7656 13308
rect 7055 13277 7067 13280
rect 7009 13271 7067 13277
rect 7650 13268 7656 13280
rect 7708 13268 7714 13320
rect 8938 13268 8944 13320
rect 8996 13308 9002 13320
rect 9033 13311 9091 13317
rect 9033 13308 9045 13311
rect 8996 13280 9045 13308
rect 8996 13268 9002 13280
rect 9033 13277 9045 13280
rect 9079 13277 9091 13311
rect 9306 13308 9312 13320
rect 9267 13280 9312 13308
rect 9033 13271 9091 13277
rect 9306 13268 9312 13280
rect 9364 13268 9370 13320
rect 10502 13308 10508 13320
rect 10463 13280 10508 13308
rect 10502 13268 10508 13280
rect 10560 13268 10566 13320
rect 13096 13240 13124 13475
rect 13814 13472 13820 13484
rect 13872 13512 13878 13524
rect 14918 13512 14924 13524
rect 13872 13484 14924 13512
rect 13872 13472 13878 13484
rect 14918 13472 14924 13484
rect 14976 13512 14982 13524
rect 14976 13484 16160 13512
rect 14976 13472 14982 13484
rect 15010 13444 15016 13456
rect 14971 13416 15016 13444
rect 15010 13404 15016 13416
rect 15068 13404 15074 13456
rect 16132 13444 16160 13484
rect 16206 13472 16212 13524
rect 16264 13512 16270 13524
rect 16301 13515 16359 13521
rect 16301 13512 16313 13515
rect 16264 13484 16313 13512
rect 16264 13472 16270 13484
rect 16301 13481 16313 13484
rect 16347 13481 16359 13515
rect 16301 13475 16359 13481
rect 16574 13444 16580 13456
rect 16132 13416 16580 13444
rect 16574 13404 16580 13416
rect 16632 13444 16638 13456
rect 17773 13447 17831 13453
rect 17773 13444 17785 13447
rect 16632 13416 17785 13444
rect 16632 13404 16638 13416
rect 17773 13413 17785 13416
rect 17819 13413 17831 13447
rect 17773 13407 17831 13413
rect 14366 13376 14372 13388
rect 14327 13348 14372 13376
rect 14366 13336 14372 13348
rect 14424 13336 14430 13388
rect 17678 13376 17684 13388
rect 17639 13348 17684 13376
rect 17678 13336 17684 13348
rect 17736 13336 17742 13388
rect 17586 13268 17592 13320
rect 17644 13308 17650 13320
rect 17865 13311 17923 13317
rect 17865 13308 17877 13311
rect 17644 13280 17877 13308
rect 17644 13268 17650 13280
rect 17865 13277 17877 13280
rect 17911 13277 17923 13311
rect 17865 13271 17923 13277
rect 11532 13212 13124 13240
rect 10226 13132 10232 13184
rect 10284 13172 10290 13184
rect 11532 13172 11560 13212
rect 10284 13144 11560 13172
rect 11977 13175 12035 13181
rect 10284 13132 10290 13144
rect 11977 13141 11989 13175
rect 12023 13172 12035 13175
rect 12434 13172 12440 13184
rect 12023 13144 12440 13172
rect 12023 13141 12035 13144
rect 11977 13135 12035 13141
rect 12434 13132 12440 13144
rect 12492 13172 12498 13184
rect 14734 13172 14740 13184
rect 12492 13144 14740 13172
rect 12492 13132 12498 13144
rect 14734 13132 14740 13144
rect 14792 13132 14798 13184
rect 17313 13175 17371 13181
rect 17313 13141 17325 13175
rect 17359 13172 17371 13175
rect 17402 13172 17408 13184
rect 17359 13144 17408 13172
rect 17359 13141 17371 13144
rect 17313 13135 17371 13141
rect 17402 13132 17408 13144
rect 17460 13132 17466 13184
rect 184 13082 18860 13104
rect 184 13030 1556 13082
rect 1608 13030 1620 13082
rect 1672 13030 1684 13082
rect 1736 13030 1748 13082
rect 1800 13030 1812 13082
rect 1864 13030 4656 13082
rect 4708 13030 4720 13082
rect 4772 13030 4784 13082
rect 4836 13030 4848 13082
rect 4900 13030 4912 13082
rect 4964 13030 7756 13082
rect 7808 13030 7820 13082
rect 7872 13030 7884 13082
rect 7936 13030 7948 13082
rect 8000 13030 8012 13082
rect 8064 13030 10856 13082
rect 10908 13030 10920 13082
rect 10972 13030 10984 13082
rect 11036 13030 11048 13082
rect 11100 13030 11112 13082
rect 11164 13030 13956 13082
rect 14008 13030 14020 13082
rect 14072 13030 14084 13082
rect 14136 13030 14148 13082
rect 14200 13030 14212 13082
rect 14264 13030 17056 13082
rect 17108 13030 17120 13082
rect 17172 13030 17184 13082
rect 17236 13030 17248 13082
rect 17300 13030 17312 13082
rect 17364 13030 18860 13082
rect 184 13008 18860 13030
rect 934 12928 940 12980
rect 992 12968 998 12980
rect 1581 12971 1639 12977
rect 1581 12968 1593 12971
rect 992 12940 1593 12968
rect 992 12928 998 12940
rect 1581 12937 1593 12940
rect 1627 12937 1639 12971
rect 1581 12931 1639 12937
rect 11241 12971 11299 12977
rect 11241 12937 11253 12971
rect 11287 12968 11299 12971
rect 11330 12968 11336 12980
rect 11287 12940 11336 12968
rect 11287 12937 11299 12940
rect 11241 12931 11299 12937
rect 11330 12928 11336 12940
rect 11388 12928 11394 12980
rect 15930 12928 15936 12980
rect 15988 12968 15994 12980
rect 16390 12968 16396 12980
rect 15988 12940 16396 12968
rect 15988 12928 15994 12940
rect 16390 12928 16396 12940
rect 16448 12928 16454 12980
rect 16482 12928 16488 12980
rect 16540 12968 16546 12980
rect 16761 12971 16819 12977
rect 16761 12968 16773 12971
rect 16540 12940 16773 12968
rect 16540 12928 16546 12940
rect 16761 12937 16773 12940
rect 16807 12937 16819 12971
rect 16761 12931 16819 12937
rect 16942 12928 16948 12980
rect 17000 12968 17006 12980
rect 17957 12971 18015 12977
rect 17957 12968 17969 12971
rect 17000 12940 17969 12968
rect 17000 12928 17006 12940
rect 17957 12937 17969 12940
rect 18003 12937 18015 12971
rect 17957 12931 18015 12937
rect 8938 12860 8944 12912
rect 8996 12900 9002 12912
rect 12526 12900 12532 12912
rect 8996 12872 12532 12900
rect 8996 12860 9002 12872
rect 12526 12860 12532 12872
rect 12584 12860 12590 12912
rect 12710 12860 12716 12912
rect 12768 12900 12774 12912
rect 18138 12900 18144 12912
rect 12768 12872 18144 12900
rect 12768 12860 12774 12872
rect 18138 12860 18144 12872
rect 18196 12860 18202 12912
rect 2130 12832 2136 12844
rect 2091 12804 2136 12832
rect 2130 12792 2136 12804
rect 2188 12792 2194 12844
rect 2958 12792 2964 12844
rect 3016 12832 3022 12844
rect 3237 12835 3295 12841
rect 3237 12832 3249 12835
rect 3016 12804 3249 12832
rect 3016 12792 3022 12804
rect 3237 12801 3249 12804
rect 3283 12801 3295 12835
rect 3237 12795 3295 12801
rect 3421 12835 3479 12841
rect 3421 12801 3433 12835
rect 3467 12832 3479 12835
rect 3510 12832 3516 12844
rect 3467 12804 3516 12832
rect 3467 12801 3479 12804
rect 3421 12795 3479 12801
rect 3510 12792 3516 12804
rect 3568 12792 3574 12844
rect 7466 12792 7472 12844
rect 7524 12832 7530 12844
rect 7561 12835 7619 12841
rect 7561 12832 7573 12835
rect 7524 12804 7573 12832
rect 7524 12792 7530 12804
rect 7561 12801 7573 12804
rect 7607 12801 7619 12835
rect 7561 12795 7619 12801
rect 7650 12792 7656 12844
rect 7708 12832 7714 12844
rect 7745 12835 7803 12841
rect 7745 12832 7757 12835
rect 7708 12804 7757 12832
rect 7708 12792 7714 12804
rect 7745 12801 7757 12804
rect 7791 12801 7803 12835
rect 7745 12795 7803 12801
rect 11425 12835 11483 12841
rect 11425 12801 11437 12835
rect 11471 12832 11483 12835
rect 12345 12835 12403 12841
rect 12345 12832 12357 12835
rect 11471 12804 12357 12832
rect 11471 12801 11483 12804
rect 11425 12795 11483 12801
rect 12345 12801 12357 12804
rect 12391 12801 12403 12835
rect 12345 12795 12403 12801
rect 12434 12792 12440 12844
rect 12492 12832 12498 12844
rect 12492 12804 12664 12832
rect 12492 12792 12498 12804
rect 2041 12767 2099 12773
rect 2041 12733 2053 12767
rect 2087 12764 2099 12767
rect 2222 12764 2228 12776
rect 2087 12736 2228 12764
rect 2087 12733 2099 12736
rect 2041 12727 2099 12733
rect 2222 12724 2228 12736
rect 2280 12724 2286 12776
rect 4433 12767 4491 12773
rect 4433 12733 4445 12767
rect 4479 12764 4491 12767
rect 5166 12764 5172 12776
rect 4479 12736 5172 12764
rect 4479 12733 4491 12736
rect 4433 12727 4491 12733
rect 5166 12724 5172 12736
rect 5224 12724 5230 12776
rect 7006 12724 7012 12776
rect 7064 12764 7070 12776
rect 7837 12767 7895 12773
rect 7837 12764 7849 12767
rect 7064 12736 7849 12764
rect 7064 12724 7070 12736
rect 7837 12733 7849 12736
rect 7883 12733 7895 12767
rect 11146 12764 11152 12776
rect 11107 12736 11152 12764
rect 7837 12727 7895 12733
rect 11146 12724 11152 12736
rect 11204 12724 11210 12776
rect 12526 12764 12532 12776
rect 12487 12736 12532 12764
rect 12526 12724 12532 12736
rect 12584 12724 12590 12776
rect 12636 12773 12664 12804
rect 12986 12792 12992 12844
rect 13044 12832 13050 12844
rect 13909 12835 13967 12841
rect 13909 12832 13921 12835
rect 13044 12804 13921 12832
rect 13044 12792 13050 12804
rect 13909 12801 13921 12804
rect 13955 12801 13967 12835
rect 13909 12795 13967 12801
rect 17221 12835 17279 12841
rect 17221 12801 17233 12835
rect 17267 12832 17279 12835
rect 17402 12832 17408 12844
rect 17267 12804 17408 12832
rect 17267 12801 17279 12804
rect 17221 12795 17279 12801
rect 17402 12792 17408 12804
rect 17460 12792 17466 12844
rect 12621 12767 12679 12773
rect 12621 12733 12633 12767
rect 12667 12733 12679 12767
rect 12621 12727 12679 12733
rect 12713 12767 12771 12773
rect 12713 12733 12725 12767
rect 12759 12764 12771 12767
rect 12894 12764 12900 12776
rect 12759 12736 12900 12764
rect 12759 12733 12771 12736
rect 12713 12727 12771 12733
rect 12894 12724 12900 12736
rect 12952 12724 12958 12776
rect 13998 12724 14004 12776
rect 14056 12764 14062 12776
rect 14185 12767 14243 12773
rect 14185 12764 14197 12767
rect 14056 12736 14197 12764
rect 14056 12724 14062 12736
rect 14185 12733 14197 12736
rect 14231 12733 14243 12767
rect 14642 12764 14648 12776
rect 14603 12736 14648 12764
rect 14185 12727 14243 12733
rect 14642 12724 14648 12736
rect 14700 12724 14706 12776
rect 14826 12764 14832 12776
rect 14787 12736 14832 12764
rect 14826 12724 14832 12736
rect 14884 12724 14890 12776
rect 15289 12767 15347 12773
rect 15289 12733 15301 12767
rect 15335 12764 15347 12767
rect 15930 12764 15936 12776
rect 15335 12736 15936 12764
rect 15335 12733 15347 12736
rect 15289 12727 15347 12733
rect 15930 12724 15936 12736
rect 15988 12724 15994 12776
rect 16025 12767 16083 12773
rect 16025 12733 16037 12767
rect 16071 12733 16083 12767
rect 16025 12727 16083 12733
rect 1949 12699 2007 12705
rect 1949 12665 1961 12699
rect 1995 12696 2007 12699
rect 3145 12699 3203 12705
rect 1995 12668 2820 12696
rect 1995 12665 2007 12668
rect 1949 12659 2007 12665
rect 2792 12637 2820 12668
rect 3145 12665 3157 12699
rect 3191 12696 3203 12699
rect 3694 12696 3700 12708
rect 3191 12668 3700 12696
rect 3191 12665 3203 12668
rect 3145 12659 3203 12665
rect 3694 12656 3700 12668
rect 3752 12656 3758 12708
rect 4700 12699 4758 12705
rect 4700 12665 4712 12699
rect 4746 12696 4758 12699
rect 4982 12696 4988 12708
rect 4746 12668 4988 12696
rect 4746 12665 4758 12668
rect 4700 12659 4758 12665
rect 4982 12656 4988 12668
rect 5040 12656 5046 12708
rect 6730 12656 6736 12708
rect 6788 12696 6794 12708
rect 7193 12699 7251 12705
rect 7193 12696 7205 12699
rect 6788 12668 7205 12696
rect 6788 12656 6794 12668
rect 7193 12665 7205 12668
rect 7239 12696 7251 12699
rect 7239 12668 8800 12696
rect 7239 12665 7251 12668
rect 7193 12659 7251 12665
rect 2777 12631 2835 12637
rect 2777 12597 2789 12631
rect 2823 12597 2835 12631
rect 5810 12628 5816 12640
rect 5771 12600 5816 12628
rect 2777 12591 2835 12597
rect 5810 12588 5816 12600
rect 5868 12588 5874 12640
rect 8110 12588 8116 12640
rect 8168 12628 8174 12640
rect 8205 12631 8263 12637
rect 8205 12628 8217 12631
rect 8168 12600 8217 12628
rect 8168 12588 8174 12600
rect 8205 12597 8217 12600
rect 8251 12597 8263 12631
rect 8772 12628 8800 12668
rect 10502 12656 10508 12708
rect 10560 12696 10566 12708
rect 11425 12699 11483 12705
rect 11425 12696 11437 12699
rect 10560 12668 11437 12696
rect 10560 12656 10566 12668
rect 11425 12665 11437 12668
rect 11471 12665 11483 12699
rect 16040 12696 16068 12727
rect 16114 12724 16120 12776
rect 16172 12764 16178 12776
rect 16209 12767 16267 12773
rect 16209 12764 16221 12767
rect 16172 12736 16221 12764
rect 16172 12724 16178 12736
rect 16209 12733 16221 12736
rect 16255 12733 16267 12767
rect 16209 12727 16267 12733
rect 16298 12724 16304 12776
rect 16356 12764 16362 12776
rect 16393 12767 16451 12773
rect 16393 12764 16405 12767
rect 16356 12736 16405 12764
rect 16356 12724 16362 12736
rect 16393 12733 16405 12736
rect 16439 12733 16451 12767
rect 17494 12764 17500 12776
rect 17455 12736 17500 12764
rect 16393 12727 16451 12733
rect 17494 12724 17500 12736
rect 17552 12724 17558 12776
rect 16666 12696 16672 12708
rect 11425 12659 11483 12665
rect 12406 12668 15332 12696
rect 16040 12668 16672 12696
rect 12406 12628 12434 12668
rect 8772 12600 12434 12628
rect 8205 12591 8263 12597
rect 12526 12588 12532 12640
rect 12584 12628 12590 12640
rect 12802 12628 12808 12640
rect 12584 12600 12808 12628
rect 12584 12588 12590 12600
rect 12802 12588 12808 12600
rect 12860 12628 12866 12640
rect 12986 12628 12992 12640
rect 12860 12600 12992 12628
rect 12860 12588 12866 12600
rect 12986 12588 12992 12600
rect 13044 12588 13050 12640
rect 15304 12628 15332 12668
rect 16666 12656 16672 12668
rect 16724 12656 16730 12708
rect 16761 12699 16819 12705
rect 16761 12665 16773 12699
rect 16807 12696 16819 12699
rect 17313 12699 17371 12705
rect 17313 12696 17325 12699
rect 16807 12668 17325 12696
rect 16807 12665 16819 12668
rect 16761 12659 16819 12665
rect 17313 12665 17325 12668
rect 17359 12665 17371 12699
rect 18322 12696 18328 12708
rect 17313 12659 17371 12665
rect 17420 12668 18328 12696
rect 17420 12628 17448 12668
rect 18322 12656 18328 12668
rect 18380 12656 18386 12708
rect 15304 12600 17448 12628
rect 184 12538 18920 12560
rect 184 12486 3106 12538
rect 3158 12486 3170 12538
rect 3222 12486 3234 12538
rect 3286 12486 3298 12538
rect 3350 12486 3362 12538
rect 3414 12486 6206 12538
rect 6258 12486 6270 12538
rect 6322 12486 6334 12538
rect 6386 12486 6398 12538
rect 6450 12486 6462 12538
rect 6514 12486 9306 12538
rect 9358 12486 9370 12538
rect 9422 12486 9434 12538
rect 9486 12486 9498 12538
rect 9550 12486 9562 12538
rect 9614 12486 12406 12538
rect 12458 12486 12470 12538
rect 12522 12486 12534 12538
rect 12586 12486 12598 12538
rect 12650 12486 12662 12538
rect 12714 12486 15506 12538
rect 15558 12486 15570 12538
rect 15622 12486 15634 12538
rect 15686 12486 15698 12538
rect 15750 12486 15762 12538
rect 15814 12486 18606 12538
rect 18658 12486 18670 12538
rect 18722 12486 18734 12538
rect 18786 12486 18798 12538
rect 18850 12486 18862 12538
rect 18914 12486 18920 12538
rect 184 12464 18920 12486
rect 8018 12384 8024 12436
rect 8076 12424 8082 12436
rect 9490 12424 9496 12436
rect 8076 12396 9496 12424
rect 8076 12384 8082 12396
rect 9490 12384 9496 12396
rect 9548 12384 9554 12436
rect 12894 12424 12900 12436
rect 11164 12396 12900 12424
rect 3620 12328 5396 12356
rect 3620 12300 3648 12328
rect 2041 12291 2099 12297
rect 2041 12257 2053 12291
rect 2087 12288 2099 12291
rect 2774 12288 2780 12300
rect 2087 12260 2780 12288
rect 2087 12257 2099 12260
rect 2041 12251 2099 12257
rect 2774 12248 2780 12260
rect 2832 12288 2838 12300
rect 3602 12297 3608 12300
rect 3329 12291 3387 12297
rect 3329 12288 3341 12291
rect 2832 12260 3341 12288
rect 2832 12248 2838 12260
rect 3329 12257 3341 12260
rect 3375 12257 3387 12291
rect 3596 12288 3608 12297
rect 3563 12260 3608 12288
rect 3329 12251 3387 12257
rect 3596 12251 3608 12260
rect 3602 12248 3608 12251
rect 3660 12248 3666 12300
rect 5258 12288 5264 12300
rect 4724 12260 5264 12288
rect 4724 12161 4752 12260
rect 5258 12248 5264 12260
rect 5316 12248 5322 12300
rect 5368 12297 5396 12328
rect 5810 12316 5816 12368
rect 5868 12356 5874 12368
rect 11164 12365 11192 12396
rect 12894 12384 12900 12396
rect 12952 12424 12958 12436
rect 14182 12424 14188 12436
rect 12952 12396 14188 12424
rect 12952 12384 12958 12396
rect 14182 12384 14188 12396
rect 14240 12384 14246 12436
rect 14277 12427 14335 12433
rect 14277 12393 14289 12427
rect 14323 12424 14335 12427
rect 14642 12424 14648 12436
rect 14323 12396 14648 12424
rect 14323 12393 14335 12396
rect 14277 12387 14335 12393
rect 14642 12384 14648 12396
rect 14700 12384 14706 12436
rect 15562 12384 15568 12436
rect 15620 12424 15626 12436
rect 15657 12427 15715 12433
rect 15657 12424 15669 12427
rect 15620 12396 15669 12424
rect 15620 12384 15626 12396
rect 15657 12393 15669 12396
rect 15703 12424 15715 12427
rect 18506 12424 18512 12436
rect 15703 12396 18512 12424
rect 15703 12393 15715 12396
rect 15657 12387 15715 12393
rect 18506 12384 18512 12396
rect 18564 12384 18570 12436
rect 5905 12359 5963 12365
rect 5905 12356 5917 12359
rect 5868 12328 5917 12356
rect 5868 12316 5874 12328
rect 5905 12325 5917 12328
rect 5951 12325 5963 12359
rect 11149 12359 11207 12365
rect 5905 12319 5963 12325
rect 5354 12291 5412 12297
rect 5354 12257 5366 12291
rect 5400 12257 5412 12291
rect 5354 12251 5412 12257
rect 5629 12291 5687 12297
rect 5629 12257 5641 12291
rect 5675 12288 5687 12291
rect 6089 12291 6147 12297
rect 6089 12288 6101 12291
rect 5675 12260 6101 12288
rect 5675 12257 5687 12260
rect 5629 12251 5687 12257
rect 6089 12257 6101 12260
rect 6135 12257 6147 12291
rect 6089 12251 6147 12257
rect 6181 12291 6239 12297
rect 6181 12257 6193 12291
rect 6227 12257 6239 12291
rect 6181 12251 6239 12257
rect 5534 12180 5540 12232
rect 5592 12220 5598 12232
rect 6196 12220 6224 12251
rect 5592 12192 6224 12220
rect 7193 12223 7251 12229
rect 5592 12180 5598 12192
rect 7193 12189 7205 12223
rect 7239 12220 7251 12223
rect 8496 12220 8524 12342
rect 11149 12325 11161 12359
rect 11195 12325 11207 12359
rect 11149 12319 11207 12325
rect 11333 12359 11391 12365
rect 11333 12325 11345 12359
rect 11379 12356 11391 12359
rect 11882 12356 11888 12368
rect 11379 12328 11888 12356
rect 11379 12325 11391 12328
rect 11333 12319 11391 12325
rect 11882 12316 11888 12328
rect 11940 12356 11946 12368
rect 13909 12359 13967 12365
rect 13909 12356 13921 12359
rect 11940 12328 13921 12356
rect 11940 12316 11946 12328
rect 13909 12325 13921 12328
rect 13955 12356 13967 12359
rect 13998 12356 14004 12368
rect 13955 12328 14004 12356
rect 13955 12325 13967 12328
rect 13909 12319 13967 12325
rect 13998 12316 14004 12328
rect 14056 12356 14062 12368
rect 15010 12356 15016 12368
rect 14056 12328 15016 12356
rect 14056 12316 14062 12328
rect 15010 12316 15016 12328
rect 15068 12316 15074 12368
rect 16298 12356 16304 12368
rect 16259 12328 16304 12356
rect 16298 12316 16304 12328
rect 16356 12316 16362 12368
rect 16666 12356 16672 12368
rect 16627 12328 16672 12356
rect 16666 12316 16672 12328
rect 16724 12316 16730 12368
rect 16942 12316 16948 12368
rect 17000 12356 17006 12368
rect 17129 12359 17187 12365
rect 17129 12356 17141 12359
rect 17000 12328 17141 12356
rect 17000 12316 17006 12328
rect 17129 12325 17141 12328
rect 17175 12325 17187 12359
rect 17586 12356 17592 12368
rect 17547 12328 17592 12356
rect 17129 12319 17187 12325
rect 17586 12316 17592 12328
rect 17644 12316 17650 12368
rect 9122 12248 9128 12300
rect 9180 12288 9186 12300
rect 9217 12291 9275 12297
rect 9217 12288 9229 12291
rect 9180 12260 9229 12288
rect 9180 12248 9186 12260
rect 9217 12257 9229 12260
rect 9263 12257 9275 12291
rect 9217 12251 9275 12257
rect 9306 12248 9312 12300
rect 9364 12288 9370 12300
rect 9585 12291 9643 12297
rect 9585 12288 9597 12291
rect 9364 12260 9597 12288
rect 9364 12248 9370 12260
rect 9585 12257 9597 12260
rect 9631 12257 9643 12291
rect 9585 12251 9643 12257
rect 11425 12291 11483 12297
rect 11425 12257 11437 12291
rect 11471 12257 11483 12291
rect 11425 12251 11483 12257
rect 12529 12291 12587 12297
rect 12529 12257 12541 12291
rect 12575 12288 12587 12291
rect 12802 12288 12808 12300
rect 12575 12260 12808 12288
rect 12575 12257 12587 12260
rect 12529 12251 12587 12257
rect 9674 12220 9680 12232
rect 7239 12192 9680 12220
rect 7239 12189 7251 12192
rect 7193 12183 7251 12189
rect 9674 12180 9680 12192
rect 9732 12180 9738 12232
rect 11440 12220 11468 12251
rect 12802 12248 12808 12260
rect 12860 12248 12866 12300
rect 13722 12288 13728 12300
rect 13635 12260 13728 12288
rect 13722 12248 13728 12260
rect 13780 12288 13786 12300
rect 14108 12288 14320 12292
rect 15105 12291 15163 12297
rect 15105 12288 15117 12291
rect 13780 12264 15117 12288
rect 13780 12260 14136 12264
rect 14292 12260 15117 12264
rect 13780 12248 13786 12260
rect 15105 12257 15117 12260
rect 15151 12257 15163 12291
rect 15105 12251 15163 12257
rect 16117 12291 16175 12297
rect 16117 12257 16129 12291
rect 16163 12288 16175 12291
rect 16206 12288 16212 12300
rect 16163 12260 16212 12288
rect 16163 12257 16175 12260
rect 16117 12251 16175 12257
rect 16206 12248 16212 12260
rect 16264 12288 16270 12300
rect 16577 12291 16635 12297
rect 16577 12288 16589 12291
rect 16264 12260 16589 12288
rect 16264 12248 16270 12260
rect 16577 12257 16589 12260
rect 16623 12257 16635 12291
rect 16577 12251 16635 12257
rect 16761 12291 16819 12297
rect 16761 12257 16773 12291
rect 16807 12257 16819 12291
rect 16761 12251 16819 12257
rect 17497 12291 17555 12297
rect 17497 12257 17509 12291
rect 17543 12257 17555 12291
rect 17497 12251 17555 12257
rect 17681 12291 17739 12297
rect 17681 12257 17693 12291
rect 17727 12288 17739 12291
rect 17862 12288 17868 12300
rect 17727 12260 17868 12288
rect 17727 12257 17739 12260
rect 17681 12251 17739 12257
rect 13998 12220 14004 12232
rect 11440 12192 14004 12220
rect 13998 12180 14004 12192
rect 14056 12180 14062 12232
rect 14090 12223 14148 12229
rect 14090 12189 14102 12223
rect 14136 12189 14148 12223
rect 14090 12183 14148 12189
rect 4709 12155 4767 12161
rect 4709 12121 4721 12155
rect 4755 12121 4767 12155
rect 4709 12115 4767 12121
rect 11149 12155 11207 12161
rect 11149 12121 11161 12155
rect 11195 12152 11207 12155
rect 11330 12152 11336 12164
rect 11195 12124 11336 12152
rect 11195 12121 11207 12124
rect 11149 12115 11207 12121
rect 11330 12112 11336 12124
rect 11388 12112 11394 12164
rect 14108 12152 14136 12183
rect 14182 12180 14188 12232
rect 14240 12220 14246 12232
rect 14921 12223 14979 12229
rect 14240 12192 14284 12220
rect 14240 12180 14246 12192
rect 14921 12189 14933 12223
rect 14967 12189 14979 12223
rect 14921 12183 14979 12189
rect 14274 12152 14280 12164
rect 14108 12124 14280 12152
rect 14274 12112 14280 12124
rect 14332 12112 14338 12164
rect 14936 12152 14964 12183
rect 15010 12180 15016 12232
rect 15068 12220 15074 12232
rect 15068 12192 15113 12220
rect 15068 12180 15074 12192
rect 15194 12180 15200 12232
rect 15252 12220 15258 12232
rect 15930 12220 15936 12232
rect 15252 12192 15297 12220
rect 15891 12192 15936 12220
rect 15252 12180 15258 12192
rect 15930 12180 15936 12192
rect 15988 12180 15994 12232
rect 15102 12152 15108 12164
rect 14384 12124 15108 12152
rect 1946 12084 1952 12096
rect 1907 12056 1952 12084
rect 1946 12044 1952 12056
rect 2004 12044 2010 12096
rect 6181 12087 6239 12093
rect 6181 12053 6193 12087
rect 6227 12084 6239 12087
rect 6730 12084 6736 12096
rect 6227 12056 6736 12084
rect 6227 12053 6239 12056
rect 6181 12047 6239 12053
rect 6730 12044 6736 12056
rect 6788 12044 6794 12096
rect 7791 12087 7849 12093
rect 7791 12053 7803 12087
rect 7837 12084 7849 12087
rect 8846 12084 8852 12096
rect 7837 12056 8852 12084
rect 7837 12053 7849 12056
rect 7791 12047 7849 12053
rect 8846 12044 8852 12056
rect 8904 12044 8910 12096
rect 12621 12087 12679 12093
rect 12621 12053 12633 12087
rect 12667 12084 12679 12087
rect 12894 12084 12900 12096
rect 12667 12056 12900 12084
rect 12667 12053 12679 12056
rect 12621 12047 12679 12053
rect 12894 12044 12900 12056
rect 12952 12044 12958 12096
rect 13998 12044 14004 12096
rect 14056 12084 14062 12096
rect 14384 12084 14412 12124
rect 15102 12112 15108 12124
rect 15160 12112 15166 12164
rect 15948 12152 15976 12180
rect 16776 12152 16804 12251
rect 15948 12124 16804 12152
rect 14056 12056 14412 12084
rect 14056 12044 14062 12056
rect 14458 12044 14464 12096
rect 14516 12084 14522 12096
rect 14737 12087 14795 12093
rect 14737 12084 14749 12087
rect 14516 12056 14749 12084
rect 14516 12044 14522 12056
rect 14737 12053 14749 12056
rect 14783 12053 14795 12087
rect 14737 12047 14795 12053
rect 16390 12044 16396 12096
rect 16448 12084 16454 12096
rect 17512 12084 17540 12251
rect 17862 12248 17868 12260
rect 17920 12248 17926 12300
rect 18414 12288 18420 12300
rect 18375 12260 18420 12288
rect 18414 12248 18420 12260
rect 18472 12248 18478 12300
rect 18230 12152 18236 12164
rect 18191 12124 18236 12152
rect 18230 12112 18236 12124
rect 18288 12112 18294 12164
rect 16448 12056 17540 12084
rect 16448 12044 16454 12056
rect 184 11994 18860 12016
rect 184 11942 1556 11994
rect 1608 11942 1620 11994
rect 1672 11942 1684 11994
rect 1736 11942 1748 11994
rect 1800 11942 1812 11994
rect 1864 11942 4656 11994
rect 4708 11942 4720 11994
rect 4772 11942 4784 11994
rect 4836 11942 4848 11994
rect 4900 11942 4912 11994
rect 4964 11942 7756 11994
rect 7808 11942 7820 11994
rect 7872 11942 7884 11994
rect 7936 11942 7948 11994
rect 8000 11942 8012 11994
rect 8064 11942 10856 11994
rect 10908 11942 10920 11994
rect 10972 11942 10984 11994
rect 11036 11942 11048 11994
rect 11100 11942 11112 11994
rect 11164 11942 13956 11994
rect 14008 11942 14020 11994
rect 14072 11942 14084 11994
rect 14136 11942 14148 11994
rect 14200 11942 14212 11994
rect 14264 11942 17056 11994
rect 17108 11942 17120 11994
rect 17172 11942 17184 11994
rect 17236 11942 17248 11994
rect 17300 11942 17312 11994
rect 17364 11942 18860 11994
rect 184 11920 18860 11942
rect 1946 11880 1952 11892
rect 1596 11852 1952 11880
rect 1596 11753 1624 11852
rect 1946 11840 1952 11852
rect 2004 11840 2010 11892
rect 7558 11840 7564 11892
rect 7616 11880 7622 11892
rect 7745 11883 7803 11889
rect 7745 11880 7757 11883
rect 7616 11852 7757 11880
rect 7616 11840 7622 11852
rect 7745 11849 7757 11852
rect 7791 11849 7803 11883
rect 7745 11843 7803 11849
rect 14274 11840 14280 11892
rect 14332 11880 14338 11892
rect 15194 11880 15200 11892
rect 14332 11852 15200 11880
rect 14332 11840 14338 11852
rect 15194 11840 15200 11852
rect 15252 11840 15258 11892
rect 7466 11772 7472 11824
rect 7524 11812 7530 11824
rect 8021 11815 8079 11821
rect 8021 11812 8033 11815
rect 7524 11784 8033 11812
rect 7524 11772 7530 11784
rect 8021 11781 8033 11784
rect 8067 11781 8079 11815
rect 8021 11775 8079 11781
rect 1581 11747 1639 11753
rect 1581 11713 1593 11747
rect 1627 11713 1639 11747
rect 6457 11747 6515 11753
rect 6457 11744 6469 11747
rect 1581 11707 1639 11713
rect 6012 11716 6469 11744
rect 1949 11679 2007 11685
rect 1949 11645 1961 11679
rect 1995 11676 2007 11679
rect 2038 11676 2044 11688
rect 1995 11648 2044 11676
rect 1995 11645 2007 11648
rect 1949 11639 2007 11645
rect 2038 11636 2044 11648
rect 2096 11636 2102 11688
rect 6012 11685 6040 11716
rect 6457 11713 6469 11716
rect 6503 11744 6515 11747
rect 12894 11744 12900 11756
rect 6503 11716 12434 11744
rect 12855 11716 12900 11744
rect 6503 11713 6515 11716
rect 6457 11707 6515 11713
rect 5997 11679 6055 11685
rect 5997 11645 6009 11679
rect 6043 11645 6055 11679
rect 7098 11676 7104 11688
rect 7059 11648 7104 11676
rect 5997 11639 6055 11645
rect 7098 11636 7104 11648
rect 7156 11636 7162 11688
rect 7193 11679 7251 11685
rect 7193 11645 7205 11679
rect 7239 11645 7251 11679
rect 7374 11676 7380 11688
rect 7335 11648 7380 11676
rect 7193 11639 7251 11645
rect 2314 11568 2320 11620
rect 2372 11568 2378 11620
rect 7208 11608 7236 11639
rect 7374 11636 7380 11648
rect 7432 11636 7438 11688
rect 8018 11676 8024 11688
rect 7979 11648 8024 11676
rect 8018 11636 8024 11648
rect 8076 11636 8082 11688
rect 8202 11676 8208 11688
rect 8115 11648 8208 11676
rect 8202 11636 8208 11648
rect 8260 11636 8266 11688
rect 8294 11636 8300 11688
rect 8352 11676 8358 11688
rect 8757 11679 8815 11685
rect 8757 11676 8769 11679
rect 8352 11648 8769 11676
rect 8352 11636 8358 11648
rect 8757 11645 8769 11648
rect 8803 11645 8815 11679
rect 8757 11639 8815 11645
rect 7466 11608 7472 11620
rect 7208 11580 7472 11608
rect 7466 11568 7472 11580
rect 7524 11568 7530 11620
rect 7650 11568 7656 11620
rect 7708 11608 7714 11620
rect 7745 11611 7803 11617
rect 7745 11608 7757 11611
rect 7708 11580 7757 11608
rect 7708 11568 7714 11580
rect 7745 11577 7757 11580
rect 7791 11577 7803 11611
rect 7745 11571 7803 11577
rect 1670 11500 1676 11552
rect 1728 11540 1734 11552
rect 2222 11540 2228 11552
rect 1728 11512 2228 11540
rect 1728 11500 1734 11512
rect 2222 11500 2228 11512
rect 2280 11540 2286 11552
rect 3375 11543 3433 11549
rect 3375 11540 3387 11543
rect 2280 11512 3387 11540
rect 2280 11500 2286 11512
rect 3375 11509 3387 11512
rect 3421 11509 3433 11543
rect 4522 11540 4528 11552
rect 4483 11512 4528 11540
rect 3375 11503 3433 11509
rect 4522 11500 4528 11512
rect 4580 11500 4586 11552
rect 7006 11500 7012 11552
rect 7064 11540 7070 11552
rect 8220 11540 8248 11636
rect 7064 11512 8248 11540
rect 8772 11540 8800 11639
rect 8846 11636 8852 11688
rect 8904 11676 8910 11688
rect 9125 11679 9183 11685
rect 9125 11676 9137 11679
rect 8904 11648 9137 11676
rect 8904 11636 8910 11648
rect 9125 11645 9137 11648
rect 9171 11645 9183 11679
rect 9125 11639 9183 11645
rect 9490 11568 9496 11620
rect 9548 11568 9554 11620
rect 12406 11608 12434 11716
rect 12894 11704 12900 11716
rect 12952 11704 12958 11756
rect 16574 11744 16580 11756
rect 16316 11716 16580 11744
rect 12802 11676 12808 11688
rect 12763 11648 12808 11676
rect 12802 11636 12808 11648
rect 12860 11636 12866 11688
rect 14182 11636 14188 11688
rect 14240 11676 14246 11688
rect 15286 11676 15292 11688
rect 14240 11648 15292 11676
rect 14240 11636 14246 11648
rect 15286 11636 15292 11648
rect 15344 11636 15350 11688
rect 15562 11676 15568 11688
rect 15523 11648 15568 11676
rect 15562 11636 15568 11648
rect 15620 11636 15626 11688
rect 16316 11685 16344 11716
rect 16574 11704 16580 11716
rect 16632 11704 16638 11756
rect 16301 11679 16359 11685
rect 16301 11645 16313 11679
rect 16347 11645 16359 11679
rect 16301 11639 16359 11645
rect 15378 11608 15384 11620
rect 12406 11580 15384 11608
rect 15378 11568 15384 11580
rect 15436 11568 15442 11620
rect 16844 11611 16902 11617
rect 16844 11577 16856 11611
rect 16890 11608 16902 11611
rect 16942 11608 16948 11620
rect 16890 11580 16948 11608
rect 16890 11577 16902 11580
rect 16844 11571 16902 11577
rect 16942 11568 16948 11580
rect 17000 11568 17006 11620
rect 9214 11540 9220 11552
rect 8772 11512 9220 11540
rect 7064 11500 7070 11512
rect 9214 11500 9220 11512
rect 9272 11500 9278 11552
rect 9766 11500 9772 11552
rect 9824 11540 9830 11552
rect 10551 11543 10609 11549
rect 10551 11540 10563 11543
rect 9824 11512 10563 11540
rect 9824 11500 9830 11512
rect 10551 11509 10563 11512
rect 10597 11509 10609 11543
rect 10551 11503 10609 11509
rect 11790 11500 11796 11552
rect 11848 11540 11854 11552
rect 12345 11543 12403 11549
rect 12345 11540 12357 11543
rect 11848 11512 12357 11540
rect 11848 11500 11854 11512
rect 12345 11509 12357 11512
rect 12391 11509 12403 11543
rect 12345 11503 12403 11509
rect 12713 11543 12771 11549
rect 12713 11509 12725 11543
rect 12759 11540 12771 11543
rect 14182 11540 14188 11552
rect 12759 11512 14188 11540
rect 12759 11509 12771 11512
rect 12713 11503 12771 11509
rect 14182 11500 14188 11512
rect 14240 11500 14246 11552
rect 14277 11543 14335 11549
rect 14277 11509 14289 11543
rect 14323 11540 14335 11543
rect 14366 11540 14372 11552
rect 14323 11512 14372 11540
rect 14323 11509 14335 11512
rect 14277 11503 14335 11509
rect 14366 11500 14372 11512
rect 14424 11500 14430 11552
rect 14734 11500 14740 11552
rect 14792 11540 14798 11552
rect 16025 11543 16083 11549
rect 16025 11540 16037 11543
rect 14792 11512 16037 11540
rect 14792 11500 14798 11512
rect 16025 11509 16037 11512
rect 16071 11509 16083 11543
rect 16025 11503 16083 11509
rect 17770 11500 17776 11552
rect 17828 11540 17834 11552
rect 17957 11543 18015 11549
rect 17957 11540 17969 11543
rect 17828 11512 17969 11540
rect 17828 11500 17834 11512
rect 17957 11509 17969 11512
rect 18003 11509 18015 11543
rect 18414 11540 18420 11552
rect 18375 11512 18420 11540
rect 17957 11503 18015 11509
rect 18414 11500 18420 11512
rect 18472 11500 18478 11552
rect 184 11450 18920 11472
rect 184 11398 3106 11450
rect 3158 11398 3170 11450
rect 3222 11398 3234 11450
rect 3286 11398 3298 11450
rect 3350 11398 3362 11450
rect 3414 11398 6206 11450
rect 6258 11398 6270 11450
rect 6322 11398 6334 11450
rect 6386 11398 6398 11450
rect 6450 11398 6462 11450
rect 6514 11398 9306 11450
rect 9358 11398 9370 11450
rect 9422 11398 9434 11450
rect 9486 11398 9498 11450
rect 9550 11398 9562 11450
rect 9614 11398 12406 11450
rect 12458 11398 12470 11450
rect 12522 11398 12534 11450
rect 12586 11398 12598 11450
rect 12650 11398 12662 11450
rect 12714 11398 15506 11450
rect 15558 11398 15570 11450
rect 15622 11398 15634 11450
rect 15686 11398 15698 11450
rect 15750 11398 15762 11450
rect 15814 11398 18606 11450
rect 18658 11398 18670 11450
rect 18722 11398 18734 11450
rect 18786 11398 18798 11450
rect 18850 11398 18862 11450
rect 18914 11398 18920 11450
rect 184 11376 18920 11398
rect 1670 11336 1676 11348
rect 1631 11308 1676 11336
rect 1670 11296 1676 11308
rect 1728 11296 1734 11348
rect 2038 11336 2044 11348
rect 1999 11308 2044 11336
rect 2038 11296 2044 11308
rect 2096 11296 2102 11348
rect 5534 11336 5540 11348
rect 5495 11308 5540 11336
rect 5534 11296 5540 11308
rect 5592 11296 5598 11348
rect 8294 11336 8300 11348
rect 8255 11308 8300 11336
rect 8294 11296 8300 11308
rect 8352 11296 8358 11348
rect 8018 11268 8024 11280
rect 5184 11240 8024 11268
rect 3786 11200 3792 11212
rect 3747 11172 3792 11200
rect 3786 11160 3792 11172
rect 3844 11160 3850 11212
rect 3973 11203 4031 11209
rect 3973 11169 3985 11203
rect 4019 11200 4031 11203
rect 4062 11200 4068 11212
rect 4019 11172 4068 11200
rect 4019 11169 4031 11172
rect 3973 11163 4031 11169
rect 4062 11160 4068 11172
rect 4120 11160 4126 11212
rect 5184 11209 5212 11240
rect 8018 11228 8024 11240
rect 8076 11228 8082 11280
rect 9030 11228 9036 11280
rect 9088 11268 9094 11280
rect 9585 11271 9643 11277
rect 9585 11268 9597 11271
rect 9088 11240 9597 11268
rect 9088 11228 9094 11240
rect 9585 11237 9597 11240
rect 9631 11237 9643 11271
rect 11606 11268 11612 11280
rect 11454 11240 11612 11268
rect 9585 11231 9643 11237
rect 11606 11228 11612 11240
rect 11664 11228 11670 11280
rect 14642 11268 14648 11280
rect 14016 11240 14648 11268
rect 5169 11203 5227 11209
rect 5169 11169 5181 11203
rect 5215 11169 5227 11203
rect 5169 11163 5227 11169
rect 1489 11135 1547 11141
rect 1489 11101 1501 11135
rect 1535 11101 1547 11135
rect 1489 11095 1547 11101
rect 1581 11135 1639 11141
rect 1581 11101 1593 11135
rect 1627 11132 1639 11135
rect 2682 11132 2688 11144
rect 1627 11104 2688 11132
rect 1627 11101 1639 11104
rect 1581 11095 1639 11101
rect 1504 11064 1532 11095
rect 2682 11092 2688 11104
rect 2740 11092 2746 11144
rect 3602 11092 3608 11144
rect 3660 11132 3666 11144
rect 5184 11132 5212 11163
rect 5258 11160 5264 11212
rect 5316 11200 5322 11212
rect 8036 11200 8064 11228
rect 9766 11200 9772 11212
rect 5316 11172 5361 11200
rect 8036 11172 9772 11200
rect 5316 11160 5322 11172
rect 9766 11160 9772 11172
rect 9824 11160 9830 11212
rect 9950 11200 9956 11212
rect 9911 11172 9956 11200
rect 9950 11160 9956 11172
rect 10008 11160 10014 11212
rect 14016 11209 14044 11240
rect 14642 11228 14648 11240
rect 14700 11228 14706 11280
rect 16114 11228 16120 11280
rect 16172 11228 16178 11280
rect 14001 11203 14059 11209
rect 14001 11169 14013 11203
rect 14047 11169 14059 11203
rect 14001 11163 14059 11169
rect 14185 11203 14243 11209
rect 14185 11169 14197 11203
rect 14231 11200 14243 11203
rect 14458 11200 14464 11212
rect 14231 11172 14464 11200
rect 14231 11169 14243 11172
rect 14185 11163 14243 11169
rect 14458 11160 14464 11172
rect 14516 11160 14522 11212
rect 14734 11200 14740 11212
rect 14695 11172 14740 11200
rect 14734 11160 14740 11172
rect 14792 11160 14798 11212
rect 16942 11160 16948 11212
rect 17000 11200 17006 11212
rect 17129 11203 17187 11209
rect 17129 11200 17141 11203
rect 17000 11172 17141 11200
rect 17000 11160 17006 11172
rect 17129 11169 17141 11172
rect 17175 11169 17187 11203
rect 17129 11163 17187 11169
rect 17283 11203 17341 11209
rect 17283 11169 17295 11203
rect 17329 11200 17341 11203
rect 17770 11200 17776 11212
rect 17329 11172 17776 11200
rect 17329 11169 17341 11172
rect 17283 11163 17341 11169
rect 10226 11132 10232 11144
rect 3660 11104 5212 11132
rect 10187 11104 10232 11132
rect 3660 11092 3666 11104
rect 10226 11092 10232 11104
rect 10284 11092 10290 11144
rect 14093 11135 14151 11141
rect 14093 11101 14105 11135
rect 14139 11132 14151 11135
rect 15105 11135 15163 11141
rect 15105 11132 15117 11135
rect 14139 11104 15117 11132
rect 14139 11101 14151 11104
rect 14093 11095 14151 11101
rect 15105 11101 15117 11104
rect 15151 11101 15163 11135
rect 17144 11132 17172 11163
rect 17770 11160 17776 11172
rect 17828 11160 17834 11212
rect 17866 11203 17924 11209
rect 17866 11169 17878 11203
rect 17912 11169 17924 11203
rect 17866 11163 17924 11169
rect 17880 11132 17908 11163
rect 17144 11104 17908 11132
rect 15105 11095 15163 11101
rect 2130 11064 2136 11076
rect 1504 11036 2136 11064
rect 2130 11024 2136 11036
rect 2188 11024 2194 11076
rect 17494 11024 17500 11076
rect 17552 11064 17558 11076
rect 18141 11067 18199 11073
rect 18141 11064 18153 11067
rect 17552 11036 18153 11064
rect 17552 11024 17558 11036
rect 18141 11033 18153 11036
rect 18187 11033 18199 11067
rect 18141 11027 18199 11033
rect 3142 10956 3148 11008
rect 3200 10996 3206 11008
rect 3973 10999 4031 11005
rect 3973 10996 3985 10999
rect 3200 10968 3985 10996
rect 3200 10956 3206 10968
rect 3973 10965 3985 10968
rect 4019 10965 4031 10999
rect 3973 10959 4031 10965
rect 11514 10956 11520 11008
rect 11572 10996 11578 11008
rect 11701 10999 11759 11005
rect 11701 10996 11713 10999
rect 11572 10968 11713 10996
rect 11572 10956 11578 10968
rect 11701 10965 11713 10968
rect 11747 10965 11759 10999
rect 11701 10959 11759 10965
rect 15562 10956 15568 11008
rect 15620 10996 15626 11008
rect 15930 10996 15936 11008
rect 15620 10968 15936 10996
rect 15620 10956 15626 10968
rect 15930 10956 15936 10968
rect 15988 10996 15994 11008
rect 16531 10999 16589 11005
rect 16531 10996 16543 10999
rect 15988 10968 16543 10996
rect 15988 10956 15994 10968
rect 16531 10965 16543 10968
rect 16577 10965 16589 10999
rect 16531 10959 16589 10965
rect 17313 10999 17371 11005
rect 17313 10965 17325 10999
rect 17359 10996 17371 10999
rect 17402 10996 17408 11008
rect 17359 10968 17408 10996
rect 17359 10965 17371 10968
rect 17313 10959 17371 10965
rect 17402 10956 17408 10968
rect 17460 10956 17466 11008
rect 184 10906 18860 10928
rect 184 10854 1556 10906
rect 1608 10854 1620 10906
rect 1672 10854 1684 10906
rect 1736 10854 1748 10906
rect 1800 10854 1812 10906
rect 1864 10854 4656 10906
rect 4708 10854 4720 10906
rect 4772 10854 4784 10906
rect 4836 10854 4848 10906
rect 4900 10854 4912 10906
rect 4964 10854 7756 10906
rect 7808 10854 7820 10906
rect 7872 10854 7884 10906
rect 7936 10854 7948 10906
rect 8000 10854 8012 10906
rect 8064 10854 10856 10906
rect 10908 10854 10920 10906
rect 10972 10854 10984 10906
rect 11036 10854 11048 10906
rect 11100 10854 11112 10906
rect 11164 10854 13956 10906
rect 14008 10854 14020 10906
rect 14072 10854 14084 10906
rect 14136 10854 14148 10906
rect 14200 10854 14212 10906
rect 14264 10854 17056 10906
rect 17108 10854 17120 10906
rect 17172 10854 17184 10906
rect 17236 10854 17248 10906
rect 17300 10854 17312 10906
rect 17364 10854 18860 10906
rect 184 10832 18860 10854
rect 2682 10792 2688 10804
rect 2643 10764 2688 10792
rect 2682 10752 2688 10764
rect 2740 10752 2746 10804
rect 6457 10795 6515 10801
rect 6457 10761 6469 10795
rect 6503 10792 6515 10795
rect 6638 10792 6644 10804
rect 6503 10764 6644 10792
rect 6503 10761 6515 10764
rect 6457 10755 6515 10761
rect 6638 10752 6644 10764
rect 6696 10752 6702 10804
rect 7650 10752 7656 10804
rect 7708 10792 7714 10804
rect 7745 10795 7803 10801
rect 7745 10792 7757 10795
rect 7708 10764 7757 10792
rect 7708 10752 7714 10764
rect 7745 10761 7757 10764
rect 7791 10761 7803 10795
rect 7745 10755 7803 10761
rect 10226 10752 10232 10804
rect 10284 10792 10290 10804
rect 11149 10795 11207 10801
rect 11149 10792 11161 10795
rect 10284 10764 11161 10792
rect 10284 10752 10290 10764
rect 11149 10761 11161 10764
rect 11195 10761 11207 10795
rect 11149 10755 11207 10761
rect 15194 10752 15200 10804
rect 15252 10792 15258 10804
rect 15473 10795 15531 10801
rect 15473 10792 15485 10795
rect 15252 10764 15485 10792
rect 15252 10752 15258 10764
rect 15473 10761 15485 10764
rect 15519 10761 15531 10795
rect 16942 10792 16948 10804
rect 16903 10764 16948 10792
rect 15473 10755 15531 10761
rect 16942 10752 16948 10764
rect 17000 10792 17006 10804
rect 17589 10795 17647 10801
rect 17589 10792 17601 10795
rect 17000 10764 17601 10792
rect 17000 10752 17006 10764
rect 17589 10761 17601 10764
rect 17635 10761 17647 10795
rect 17589 10755 17647 10761
rect 3694 10684 3700 10736
rect 3752 10724 3758 10736
rect 3752 10696 4568 10724
rect 3752 10684 3758 10696
rect 2133 10659 2191 10665
rect 2133 10625 2145 10659
rect 2179 10656 2191 10659
rect 2590 10656 2596 10668
rect 2179 10628 2596 10656
rect 2179 10625 2191 10628
rect 2133 10619 2191 10625
rect 2590 10616 2596 10628
rect 2648 10616 2654 10668
rect 3142 10656 3148 10668
rect 3103 10628 3148 10656
rect 3142 10616 3148 10628
rect 3200 10616 3206 10668
rect 3329 10659 3387 10665
rect 3329 10625 3341 10659
rect 3375 10625 3387 10659
rect 3329 10619 3387 10625
rect 2041 10591 2099 10597
rect 2041 10557 2053 10591
rect 2087 10588 2099 10591
rect 2222 10588 2228 10600
rect 2087 10560 2228 10588
rect 2087 10557 2099 10560
rect 2041 10551 2099 10557
rect 2222 10548 2228 10560
rect 2280 10588 2286 10600
rect 2682 10588 2688 10600
rect 2280 10560 2688 10588
rect 2280 10548 2286 10560
rect 2682 10548 2688 10560
rect 2740 10548 2746 10600
rect 3053 10523 3111 10529
rect 3053 10520 3065 10523
rect 2424 10492 3065 10520
rect 2424 10461 2452 10492
rect 3053 10489 3065 10492
rect 3099 10489 3111 10523
rect 3344 10520 3372 10619
rect 3878 10616 3884 10668
rect 3936 10656 3942 10668
rect 4540 10665 4568 10696
rect 4982 10684 4988 10736
rect 5040 10724 5046 10736
rect 5040 10696 7696 10724
rect 5040 10684 5046 10696
rect 4433 10659 4491 10665
rect 4433 10656 4445 10659
rect 3936 10628 4445 10656
rect 3936 10616 3942 10628
rect 4433 10625 4445 10628
rect 4479 10625 4491 10659
rect 4433 10619 4491 10625
rect 4525 10659 4583 10665
rect 4525 10625 4537 10659
rect 4571 10656 4583 10659
rect 6914 10656 6920 10668
rect 4571 10628 6920 10656
rect 4571 10625 4583 10628
rect 4525 10619 4583 10625
rect 6914 10616 6920 10628
rect 6972 10616 6978 10668
rect 4246 10588 4252 10600
rect 4207 10560 4252 10588
rect 4246 10548 4252 10560
rect 4304 10548 4310 10600
rect 6365 10591 6423 10597
rect 6365 10557 6377 10591
rect 6411 10557 6423 10591
rect 6365 10551 6423 10557
rect 4338 10520 4344 10532
rect 3344 10492 4344 10520
rect 3053 10483 3111 10489
rect 4338 10480 4344 10492
rect 4396 10520 4402 10532
rect 6380 10520 6408 10551
rect 6546 10548 6552 10600
rect 6604 10588 6610 10600
rect 6641 10591 6699 10597
rect 6641 10588 6653 10591
rect 6604 10560 6653 10588
rect 6604 10548 6610 10560
rect 6641 10557 6653 10560
rect 6687 10557 6699 10591
rect 6641 10551 6699 10557
rect 6730 10548 6736 10600
rect 6788 10588 6794 10600
rect 7668 10597 7696 10696
rect 11790 10656 11796 10668
rect 11751 10628 11796 10656
rect 11790 10616 11796 10628
rect 11848 10616 11854 10668
rect 12802 10656 12808 10668
rect 12763 10628 12808 10656
rect 12802 10616 12808 10628
rect 12860 10616 12866 10668
rect 7653 10591 7711 10597
rect 6788 10560 6833 10588
rect 6788 10548 6794 10560
rect 7653 10557 7665 10591
rect 7699 10557 7711 10591
rect 8110 10588 8116 10600
rect 8071 10560 8116 10588
rect 7653 10551 7711 10557
rect 8110 10548 8116 10560
rect 8168 10548 8174 10600
rect 11514 10588 11520 10600
rect 11475 10560 11520 10588
rect 11514 10548 11520 10560
rect 11572 10548 11578 10600
rect 15562 10588 15568 10600
rect 15523 10560 15568 10588
rect 15562 10548 15568 10560
rect 15620 10548 15626 10600
rect 8570 10520 8576 10532
rect 4396 10492 8576 10520
rect 4396 10480 4402 10492
rect 8570 10480 8576 10492
rect 8628 10480 8634 10532
rect 12529 10523 12587 10529
rect 12529 10489 12541 10523
rect 12575 10520 12587 10523
rect 12802 10520 12808 10532
rect 12575 10492 12808 10520
rect 12575 10489 12587 10492
rect 12529 10483 12587 10489
rect 12802 10480 12808 10492
rect 12860 10480 12866 10532
rect 2409 10455 2467 10461
rect 2409 10421 2421 10455
rect 2455 10421 2467 10455
rect 4062 10452 4068 10464
rect 4023 10424 4068 10452
rect 2409 10415 2467 10421
rect 4062 10412 4068 10424
rect 4120 10412 4126 10464
rect 6917 10455 6975 10461
rect 6917 10421 6929 10455
rect 6963 10452 6975 10455
rect 8110 10452 8116 10464
rect 6963 10424 8116 10452
rect 6963 10421 6975 10424
rect 6917 10415 6975 10421
rect 8110 10412 8116 10424
rect 8168 10412 8174 10464
rect 11609 10455 11667 10461
rect 11609 10421 11621 10455
rect 11655 10452 11667 10455
rect 12161 10455 12219 10461
rect 12161 10452 12173 10455
rect 11655 10424 12173 10452
rect 11655 10421 11667 10424
rect 11609 10415 11667 10421
rect 12161 10421 12173 10424
rect 12207 10421 12219 10455
rect 12161 10415 12219 10421
rect 12621 10455 12679 10461
rect 12621 10421 12633 10455
rect 12667 10452 12679 10455
rect 13170 10452 13176 10464
rect 12667 10424 13176 10452
rect 12667 10421 12679 10424
rect 12621 10415 12679 10421
rect 13170 10412 13176 10424
rect 13228 10412 13234 10464
rect 184 10362 18920 10384
rect 184 10310 3106 10362
rect 3158 10310 3170 10362
rect 3222 10310 3234 10362
rect 3286 10310 3298 10362
rect 3350 10310 3362 10362
rect 3414 10310 6206 10362
rect 6258 10310 6270 10362
rect 6322 10310 6334 10362
rect 6386 10310 6398 10362
rect 6450 10310 6462 10362
rect 6514 10310 9306 10362
rect 9358 10310 9370 10362
rect 9422 10310 9434 10362
rect 9486 10310 9498 10362
rect 9550 10310 9562 10362
rect 9614 10310 12406 10362
rect 12458 10310 12470 10362
rect 12522 10310 12534 10362
rect 12586 10310 12598 10362
rect 12650 10310 12662 10362
rect 12714 10310 15506 10362
rect 15558 10310 15570 10362
rect 15622 10310 15634 10362
rect 15686 10310 15698 10362
rect 15750 10310 15762 10362
rect 15814 10310 18606 10362
rect 18658 10310 18670 10362
rect 18722 10310 18734 10362
rect 18786 10310 18798 10362
rect 18850 10310 18862 10362
rect 18914 10310 18920 10362
rect 184 10288 18920 10310
rect 753 10251 811 10257
rect 753 10217 765 10251
rect 799 10248 811 10251
rect 1394 10248 1400 10260
rect 799 10220 1400 10248
rect 799 10217 811 10220
rect 753 10211 811 10217
rect 1394 10208 1400 10220
rect 1452 10208 1458 10260
rect 3786 10248 3792 10260
rect 3747 10220 3792 10248
rect 3786 10208 3792 10220
rect 3844 10208 3850 10260
rect 6546 10248 6552 10260
rect 6507 10220 6552 10248
rect 6546 10208 6552 10220
rect 6604 10208 6610 10260
rect 7193 10251 7251 10257
rect 7193 10217 7205 10251
rect 7239 10248 7251 10251
rect 7374 10248 7380 10260
rect 7239 10220 7380 10248
rect 7239 10217 7251 10220
rect 7193 10211 7251 10217
rect 7374 10208 7380 10220
rect 7432 10208 7438 10260
rect 11882 10248 11888 10260
rect 11843 10220 11888 10248
rect 11882 10208 11888 10220
rect 11940 10248 11946 10260
rect 12342 10248 12348 10260
rect 11940 10220 12348 10248
rect 11940 10208 11946 10220
rect 12342 10208 12348 10220
rect 12400 10208 12406 10260
rect 12802 10248 12808 10260
rect 12763 10220 12808 10248
rect 12802 10208 12808 10220
rect 12860 10208 12866 10260
rect 5261 10183 5319 10189
rect 5261 10149 5273 10183
rect 5307 10180 5319 10183
rect 8110 10180 8116 10192
rect 5307 10152 6316 10180
rect 8071 10152 8116 10180
rect 5307 10149 5319 10152
rect 5261 10143 5319 10149
rect 569 10115 627 10121
rect 569 10081 581 10115
rect 615 10112 627 10115
rect 934 10112 940 10124
rect 615 10084 940 10112
rect 615 10081 627 10084
rect 569 10075 627 10081
rect 934 10072 940 10084
rect 992 10112 998 10124
rect 1029 10115 1087 10121
rect 1029 10112 1041 10115
rect 992 10084 1041 10112
rect 992 10072 998 10084
rect 1029 10081 1041 10084
rect 1075 10081 1087 10115
rect 3786 10112 3792 10124
rect 3747 10084 3792 10112
rect 1029 10075 1087 10081
rect 3786 10072 3792 10084
rect 3844 10072 3850 10124
rect 5169 10115 5227 10121
rect 5169 10081 5181 10115
rect 5215 10081 5227 10115
rect 5350 10112 5356 10124
rect 5311 10084 5356 10112
rect 5169 10075 5227 10081
rect 3694 10004 3700 10056
rect 3752 10044 3758 10056
rect 3881 10047 3939 10053
rect 3881 10044 3893 10047
rect 3752 10016 3893 10044
rect 3752 10004 3758 10016
rect 3881 10013 3893 10016
rect 3927 10013 3939 10047
rect 3881 10007 3939 10013
rect 4065 10047 4123 10053
rect 4065 10013 4077 10047
rect 4111 10044 4123 10047
rect 4246 10044 4252 10056
rect 4111 10016 4252 10044
rect 4111 10013 4123 10016
rect 4065 10007 4123 10013
rect 4246 10004 4252 10016
rect 4304 10044 4310 10056
rect 5184 10044 5212 10075
rect 5350 10072 5356 10084
rect 5408 10112 5414 10124
rect 6288 10121 6316 10152
rect 8110 10140 8116 10152
rect 8168 10140 8174 10192
rect 8662 10140 8668 10192
rect 8720 10140 8726 10192
rect 11333 10183 11391 10189
rect 11333 10149 11345 10183
rect 11379 10180 11391 10183
rect 17494 10180 17500 10192
rect 11379 10152 12664 10180
rect 17455 10152 17500 10180
rect 11379 10149 11391 10152
rect 11333 10143 11391 10149
rect 5813 10115 5871 10121
rect 5813 10112 5825 10115
rect 5408 10084 5825 10112
rect 5408 10072 5414 10084
rect 5813 10081 5825 10084
rect 5859 10081 5871 10115
rect 5813 10075 5871 10081
rect 6273 10115 6331 10121
rect 6273 10081 6285 10115
rect 6319 10081 6331 10115
rect 6273 10075 6331 10081
rect 7009 10115 7067 10121
rect 7009 10081 7021 10115
rect 7055 10112 7067 10115
rect 7190 10112 7196 10124
rect 7055 10084 7196 10112
rect 7055 10081 7067 10084
rect 7009 10075 7067 10081
rect 7190 10072 7196 10084
rect 7248 10072 7254 10124
rect 11149 10115 11207 10121
rect 11149 10081 11161 10115
rect 11195 10112 11207 10115
rect 11514 10112 11520 10124
rect 11195 10084 11520 10112
rect 11195 10081 11207 10084
rect 11149 10075 11207 10081
rect 11514 10072 11520 10084
rect 11572 10112 11578 10124
rect 11701 10115 11759 10121
rect 11701 10112 11713 10115
rect 11572 10084 11713 10112
rect 11572 10072 11578 10084
rect 11701 10081 11713 10084
rect 11747 10081 11759 10115
rect 11701 10075 11759 10081
rect 11885 10115 11943 10121
rect 11885 10081 11897 10115
rect 11931 10081 11943 10115
rect 12342 10112 12348 10124
rect 12303 10084 12348 10112
rect 11885 10075 11943 10081
rect 5629 10047 5687 10053
rect 5629 10044 5641 10047
rect 4304 10016 5641 10044
rect 4304 10004 4310 10016
rect 5629 10013 5641 10016
rect 5675 10013 5687 10047
rect 6546 10044 6552 10056
rect 6507 10016 6552 10044
rect 5629 10007 5687 10013
rect 5644 9976 5672 10007
rect 6546 10004 6552 10016
rect 6604 10004 6610 10056
rect 6822 10044 6828 10056
rect 6783 10016 6828 10044
rect 6822 10004 6828 10016
rect 6880 10004 6886 10056
rect 7558 10004 7564 10056
rect 7616 10044 7622 10056
rect 7837 10047 7895 10053
rect 7837 10044 7849 10047
rect 7616 10016 7849 10044
rect 7616 10004 7622 10016
rect 7837 10013 7849 10016
rect 7883 10013 7895 10047
rect 7837 10007 7895 10013
rect 10873 10047 10931 10053
rect 10873 10013 10885 10047
rect 10919 10044 10931 10047
rect 11900 10044 11928 10075
rect 12342 10072 12348 10084
rect 12400 10072 12406 10124
rect 12636 10121 12664 10152
rect 17494 10140 17500 10152
rect 17552 10140 17558 10192
rect 12437 10115 12495 10121
rect 12437 10081 12449 10115
rect 12483 10081 12495 10115
rect 12437 10075 12495 10081
rect 12621 10115 12679 10121
rect 12621 10081 12633 10115
rect 12667 10081 12679 10115
rect 13262 10112 13268 10124
rect 13223 10084 13268 10112
rect 12621 10075 12679 10081
rect 11974 10044 11980 10056
rect 10919 10016 11980 10044
rect 10919 10013 10931 10016
rect 10873 10007 10931 10013
rect 11974 10004 11980 10016
rect 12032 10004 12038 10056
rect 12452 10044 12480 10075
rect 13262 10072 13268 10084
rect 13320 10072 13326 10124
rect 13541 10115 13599 10121
rect 13541 10081 13553 10115
rect 13587 10112 13599 10115
rect 13630 10112 13636 10124
rect 13587 10084 13636 10112
rect 13587 10081 13599 10084
rect 13541 10075 13599 10081
rect 13630 10072 13636 10084
rect 13688 10072 13694 10124
rect 17402 10112 17408 10124
rect 17363 10084 17408 10112
rect 17402 10072 17408 10084
rect 17460 10072 17466 10124
rect 17681 10115 17739 10121
rect 17681 10081 17693 10115
rect 17727 10112 17739 10115
rect 17954 10112 17960 10124
rect 17727 10084 17960 10112
rect 17727 10081 17739 10084
rect 17681 10075 17739 10081
rect 17954 10072 17960 10084
rect 18012 10072 18018 10124
rect 12894 10044 12900 10056
rect 12452 10016 12900 10044
rect 12894 10004 12900 10016
rect 12952 10004 12958 10056
rect 13449 10047 13507 10053
rect 13449 10013 13461 10047
rect 13495 10044 13507 10047
rect 13722 10044 13728 10056
rect 13495 10016 13728 10044
rect 13495 10013 13507 10016
rect 13449 10007 13507 10013
rect 13722 10004 13728 10016
rect 13780 10044 13786 10056
rect 14550 10044 14556 10056
rect 13780 10016 14556 10044
rect 13780 10004 13786 10016
rect 14550 10004 14556 10016
rect 14608 10004 14614 10056
rect 7374 9976 7380 9988
rect 5644 9948 7380 9976
rect 7374 9936 7380 9948
rect 7432 9936 7438 9988
rect 5997 9911 6055 9917
rect 5997 9877 6009 9911
rect 6043 9908 6055 9911
rect 6365 9911 6423 9917
rect 6365 9908 6377 9911
rect 6043 9880 6377 9908
rect 6043 9877 6055 9880
rect 5997 9871 6055 9877
rect 6365 9877 6377 9880
rect 6411 9877 6423 9911
rect 6365 9871 6423 9877
rect 9122 9868 9128 9920
rect 9180 9908 9186 9920
rect 9585 9911 9643 9917
rect 9585 9908 9597 9911
rect 9180 9880 9597 9908
rect 9180 9868 9186 9880
rect 9585 9877 9597 9880
rect 9631 9877 9643 9911
rect 9585 9871 9643 9877
rect 10778 9868 10784 9920
rect 10836 9908 10842 9920
rect 10965 9911 11023 9917
rect 10965 9908 10977 9911
rect 10836 9880 10977 9908
rect 10836 9868 10842 9880
rect 10965 9877 10977 9880
rect 11011 9877 11023 9911
rect 10965 9871 11023 9877
rect 13081 9911 13139 9917
rect 13081 9877 13093 9911
rect 13127 9908 13139 9911
rect 13170 9908 13176 9920
rect 13127 9880 13176 9908
rect 13127 9877 13139 9880
rect 13081 9871 13139 9877
rect 13170 9868 13176 9880
rect 13228 9868 13234 9920
rect 16666 9868 16672 9920
rect 16724 9908 16730 9920
rect 17405 9911 17463 9917
rect 17405 9908 17417 9911
rect 16724 9880 17417 9908
rect 16724 9868 16730 9880
rect 17405 9877 17417 9880
rect 17451 9877 17463 9911
rect 17405 9871 17463 9877
rect 184 9818 18860 9840
rect 184 9766 1556 9818
rect 1608 9766 1620 9818
rect 1672 9766 1684 9818
rect 1736 9766 1748 9818
rect 1800 9766 1812 9818
rect 1864 9766 4656 9818
rect 4708 9766 4720 9818
rect 4772 9766 4784 9818
rect 4836 9766 4848 9818
rect 4900 9766 4912 9818
rect 4964 9766 7756 9818
rect 7808 9766 7820 9818
rect 7872 9766 7884 9818
rect 7936 9766 7948 9818
rect 8000 9766 8012 9818
rect 8064 9766 10856 9818
rect 10908 9766 10920 9818
rect 10972 9766 10984 9818
rect 11036 9766 11048 9818
rect 11100 9766 11112 9818
rect 11164 9766 13956 9818
rect 14008 9766 14020 9818
rect 14072 9766 14084 9818
rect 14136 9766 14148 9818
rect 14200 9766 14212 9818
rect 14264 9766 17056 9818
rect 17108 9766 17120 9818
rect 17172 9766 17184 9818
rect 17236 9766 17248 9818
rect 17300 9766 17312 9818
rect 17364 9766 18860 9818
rect 184 9744 18860 9766
rect 10778 9664 10784 9716
rect 10836 9704 10842 9716
rect 12989 9707 13047 9713
rect 10836 9676 11008 9704
rect 10836 9664 10842 9676
rect 4338 9596 4344 9648
rect 4396 9636 4402 9648
rect 4396 9608 4568 9636
rect 4396 9596 4402 9608
rect 2130 9568 2136 9580
rect 2091 9540 2136 9568
rect 2130 9528 2136 9540
rect 2188 9528 2194 9580
rect 2240 9540 3096 9568
rect 1949 9503 2007 9509
rect 1949 9469 1961 9503
rect 1995 9500 2007 9503
rect 2240 9500 2268 9540
rect 2314 9500 2320 9512
rect 1995 9472 2320 9500
rect 1995 9469 2007 9472
rect 1949 9463 2007 9469
rect 2314 9460 2320 9472
rect 2372 9460 2378 9512
rect 2682 9460 2688 9512
rect 2740 9500 2746 9512
rect 3068 9509 3096 9540
rect 4062 9528 4068 9580
rect 4120 9568 4126 9580
rect 4540 9577 4568 9608
rect 8202 9596 8208 9648
rect 8260 9636 8266 9648
rect 8757 9639 8815 9645
rect 8757 9636 8769 9639
rect 8260 9608 8769 9636
rect 8260 9596 8266 9608
rect 8757 9605 8769 9608
rect 8803 9605 8815 9639
rect 10980 9636 11008 9676
rect 12989 9673 13001 9707
rect 13035 9704 13047 9707
rect 13262 9704 13268 9716
rect 13035 9676 13268 9704
rect 13035 9673 13047 9676
rect 12989 9667 13047 9673
rect 13262 9664 13268 9676
rect 13320 9664 13326 9716
rect 15933 9639 15991 9645
rect 15933 9636 15945 9639
rect 10980 9608 11928 9636
rect 8757 9599 8815 9605
rect 4433 9571 4491 9577
rect 4433 9568 4445 9571
rect 4120 9540 4445 9568
rect 4120 9528 4126 9540
rect 4433 9537 4445 9540
rect 4479 9537 4491 9571
rect 4433 9531 4491 9537
rect 4525 9571 4583 9577
rect 4525 9537 4537 9571
rect 4571 9537 4583 9571
rect 7098 9568 7104 9580
rect 7059 9540 7104 9568
rect 4525 9531 4583 9537
rect 7098 9528 7104 9540
rect 7156 9528 7162 9580
rect 11900 9577 11928 9608
rect 15028 9608 15945 9636
rect 15028 9577 15056 9608
rect 15933 9605 15945 9608
rect 15979 9605 15991 9639
rect 17954 9636 17960 9648
rect 17915 9608 17960 9636
rect 15933 9599 15991 9605
rect 17954 9596 17960 9608
rect 18012 9596 18018 9648
rect 11885 9571 11943 9577
rect 11885 9537 11897 9571
rect 11931 9537 11943 9571
rect 11885 9531 11943 9537
rect 15013 9571 15071 9577
rect 15013 9537 15025 9571
rect 15059 9537 15071 9571
rect 15013 9531 15071 9537
rect 2869 9503 2927 9509
rect 2869 9500 2881 9503
rect 2740 9472 2881 9500
rect 2740 9460 2746 9472
rect 2869 9469 2881 9472
rect 2915 9469 2927 9503
rect 2869 9463 2927 9469
rect 3053 9503 3111 9509
rect 3053 9469 3065 9503
rect 3099 9469 3111 9503
rect 3053 9463 3111 9469
rect 6822 9460 6828 9512
rect 6880 9500 6886 9512
rect 7009 9503 7067 9509
rect 7009 9500 7021 9503
rect 6880 9472 7021 9500
rect 6880 9460 6886 9472
rect 7009 9469 7021 9472
rect 7055 9469 7067 9503
rect 7190 9500 7196 9512
rect 7151 9472 7196 9500
rect 7009 9463 7067 9469
rect 7190 9460 7196 9472
rect 7248 9500 7254 9512
rect 9033 9503 9091 9509
rect 9033 9500 9045 9503
rect 7248 9472 9045 9500
rect 7248 9460 7254 9472
rect 9033 9469 9045 9472
rect 9079 9500 9091 9503
rect 9214 9500 9220 9512
rect 9079 9472 9220 9500
rect 9079 9469 9091 9472
rect 9033 9463 9091 9469
rect 9214 9460 9220 9472
rect 9272 9460 9278 9512
rect 10134 9500 10140 9512
rect 10095 9472 10140 9500
rect 10134 9460 10140 9472
rect 10192 9460 10198 9512
rect 11974 9500 11980 9512
rect 11935 9472 11980 9500
rect 11974 9460 11980 9472
rect 12032 9460 12038 9512
rect 15194 9500 15200 9512
rect 15155 9472 15200 9500
rect 15194 9460 15200 9472
rect 15252 9460 15258 9512
rect 15289 9503 15347 9509
rect 15289 9469 15301 9503
rect 15335 9500 15347 9503
rect 16206 9500 16212 9512
rect 15335 9472 16212 9500
rect 15335 9469 15347 9472
rect 15289 9463 15347 9469
rect 16206 9460 16212 9472
rect 16264 9460 16270 9512
rect 16298 9460 16304 9512
rect 16356 9500 16362 9512
rect 16850 9509 16856 9512
rect 16577 9503 16635 9509
rect 16577 9500 16589 9503
rect 16356 9472 16589 9500
rect 16356 9460 16362 9472
rect 16577 9469 16589 9472
rect 16623 9469 16635 9503
rect 16844 9500 16856 9509
rect 16811 9472 16856 9500
rect 16577 9463 16635 9469
rect 16844 9463 16856 9472
rect 16850 9460 16856 9463
rect 16908 9460 16914 9512
rect 2041 9435 2099 9441
rect 2041 9401 2053 9435
rect 2087 9432 2099 9435
rect 2087 9404 4016 9432
rect 2087 9401 2099 9404
rect 2041 9395 2099 9401
rect 842 9324 848 9376
rect 900 9364 906 9376
rect 1581 9367 1639 9373
rect 1581 9364 1593 9367
rect 900 9336 1593 9364
rect 900 9324 906 9336
rect 1581 9333 1593 9336
rect 1627 9333 1639 9367
rect 2958 9364 2964 9376
rect 2919 9336 2964 9364
rect 1581 9327 1639 9333
rect 2958 9324 2964 9336
rect 3016 9324 3022 9376
rect 3988 9373 4016 9404
rect 8570 9392 8576 9444
rect 8628 9432 8634 9444
rect 8757 9435 8815 9441
rect 8757 9432 8769 9435
rect 8628 9404 8769 9432
rect 8628 9392 8634 9404
rect 8757 9401 8769 9404
rect 8803 9401 8815 9435
rect 15930 9432 15936 9444
rect 15891 9404 15936 9432
rect 8757 9395 8815 9401
rect 15930 9392 15936 9404
rect 15988 9392 15994 9444
rect 3973 9367 4031 9373
rect 3973 9333 3985 9367
rect 4019 9333 4031 9367
rect 4338 9364 4344 9376
rect 4299 9336 4344 9364
rect 3973 9327 4031 9333
rect 4338 9324 4344 9336
rect 4396 9324 4402 9376
rect 7282 9324 7288 9376
rect 7340 9364 7346 9376
rect 7745 9367 7803 9373
rect 7745 9364 7757 9367
rect 7340 9336 7757 9364
rect 7340 9324 7346 9336
rect 7745 9333 7757 9336
rect 7791 9364 7803 9367
rect 8662 9364 8668 9376
rect 7791 9336 8668 9364
rect 7791 9333 7803 9336
rect 7745 9327 7803 9333
rect 8662 9324 8668 9336
rect 8720 9324 8726 9376
rect 8938 9364 8944 9376
rect 8899 9336 8944 9364
rect 8938 9324 8944 9336
rect 8996 9324 9002 9376
rect 9950 9324 9956 9376
rect 10008 9364 10014 9376
rect 10137 9367 10195 9373
rect 10137 9364 10149 9367
rect 10008 9336 10149 9364
rect 10008 9324 10014 9336
rect 10137 9333 10149 9336
rect 10183 9333 10195 9367
rect 10137 9327 10195 9333
rect 12345 9367 12403 9373
rect 12345 9333 12357 9367
rect 12391 9364 12403 9367
rect 12802 9364 12808 9376
rect 12391 9336 12808 9364
rect 12391 9333 12403 9336
rect 12345 9327 12403 9333
rect 12802 9324 12808 9336
rect 12860 9324 12866 9376
rect 15013 9367 15071 9373
rect 15013 9333 15025 9367
rect 15059 9364 15071 9367
rect 15102 9364 15108 9376
rect 15059 9336 15108 9364
rect 15059 9333 15071 9336
rect 15013 9327 15071 9333
rect 15102 9324 15108 9336
rect 15160 9324 15166 9376
rect 15286 9324 15292 9376
rect 15344 9364 15350 9376
rect 16117 9367 16175 9373
rect 16117 9364 16129 9367
rect 15344 9336 16129 9364
rect 15344 9324 15350 9336
rect 16117 9333 16129 9336
rect 16163 9333 16175 9367
rect 16117 9327 16175 9333
rect 184 9274 18920 9296
rect 184 9222 3106 9274
rect 3158 9222 3170 9274
rect 3222 9222 3234 9274
rect 3286 9222 3298 9274
rect 3350 9222 3362 9274
rect 3414 9222 6206 9274
rect 6258 9222 6270 9274
rect 6322 9222 6334 9274
rect 6386 9222 6398 9274
rect 6450 9222 6462 9274
rect 6514 9222 9306 9274
rect 9358 9222 9370 9274
rect 9422 9222 9434 9274
rect 9486 9222 9498 9274
rect 9550 9222 9562 9274
rect 9614 9222 12406 9274
rect 12458 9222 12470 9274
rect 12522 9222 12534 9274
rect 12586 9222 12598 9274
rect 12650 9222 12662 9274
rect 12714 9222 15506 9274
rect 15558 9222 15570 9274
rect 15622 9222 15634 9274
rect 15686 9222 15698 9274
rect 15750 9222 15762 9274
rect 15814 9222 18606 9274
rect 18658 9222 18670 9274
rect 18722 9222 18734 9274
rect 18786 9222 18798 9274
rect 18850 9222 18862 9274
rect 18914 9222 18920 9274
rect 184 9200 18920 9222
rect 2314 9160 2320 9172
rect 2275 9132 2320 9160
rect 2314 9120 2320 9132
rect 2372 9120 2378 9172
rect 3605 9163 3663 9169
rect 3605 9129 3617 9163
rect 3651 9160 3663 9163
rect 4338 9160 4344 9172
rect 3651 9132 4344 9160
rect 3651 9129 3663 9132
rect 3605 9123 3663 9129
rect 4338 9120 4344 9132
rect 4396 9120 4402 9172
rect 5169 9163 5227 9169
rect 5169 9129 5181 9163
rect 5215 9160 5227 9163
rect 5350 9160 5356 9172
rect 5215 9132 5356 9160
rect 5215 9129 5227 9132
rect 5169 9123 5227 9129
rect 5350 9120 5356 9132
rect 5408 9120 5414 9172
rect 7193 9163 7251 9169
rect 7193 9129 7205 9163
rect 7239 9160 7251 9163
rect 7282 9160 7288 9172
rect 7239 9132 7288 9160
rect 7239 9129 7251 9132
rect 7193 9123 7251 9129
rect 7282 9120 7288 9132
rect 7340 9120 7346 9172
rect 9214 9120 9220 9172
rect 9272 9160 9278 9172
rect 9355 9163 9413 9169
rect 9355 9160 9367 9163
rect 9272 9132 9367 9160
rect 9272 9120 9278 9132
rect 9355 9129 9367 9132
rect 9401 9129 9413 9163
rect 9355 9123 9413 9129
rect 11747 9163 11805 9169
rect 11747 9129 11759 9163
rect 11793 9160 11805 9163
rect 11974 9160 11980 9172
rect 11793 9132 11980 9160
rect 11793 9129 11805 9132
rect 11747 9123 11805 9129
rect 11974 9120 11980 9132
rect 12032 9120 12038 9172
rect 12802 9120 12808 9172
rect 12860 9160 12866 9172
rect 12989 9163 13047 9169
rect 12989 9160 13001 9163
rect 12860 9132 13001 9160
rect 12860 9120 12866 9132
rect 12989 9129 13001 9132
rect 13035 9129 13047 9163
rect 12989 9123 13047 9129
rect 18138 9120 18144 9172
rect 18196 9160 18202 9172
rect 18233 9163 18291 9169
rect 18233 9160 18245 9163
rect 18196 9132 18245 9160
rect 18196 9120 18202 9132
rect 18233 9129 18245 9132
rect 18279 9129 18291 9163
rect 18233 9123 18291 9129
rect 842 9092 848 9104
rect 803 9064 848 9092
rect 842 9052 848 9064
rect 900 9052 906 9104
rect 2866 9092 2872 9104
rect 2070 9064 2872 9092
rect 2866 9052 2872 9064
rect 2924 9052 2930 9104
rect 8662 9052 8668 9104
rect 8720 9052 8726 9104
rect 11238 9052 11244 9104
rect 11296 9052 11302 9104
rect 13262 9052 13268 9104
rect 13320 9092 13326 9104
rect 13538 9092 13544 9104
rect 13320 9064 13544 9092
rect 13320 9052 13326 9064
rect 13538 9052 13544 9064
rect 13596 9092 13602 9104
rect 13909 9095 13967 9101
rect 13909 9092 13921 9095
rect 13596 9064 13921 9092
rect 13596 9052 13602 9064
rect 13909 9061 13921 9064
rect 13955 9092 13967 9095
rect 14185 9095 14243 9101
rect 14185 9092 14197 9095
rect 13955 9064 14197 9092
rect 13955 9061 13967 9064
rect 13909 9055 13967 9061
rect 14185 9061 14197 9064
rect 14231 9061 14243 9095
rect 14185 9055 14243 9061
rect 16114 9052 16120 9104
rect 16172 9092 16178 9104
rect 16482 9092 16488 9104
rect 16172 9064 16488 9092
rect 16172 9052 16178 9064
rect 16482 9052 16488 9064
rect 16540 9052 16546 9104
rect 2958 8984 2964 9036
rect 3016 9024 3022 9036
rect 3145 9027 3203 9033
rect 3145 9024 3157 9027
rect 3016 8996 3157 9024
rect 3016 8984 3022 8996
rect 3145 8993 3157 8996
rect 3191 8993 3203 9027
rect 3145 8987 3203 8993
rect 3237 9027 3295 9033
rect 3237 8993 3249 9027
rect 3283 8993 3295 9027
rect 3418 9024 3424 9036
rect 3379 8996 3424 9024
rect 3237 8987 3295 8993
rect 566 8956 572 8968
rect 527 8928 572 8956
rect 566 8916 572 8928
rect 624 8916 630 8968
rect 3160 8888 3188 8987
rect 3252 8956 3280 8987
rect 3418 8984 3424 8996
rect 3476 8984 3482 9036
rect 6293 9027 6351 9033
rect 6293 8993 6305 9027
rect 6339 9024 6351 9027
rect 7006 9024 7012 9036
rect 6339 8996 7012 9024
rect 6339 8993 6351 8996
rect 6293 8987 6351 8993
rect 7006 8984 7012 8996
rect 7064 8984 7070 9036
rect 9950 9024 9956 9036
rect 9911 8996 9956 9024
rect 9950 8984 9956 8996
rect 10008 8984 10014 9036
rect 13633 9027 13691 9033
rect 13633 8993 13645 9027
rect 13679 9024 13691 9027
rect 13722 9024 13728 9036
rect 13679 8996 13728 9024
rect 13679 8993 13691 8996
rect 13633 8987 13691 8993
rect 13722 8984 13728 8996
rect 13780 8984 13786 9036
rect 13814 8984 13820 9036
rect 13872 9024 13878 9036
rect 14737 9027 14795 9033
rect 14737 9024 14749 9027
rect 13872 8996 14749 9024
rect 13872 8984 13878 8996
rect 14737 8993 14749 8996
rect 14783 8993 14795 9027
rect 15102 9024 15108 9036
rect 15063 8996 15108 9024
rect 14737 8987 14795 8993
rect 15102 8984 15108 8996
rect 15160 8984 15166 9036
rect 17957 9027 18015 9033
rect 17957 8993 17969 9027
rect 18003 9024 18015 9027
rect 18414 9024 18420 9036
rect 18003 8996 18420 9024
rect 18003 8993 18015 8996
rect 17957 8987 18015 8993
rect 18414 8984 18420 8996
rect 18472 8984 18478 9036
rect 4338 8956 4344 8968
rect 3252 8928 4344 8956
rect 4338 8916 4344 8928
rect 4396 8916 4402 8968
rect 6549 8959 6607 8965
rect 6549 8925 6561 8959
rect 6595 8956 6607 8959
rect 7558 8956 7564 8968
rect 6595 8928 7564 8956
rect 6595 8925 6607 8928
rect 6549 8919 6607 8925
rect 4430 8888 4436 8900
rect 3160 8860 4436 8888
rect 4430 8848 4436 8860
rect 4488 8848 4494 8900
rect 2866 8820 2872 8832
rect 2827 8792 2872 8820
rect 2866 8780 2872 8792
rect 2924 8780 2930 8832
rect 5534 8780 5540 8832
rect 5592 8820 5598 8832
rect 6564 8820 6592 8919
rect 7558 8916 7564 8928
rect 7616 8916 7622 8968
rect 7929 8959 7987 8965
rect 7929 8925 7941 8959
rect 7975 8956 7987 8959
rect 8110 8956 8116 8968
rect 7975 8928 8116 8956
rect 7975 8925 7987 8928
rect 7929 8919 7987 8925
rect 8110 8916 8116 8928
rect 8168 8916 8174 8968
rect 10318 8956 10324 8968
rect 10279 8928 10324 8956
rect 10318 8916 10324 8928
rect 10376 8916 10382 8968
rect 13078 8956 13084 8968
rect 13039 8928 13084 8956
rect 13078 8916 13084 8928
rect 13136 8916 13142 8968
rect 13262 8956 13268 8968
rect 13223 8928 13268 8956
rect 13262 8916 13268 8928
rect 13320 8916 13326 8968
rect 16206 8916 16212 8968
rect 16264 8956 16270 8968
rect 16531 8959 16589 8965
rect 16531 8956 16543 8959
rect 16264 8928 16543 8956
rect 16264 8916 16270 8928
rect 16531 8925 16543 8928
rect 16577 8925 16589 8959
rect 16531 8919 16589 8925
rect 13725 8891 13783 8897
rect 13725 8857 13737 8891
rect 13771 8888 13783 8891
rect 13814 8888 13820 8900
rect 13771 8860 13820 8888
rect 13771 8857 13783 8860
rect 13725 8851 13783 8857
rect 13814 8848 13820 8860
rect 13872 8888 13878 8900
rect 14734 8888 14740 8900
rect 13872 8860 14740 8888
rect 13872 8848 13878 8860
rect 14734 8848 14740 8860
rect 14792 8848 14798 8900
rect 12618 8820 12624 8832
rect 5592 8792 6592 8820
rect 12579 8792 12624 8820
rect 5592 8780 5598 8792
rect 12618 8780 12624 8792
rect 12676 8780 12682 8832
rect 13630 8820 13636 8832
rect 13591 8792 13636 8820
rect 13630 8780 13636 8792
rect 13688 8780 13694 8832
rect 184 8730 18860 8752
rect 184 8678 1556 8730
rect 1608 8678 1620 8730
rect 1672 8678 1684 8730
rect 1736 8678 1748 8730
rect 1800 8678 1812 8730
rect 1864 8678 4656 8730
rect 4708 8678 4720 8730
rect 4772 8678 4784 8730
rect 4836 8678 4848 8730
rect 4900 8678 4912 8730
rect 4964 8678 7756 8730
rect 7808 8678 7820 8730
rect 7872 8678 7884 8730
rect 7936 8678 7948 8730
rect 8000 8678 8012 8730
rect 8064 8678 10856 8730
rect 10908 8678 10920 8730
rect 10972 8678 10984 8730
rect 11036 8678 11048 8730
rect 11100 8678 11112 8730
rect 11164 8678 13956 8730
rect 14008 8678 14020 8730
rect 14072 8678 14084 8730
rect 14136 8678 14148 8730
rect 14200 8678 14212 8730
rect 14264 8678 17056 8730
rect 17108 8678 17120 8730
rect 17172 8678 17184 8730
rect 17236 8678 17248 8730
rect 17300 8678 17312 8730
rect 17364 8678 18860 8730
rect 184 8656 18860 8678
rect 2590 8616 2596 8628
rect 2551 8588 2596 8616
rect 2590 8576 2596 8588
rect 2648 8576 2654 8628
rect 2961 8619 3019 8625
rect 2961 8585 2973 8619
rect 3007 8616 3019 8619
rect 3418 8616 3424 8628
rect 3007 8588 3424 8616
rect 3007 8585 3019 8588
rect 2961 8579 3019 8585
rect 3418 8576 3424 8588
rect 3476 8576 3482 8628
rect 6914 8616 6920 8628
rect 6875 8588 6920 8616
rect 6914 8576 6920 8588
rect 6972 8576 6978 8628
rect 8110 8616 8116 8628
rect 8071 8588 8116 8616
rect 8110 8576 8116 8588
rect 8168 8576 8174 8628
rect 8570 8576 8576 8628
rect 8628 8616 8634 8628
rect 8849 8619 8907 8625
rect 8849 8616 8861 8619
rect 8628 8588 8861 8616
rect 8628 8576 8634 8588
rect 8849 8585 8861 8588
rect 8895 8585 8907 8619
rect 8849 8579 8907 8585
rect 10318 8576 10324 8628
rect 10376 8616 10382 8628
rect 11149 8619 11207 8625
rect 11149 8616 11161 8619
rect 10376 8588 11161 8616
rect 10376 8576 10382 8588
rect 11149 8585 11161 8588
rect 11195 8585 11207 8619
rect 11149 8579 11207 8585
rect 13078 8576 13084 8628
rect 13136 8616 13142 8628
rect 13541 8619 13599 8625
rect 13541 8616 13553 8619
rect 13136 8588 13553 8616
rect 13136 8576 13142 8588
rect 13541 8585 13553 8588
rect 13587 8585 13599 8619
rect 13541 8579 13599 8585
rect 13814 8576 13820 8628
rect 13872 8616 13878 8628
rect 14001 8619 14059 8625
rect 14001 8616 14013 8619
rect 13872 8588 14013 8616
rect 13872 8576 13878 8588
rect 14001 8585 14013 8588
rect 14047 8585 14059 8619
rect 14001 8579 14059 8585
rect 17678 8576 17684 8628
rect 17736 8616 17742 8628
rect 17911 8619 17969 8625
rect 17911 8616 17923 8619
rect 17736 8588 17923 8616
rect 17736 8576 17742 8588
rect 17911 8585 17923 8588
rect 17957 8585 17969 8619
rect 17911 8579 17969 8585
rect 2608 8548 2636 8576
rect 8021 8551 8079 8557
rect 2608 8520 3280 8548
rect 2314 8440 2320 8492
rect 2372 8480 2378 8492
rect 2372 8452 2820 8480
rect 2372 8440 2378 8452
rect 2792 8421 2820 8452
rect 3252 8421 3280 8520
rect 8021 8517 8033 8551
rect 8067 8548 8079 8551
rect 8938 8548 8944 8560
rect 8067 8520 8944 8548
rect 8067 8517 8079 8520
rect 8021 8511 8079 8517
rect 8938 8508 8944 8520
rect 8996 8508 9002 8560
rect 12618 8548 12624 8560
rect 11624 8520 12624 8548
rect 8202 8480 8208 8492
rect 6748 8452 8064 8480
rect 8163 8452 8208 8480
rect 2501 8415 2559 8421
rect 2501 8381 2513 8415
rect 2547 8381 2559 8415
rect 2501 8375 2559 8381
rect 2777 8415 2835 8421
rect 2777 8381 2789 8415
rect 2823 8381 2835 8415
rect 2777 8375 2835 8381
rect 3237 8415 3295 8421
rect 3237 8381 3249 8415
rect 3283 8381 3295 8415
rect 5534 8412 5540 8424
rect 5495 8384 5540 8412
rect 3237 8375 3295 8381
rect 2516 8344 2544 8375
rect 5534 8372 5540 8384
rect 5592 8372 5598 8424
rect 6748 8421 6776 8452
rect 6733 8415 6791 8421
rect 6733 8381 6745 8415
rect 6779 8381 6791 8415
rect 6733 8375 6791 8381
rect 7006 8372 7012 8424
rect 7064 8412 7070 8424
rect 7064 8384 7157 8412
rect 7064 8372 7070 8384
rect 7190 8372 7196 8424
rect 7248 8412 7254 8424
rect 7929 8415 7987 8421
rect 7929 8412 7941 8415
rect 7248 8384 7941 8412
rect 7248 8372 7254 8384
rect 7929 8381 7941 8384
rect 7975 8381 7987 8415
rect 8036 8412 8064 8452
rect 8202 8440 8208 8452
rect 8260 8440 8266 8492
rect 11624 8489 11652 8520
rect 12618 8508 12624 8520
rect 12676 8508 12682 8560
rect 11609 8483 11667 8489
rect 11609 8449 11621 8483
rect 11655 8449 11667 8483
rect 11790 8480 11796 8492
rect 11751 8452 11796 8480
rect 11609 8443 11667 8449
rect 11790 8440 11796 8452
rect 11848 8440 11854 8492
rect 16117 8483 16175 8489
rect 16117 8449 16129 8483
rect 16163 8480 16175 8483
rect 16298 8480 16304 8492
rect 16163 8452 16304 8480
rect 16163 8449 16175 8452
rect 16117 8443 16175 8449
rect 16298 8440 16304 8452
rect 16356 8440 16362 8492
rect 8386 8412 8392 8424
rect 8036 8384 8392 8412
rect 7929 8375 7987 8381
rect 8386 8372 8392 8384
rect 8444 8372 8450 8424
rect 9122 8412 9128 8424
rect 9083 8384 9128 8412
rect 9122 8372 9128 8384
rect 9180 8372 9186 8424
rect 11517 8415 11575 8421
rect 11517 8381 11529 8415
rect 11563 8412 11575 8415
rect 11974 8412 11980 8424
rect 11563 8384 11980 8412
rect 11563 8381 11575 8384
rect 11517 8375 11575 8381
rect 11974 8372 11980 8384
rect 12032 8372 12038 8424
rect 13170 8372 13176 8424
rect 13228 8412 13234 8424
rect 13541 8415 13599 8421
rect 13541 8412 13553 8415
rect 13228 8384 13553 8412
rect 13228 8372 13234 8384
rect 13541 8381 13553 8384
rect 13587 8381 13599 8415
rect 13541 8375 13599 8381
rect 13630 8372 13636 8424
rect 13688 8412 13694 8424
rect 13725 8415 13783 8421
rect 13725 8412 13737 8415
rect 13688 8384 13737 8412
rect 13688 8372 13694 8384
rect 13725 8381 13737 8384
rect 13771 8381 13783 8415
rect 13725 8375 13783 8381
rect 16485 8415 16543 8421
rect 16485 8381 16497 8415
rect 16531 8412 16543 8415
rect 16574 8412 16580 8424
rect 16531 8384 16580 8412
rect 16531 8381 16543 8384
rect 16485 8375 16543 8381
rect 16574 8372 16580 8384
rect 16632 8372 16638 8424
rect 2682 8344 2688 8356
rect 2516 8316 2688 8344
rect 2682 8304 2688 8316
rect 2740 8304 2746 8356
rect 3329 8347 3387 8353
rect 3329 8313 3341 8347
rect 3375 8344 3387 8347
rect 4338 8344 4344 8356
rect 3375 8316 4344 8344
rect 3375 8313 3387 8316
rect 3329 8307 3387 8313
rect 4338 8304 4344 8316
rect 4396 8304 4402 8356
rect 5258 8344 5264 8356
rect 5219 8316 5264 8344
rect 5258 8304 5264 8316
rect 5316 8304 5322 8356
rect 6546 8344 6552 8356
rect 6507 8316 6552 8344
rect 6546 8304 6552 8316
rect 6604 8304 6610 8356
rect 7024 8344 7052 8372
rect 9950 8344 9956 8356
rect 7024 8316 9956 8344
rect 9950 8304 9956 8316
rect 10008 8304 10014 8356
rect 16776 8316 16882 8344
rect 9674 8236 9680 8288
rect 9732 8276 9738 8288
rect 10781 8279 10839 8285
rect 10781 8276 10793 8279
rect 9732 8248 10793 8276
rect 9732 8236 9738 8248
rect 10781 8245 10793 8248
rect 10827 8276 10839 8279
rect 10870 8276 10876 8288
rect 10827 8248 10876 8276
rect 10827 8245 10839 8248
rect 10781 8239 10839 8245
rect 10870 8236 10876 8248
rect 10928 8236 10934 8288
rect 16482 8236 16488 8288
rect 16540 8276 16546 8288
rect 16776 8276 16804 8316
rect 16540 8248 16804 8276
rect 16540 8236 16546 8248
rect 184 8186 18920 8208
rect 184 8134 3106 8186
rect 3158 8134 3170 8186
rect 3222 8134 3234 8186
rect 3286 8134 3298 8186
rect 3350 8134 3362 8186
rect 3414 8134 6206 8186
rect 6258 8134 6270 8186
rect 6322 8134 6334 8186
rect 6386 8134 6398 8186
rect 6450 8134 6462 8186
rect 6514 8134 9306 8186
rect 9358 8134 9370 8186
rect 9422 8134 9434 8186
rect 9486 8134 9498 8186
rect 9550 8134 9562 8186
rect 9614 8134 12406 8186
rect 12458 8134 12470 8186
rect 12522 8134 12534 8186
rect 12586 8134 12598 8186
rect 12650 8134 12662 8186
rect 12714 8134 15506 8186
rect 15558 8134 15570 8186
rect 15622 8134 15634 8186
rect 15686 8134 15698 8186
rect 15750 8134 15762 8186
rect 15814 8134 18606 8186
rect 18658 8134 18670 8186
rect 18722 8134 18734 8186
rect 18786 8134 18798 8186
rect 18850 8134 18862 8186
rect 18914 8134 18920 8186
rect 184 8112 18920 8134
rect 2409 8075 2467 8081
rect 2409 8041 2421 8075
rect 2455 8072 2467 8075
rect 2590 8072 2596 8084
rect 2455 8044 2596 8072
rect 2455 8041 2467 8044
rect 2409 8035 2467 8041
rect 2590 8032 2596 8044
rect 2648 8032 2654 8084
rect 3237 8075 3295 8081
rect 3237 8041 3249 8075
rect 3283 8072 3295 8075
rect 5442 8072 5448 8084
rect 3283 8044 5448 8072
rect 3283 8041 3295 8044
rect 3237 8035 3295 8041
rect 5442 8032 5448 8044
rect 5500 8032 5506 8084
rect 13262 8032 13268 8084
rect 13320 8072 13326 8084
rect 15930 8072 15936 8084
rect 13320 8044 15936 8072
rect 13320 8032 13326 8044
rect 2866 8004 2872 8016
rect 2162 7976 2872 8004
rect 2866 7964 2872 7976
rect 2924 7964 2930 8016
rect 4522 8004 4528 8016
rect 4483 7976 4528 8004
rect 4522 7964 4528 7976
rect 4580 7964 4586 8016
rect 7282 8004 7288 8016
rect 6578 7976 7288 8004
rect 7282 7964 7288 7976
rect 7340 7964 7346 8016
rect 9766 7964 9772 8016
rect 9824 8004 9830 8016
rect 10321 8007 10379 8013
rect 10321 8004 10333 8007
rect 9824 7976 10333 8004
rect 9824 7964 9830 7976
rect 10321 7973 10333 7976
rect 10367 7973 10379 8007
rect 10321 7967 10379 7973
rect 11149 8007 11207 8013
rect 11149 7973 11161 8007
rect 11195 8004 11207 8007
rect 11238 8004 11244 8016
rect 11195 7976 11244 8004
rect 11195 7973 11207 7976
rect 11149 7967 11207 7973
rect 11238 7964 11244 7976
rect 11296 7964 11302 8016
rect 14366 8004 14372 8016
rect 14327 7976 14372 8004
rect 14366 7964 14372 7976
rect 14424 7964 14430 8016
rect 5169 7939 5227 7945
rect 5169 7905 5181 7939
rect 5215 7936 5227 7939
rect 5258 7936 5264 7948
rect 5215 7908 5264 7936
rect 5215 7905 5227 7908
rect 5169 7899 5227 7905
rect 5258 7896 5264 7908
rect 5316 7896 5322 7948
rect 6914 7896 6920 7948
rect 6972 7936 6978 7948
rect 7929 7939 7987 7945
rect 7929 7936 7941 7939
rect 6972 7908 7941 7936
rect 6972 7896 6978 7908
rect 7929 7905 7941 7908
rect 7975 7936 7987 7939
rect 8297 7939 8355 7945
rect 7975 7908 8248 7936
rect 7975 7905 7987 7908
rect 7929 7899 7987 7905
rect 566 7828 572 7880
rect 624 7868 630 7880
rect 661 7871 719 7877
rect 661 7868 673 7871
rect 624 7840 673 7868
rect 624 7828 630 7840
rect 661 7837 673 7840
rect 707 7837 719 7871
rect 934 7868 940 7880
rect 895 7840 940 7868
rect 661 7831 719 7837
rect 934 7828 940 7840
rect 992 7828 998 7880
rect 5537 7871 5595 7877
rect 5537 7837 5549 7871
rect 5583 7868 5595 7871
rect 5718 7868 5724 7880
rect 5583 7840 5724 7868
rect 5583 7837 5595 7840
rect 5537 7831 5595 7837
rect 5718 7828 5724 7840
rect 5776 7828 5782 7880
rect 7374 7828 7380 7880
rect 7432 7868 7438 7880
rect 8110 7868 8116 7880
rect 7432 7840 8116 7868
rect 7432 7828 7438 7840
rect 8110 7828 8116 7840
rect 8168 7828 8174 7880
rect 7466 7760 7472 7812
rect 7524 7800 7530 7812
rect 7650 7800 7656 7812
rect 7524 7772 7656 7800
rect 7524 7760 7530 7772
rect 7650 7760 7656 7772
rect 7708 7800 7714 7812
rect 7929 7803 7987 7809
rect 7929 7800 7941 7803
rect 7708 7772 7941 7800
rect 7708 7760 7714 7772
rect 7929 7769 7941 7772
rect 7975 7769 7987 7803
rect 8220 7800 8248 7908
rect 8297 7905 8309 7939
rect 8343 7936 8355 7939
rect 8386 7936 8392 7948
rect 8343 7908 8392 7936
rect 8343 7905 8355 7908
rect 8297 7899 8355 7905
rect 8386 7896 8392 7908
rect 8444 7896 8450 7948
rect 8754 7896 8760 7948
rect 8812 7936 8818 7948
rect 9033 7939 9091 7945
rect 9033 7936 9045 7939
rect 8812 7908 9045 7936
rect 8812 7896 8818 7908
rect 9033 7905 9045 7908
rect 9079 7905 9091 7939
rect 10870 7936 10876 7948
rect 10831 7908 10876 7936
rect 9033 7899 9091 7905
rect 10870 7896 10876 7908
rect 10928 7896 10934 7948
rect 14921 7939 14979 7945
rect 14921 7905 14933 7939
rect 14967 7905 14979 7939
rect 14921 7899 14979 7905
rect 15013 7939 15071 7945
rect 15013 7905 15025 7939
rect 15059 7936 15071 7939
rect 15194 7936 15200 7948
rect 15059 7908 15200 7936
rect 15059 7905 15071 7908
rect 15013 7899 15071 7905
rect 8404 7868 8432 7896
rect 8849 7871 8907 7877
rect 8849 7868 8861 7871
rect 8404 7840 8861 7868
rect 8849 7837 8861 7840
rect 8895 7837 8907 7871
rect 14936 7868 14964 7899
rect 15194 7896 15200 7908
rect 15252 7896 15258 7948
rect 15304 7945 15332 8044
rect 15930 8032 15936 8044
rect 15988 8032 15994 8084
rect 16574 8072 16580 8084
rect 16535 8044 16580 8072
rect 16574 8032 16580 8044
rect 16632 8032 16638 8084
rect 17678 8032 17684 8084
rect 17736 8072 17742 8084
rect 17773 8075 17831 8081
rect 17773 8072 17785 8075
rect 17736 8044 17785 8072
rect 17736 8032 17742 8044
rect 17773 8041 17785 8044
rect 17819 8041 17831 8075
rect 17773 8035 17831 8041
rect 15657 8007 15715 8013
rect 15657 7973 15669 8007
rect 15703 8004 15715 8007
rect 15838 8004 15844 8016
rect 15703 7976 15844 8004
rect 15703 7973 15715 7976
rect 15657 7967 15715 7973
rect 15838 7964 15844 7976
rect 15896 7964 15902 8016
rect 15289 7939 15347 7945
rect 15289 7905 15301 7939
rect 15335 7905 15347 7939
rect 16574 7936 16580 7948
rect 16535 7908 16580 7936
rect 15289 7899 15347 7905
rect 16574 7896 16580 7908
rect 16632 7896 16638 7948
rect 16761 7939 16819 7945
rect 16761 7905 16773 7939
rect 16807 7936 16819 7939
rect 17129 7939 17187 7945
rect 17129 7936 17141 7939
rect 16807 7908 17141 7936
rect 16807 7905 16819 7908
rect 16761 7899 16819 7905
rect 17129 7905 17141 7908
rect 17175 7905 17187 7939
rect 17129 7899 17187 7905
rect 16666 7868 16672 7880
rect 14936 7840 16672 7868
rect 8849 7831 8907 7837
rect 16666 7828 16672 7840
rect 16724 7828 16730 7880
rect 17310 7868 17316 7880
rect 17271 7840 17316 7868
rect 17310 7828 17316 7840
rect 17368 7828 17374 7880
rect 17405 7871 17463 7877
rect 17405 7837 17417 7871
rect 17451 7868 17463 7871
rect 17770 7868 17776 7880
rect 17451 7840 17776 7868
rect 17451 7837 17463 7840
rect 17405 7831 17463 7837
rect 17770 7828 17776 7840
rect 17828 7828 17834 7880
rect 9214 7800 9220 7812
rect 8220 7772 9220 7800
rect 7929 7763 7987 7769
rect 9214 7760 9220 7772
rect 9272 7800 9278 7812
rect 10045 7803 10103 7809
rect 10045 7800 10057 7803
rect 9272 7772 10057 7800
rect 9272 7760 9278 7772
rect 10045 7769 10057 7772
rect 10091 7769 10103 7803
rect 10045 7763 10103 7769
rect 15197 7803 15255 7809
rect 15197 7769 15209 7803
rect 15243 7800 15255 7803
rect 15378 7800 15384 7812
rect 15243 7772 15384 7800
rect 15243 7769 15255 7772
rect 15197 7763 15255 7769
rect 15378 7760 15384 7772
rect 15436 7760 15442 7812
rect 6822 7692 6828 7744
rect 6880 7732 6886 7744
rect 6963 7735 7021 7741
rect 6963 7732 6975 7735
rect 6880 7704 6975 7732
rect 6880 7692 6886 7704
rect 6963 7701 6975 7704
rect 7009 7701 7021 7735
rect 6963 7695 7021 7701
rect 13081 7735 13139 7741
rect 13081 7701 13093 7735
rect 13127 7732 13139 7735
rect 13814 7732 13820 7744
rect 13127 7704 13820 7732
rect 13127 7701 13139 7704
rect 13081 7695 13139 7701
rect 13814 7692 13820 7704
rect 13872 7692 13878 7744
rect 14734 7732 14740 7744
rect 14695 7704 14740 7732
rect 14734 7692 14740 7704
rect 14792 7692 14798 7744
rect 184 7642 18860 7664
rect 184 7590 1556 7642
rect 1608 7590 1620 7642
rect 1672 7590 1684 7642
rect 1736 7590 1748 7642
rect 1800 7590 1812 7642
rect 1864 7590 4656 7642
rect 4708 7590 4720 7642
rect 4772 7590 4784 7642
rect 4836 7590 4848 7642
rect 4900 7590 4912 7642
rect 4964 7590 7756 7642
rect 7808 7590 7820 7642
rect 7872 7590 7884 7642
rect 7936 7590 7948 7642
rect 8000 7590 8012 7642
rect 8064 7590 10856 7642
rect 10908 7590 10920 7642
rect 10972 7590 10984 7642
rect 11036 7590 11048 7642
rect 11100 7590 11112 7642
rect 11164 7590 13956 7642
rect 14008 7590 14020 7642
rect 14072 7590 14084 7642
rect 14136 7590 14148 7642
rect 14200 7590 14212 7642
rect 14264 7590 17056 7642
rect 17108 7590 17120 7642
rect 17172 7590 17184 7642
rect 17236 7590 17248 7642
rect 17300 7590 17312 7642
rect 17364 7590 18860 7642
rect 184 7568 18860 7590
rect 934 7488 940 7540
rect 992 7528 998 7540
rect 1581 7531 1639 7537
rect 1581 7528 1593 7531
rect 992 7500 1593 7528
rect 992 7488 998 7500
rect 1581 7497 1593 7500
rect 1627 7497 1639 7531
rect 1581 7491 1639 7497
rect 4246 7488 4252 7540
rect 4304 7528 4310 7540
rect 4304 7500 4568 7528
rect 4304 7488 4310 7500
rect 3605 7463 3663 7469
rect 3605 7429 3617 7463
rect 3651 7460 3663 7463
rect 3651 7432 4476 7460
rect 3651 7429 3663 7432
rect 3605 7423 3663 7429
rect 2130 7392 2136 7404
rect 2091 7364 2136 7392
rect 2130 7352 2136 7364
rect 2188 7352 2194 7404
rect 2774 7352 2780 7404
rect 2832 7392 2838 7404
rect 3145 7395 3203 7401
rect 3145 7392 3157 7395
rect 2832 7364 3157 7392
rect 2832 7352 2838 7364
rect 3145 7361 3157 7364
rect 3191 7392 3203 7395
rect 3786 7392 3792 7404
rect 3191 7364 3792 7392
rect 3191 7361 3203 7364
rect 3145 7355 3203 7361
rect 3786 7352 3792 7364
rect 3844 7352 3850 7404
rect 4448 7401 4476 7432
rect 4540 7401 4568 7500
rect 8110 7488 8116 7540
rect 8168 7528 8174 7540
rect 9861 7531 9919 7537
rect 8168 7500 9352 7528
rect 8168 7488 8174 7500
rect 8938 7460 8944 7472
rect 8899 7432 8944 7460
rect 8938 7420 8944 7432
rect 8996 7420 9002 7472
rect 9214 7460 9220 7472
rect 9175 7432 9220 7460
rect 9214 7420 9220 7432
rect 9272 7420 9278 7472
rect 4433 7395 4491 7401
rect 4433 7361 4445 7395
rect 4479 7361 4491 7395
rect 4433 7355 4491 7361
rect 4525 7395 4583 7401
rect 4525 7361 4537 7395
rect 4571 7361 4583 7395
rect 4525 7355 4583 7361
rect 8386 7352 8392 7404
rect 8444 7392 8450 7404
rect 9324 7401 9352 7500
rect 9861 7497 9873 7531
rect 9907 7528 9919 7531
rect 10410 7528 10416 7540
rect 9907 7500 10416 7528
rect 9907 7497 9919 7500
rect 9861 7491 9919 7497
rect 9033 7395 9091 7401
rect 9033 7392 9045 7395
rect 8444 7364 9045 7392
rect 8444 7352 8450 7364
rect 9033 7361 9045 7364
rect 9079 7361 9091 7395
rect 9033 7355 9091 7361
rect 9309 7395 9367 7401
rect 9309 7361 9321 7395
rect 9355 7392 9367 7395
rect 9876 7392 9904 7491
rect 10410 7488 10416 7500
rect 10468 7488 10474 7540
rect 11238 7488 11244 7540
rect 11296 7528 11302 7540
rect 12250 7528 12256 7540
rect 11296 7500 12256 7528
rect 11296 7488 11302 7500
rect 12250 7488 12256 7500
rect 12308 7528 12314 7540
rect 15565 7531 15623 7537
rect 12308 7500 15332 7528
rect 12308 7488 12314 7500
rect 11790 7392 11796 7404
rect 9355 7364 9904 7392
rect 11751 7364 11796 7392
rect 9355 7361 9367 7364
rect 9309 7355 9367 7361
rect 11790 7352 11796 7364
rect 11848 7352 11854 7404
rect 12805 7395 12863 7401
rect 12805 7361 12817 7395
rect 12851 7392 12863 7395
rect 13262 7392 13268 7404
rect 12851 7364 13268 7392
rect 12851 7361 12863 7364
rect 12805 7355 12863 7361
rect 13262 7352 13268 7364
rect 13320 7352 13326 7404
rect 14093 7395 14151 7401
rect 14093 7361 14105 7395
rect 14139 7392 14151 7395
rect 14734 7392 14740 7404
rect 14139 7364 14740 7392
rect 14139 7361 14151 7364
rect 14093 7355 14151 7361
rect 14734 7352 14740 7364
rect 14792 7352 14798 7404
rect 1949 7327 2007 7333
rect 1949 7293 1961 7327
rect 1995 7324 2007 7327
rect 2590 7324 2596 7336
rect 1995 7296 2596 7324
rect 1995 7293 2007 7296
rect 1949 7287 2007 7293
rect 2590 7284 2596 7296
rect 2648 7284 2654 7336
rect 3237 7327 3295 7333
rect 3237 7293 3249 7327
rect 3283 7324 3295 7327
rect 3602 7324 3608 7336
rect 3283 7296 3608 7324
rect 3283 7293 3295 7296
rect 3237 7287 3295 7293
rect 3602 7284 3608 7296
rect 3660 7284 3666 7336
rect 4338 7324 4344 7336
rect 4299 7296 4344 7324
rect 4338 7284 4344 7296
rect 4396 7284 4402 7336
rect 6822 7324 6828 7336
rect 6783 7296 6828 7324
rect 6822 7284 6828 7296
rect 6880 7284 6886 7336
rect 8294 7284 8300 7336
rect 8352 7324 8358 7336
rect 8849 7327 8907 7333
rect 8849 7324 8861 7327
rect 8352 7296 8861 7324
rect 8352 7284 8358 7296
rect 8849 7293 8861 7296
rect 8895 7293 8907 7327
rect 9950 7324 9956 7336
rect 9911 7296 9956 7324
rect 8849 7287 8907 7293
rect 9950 7284 9956 7296
rect 10008 7284 10014 7336
rect 10778 7324 10784 7336
rect 10739 7296 10784 7324
rect 10778 7284 10784 7296
rect 10836 7324 10842 7336
rect 11517 7327 11575 7333
rect 11517 7324 11529 7327
rect 10836 7296 11529 7324
rect 10836 7284 10842 7296
rect 11517 7293 11529 7296
rect 11563 7324 11575 7327
rect 11882 7324 11888 7336
rect 11563 7296 11888 7324
rect 11563 7293 11575 7296
rect 11517 7287 11575 7293
rect 11882 7284 11888 7296
rect 11940 7284 11946 7336
rect 12529 7327 12587 7333
rect 12529 7324 12541 7327
rect 12406 7296 12541 7324
rect 2041 7259 2099 7265
rect 2041 7225 2053 7259
rect 2087 7256 2099 7259
rect 2087 7228 4016 7256
rect 2087 7225 2099 7228
rect 2041 7219 2099 7225
rect 2685 7191 2743 7197
rect 2685 7157 2697 7191
rect 2731 7188 2743 7191
rect 2866 7188 2872 7200
rect 2731 7160 2872 7188
rect 2731 7157 2743 7160
rect 2685 7151 2743 7157
rect 2866 7148 2872 7160
rect 2924 7148 2930 7200
rect 3988 7197 4016 7228
rect 5810 7216 5816 7268
rect 5868 7256 5874 7268
rect 6365 7259 6423 7265
rect 6365 7256 6377 7259
rect 5868 7228 6377 7256
rect 5868 7216 5874 7228
rect 6365 7225 6377 7228
rect 6411 7225 6423 7259
rect 6365 7219 6423 7225
rect 8941 7259 8999 7265
rect 8941 7225 8953 7259
rect 8987 7256 8999 7259
rect 10689 7259 10747 7265
rect 8987 7228 9904 7256
rect 8987 7225 8999 7228
rect 8941 7219 8999 7225
rect 3973 7191 4031 7197
rect 3973 7157 3985 7191
rect 4019 7157 4031 7191
rect 3973 7151 4031 7157
rect 5077 7191 5135 7197
rect 5077 7157 5089 7191
rect 5123 7188 5135 7191
rect 5902 7188 5908 7200
rect 5123 7160 5908 7188
rect 5123 7157 5135 7160
rect 5077 7151 5135 7157
rect 5902 7148 5908 7160
rect 5960 7148 5966 7200
rect 9876 7188 9904 7228
rect 10689 7225 10701 7259
rect 10735 7256 10747 7259
rect 12406 7256 12434 7296
rect 12529 7293 12541 7296
rect 12575 7324 12587 7327
rect 12894 7324 12900 7336
rect 12575 7296 12900 7324
rect 12575 7293 12587 7296
rect 12529 7287 12587 7293
rect 12894 7284 12900 7296
rect 12952 7284 12958 7336
rect 13814 7324 13820 7336
rect 13775 7296 13820 7324
rect 13814 7284 13820 7296
rect 13872 7284 13878 7336
rect 10735 7228 12434 7256
rect 15304 7256 15332 7500
rect 15565 7497 15577 7531
rect 15611 7528 15623 7531
rect 15838 7528 15844 7540
rect 15611 7500 15844 7528
rect 15611 7497 15623 7500
rect 15565 7491 15623 7497
rect 15838 7488 15844 7500
rect 15896 7488 15902 7540
rect 16574 7488 16580 7540
rect 16632 7528 16638 7540
rect 17221 7531 17279 7537
rect 17221 7528 17233 7531
rect 16632 7500 17233 7528
rect 16632 7488 16638 7500
rect 17221 7497 17233 7500
rect 17267 7497 17279 7531
rect 17221 7491 17279 7497
rect 15838 7352 15844 7404
rect 15896 7392 15902 7404
rect 15896 7364 16160 7392
rect 15896 7352 15902 7364
rect 15930 7324 15936 7336
rect 15891 7296 15936 7324
rect 15930 7284 15936 7296
rect 15988 7284 15994 7336
rect 16132 7333 16160 7364
rect 16117 7327 16175 7333
rect 16117 7293 16129 7327
rect 16163 7324 16175 7327
rect 16393 7327 16451 7333
rect 16393 7324 16405 7327
rect 16163 7296 16405 7324
rect 16163 7293 16175 7296
rect 16117 7287 16175 7293
rect 16393 7293 16405 7296
rect 16439 7293 16451 7327
rect 17402 7324 17408 7336
rect 17363 7296 17408 7324
rect 16393 7287 16451 7293
rect 17402 7284 17408 7296
rect 17460 7284 17466 7336
rect 17497 7327 17555 7333
rect 17497 7293 17509 7327
rect 17543 7293 17555 7327
rect 17497 7287 17555 7293
rect 17589 7327 17647 7333
rect 17589 7293 17601 7327
rect 17635 7324 17647 7327
rect 17678 7324 17684 7336
rect 17635 7296 17684 7324
rect 17635 7293 17647 7296
rect 17589 7287 17647 7293
rect 16482 7256 16488 7268
rect 15304 7242 16488 7256
rect 15318 7228 16488 7242
rect 10735 7225 10747 7228
rect 10689 7219 10747 7225
rect 16482 7216 16488 7228
rect 16540 7216 16546 7268
rect 17512 7256 17540 7287
rect 17678 7284 17684 7296
rect 17736 7284 17742 7336
rect 17770 7256 17776 7268
rect 17512 7228 17776 7256
rect 17770 7216 17776 7228
rect 17828 7216 17834 7268
rect 10778 7188 10784 7200
rect 9876 7160 10784 7188
rect 10778 7148 10784 7160
rect 10836 7148 10842 7200
rect 11146 7188 11152 7200
rect 11107 7160 11152 7188
rect 11146 7148 11152 7160
rect 11204 7148 11210 7200
rect 11609 7191 11667 7197
rect 11609 7157 11621 7191
rect 11655 7188 11667 7191
rect 12161 7191 12219 7197
rect 12161 7188 12173 7191
rect 11655 7160 12173 7188
rect 11655 7157 11667 7160
rect 11609 7151 11667 7157
rect 12161 7157 12173 7160
rect 12207 7157 12219 7191
rect 12161 7151 12219 7157
rect 12621 7191 12679 7197
rect 12621 7157 12633 7191
rect 12667 7188 12679 7191
rect 12802 7188 12808 7200
rect 12667 7160 12808 7188
rect 12667 7157 12679 7160
rect 12621 7151 12679 7157
rect 12802 7148 12808 7160
rect 12860 7148 12866 7200
rect 15010 7148 15016 7200
rect 15068 7188 15074 7200
rect 15838 7188 15844 7200
rect 15068 7160 15844 7188
rect 15068 7148 15074 7160
rect 15838 7148 15844 7160
rect 15896 7148 15902 7200
rect 16022 7188 16028 7200
rect 15983 7160 16028 7188
rect 16022 7148 16028 7160
rect 16080 7148 16086 7200
rect 184 7098 18920 7120
rect 184 7046 3106 7098
rect 3158 7046 3170 7098
rect 3222 7046 3234 7098
rect 3286 7046 3298 7098
rect 3350 7046 3362 7098
rect 3414 7046 6206 7098
rect 6258 7046 6270 7098
rect 6322 7046 6334 7098
rect 6386 7046 6398 7098
rect 6450 7046 6462 7098
rect 6514 7046 9306 7098
rect 9358 7046 9370 7098
rect 9422 7046 9434 7098
rect 9486 7046 9498 7098
rect 9550 7046 9562 7098
rect 9614 7046 12406 7098
rect 12458 7046 12470 7098
rect 12522 7046 12534 7098
rect 12586 7046 12598 7098
rect 12650 7046 12662 7098
rect 12714 7046 15506 7098
rect 15558 7046 15570 7098
rect 15622 7046 15634 7098
rect 15686 7046 15698 7098
rect 15750 7046 15762 7098
rect 15814 7046 18606 7098
rect 18658 7046 18670 7098
rect 18722 7046 18734 7098
rect 18786 7046 18798 7098
rect 18850 7046 18862 7098
rect 18914 7046 18920 7098
rect 184 7024 18920 7046
rect 11882 6984 11888 6996
rect 11843 6956 11888 6984
rect 11882 6944 11888 6956
rect 11940 6944 11946 6996
rect 15194 6944 15200 6996
rect 15252 6984 15258 6996
rect 15381 6987 15439 6993
rect 15381 6984 15393 6987
rect 15252 6956 15393 6984
rect 15252 6944 15258 6956
rect 15381 6953 15393 6956
rect 15427 6953 15439 6987
rect 15381 6947 15439 6953
rect 566 6876 572 6928
rect 624 6916 630 6928
rect 4246 6916 4252 6928
rect 624 6888 4252 6916
rect 624 6876 630 6888
rect 2056 6857 2084 6888
rect 4246 6876 4252 6888
rect 4304 6876 4310 6928
rect 11422 6876 11428 6928
rect 11480 6876 11486 6928
rect 13814 6916 13820 6928
rect 12544 6888 13820 6916
rect 2041 6851 2099 6857
rect 2041 6817 2053 6851
rect 2087 6848 2099 6851
rect 2087 6820 2121 6848
rect 2087 6817 2099 6820
rect 2041 6811 2099 6817
rect 4154 6808 4160 6860
rect 4212 6848 4218 6860
rect 5169 6851 5227 6857
rect 5169 6848 5181 6851
rect 4212 6820 5181 6848
rect 4212 6808 4218 6820
rect 5169 6817 5181 6820
rect 5215 6817 5227 6851
rect 5169 6811 5227 6817
rect 5258 6808 5264 6860
rect 5316 6848 5322 6860
rect 5721 6851 5779 6857
rect 5316 6820 5361 6848
rect 5316 6808 5322 6820
rect 5721 6817 5733 6851
rect 5767 6848 5779 6851
rect 5810 6848 5816 6860
rect 5767 6820 5816 6848
rect 5767 6817 5779 6820
rect 5721 6811 5779 6817
rect 5810 6808 5816 6820
rect 5868 6808 5874 6860
rect 10134 6848 10140 6860
rect 10095 6820 10140 6848
rect 10134 6808 10140 6820
rect 10192 6808 10198 6860
rect 12544 6857 12572 6888
rect 13814 6876 13820 6888
rect 13872 6876 13878 6928
rect 15930 6916 15936 6928
rect 15212 6888 15936 6916
rect 12529 6851 12587 6857
rect 12529 6848 12541 6851
rect 12406 6820 12541 6848
rect 10152 6780 10180 6808
rect 12406 6780 12434 6820
rect 12529 6817 12541 6820
rect 12575 6817 12587 6851
rect 12529 6811 12587 6817
rect 12796 6851 12854 6857
rect 12796 6817 12808 6851
rect 12842 6848 12854 6851
rect 13538 6848 13544 6860
rect 12842 6820 13544 6848
rect 12842 6817 12854 6820
rect 12796 6811 12854 6817
rect 13538 6808 13544 6820
rect 13596 6808 13602 6860
rect 14921 6851 14979 6857
rect 14921 6848 14933 6851
rect 13924 6820 14933 6848
rect 10152 6752 12434 6780
rect 5537 6715 5595 6721
rect 5537 6681 5549 6715
rect 5583 6712 5595 6715
rect 5718 6712 5724 6724
rect 5583 6684 5724 6712
rect 5583 6681 5595 6684
rect 5537 6675 5595 6681
rect 5718 6672 5724 6684
rect 5776 6672 5782 6724
rect 13924 6721 13952 6820
rect 14921 6817 14933 6820
rect 14967 6848 14979 6851
rect 15212 6848 15240 6888
rect 15930 6876 15936 6888
rect 15988 6876 15994 6928
rect 14967 6820 15240 6848
rect 15657 6851 15715 6857
rect 14967 6817 14979 6820
rect 14921 6811 14979 6817
rect 15657 6817 15669 6851
rect 15703 6848 15715 6851
rect 16022 6848 16028 6860
rect 15703 6820 16028 6848
rect 15703 6817 15715 6820
rect 15657 6811 15715 6817
rect 16022 6808 16028 6820
rect 16080 6808 16086 6860
rect 17957 6851 18015 6857
rect 17957 6817 17969 6851
rect 18003 6848 18015 6851
rect 18414 6848 18420 6860
rect 18003 6820 18420 6848
rect 18003 6817 18015 6820
rect 17957 6811 18015 6817
rect 18414 6808 18420 6820
rect 18472 6808 18478 6860
rect 14550 6780 14556 6792
rect 14200 6752 14556 6780
rect 13909 6715 13967 6721
rect 13909 6681 13921 6715
rect 13955 6681 13967 6715
rect 13909 6675 13967 6681
rect 1946 6644 1952 6656
rect 1907 6616 1952 6644
rect 1946 6604 1952 6616
rect 2004 6604 2010 6656
rect 5626 6644 5632 6656
rect 5587 6616 5632 6644
rect 5626 6604 5632 6616
rect 5684 6604 5690 6656
rect 10400 6647 10458 6653
rect 10400 6613 10412 6647
rect 10446 6644 10458 6647
rect 11146 6644 11152 6656
rect 10446 6616 11152 6644
rect 10446 6613 10458 6616
rect 10400 6607 10458 6613
rect 11146 6604 11152 6616
rect 11204 6604 11210 6656
rect 13538 6604 13544 6656
rect 13596 6644 13602 6656
rect 14200 6653 14228 6752
rect 14550 6740 14556 6752
rect 14608 6780 14614 6792
rect 14737 6783 14795 6789
rect 14737 6780 14749 6783
rect 14608 6752 14749 6780
rect 14608 6740 14614 6752
rect 14737 6749 14749 6752
rect 14783 6780 14795 6783
rect 15010 6780 15016 6792
rect 14783 6752 15016 6780
rect 14783 6749 14795 6752
rect 14737 6743 14795 6749
rect 15010 6740 15016 6752
rect 15068 6740 15074 6792
rect 15378 6780 15384 6792
rect 15339 6752 15384 6780
rect 15378 6740 15384 6752
rect 15436 6740 15442 6792
rect 15105 6715 15163 6721
rect 15105 6681 15117 6715
rect 15151 6712 15163 6715
rect 15565 6715 15623 6721
rect 15565 6712 15577 6715
rect 15151 6684 15577 6712
rect 15151 6681 15163 6684
rect 15105 6675 15163 6681
rect 15565 6681 15577 6684
rect 15611 6681 15623 6715
rect 15565 6675 15623 6681
rect 14185 6647 14243 6653
rect 14185 6644 14197 6647
rect 13596 6616 14197 6644
rect 13596 6604 13602 6616
rect 14185 6613 14197 6616
rect 14231 6613 14243 6647
rect 14185 6607 14243 6613
rect 15286 6604 15292 6656
rect 15344 6644 15350 6656
rect 18233 6647 18291 6653
rect 18233 6644 18245 6647
rect 15344 6616 18245 6644
rect 15344 6604 15350 6616
rect 18233 6613 18245 6616
rect 18279 6613 18291 6647
rect 18233 6607 18291 6613
rect 184 6554 18860 6576
rect 184 6502 1556 6554
rect 1608 6502 1620 6554
rect 1672 6502 1684 6554
rect 1736 6502 1748 6554
rect 1800 6502 1812 6554
rect 1864 6502 4656 6554
rect 4708 6502 4720 6554
rect 4772 6502 4784 6554
rect 4836 6502 4848 6554
rect 4900 6502 4912 6554
rect 4964 6502 7756 6554
rect 7808 6502 7820 6554
rect 7872 6502 7884 6554
rect 7936 6502 7948 6554
rect 8000 6502 8012 6554
rect 8064 6502 10856 6554
rect 10908 6502 10920 6554
rect 10972 6502 10984 6554
rect 11036 6502 11048 6554
rect 11100 6502 11112 6554
rect 11164 6502 13956 6554
rect 14008 6502 14020 6554
rect 14072 6502 14084 6554
rect 14136 6502 14148 6554
rect 14200 6502 14212 6554
rect 14264 6502 17056 6554
rect 17108 6502 17120 6554
rect 17172 6502 17184 6554
rect 17236 6502 17248 6554
rect 17300 6502 17312 6554
rect 17364 6502 18860 6554
rect 184 6480 18860 6502
rect 1946 6440 1952 6452
rect 1596 6412 1952 6440
rect 1596 6313 1624 6412
rect 1946 6400 1952 6412
rect 2004 6400 2010 6452
rect 9030 6400 9036 6452
rect 9088 6440 9094 6452
rect 12621 6443 12679 6449
rect 9088 6412 12434 6440
rect 9088 6400 9094 6412
rect 12406 6372 12434 6412
rect 12621 6409 12633 6443
rect 12667 6440 12679 6443
rect 12802 6440 12808 6452
rect 12667 6412 12808 6440
rect 12667 6409 12679 6412
rect 12621 6403 12679 6409
rect 12802 6400 12808 6412
rect 12860 6400 12866 6452
rect 13633 6443 13691 6449
rect 13633 6409 13645 6443
rect 13679 6440 13691 6443
rect 13722 6440 13728 6452
rect 13679 6412 13728 6440
rect 13679 6409 13691 6412
rect 13633 6403 13691 6409
rect 13722 6400 13728 6412
rect 13780 6400 13786 6452
rect 14550 6440 14556 6452
rect 14511 6412 14556 6440
rect 14550 6400 14556 6412
rect 14608 6400 14614 6452
rect 16850 6440 16856 6452
rect 15856 6412 16856 6440
rect 15286 6372 15292 6384
rect 12406 6344 15292 6372
rect 15286 6332 15292 6344
rect 15344 6332 15350 6384
rect 1581 6307 1639 6313
rect 1581 6273 1593 6307
rect 1627 6273 1639 6307
rect 1581 6267 1639 6273
rect 1949 6307 2007 6313
rect 1949 6273 1961 6307
rect 1995 6304 2007 6307
rect 2958 6304 2964 6316
rect 1995 6276 2964 6304
rect 1995 6273 2007 6276
rect 1949 6267 2007 6273
rect 2958 6264 2964 6276
rect 3016 6264 3022 6316
rect 4246 6304 4252 6316
rect 4159 6276 4252 6304
rect 4246 6264 4252 6276
rect 4304 6304 4310 6316
rect 5534 6304 5540 6316
rect 4304 6276 5540 6304
rect 4304 6264 4310 6276
rect 5534 6264 5540 6276
rect 5592 6304 5598 6316
rect 6365 6307 6423 6313
rect 6365 6304 6377 6307
rect 5592 6276 6377 6304
rect 5592 6264 5598 6276
rect 6365 6273 6377 6276
rect 6411 6304 6423 6307
rect 12989 6307 13047 6313
rect 6411 6276 8800 6304
rect 6411 6273 6423 6276
rect 6365 6267 6423 6273
rect 8772 6248 8800 6276
rect 12989 6273 13001 6307
rect 13035 6304 13047 6307
rect 15856 6304 15884 6412
rect 16850 6400 16856 6412
rect 16908 6400 16914 6452
rect 13035 6276 15884 6304
rect 15933 6307 15991 6313
rect 13035 6273 13047 6276
rect 12989 6267 13047 6273
rect 15933 6273 15945 6307
rect 15979 6304 15991 6307
rect 16206 6304 16212 6316
rect 15979 6276 16212 6304
rect 15979 6273 15991 6276
rect 15933 6267 15991 6273
rect 16206 6264 16212 6276
rect 16264 6264 16270 6316
rect 6730 6236 6736 6248
rect 6691 6208 6736 6236
rect 6730 6196 6736 6208
rect 6788 6196 6794 6248
rect 8754 6236 8760 6248
rect 8715 6208 8760 6236
rect 8754 6196 8760 6208
rect 8812 6196 8818 6248
rect 12897 6239 12955 6245
rect 12897 6205 12909 6239
rect 12943 6236 12955 6239
rect 13722 6236 13728 6248
rect 12943 6208 13728 6236
rect 12943 6205 12955 6208
rect 12897 6199 12955 6205
rect 13722 6196 13728 6208
rect 13780 6236 13786 6248
rect 14734 6236 14740 6248
rect 13780 6208 14740 6236
rect 13780 6196 13786 6208
rect 14734 6196 14740 6208
rect 14792 6196 14798 6248
rect 16298 6236 16304 6248
rect 16259 6208 16304 6236
rect 16298 6196 16304 6208
rect 16356 6196 16362 6248
rect 2866 6128 2872 6180
rect 2924 6128 2930 6180
rect 3421 6171 3479 6177
rect 3421 6137 3433 6171
rect 3467 6168 3479 6171
rect 3510 6168 3516 6180
rect 3467 6140 3516 6168
rect 3467 6137 3479 6140
rect 3421 6131 3479 6137
rect 3510 6128 3516 6140
rect 3568 6128 3574 6180
rect 4522 6168 4528 6180
rect 4483 6140 4528 6168
rect 4522 6128 4528 6140
rect 4580 6128 4586 6180
rect 5902 6168 5908 6180
rect 5750 6140 5908 6168
rect 5902 6128 5908 6140
rect 5960 6128 5966 6180
rect 7282 6128 7288 6180
rect 7340 6128 7346 6180
rect 8110 6128 8116 6180
rect 8168 6168 8174 6180
rect 8205 6171 8263 6177
rect 8205 6168 8217 6171
rect 8168 6140 8217 6168
rect 8168 6128 8174 6140
rect 8205 6137 8217 6140
rect 8251 6137 8263 6171
rect 8205 6131 8263 6137
rect 8938 6128 8944 6180
rect 8996 6168 9002 6180
rect 9033 6171 9091 6177
rect 9033 6168 9045 6171
rect 8996 6140 9045 6168
rect 8996 6128 9002 6140
rect 9033 6137 9045 6140
rect 9079 6137 9091 6171
rect 9033 6131 9091 6137
rect 9122 6128 9128 6180
rect 9180 6168 9186 6180
rect 10778 6168 10784 6180
rect 9180 6140 9522 6168
rect 10739 6140 10784 6168
rect 9180 6128 9186 6140
rect 4798 6060 4804 6112
rect 4856 6100 4862 6112
rect 5997 6103 6055 6109
rect 5997 6100 6009 6103
rect 4856 6072 6009 6100
rect 4856 6060 4862 6072
rect 5997 6069 6009 6072
rect 6043 6069 6055 6103
rect 9416 6100 9444 6140
rect 10778 6128 10784 6140
rect 10836 6128 10842 6180
rect 16666 6128 16672 6180
rect 16724 6128 16730 6180
rect 17770 6168 17776 6180
rect 17731 6140 17776 6168
rect 17770 6128 17776 6140
rect 17828 6128 17834 6180
rect 9674 6100 9680 6112
rect 9416 6072 9680 6100
rect 5997 6063 6055 6069
rect 9674 6060 9680 6072
rect 9732 6060 9738 6112
rect 184 6010 18920 6032
rect 184 5958 3106 6010
rect 3158 5958 3170 6010
rect 3222 5958 3234 6010
rect 3286 5958 3298 6010
rect 3350 5958 3362 6010
rect 3414 5958 6206 6010
rect 6258 5958 6270 6010
rect 6322 5958 6334 6010
rect 6386 5958 6398 6010
rect 6450 5958 6462 6010
rect 6514 5958 9306 6010
rect 9358 5958 9370 6010
rect 9422 5958 9434 6010
rect 9486 5958 9498 6010
rect 9550 5958 9562 6010
rect 9614 5958 12406 6010
rect 12458 5958 12470 6010
rect 12522 5958 12534 6010
rect 12586 5958 12598 6010
rect 12650 5958 12662 6010
rect 12714 5958 15506 6010
rect 15558 5958 15570 6010
rect 15622 5958 15634 6010
rect 15686 5958 15698 6010
rect 15750 5958 15762 6010
rect 15814 5958 18606 6010
rect 18658 5958 18670 6010
rect 18722 5958 18734 6010
rect 18786 5958 18798 6010
rect 18850 5958 18862 6010
rect 18914 5958 18920 6010
rect 184 5936 18920 5958
rect 2314 5896 2320 5908
rect 2227 5868 2320 5896
rect 2314 5856 2320 5868
rect 2372 5896 2378 5908
rect 5169 5899 5227 5905
rect 2372 5868 4108 5896
rect 2372 5856 2378 5868
rect 2866 5828 2872 5840
rect 2070 5800 2872 5828
rect 2866 5788 2872 5800
rect 2924 5788 2930 5840
rect 4080 5828 4108 5868
rect 5169 5865 5181 5899
rect 5215 5896 5227 5899
rect 5258 5896 5264 5908
rect 5215 5868 5264 5896
rect 5215 5865 5227 5868
rect 5169 5859 5227 5865
rect 5258 5856 5264 5868
rect 5316 5856 5322 5908
rect 5902 5856 5908 5908
rect 5960 5896 5966 5908
rect 6273 5899 6331 5905
rect 6273 5896 6285 5899
rect 5960 5868 6285 5896
rect 5960 5856 5966 5868
rect 6273 5865 6285 5868
rect 6319 5896 6331 5899
rect 7282 5896 7288 5908
rect 6319 5868 7288 5896
rect 6319 5865 6331 5868
rect 6273 5859 6331 5865
rect 7282 5856 7288 5868
rect 7340 5896 7346 5908
rect 8573 5899 8631 5905
rect 8573 5896 8585 5899
rect 7340 5868 8585 5896
rect 7340 5856 7346 5868
rect 8573 5865 8585 5868
rect 8619 5896 8631 5899
rect 8941 5899 8999 5905
rect 8941 5896 8953 5899
rect 8619 5868 8953 5896
rect 8619 5865 8631 5868
rect 8573 5859 8631 5865
rect 8941 5865 8953 5868
rect 8987 5896 8999 5899
rect 9122 5896 9128 5908
rect 8987 5868 9128 5896
rect 8987 5865 8999 5868
rect 8941 5859 8999 5865
rect 9122 5856 9128 5868
rect 9180 5856 9186 5908
rect 13538 5856 13544 5908
rect 13596 5896 13602 5908
rect 13814 5896 13820 5908
rect 13596 5868 13820 5896
rect 13596 5856 13602 5868
rect 13814 5856 13820 5868
rect 13872 5896 13878 5908
rect 16206 5896 16212 5908
rect 13872 5868 16212 5896
rect 13872 5856 13878 5868
rect 4080 5800 5396 5828
rect 566 5760 572 5772
rect 527 5732 572 5760
rect 566 5720 572 5732
rect 624 5720 630 5772
rect 3510 5720 3516 5772
rect 3568 5760 3574 5772
rect 4617 5763 4675 5769
rect 4617 5760 4629 5763
rect 3568 5732 4629 5760
rect 3568 5720 3574 5732
rect 4617 5729 4629 5732
rect 4663 5729 4675 5763
rect 4798 5760 4804 5772
rect 4759 5732 4804 5760
rect 4617 5723 4675 5729
rect 4798 5720 4804 5732
rect 4856 5720 4862 5772
rect 5368 5769 5396 5800
rect 5353 5763 5411 5769
rect 5353 5729 5365 5763
rect 5399 5729 5411 5763
rect 5353 5723 5411 5729
rect 5445 5763 5503 5769
rect 5445 5729 5457 5763
rect 5491 5760 5503 5763
rect 5810 5760 5816 5772
rect 5491 5732 5816 5760
rect 5491 5729 5503 5732
rect 5445 5723 5503 5729
rect 5810 5720 5816 5732
rect 5868 5720 5874 5772
rect 8110 5760 8116 5772
rect 8071 5732 8116 5760
rect 8110 5720 8116 5732
rect 8168 5720 8174 5772
rect 8297 5763 8355 5769
rect 8297 5729 8309 5763
rect 8343 5760 8355 5763
rect 8478 5760 8484 5772
rect 8343 5732 8484 5760
rect 8343 5729 8355 5732
rect 8297 5723 8355 5729
rect 8478 5720 8484 5732
rect 8536 5720 8542 5772
rect 15028 5769 15056 5868
rect 16206 5856 16212 5868
rect 16264 5856 16270 5908
rect 17402 5856 17408 5908
rect 17460 5896 17466 5908
rect 17681 5899 17739 5905
rect 17681 5896 17693 5899
rect 17460 5868 17693 5896
rect 17460 5856 17466 5868
rect 17681 5865 17693 5868
rect 17727 5865 17739 5899
rect 17681 5859 17739 5865
rect 16666 5828 16672 5840
rect 16514 5800 16672 5828
rect 16666 5788 16672 5800
rect 16724 5788 16730 5840
rect 15013 5763 15071 5769
rect 15013 5729 15025 5763
rect 15059 5729 15071 5763
rect 15013 5723 15071 5729
rect 16850 5720 16856 5772
rect 16908 5760 16914 5772
rect 17405 5763 17463 5769
rect 17405 5760 17417 5763
rect 16908 5732 17417 5760
rect 16908 5720 16914 5732
rect 17405 5729 17417 5732
rect 17451 5729 17463 5763
rect 17405 5723 17463 5729
rect 17494 5720 17500 5772
rect 17552 5760 17558 5772
rect 17681 5763 17739 5769
rect 17681 5760 17693 5763
rect 17552 5732 17693 5760
rect 17552 5720 17558 5732
rect 17681 5729 17693 5732
rect 17727 5729 17739 5763
rect 17681 5723 17739 5729
rect 845 5695 903 5701
rect 845 5661 857 5695
rect 891 5692 903 5695
rect 934 5692 940 5704
rect 891 5664 940 5692
rect 891 5661 903 5664
rect 845 5655 903 5661
rect 934 5652 940 5664
rect 992 5652 998 5704
rect 4246 5652 4252 5704
rect 4304 5692 4310 5704
rect 4816 5692 4844 5720
rect 4304 5664 4844 5692
rect 5537 5695 5595 5701
rect 4304 5652 4310 5664
rect 5537 5661 5549 5695
rect 5583 5661 5595 5695
rect 5537 5655 5595 5661
rect 5629 5695 5687 5701
rect 5629 5661 5641 5695
rect 5675 5692 5687 5695
rect 5718 5692 5724 5704
rect 5675 5664 5724 5692
rect 5675 5661 5687 5664
rect 5629 5655 5687 5661
rect 4801 5627 4859 5633
rect 4801 5593 4813 5627
rect 4847 5624 4859 5627
rect 5552 5624 5580 5655
rect 5718 5652 5724 5664
rect 5776 5652 5782 5704
rect 15289 5695 15347 5701
rect 15289 5661 15301 5695
rect 15335 5692 15347 5695
rect 16942 5692 16948 5704
rect 15335 5664 16948 5692
rect 15335 5661 15347 5664
rect 15289 5655 15347 5661
rect 16942 5652 16948 5664
rect 17000 5652 17006 5704
rect 8294 5624 8300 5636
rect 4847 5596 5580 5624
rect 8255 5596 8300 5624
rect 4847 5593 4859 5596
rect 4801 5587 4859 5593
rect 8294 5584 8300 5596
rect 8352 5584 8358 5636
rect 16761 5627 16819 5633
rect 16761 5593 16773 5627
rect 16807 5624 16819 5627
rect 17586 5624 17592 5636
rect 16807 5596 17592 5624
rect 16807 5593 16819 5596
rect 16761 5587 16819 5593
rect 17586 5584 17592 5596
rect 17644 5584 17650 5636
rect 2866 5556 2872 5568
rect 2779 5528 2872 5556
rect 2866 5516 2872 5528
rect 2924 5556 2930 5568
rect 3605 5559 3663 5565
rect 3605 5556 3617 5559
rect 2924 5528 3617 5556
rect 2924 5516 2930 5528
rect 3605 5525 3617 5528
rect 3651 5556 3663 5559
rect 4157 5559 4215 5565
rect 4157 5556 4169 5559
rect 3651 5528 4169 5556
rect 3651 5525 3663 5528
rect 3605 5519 3663 5525
rect 4157 5525 4169 5528
rect 4203 5556 4215 5559
rect 5902 5556 5908 5568
rect 4203 5528 5908 5556
rect 4203 5525 4215 5528
rect 4157 5519 4215 5525
rect 5902 5516 5908 5528
rect 5960 5516 5966 5568
rect 184 5466 18860 5488
rect 184 5414 1556 5466
rect 1608 5414 1620 5466
rect 1672 5414 1684 5466
rect 1736 5414 1748 5466
rect 1800 5414 1812 5466
rect 1864 5414 4656 5466
rect 4708 5414 4720 5466
rect 4772 5414 4784 5466
rect 4836 5414 4848 5466
rect 4900 5414 4912 5466
rect 4964 5414 7756 5466
rect 7808 5414 7820 5466
rect 7872 5414 7884 5466
rect 7936 5414 7948 5466
rect 8000 5414 8012 5466
rect 8064 5414 10856 5466
rect 10908 5414 10920 5466
rect 10972 5414 10984 5466
rect 11036 5414 11048 5466
rect 11100 5414 11112 5466
rect 11164 5414 13956 5466
rect 14008 5414 14020 5466
rect 14072 5414 14084 5466
rect 14136 5414 14148 5466
rect 14200 5414 14212 5466
rect 14264 5414 17056 5466
rect 17108 5414 17120 5466
rect 17172 5414 17184 5466
rect 17236 5414 17248 5466
rect 17300 5414 17312 5466
rect 17364 5414 18860 5466
rect 184 5392 18860 5414
rect 1673 5355 1731 5361
rect 1673 5321 1685 5355
rect 1719 5352 1731 5355
rect 2130 5352 2136 5364
rect 1719 5324 2136 5352
rect 1719 5321 1731 5324
rect 1673 5315 1731 5321
rect 2130 5312 2136 5324
rect 2188 5312 2194 5364
rect 6549 5355 6607 5361
rect 6549 5321 6561 5355
rect 6595 5352 6607 5355
rect 6730 5352 6736 5364
rect 6595 5324 6736 5352
rect 6595 5321 6607 5324
rect 6549 5315 6607 5321
rect 6730 5312 6736 5324
rect 6788 5312 6794 5364
rect 7466 5312 7472 5364
rect 7524 5352 7530 5364
rect 8662 5352 8668 5364
rect 7524 5324 8668 5352
rect 7524 5312 7530 5324
rect 8662 5312 8668 5324
rect 8720 5312 8726 5364
rect 7558 5284 7564 5296
rect 6748 5256 7564 5284
rect 1946 5176 1952 5228
rect 2004 5216 2010 5228
rect 2225 5219 2283 5225
rect 2225 5216 2237 5219
rect 2004 5188 2237 5216
rect 2004 5176 2010 5188
rect 2225 5185 2237 5188
rect 2271 5185 2283 5219
rect 2225 5179 2283 5185
rect 5718 5108 5724 5160
rect 5776 5148 5782 5160
rect 6748 5157 6776 5256
rect 7558 5244 7564 5256
rect 7616 5284 7622 5296
rect 7653 5287 7711 5293
rect 7653 5284 7665 5287
rect 7616 5256 7665 5284
rect 7616 5244 7622 5256
rect 7653 5253 7665 5256
rect 7699 5253 7711 5287
rect 7653 5247 7711 5253
rect 8113 5219 8171 5225
rect 8113 5216 8125 5219
rect 6840 5188 8125 5216
rect 6840 5157 6868 5188
rect 8113 5185 8125 5188
rect 8159 5185 8171 5219
rect 8754 5216 8760 5228
rect 8715 5188 8760 5216
rect 8113 5179 8171 5185
rect 8754 5176 8760 5188
rect 8812 5176 8818 5228
rect 13081 5219 13139 5225
rect 13081 5185 13093 5219
rect 13127 5216 13139 5219
rect 13538 5216 13544 5228
rect 13127 5188 13544 5216
rect 13127 5185 13139 5188
rect 13081 5179 13139 5185
rect 13538 5176 13544 5188
rect 13596 5176 13602 5228
rect 14826 5176 14832 5228
rect 14884 5216 14890 5228
rect 15565 5219 15623 5225
rect 15565 5216 15577 5219
rect 14884 5188 15577 5216
rect 14884 5176 14890 5188
rect 15565 5185 15577 5188
rect 15611 5185 15623 5219
rect 15565 5179 15623 5185
rect 15933 5219 15991 5225
rect 15933 5185 15945 5219
rect 15979 5216 15991 5219
rect 16206 5216 16212 5228
rect 15979 5188 16212 5216
rect 15979 5185 15991 5188
rect 15933 5179 15991 5185
rect 16206 5176 16212 5188
rect 16264 5176 16270 5228
rect 6733 5151 6791 5157
rect 6733 5148 6745 5151
rect 5776 5120 6745 5148
rect 5776 5108 5782 5120
rect 6733 5117 6745 5120
rect 6779 5117 6791 5151
rect 6733 5111 6791 5117
rect 6825 5151 6883 5157
rect 6825 5117 6837 5151
rect 6871 5117 6883 5151
rect 7190 5148 7196 5160
rect 6825 5111 6883 5117
rect 6932 5120 7196 5148
rect 2041 5083 2099 5089
rect 2041 5049 2053 5083
rect 2087 5080 2099 5083
rect 6932 5080 6960 5120
rect 7190 5108 7196 5120
rect 7248 5108 7254 5160
rect 7466 5148 7472 5160
rect 7427 5120 7472 5148
rect 7466 5108 7472 5120
rect 7524 5108 7530 5160
rect 7650 5108 7656 5160
rect 7708 5148 7714 5160
rect 7834 5148 7840 5160
rect 7708 5120 7840 5148
rect 7708 5108 7714 5120
rect 7834 5108 7840 5120
rect 7892 5148 7898 5160
rect 8021 5151 8079 5157
rect 8021 5148 8033 5151
rect 7892 5120 8033 5148
rect 7892 5108 7898 5120
rect 8021 5117 8033 5120
rect 8067 5117 8079 5151
rect 8021 5111 8079 5117
rect 8205 5151 8263 5157
rect 8205 5117 8217 5151
rect 8251 5117 8263 5151
rect 8205 5111 8263 5117
rect 12713 5151 12771 5157
rect 12713 5117 12725 5151
rect 12759 5148 12771 5151
rect 12802 5148 12808 5160
rect 12759 5120 12808 5148
rect 12759 5117 12771 5120
rect 12713 5111 12771 5117
rect 7098 5080 7104 5092
rect 2087 5052 6960 5080
rect 7059 5052 7104 5080
rect 2087 5049 2099 5052
rect 2041 5043 2099 5049
rect 7098 5040 7104 5052
rect 7156 5040 7162 5092
rect 7742 5040 7748 5092
rect 7800 5080 7806 5092
rect 8110 5080 8116 5092
rect 7800 5052 8116 5080
rect 7800 5040 7806 5052
rect 8110 5040 8116 5052
rect 8168 5080 8174 5092
rect 8220 5080 8248 5111
rect 12802 5108 12808 5120
rect 12860 5108 12866 5160
rect 8168 5052 8248 5080
rect 8168 5040 8174 5052
rect 8754 5040 8760 5092
rect 8812 5080 8818 5092
rect 9033 5083 9091 5089
rect 9033 5080 9045 5083
rect 8812 5052 9045 5080
rect 8812 5040 8818 5052
rect 9033 5049 9045 5052
rect 9079 5049 9091 5083
rect 9033 5043 9091 5049
rect 9674 5040 9680 5092
rect 9732 5040 9738 5092
rect 13814 5080 13820 5092
rect 12374 5052 12480 5080
rect 13775 5052 13820 5080
rect 2130 5012 2136 5024
rect 2091 4984 2136 5012
rect 2130 4972 2136 4984
rect 2188 4972 2194 5024
rect 9766 4972 9772 5024
rect 9824 5012 9830 5024
rect 10505 5015 10563 5021
rect 10505 5012 10517 5015
rect 9824 4984 10517 5012
rect 9824 4972 9830 4984
rect 10505 4981 10517 4984
rect 10551 4981 10563 5015
rect 10505 4975 10563 4981
rect 11287 5015 11345 5021
rect 11287 4981 11299 5015
rect 11333 5012 11345 5015
rect 11882 5012 11888 5024
rect 11333 4984 11888 5012
rect 11333 4981 11345 4984
rect 11287 4975 11345 4981
rect 11882 4972 11888 4984
rect 11940 4972 11946 5024
rect 12250 4972 12256 5024
rect 12308 5012 12314 5024
rect 12452 5012 12480 5052
rect 13814 5040 13820 5052
rect 13872 5040 13878 5092
rect 16206 5080 16212 5092
rect 13924 5052 14306 5080
rect 16167 5052 16212 5080
rect 13924 5012 13952 5052
rect 16206 5040 16212 5052
rect 16264 5040 16270 5092
rect 16666 5040 16672 5092
rect 16724 5040 16730 5092
rect 12308 4984 13952 5012
rect 12308 4972 12314 4984
rect 17494 4972 17500 5024
rect 17552 5012 17558 5024
rect 17681 5015 17739 5021
rect 17681 5012 17693 5015
rect 17552 4984 17693 5012
rect 17552 4972 17558 4984
rect 17681 4981 17693 4984
rect 17727 4981 17739 5015
rect 17681 4975 17739 4981
rect 184 4922 18920 4944
rect 184 4870 3106 4922
rect 3158 4870 3170 4922
rect 3222 4870 3234 4922
rect 3286 4870 3298 4922
rect 3350 4870 3362 4922
rect 3414 4870 6206 4922
rect 6258 4870 6270 4922
rect 6322 4870 6334 4922
rect 6386 4870 6398 4922
rect 6450 4870 6462 4922
rect 6514 4870 9306 4922
rect 9358 4870 9370 4922
rect 9422 4870 9434 4922
rect 9486 4870 9498 4922
rect 9550 4870 9562 4922
rect 9614 4870 12406 4922
rect 12458 4870 12470 4922
rect 12522 4870 12534 4922
rect 12586 4870 12598 4922
rect 12650 4870 12662 4922
rect 12714 4870 15506 4922
rect 15558 4870 15570 4922
rect 15622 4870 15634 4922
rect 15686 4870 15698 4922
rect 15750 4870 15762 4922
rect 15814 4870 18606 4922
rect 18658 4870 18670 4922
rect 18722 4870 18734 4922
rect 18786 4870 18798 4922
rect 18850 4870 18862 4922
rect 18914 4870 18920 4922
rect 184 4848 18920 4870
rect 1946 4808 1952 4820
rect 1907 4780 1952 4808
rect 1946 4768 1952 4780
rect 2004 4768 2010 4820
rect 2958 4768 2964 4820
rect 3016 4808 3022 4820
rect 3053 4811 3111 4817
rect 3053 4808 3065 4811
rect 3016 4780 3065 4808
rect 3016 4768 3022 4780
rect 3053 4777 3065 4780
rect 3099 4777 3111 4811
rect 3053 4771 3111 4777
rect 3605 4811 3663 4817
rect 3605 4777 3617 4811
rect 3651 4808 3663 4811
rect 4154 4808 4160 4820
rect 3651 4780 4160 4808
rect 3651 4777 3663 4780
rect 3605 4771 3663 4777
rect 2869 4743 2927 4749
rect 2869 4709 2881 4743
rect 2915 4740 2927 4743
rect 3620 4740 3648 4771
rect 4154 4768 4160 4780
rect 4212 4768 4218 4820
rect 4522 4808 4528 4820
rect 4483 4780 4528 4808
rect 4522 4768 4528 4780
rect 4580 4768 4586 4820
rect 7190 4768 7196 4820
rect 7248 4808 7254 4820
rect 7929 4811 7987 4817
rect 7929 4808 7941 4811
rect 7248 4780 7941 4808
rect 7248 4768 7254 4780
rect 7929 4777 7941 4780
rect 7975 4808 7987 4811
rect 8846 4808 8852 4820
rect 7975 4780 8852 4808
rect 7975 4777 7987 4780
rect 7929 4771 7987 4777
rect 8846 4768 8852 4780
rect 8904 4808 8910 4820
rect 12345 4811 12403 4817
rect 8904 4780 9444 4808
rect 8904 4768 8910 4780
rect 9416 4749 9444 4780
rect 12345 4777 12357 4811
rect 12391 4808 12403 4811
rect 12802 4808 12808 4820
rect 12391 4780 12808 4808
rect 12391 4777 12403 4780
rect 12345 4771 12403 4777
rect 12802 4768 12808 4780
rect 12860 4768 12866 4820
rect 13814 4768 13820 4820
rect 13872 4808 13878 4820
rect 14001 4811 14059 4817
rect 14001 4808 14013 4811
rect 13872 4780 14013 4808
rect 13872 4768 13878 4780
rect 14001 4777 14013 4780
rect 14047 4777 14059 4811
rect 14734 4808 14740 4820
rect 14695 4780 14740 4808
rect 14001 4771 14059 4777
rect 14734 4768 14740 4780
rect 14792 4768 14798 4820
rect 15010 4768 15016 4820
rect 15068 4808 15074 4820
rect 15197 4811 15255 4817
rect 15197 4808 15209 4811
rect 15068 4780 15209 4808
rect 15068 4768 15074 4780
rect 15197 4777 15209 4780
rect 15243 4808 15255 4811
rect 15470 4808 15476 4820
rect 15243 4780 15476 4808
rect 15243 4777 15255 4780
rect 15197 4771 15255 4777
rect 15470 4768 15476 4780
rect 15528 4768 15534 4820
rect 2915 4712 3648 4740
rect 8389 4743 8447 4749
rect 2915 4709 2927 4712
rect 2869 4703 2927 4709
rect 8389 4709 8401 4743
rect 8435 4740 8447 4743
rect 9401 4743 9459 4749
rect 8435 4712 9076 4740
rect 8435 4709 8447 4712
rect 8389 4703 8447 4709
rect 1857 4675 1915 4681
rect 1857 4641 1869 4675
rect 1903 4672 1915 4675
rect 1946 4672 1952 4684
rect 1903 4644 1952 4672
rect 1903 4641 1915 4644
rect 1857 4635 1915 4641
rect 1946 4632 1952 4644
rect 2004 4632 2010 4684
rect 2774 4632 2780 4684
rect 2832 4672 2838 4684
rect 3326 4672 3332 4684
rect 2832 4644 2877 4672
rect 3287 4644 3332 4672
rect 2832 4632 2838 4644
rect 3326 4632 3332 4644
rect 3384 4632 3390 4684
rect 3878 4672 3884 4684
rect 3839 4644 3884 4672
rect 3878 4632 3884 4644
rect 3936 4632 3942 4684
rect 3973 4675 4031 4681
rect 3973 4641 3985 4675
rect 4019 4641 4031 4675
rect 3973 4635 4031 4641
rect 4801 4675 4859 4681
rect 4801 4641 4813 4675
rect 4847 4672 4859 4675
rect 5166 4672 5172 4684
rect 4847 4644 5172 4672
rect 4847 4641 4859 4644
rect 4801 4635 4859 4641
rect 3988 4604 4016 4635
rect 5166 4632 5172 4644
rect 5224 4632 5230 4684
rect 7558 4672 7564 4684
rect 7519 4644 7564 4672
rect 7558 4632 7564 4644
rect 7616 4632 7622 4684
rect 7715 4675 7773 4681
rect 7715 4641 7727 4675
rect 7761 4672 7773 4675
rect 7834 4672 7840 4684
rect 7761 4644 7840 4672
rect 7761 4641 7773 4644
rect 7715 4635 7773 4641
rect 7834 4632 7840 4644
rect 7892 4672 7898 4684
rect 8297 4675 8355 4681
rect 8297 4672 8309 4675
rect 7892 4644 8309 4672
rect 7892 4632 7898 4644
rect 8297 4641 8309 4644
rect 8343 4641 8355 4675
rect 8297 4635 8355 4641
rect 8478 4632 8484 4684
rect 8536 4672 8542 4684
rect 8536 4644 8629 4672
rect 8536 4632 8542 4644
rect 8662 4632 8668 4684
rect 8720 4672 8726 4684
rect 9048 4681 9076 4712
rect 9401 4709 9413 4743
rect 9447 4709 9459 4743
rect 12250 4740 12256 4752
rect 11730 4712 12256 4740
rect 9401 4703 9459 4709
rect 12250 4700 12256 4712
rect 12308 4700 12314 4752
rect 13262 4740 13268 4752
rect 12544 4712 13268 4740
rect 8941 4675 8999 4681
rect 8941 4672 8953 4675
rect 8720 4644 8953 4672
rect 8720 4632 8726 4644
rect 8941 4641 8953 4644
rect 8987 4641 8999 4675
rect 8941 4635 8999 4641
rect 9033 4675 9091 4681
rect 9033 4641 9045 4675
rect 9079 4641 9091 4675
rect 9033 4635 9091 4641
rect 9309 4675 9367 4681
rect 9309 4641 9321 4675
rect 9355 4672 9367 4675
rect 9950 4672 9956 4684
rect 9355 4644 9956 4672
rect 9355 4641 9367 4644
rect 9309 4635 9367 4641
rect 9950 4632 9956 4644
rect 10008 4632 10014 4684
rect 10134 4632 10140 4684
rect 10192 4672 10198 4684
rect 12544 4681 12572 4712
rect 13262 4700 13268 4712
rect 13320 4700 13326 4752
rect 14274 4700 14280 4752
rect 14332 4700 14338 4752
rect 10229 4675 10287 4681
rect 10229 4672 10241 4675
rect 10192 4644 10241 4672
rect 10192 4632 10198 4644
rect 10229 4641 10241 4644
rect 10275 4641 10287 4675
rect 10229 4635 10287 4641
rect 12529 4675 12587 4681
rect 12529 4641 12541 4675
rect 12575 4641 12587 4675
rect 12529 4635 12587 4641
rect 12710 4632 12716 4684
rect 12768 4672 12774 4684
rect 12805 4675 12863 4681
rect 12805 4672 12817 4675
rect 12768 4644 12817 4672
rect 12768 4632 12774 4644
rect 12805 4641 12817 4644
rect 12851 4641 12863 4675
rect 13722 4672 13728 4684
rect 13683 4644 13728 4672
rect 12805 4635 12863 4641
rect 13722 4632 13728 4644
rect 13780 4632 13786 4684
rect 13817 4675 13875 4681
rect 13817 4641 13829 4675
rect 13863 4672 13875 4675
rect 14292 4672 14320 4700
rect 13863 4644 14320 4672
rect 13863 4641 13875 4644
rect 13817 4635 13875 4641
rect 4522 4604 4528 4616
rect 3252 4576 4016 4604
rect 4483 4576 4528 4604
rect 2038 4428 2044 4480
rect 2096 4468 2102 4480
rect 3252 4477 3280 4576
rect 3988 4536 4016 4576
rect 4522 4564 4528 4576
rect 4580 4564 4586 4616
rect 5718 4604 5724 4616
rect 5552 4576 5724 4604
rect 5552 4548 5580 4576
rect 5718 4564 5724 4576
rect 5776 4564 5782 4616
rect 7576 4604 7604 4632
rect 8110 4604 8116 4616
rect 7576 4576 8116 4604
rect 8110 4564 8116 4576
rect 8168 4564 8174 4616
rect 4154 4536 4160 4548
rect 3988 4508 4160 4536
rect 4154 4496 4160 4508
rect 4212 4536 4218 4548
rect 5534 4536 5540 4548
rect 4212 4508 5540 4536
rect 4212 4496 4218 4508
rect 5534 4496 5540 4508
rect 5592 4496 5598 4548
rect 8496 4536 8524 4632
rect 10505 4607 10563 4613
rect 10505 4573 10517 4607
rect 10551 4604 10563 4607
rect 11238 4604 11244 4616
rect 10551 4576 11244 4604
rect 10551 4573 10563 4576
rect 10505 4567 10563 4573
rect 11238 4564 11244 4576
rect 11296 4564 11302 4616
rect 11882 4564 11888 4616
rect 11940 4604 11946 4616
rect 12621 4607 12679 4613
rect 12621 4604 12633 4607
rect 11940 4576 12633 4604
rect 11940 4564 11946 4576
rect 12621 4573 12633 4576
rect 12667 4604 12679 4607
rect 13538 4604 13544 4616
rect 12667 4576 13544 4604
rect 12667 4573 12679 4576
rect 12621 4567 12679 4573
rect 13538 4564 13544 4576
rect 13596 4564 13602 4616
rect 14001 4607 14059 4613
rect 14001 4573 14013 4607
rect 14047 4604 14059 4607
rect 14274 4604 14280 4616
rect 14047 4576 14280 4604
rect 14047 4573 14059 4576
rect 14001 4567 14059 4573
rect 14274 4564 14280 4576
rect 14332 4564 14338 4616
rect 9766 4536 9772 4548
rect 8496 4508 9772 4536
rect 9766 4496 9772 4508
rect 9824 4496 9830 4548
rect 11977 4539 12035 4545
rect 11977 4505 11989 4539
rect 12023 4536 12035 4539
rect 12713 4539 12771 4545
rect 12023 4508 12434 4536
rect 12023 4505 12035 4508
rect 11977 4499 12035 4505
rect 12406 4480 12434 4508
rect 12713 4505 12725 4539
rect 12759 4536 12771 4539
rect 14458 4536 14464 4548
rect 12759 4508 14464 4536
rect 12759 4505 12771 4508
rect 12713 4499 12771 4505
rect 14458 4496 14464 4508
rect 14516 4536 14522 4548
rect 15378 4536 15384 4548
rect 14516 4508 15384 4536
rect 14516 4496 14522 4508
rect 15378 4496 15384 4508
rect 15436 4496 15442 4548
rect 3237 4471 3295 4477
rect 3237 4468 3249 4471
rect 2096 4440 3249 4468
rect 2096 4428 2102 4440
rect 3237 4437 3249 4440
rect 3283 4437 3295 4471
rect 3237 4431 3295 4437
rect 4709 4471 4767 4477
rect 4709 4437 4721 4471
rect 4755 4468 4767 4471
rect 5718 4468 5724 4480
rect 4755 4440 5724 4468
rect 4755 4437 4767 4440
rect 4709 4431 4767 4437
rect 5718 4428 5724 4440
rect 5776 4428 5782 4480
rect 8754 4468 8760 4480
rect 8715 4440 8760 4468
rect 8754 4428 8760 4440
rect 8812 4428 8818 4480
rect 12406 4440 12440 4480
rect 12434 4428 12440 4440
rect 12492 4428 12498 4480
rect 184 4378 18860 4400
rect 184 4326 1556 4378
rect 1608 4326 1620 4378
rect 1672 4326 1684 4378
rect 1736 4326 1748 4378
rect 1800 4326 1812 4378
rect 1864 4326 4656 4378
rect 4708 4326 4720 4378
rect 4772 4326 4784 4378
rect 4836 4326 4848 4378
rect 4900 4326 4912 4378
rect 4964 4326 7756 4378
rect 7808 4326 7820 4378
rect 7872 4326 7884 4378
rect 7936 4326 7948 4378
rect 8000 4326 8012 4378
rect 8064 4326 10856 4378
rect 10908 4326 10920 4378
rect 10972 4326 10984 4378
rect 11036 4326 11048 4378
rect 11100 4326 11112 4378
rect 11164 4326 13956 4378
rect 14008 4326 14020 4378
rect 14072 4326 14084 4378
rect 14136 4326 14148 4378
rect 14200 4326 14212 4378
rect 14264 4326 17056 4378
rect 17108 4326 17120 4378
rect 17172 4326 17184 4378
rect 17236 4326 17248 4378
rect 17300 4326 17312 4378
rect 17364 4326 18860 4378
rect 184 4304 18860 4326
rect 845 4267 903 4273
rect 845 4233 857 4267
rect 891 4264 903 4267
rect 891 4236 2774 4264
rect 891 4233 903 4236
rect 845 4227 903 4233
rect 1946 4156 1952 4208
rect 2004 4156 2010 4208
rect 2746 4196 2774 4236
rect 3326 4224 3332 4276
rect 3384 4264 3390 4276
rect 3421 4267 3479 4273
rect 3421 4264 3433 4267
rect 3384 4236 3433 4264
rect 3384 4224 3390 4236
rect 3421 4233 3433 4236
rect 3467 4233 3479 4267
rect 5718 4264 5724 4276
rect 5679 4236 5724 4264
rect 3421 4227 3479 4233
rect 5718 4224 5724 4236
rect 5776 4224 5782 4276
rect 8846 4224 8852 4276
rect 8904 4264 8910 4276
rect 8941 4267 8999 4273
rect 8941 4264 8953 4267
rect 8904 4236 8953 4264
rect 8904 4224 8910 4236
rect 8941 4233 8953 4236
rect 8987 4233 8999 4267
rect 12434 4264 12440 4276
rect 8941 4227 8999 4233
rect 11440 4236 12440 4264
rect 5736 4196 5764 4224
rect 6546 4196 6552 4208
rect 2746 4168 5764 4196
rect 6012 4168 6552 4196
rect 1029 4131 1087 4137
rect 1029 4097 1041 4131
rect 1075 4128 1087 4131
rect 1581 4131 1639 4137
rect 1581 4128 1593 4131
rect 1075 4100 1593 4128
rect 1075 4097 1087 4100
rect 1029 4091 1087 4097
rect 1581 4097 1593 4100
rect 1627 4097 1639 4131
rect 1964 4128 1992 4156
rect 3878 4128 3884 4140
rect 1581 4091 1639 4097
rect 1780 4100 3884 4128
rect 750 4060 756 4072
rect 711 4032 756 4060
rect 750 4020 756 4032
rect 808 4020 814 4072
rect 1780 4069 1808 4100
rect 1765 4063 1823 4069
rect 1765 4029 1777 4063
rect 1811 4029 1823 4063
rect 1765 4023 1823 4029
rect 1857 4063 1915 4069
rect 1857 4029 1869 4063
rect 1903 4029 1915 4063
rect 1857 4023 1915 4029
rect 934 3952 940 4004
rect 992 3992 998 4004
rect 1029 3995 1087 4001
rect 1029 3992 1041 3995
rect 992 3964 1041 3992
rect 992 3952 998 3964
rect 1029 3961 1041 3964
rect 1075 3961 1087 3995
rect 1872 3992 1900 4023
rect 1946 4020 1952 4072
rect 2004 4060 2010 4072
rect 3344 4069 3372 4100
rect 3878 4088 3884 4100
rect 3936 4128 3942 4140
rect 3973 4131 4031 4137
rect 3973 4128 3985 4131
rect 3936 4100 3985 4128
rect 3936 4088 3942 4100
rect 3973 4097 3985 4100
rect 4019 4097 4031 4131
rect 4525 4131 4583 4137
rect 4525 4128 4537 4131
rect 3973 4091 4031 4097
rect 4172 4100 4537 4128
rect 3329 4063 3387 4069
rect 2004 4032 2049 4060
rect 2004 4020 2010 4032
rect 3329 4029 3341 4063
rect 3375 4029 3387 4063
rect 3510 4060 3516 4072
rect 3471 4032 3516 4060
rect 3329 4023 3387 4029
rect 3510 4020 3516 4032
rect 3568 4020 3574 4072
rect 2314 3992 2320 4004
rect 1872 3964 2320 3992
rect 1029 3955 1087 3961
rect 2314 3952 2320 3964
rect 2372 3952 2378 4004
rect 2682 3952 2688 4004
rect 2740 3992 2746 4004
rect 4172 3992 4200 4100
rect 4525 4097 4537 4100
rect 4571 4128 4583 4131
rect 5442 4128 5448 4140
rect 4571 4100 5448 4128
rect 4571 4097 4583 4100
rect 4525 4091 4583 4097
rect 5442 4088 5448 4100
rect 5500 4088 5506 4140
rect 4338 4020 4344 4072
rect 4396 4060 4402 4072
rect 5074 4060 5080 4072
rect 4396 4032 4476 4060
rect 5035 4032 5080 4060
rect 4396 4020 4402 4032
rect 2740 3964 4200 3992
rect 4448 3992 4476 4032
rect 5074 4020 5080 4032
rect 5132 4020 5138 4072
rect 5258 4060 5264 4072
rect 5219 4032 5264 4060
rect 5258 4020 5264 4032
rect 5316 4020 5322 4072
rect 5534 4020 5540 4072
rect 5592 4060 5598 4072
rect 6012 4069 6040 4168
rect 6546 4156 6552 4168
rect 6604 4196 6610 4208
rect 11440 4205 11468 4236
rect 12434 4224 12440 4236
rect 12492 4264 12498 4276
rect 12986 4264 12992 4276
rect 12492 4236 12992 4264
rect 12492 4224 12498 4236
rect 12986 4224 12992 4236
rect 13044 4224 13050 4276
rect 14274 4264 14280 4276
rect 14235 4236 14280 4264
rect 14274 4224 14280 4236
rect 14332 4224 14338 4276
rect 14734 4224 14740 4276
rect 14792 4264 14798 4276
rect 14792 4236 15424 4264
rect 14792 4224 14798 4236
rect 6917 4199 6975 4205
rect 6917 4196 6929 4199
rect 6604 4168 6929 4196
rect 6604 4156 6610 4168
rect 6917 4165 6929 4168
rect 6963 4165 6975 4199
rect 6917 4159 6975 4165
rect 11425 4199 11483 4205
rect 11425 4165 11437 4199
rect 11471 4165 11483 4199
rect 11425 4159 11483 4165
rect 12529 4199 12587 4205
rect 12529 4165 12541 4199
rect 12575 4196 12587 4199
rect 12802 4196 12808 4208
rect 12575 4168 12808 4196
rect 12575 4165 12587 4168
rect 12529 4159 12587 4165
rect 12802 4156 12808 4168
rect 12860 4156 12866 4208
rect 14185 4199 14243 4205
rect 14185 4165 14197 4199
rect 14231 4196 14243 4199
rect 14458 4196 14464 4208
rect 14231 4168 14464 4196
rect 14231 4165 14243 4168
rect 14185 4159 14243 4165
rect 7101 4131 7159 4137
rect 7101 4097 7113 4131
rect 7147 4128 7159 4131
rect 7558 4128 7564 4140
rect 7147 4100 7564 4128
rect 7147 4097 7159 4100
rect 7101 4091 7159 4097
rect 7558 4088 7564 4100
rect 7616 4088 7622 4140
rect 8757 4131 8815 4137
rect 8757 4097 8769 4131
rect 8803 4097 8815 4131
rect 8757 4091 8815 4097
rect 11149 4131 11207 4137
rect 11149 4097 11161 4131
rect 11195 4128 11207 4131
rect 11238 4128 11244 4140
rect 11195 4100 11244 4128
rect 11195 4097 11207 4100
rect 11149 4091 11207 4097
rect 5721 4063 5779 4069
rect 5721 4060 5733 4063
rect 5592 4032 5733 4060
rect 5592 4020 5598 4032
rect 5721 4029 5733 4032
rect 5767 4029 5779 4063
rect 5721 4023 5779 4029
rect 5997 4063 6055 4069
rect 5997 4029 6009 4063
rect 6043 4029 6055 4063
rect 5997 4023 6055 4029
rect 6825 4063 6883 4069
rect 6825 4029 6837 4063
rect 6871 4060 6883 4063
rect 7466 4060 7472 4072
rect 6871 4032 7472 4060
rect 6871 4029 6883 4032
rect 6825 4023 6883 4029
rect 7466 4020 7472 4032
rect 7524 4020 7530 4072
rect 5350 3992 5356 4004
rect 4448 3964 5356 3992
rect 2740 3952 2746 3964
rect 5350 3952 5356 3964
rect 5408 3992 5414 4004
rect 5905 3995 5963 4001
rect 5905 3992 5917 3995
rect 5408 3964 5917 3992
rect 5408 3952 5414 3964
rect 5905 3961 5917 3964
rect 5951 3961 5963 3995
rect 5905 3955 5963 3961
rect 7101 3995 7159 4001
rect 7101 3961 7113 3995
rect 7147 3992 7159 3995
rect 8772 3992 8800 4091
rect 11238 4088 11244 4100
rect 11296 4088 11302 4140
rect 11514 4128 11520 4140
rect 11427 4100 11520 4128
rect 11514 4088 11520 4100
rect 11572 4128 11578 4140
rect 14200 4128 14228 4159
rect 14458 4156 14464 4168
rect 14516 4196 14522 4208
rect 15396 4205 15424 4236
rect 16942 4224 16948 4276
rect 17000 4264 17006 4276
rect 17773 4267 17831 4273
rect 17773 4264 17785 4267
rect 17000 4236 17785 4264
rect 17000 4224 17006 4236
rect 17773 4233 17785 4236
rect 17819 4233 17831 4267
rect 17773 4227 17831 4233
rect 15013 4199 15071 4205
rect 15013 4196 15025 4199
rect 14516 4168 15025 4196
rect 14516 4156 14522 4168
rect 15013 4165 15025 4168
rect 15059 4165 15071 4199
rect 15013 4159 15071 4165
rect 15381 4199 15439 4205
rect 15381 4165 15393 4199
rect 15427 4165 15439 4199
rect 15381 4159 15439 4165
rect 17037 4199 17095 4205
rect 17037 4165 17049 4199
rect 17083 4196 17095 4199
rect 17586 4196 17592 4208
rect 17083 4168 17592 4196
rect 17083 4165 17095 4168
rect 17037 4159 17095 4165
rect 17586 4156 17592 4168
rect 17644 4156 17650 4208
rect 11572 4100 14228 4128
rect 14369 4131 14427 4137
rect 11572 4088 11578 4100
rect 9030 4020 9036 4072
rect 9088 4060 9094 4072
rect 11333 4063 11391 4069
rect 9088 4032 9133 4060
rect 9088 4020 9094 4032
rect 11333 4029 11345 4063
rect 11379 4029 11391 4063
rect 11333 4023 11391 4029
rect 7147 3964 8800 3992
rect 11348 3992 11376 4023
rect 11606 4020 11612 4072
rect 11664 4060 11670 4072
rect 12820 4069 12848 4100
rect 14369 4097 14381 4131
rect 14415 4128 14427 4131
rect 14734 4128 14740 4140
rect 14415 4100 14740 4128
rect 14415 4097 14427 4100
rect 14369 4091 14427 4097
rect 14734 4088 14740 4100
rect 14792 4088 14798 4140
rect 15197 4131 15255 4137
rect 15197 4097 15209 4131
rect 15243 4128 15255 4131
rect 15286 4128 15292 4140
rect 15243 4100 15292 4128
rect 15243 4097 15255 4100
rect 15197 4091 15255 4097
rect 15286 4088 15292 4100
rect 15344 4128 15350 4140
rect 16850 4128 16856 4140
rect 15344 4100 16856 4128
rect 15344 4088 15350 4100
rect 16850 4088 16856 4100
rect 16908 4128 16914 4140
rect 16945 4131 17003 4137
rect 16945 4128 16957 4131
rect 16908 4100 16957 4128
rect 16908 4088 16914 4100
rect 16945 4097 16957 4100
rect 16991 4097 17003 4131
rect 16945 4091 17003 4097
rect 17129 4131 17187 4137
rect 17129 4097 17141 4131
rect 17175 4128 17187 4131
rect 17402 4128 17408 4140
rect 17175 4100 17408 4128
rect 17175 4097 17187 4100
rect 17129 4091 17187 4097
rect 17402 4088 17408 4100
rect 17460 4088 17466 4140
rect 17770 4128 17776 4140
rect 17512 4100 17776 4128
rect 12805 4063 12863 4069
rect 11664 4032 11709 4060
rect 11664 4020 11670 4032
rect 12805 4029 12817 4063
rect 12851 4060 12863 4063
rect 12989 4063 13047 4069
rect 12851 4032 12885 4060
rect 12851 4029 12863 4032
rect 12805 4023 12863 4029
rect 12989 4029 13001 4063
rect 13035 4060 13047 4063
rect 13262 4060 13268 4072
rect 13035 4032 13268 4060
rect 13035 4029 13047 4032
rect 12989 4023 13047 4029
rect 12894 3992 12900 4004
rect 11348 3964 12900 3992
rect 7147 3961 7159 3964
rect 7101 3955 7159 3961
rect 12894 3952 12900 3964
rect 12952 3992 12958 4004
rect 13004 3992 13032 4023
rect 13262 4020 13268 4032
rect 13320 4060 13326 4072
rect 14093 4063 14151 4069
rect 14093 4060 14105 4063
rect 13320 4032 14105 4060
rect 13320 4020 13326 4032
rect 14093 4029 14105 4032
rect 14139 4029 14151 4063
rect 15470 4060 15476 4072
rect 15431 4032 15476 4060
rect 14093 4023 14151 4029
rect 15470 4020 15476 4032
rect 15528 4020 15534 4072
rect 17512 4060 17540 4100
rect 17770 4088 17776 4100
rect 17828 4088 17834 4140
rect 17328 4032 17540 4060
rect 17589 4063 17647 4069
rect 17328 4004 17356 4032
rect 17589 4029 17601 4063
rect 17635 4029 17647 4063
rect 17589 4023 17647 4029
rect 17310 3992 17316 4004
rect 12952 3964 13032 3992
rect 17271 3964 17316 3992
rect 12952 3952 12958 3964
rect 17310 3952 17316 3964
rect 17368 3952 17374 4004
rect 8757 3927 8815 3933
rect 8757 3893 8769 3927
rect 8803 3924 8815 3927
rect 8938 3924 8944 3936
rect 8803 3896 8944 3924
rect 8803 3893 8815 3896
rect 8757 3887 8815 3893
rect 8938 3884 8944 3896
rect 8996 3884 9002 3936
rect 12710 3924 12716 3936
rect 12671 3896 12716 3924
rect 12710 3884 12716 3896
rect 12768 3884 12774 3936
rect 17221 3927 17279 3933
rect 17221 3893 17233 3927
rect 17267 3924 17279 3927
rect 17604 3924 17632 4023
rect 17678 4020 17684 4072
rect 17736 4060 17742 4072
rect 17736 4032 17781 4060
rect 17736 4020 17742 4032
rect 17267 3896 17632 3924
rect 17267 3893 17279 3896
rect 17221 3887 17279 3893
rect 184 3834 18920 3856
rect 184 3782 3106 3834
rect 3158 3782 3170 3834
rect 3222 3782 3234 3834
rect 3286 3782 3298 3834
rect 3350 3782 3362 3834
rect 3414 3782 6206 3834
rect 6258 3782 6270 3834
rect 6322 3782 6334 3834
rect 6386 3782 6398 3834
rect 6450 3782 6462 3834
rect 6514 3782 9306 3834
rect 9358 3782 9370 3834
rect 9422 3782 9434 3834
rect 9486 3782 9498 3834
rect 9550 3782 9562 3834
rect 9614 3782 12406 3834
rect 12458 3782 12470 3834
rect 12522 3782 12534 3834
rect 12586 3782 12598 3834
rect 12650 3782 12662 3834
rect 12714 3782 15506 3834
rect 15558 3782 15570 3834
rect 15622 3782 15634 3834
rect 15686 3782 15698 3834
rect 15750 3782 15762 3834
rect 15814 3782 18606 3834
rect 18658 3782 18670 3834
rect 18722 3782 18734 3834
rect 18786 3782 18798 3834
rect 18850 3782 18862 3834
rect 18914 3782 18920 3834
rect 184 3760 18920 3782
rect 750 3680 756 3732
rect 808 3720 814 3732
rect 845 3723 903 3729
rect 845 3720 857 3723
rect 808 3692 857 3720
rect 808 3680 814 3692
rect 845 3689 857 3692
rect 891 3689 903 3723
rect 845 3683 903 3689
rect 3878 3680 3884 3732
rect 3936 3720 3942 3732
rect 4522 3720 4528 3732
rect 3936 3692 4384 3720
rect 4483 3692 4528 3720
rect 3936 3680 3942 3692
rect 4356 3615 4384 3692
rect 4522 3680 4528 3692
rect 4580 3680 4586 3732
rect 5442 3720 5448 3732
rect 5403 3692 5448 3720
rect 5442 3680 5448 3692
rect 5500 3680 5506 3732
rect 5626 3680 5632 3732
rect 5684 3720 5690 3732
rect 5905 3723 5963 3729
rect 5905 3720 5917 3723
rect 5684 3692 5917 3720
rect 5684 3680 5690 3692
rect 5905 3689 5917 3692
rect 5951 3689 5963 3723
rect 7558 3720 7564 3732
rect 7519 3692 7564 3720
rect 5905 3683 5963 3689
rect 7558 3680 7564 3692
rect 7616 3680 7622 3732
rect 9950 3720 9956 3732
rect 9911 3692 9956 3720
rect 9950 3680 9956 3692
rect 10008 3680 10014 3732
rect 11149 3723 11207 3729
rect 11149 3689 11161 3723
rect 11195 3720 11207 3723
rect 11606 3720 11612 3732
rect 11195 3692 11612 3720
rect 11195 3689 11207 3692
rect 11149 3683 11207 3689
rect 11606 3680 11612 3692
rect 11664 3680 11670 3732
rect 14734 3720 14740 3732
rect 14695 3692 14740 3720
rect 14734 3680 14740 3692
rect 14792 3680 14798 3732
rect 14918 3680 14924 3732
rect 14976 3720 14982 3732
rect 15197 3723 15255 3729
rect 15197 3720 15209 3723
rect 14976 3692 15209 3720
rect 14976 3680 14982 3692
rect 15197 3689 15209 3692
rect 15243 3720 15255 3723
rect 15286 3720 15292 3732
rect 15243 3692 15292 3720
rect 15243 3689 15255 3692
rect 15197 3683 15255 3689
rect 15286 3680 15292 3692
rect 15344 3680 15350 3732
rect 16025 3723 16083 3729
rect 16025 3689 16037 3723
rect 16071 3720 16083 3723
rect 16298 3720 16304 3732
rect 16071 3692 16304 3720
rect 16071 3689 16083 3692
rect 16025 3683 16083 3689
rect 16298 3680 16304 3692
rect 16356 3680 16362 3732
rect 17589 3723 17647 3729
rect 17589 3689 17601 3723
rect 17635 3720 17647 3723
rect 17678 3720 17684 3732
rect 17635 3692 17684 3720
rect 17635 3689 17647 3692
rect 17589 3683 17647 3689
rect 17678 3680 17684 3692
rect 17736 3680 17742 3732
rect 18046 3680 18052 3732
rect 18104 3720 18110 3732
rect 18233 3723 18291 3729
rect 18233 3720 18245 3723
rect 18104 3692 18245 3720
rect 18104 3680 18110 3692
rect 18233 3689 18245 3692
rect 18279 3689 18291 3723
rect 18233 3683 18291 3689
rect 11514 3652 11520 3664
rect 11256 3624 11520 3652
rect 4341 3609 4399 3615
rect 934 3584 940 3596
rect 895 3556 940 3584
rect 934 3544 940 3556
rect 992 3544 998 3596
rect 4136 3584 4142 3596
rect 4097 3556 4142 3584
rect 4136 3544 4142 3556
rect 4194 3544 4200 3596
rect 4249 3587 4307 3593
rect 4249 3553 4261 3587
rect 4295 3553 4307 3587
rect 4341 3575 4353 3609
rect 4387 3575 4399 3609
rect 5534 3584 5540 3596
rect 4341 3569 4399 3575
rect 5495 3556 5540 3584
rect 4249 3547 4307 3553
rect 4264 3516 4292 3547
rect 5534 3544 5540 3556
rect 5592 3544 5598 3596
rect 5629 3587 5687 3593
rect 5629 3553 5641 3587
rect 5675 3553 5687 3587
rect 5629 3547 5687 3553
rect 7929 3587 7987 3593
rect 7929 3553 7941 3587
rect 7975 3584 7987 3587
rect 8202 3584 8208 3596
rect 7975 3556 8208 3584
rect 7975 3553 7987 3556
rect 7929 3547 7987 3553
rect 4338 3516 4344 3528
rect 4264 3488 4344 3516
rect 4338 3476 4344 3488
rect 4396 3476 4402 3528
rect 5169 3519 5227 3525
rect 5169 3485 5181 3519
rect 5215 3516 5227 3519
rect 5258 3516 5264 3528
rect 5215 3488 5264 3516
rect 5215 3485 5227 3488
rect 5169 3479 5227 3485
rect 5184 3448 5212 3479
rect 5258 3476 5264 3488
rect 5316 3476 5322 3528
rect 5350 3476 5356 3528
rect 5408 3516 5414 3528
rect 5644 3516 5672 3547
rect 8202 3544 8208 3556
rect 8260 3544 8266 3596
rect 10226 3544 10232 3596
rect 10284 3584 10290 3596
rect 11256 3593 11284 3624
rect 11514 3612 11520 3624
rect 11572 3612 11578 3664
rect 14369 3655 14427 3661
rect 14369 3621 14381 3655
rect 14415 3652 14427 3655
rect 15010 3652 15016 3664
rect 14415 3624 15016 3652
rect 14415 3621 14427 3624
rect 14369 3615 14427 3621
rect 15010 3612 15016 3624
rect 15068 3612 15074 3664
rect 16485 3655 16543 3661
rect 16485 3621 16497 3655
rect 16531 3652 16543 3655
rect 16574 3652 16580 3664
rect 16531 3624 16580 3652
rect 16531 3621 16543 3624
rect 16485 3615 16543 3621
rect 16574 3612 16580 3624
rect 16632 3612 16638 3664
rect 10321 3587 10379 3593
rect 10321 3584 10333 3587
rect 10284 3556 10333 3584
rect 10284 3544 10290 3556
rect 10321 3553 10333 3556
rect 10367 3553 10379 3587
rect 10321 3547 10379 3553
rect 11241 3587 11299 3593
rect 11241 3553 11253 3587
rect 11287 3553 11299 3587
rect 11241 3547 11299 3553
rect 11425 3587 11483 3593
rect 11425 3553 11437 3587
rect 11471 3584 11483 3587
rect 12434 3584 12440 3596
rect 11471 3556 12440 3584
rect 11471 3553 11483 3556
rect 11425 3547 11483 3553
rect 12434 3544 12440 3556
rect 12492 3584 12498 3596
rect 12894 3584 12900 3596
rect 12492 3556 12900 3584
rect 12492 3544 12498 3556
rect 12894 3544 12900 3556
rect 12952 3544 12958 3596
rect 15105 3587 15163 3593
rect 15105 3553 15117 3587
rect 15151 3584 15163 3587
rect 15378 3584 15384 3596
rect 15151 3556 15384 3584
rect 15151 3553 15163 3556
rect 15105 3547 15163 3553
rect 15378 3544 15384 3556
rect 15436 3544 15442 3596
rect 16393 3587 16451 3593
rect 16393 3553 16405 3587
rect 16439 3584 16451 3587
rect 16850 3584 16856 3596
rect 16439 3556 16856 3584
rect 16439 3553 16451 3556
rect 16393 3547 16451 3553
rect 16850 3544 16856 3556
rect 16908 3544 16914 3596
rect 16942 3544 16948 3596
rect 17000 3584 17006 3596
rect 17129 3587 17187 3593
rect 17129 3584 17141 3587
rect 17000 3556 17141 3584
rect 17000 3544 17006 3556
rect 17129 3553 17141 3556
rect 17175 3553 17187 3587
rect 17586 3584 17592 3596
rect 17547 3556 17592 3584
rect 17129 3547 17187 3553
rect 17586 3544 17592 3556
rect 17644 3544 17650 3596
rect 17957 3587 18015 3593
rect 17957 3553 17969 3587
rect 18003 3584 18015 3587
rect 18417 3587 18475 3593
rect 18417 3584 18429 3587
rect 18003 3556 18429 3584
rect 18003 3553 18015 3556
rect 17957 3547 18015 3553
rect 18417 3553 18429 3556
rect 18463 3584 18475 3587
rect 19058 3584 19064 3596
rect 18463 3556 19064 3584
rect 18463 3553 18475 3556
rect 18417 3547 18475 3553
rect 19058 3544 19064 3556
rect 19116 3544 19122 3596
rect 5408 3488 5672 3516
rect 8021 3519 8079 3525
rect 5408 3476 5414 3488
rect 8021 3485 8033 3519
rect 8067 3485 8079 3519
rect 8021 3479 8079 3485
rect 5184 3420 5396 3448
rect 5074 3340 5080 3392
rect 5132 3380 5138 3392
rect 5258 3380 5264 3392
rect 5132 3352 5264 3380
rect 5132 3340 5138 3352
rect 5258 3340 5264 3352
rect 5316 3340 5322 3392
rect 5368 3380 5396 3420
rect 5442 3408 5448 3460
rect 5500 3448 5506 3460
rect 8036 3448 8064 3479
rect 8110 3476 8116 3528
rect 8168 3516 8174 3528
rect 10410 3516 10416 3528
rect 8168 3488 8213 3516
rect 10371 3488 10416 3516
rect 8168 3476 8174 3488
rect 10410 3476 10416 3488
rect 10468 3476 10474 3528
rect 10505 3519 10563 3525
rect 10505 3485 10517 3519
rect 10551 3485 10563 3519
rect 10505 3479 10563 3485
rect 8386 3448 8392 3460
rect 5500 3420 8392 3448
rect 5500 3408 5506 3420
rect 8386 3408 8392 3420
rect 8444 3408 8450 3460
rect 8662 3408 8668 3460
rect 8720 3448 8726 3460
rect 10520 3448 10548 3479
rect 8720 3420 10548 3448
rect 10965 3451 11023 3457
rect 8720 3408 8726 3420
rect 10965 3417 10977 3451
rect 11011 3448 11023 3451
rect 11330 3448 11336 3460
rect 11011 3420 11336 3448
rect 11011 3417 11023 3420
rect 10965 3411 11023 3417
rect 11330 3408 11336 3420
rect 11388 3408 11394 3460
rect 12912 3448 12940 3544
rect 15289 3519 15347 3525
rect 15289 3485 15301 3519
rect 15335 3485 15347 3519
rect 15289 3479 15347 3485
rect 16669 3519 16727 3525
rect 16669 3485 16681 3519
rect 16715 3516 16727 3519
rect 16960 3516 16988 3544
rect 16715 3488 16988 3516
rect 17267 3519 17325 3525
rect 16715 3485 16727 3488
rect 16669 3479 16727 3485
rect 17267 3485 17279 3519
rect 17313 3516 17325 3519
rect 17402 3516 17408 3528
rect 17313 3488 17408 3516
rect 17313 3485 17325 3488
rect 17267 3479 17325 3485
rect 15304 3448 15332 3479
rect 17402 3476 17408 3488
rect 17460 3476 17466 3528
rect 12912 3420 15332 3448
rect 6730 3380 6736 3392
rect 5368 3352 6736 3380
rect 6730 3340 6736 3352
rect 6788 3340 6794 3392
rect 16574 3340 16580 3392
rect 16632 3380 16638 3392
rect 17310 3380 17316 3392
rect 16632 3352 17316 3380
rect 16632 3340 16638 3352
rect 17310 3340 17316 3352
rect 17368 3380 17374 3392
rect 17405 3383 17463 3389
rect 17405 3380 17417 3383
rect 17368 3352 17417 3380
rect 17368 3340 17374 3352
rect 17405 3349 17417 3352
rect 17451 3349 17463 3383
rect 17405 3343 17463 3349
rect 184 3290 18860 3312
rect 184 3238 1556 3290
rect 1608 3238 1620 3290
rect 1672 3238 1684 3290
rect 1736 3238 1748 3290
rect 1800 3238 1812 3290
rect 1864 3238 4656 3290
rect 4708 3238 4720 3290
rect 4772 3238 4784 3290
rect 4836 3238 4848 3290
rect 4900 3238 4912 3290
rect 4964 3238 7756 3290
rect 7808 3238 7820 3290
rect 7872 3238 7884 3290
rect 7936 3238 7948 3290
rect 8000 3238 8012 3290
rect 8064 3238 10856 3290
rect 10908 3238 10920 3290
rect 10972 3238 10984 3290
rect 11036 3238 11048 3290
rect 11100 3238 11112 3290
rect 11164 3238 13956 3290
rect 14008 3238 14020 3290
rect 14072 3238 14084 3290
rect 14136 3238 14148 3290
rect 14200 3238 14212 3290
rect 14264 3238 17056 3290
rect 17108 3238 17120 3290
rect 17172 3238 17184 3290
rect 17236 3238 17248 3290
rect 17300 3238 17312 3290
rect 17364 3238 18860 3290
rect 184 3216 18860 3238
rect 5166 3176 5172 3188
rect 5127 3148 5172 3176
rect 5166 3136 5172 3148
rect 5224 3136 5230 3188
rect 5258 3136 5264 3188
rect 5316 3176 5322 3188
rect 6914 3176 6920 3188
rect 5316 3148 6920 3176
rect 5316 3136 5322 3148
rect 6914 3136 6920 3148
rect 6972 3136 6978 3188
rect 7009 3179 7067 3185
rect 7009 3145 7021 3179
rect 7055 3176 7067 3179
rect 7098 3176 7104 3188
rect 7055 3148 7104 3176
rect 7055 3145 7067 3148
rect 7009 3139 7067 3145
rect 7098 3136 7104 3148
rect 7156 3136 7162 3188
rect 10226 3176 10232 3188
rect 10187 3148 10232 3176
rect 10226 3136 10232 3148
rect 10284 3136 10290 3188
rect 11241 3179 11299 3185
rect 11241 3145 11253 3179
rect 11287 3176 11299 3179
rect 11330 3176 11336 3188
rect 11287 3148 11336 3176
rect 11287 3145 11299 3148
rect 11241 3139 11299 3145
rect 11330 3136 11336 3148
rect 11388 3136 11394 3188
rect 12437 3179 12495 3185
rect 12437 3145 12449 3179
rect 12483 3176 12495 3179
rect 12802 3176 12808 3188
rect 12483 3148 12808 3176
rect 12483 3145 12495 3148
rect 12437 3139 12495 3145
rect 12802 3136 12808 3148
rect 12860 3136 12866 3188
rect 14093 3179 14151 3185
rect 14093 3145 14105 3179
rect 14139 3176 14151 3179
rect 14182 3176 14188 3188
rect 14139 3148 14188 3176
rect 14139 3145 14151 3148
rect 14093 3139 14151 3145
rect 14108 3108 14136 3139
rect 14182 3136 14188 3148
rect 14240 3176 14246 3188
rect 14642 3176 14648 3188
rect 14240 3148 14648 3176
rect 14240 3136 14246 3148
rect 14642 3136 14648 3148
rect 14700 3136 14706 3188
rect 13556 3080 14136 3108
rect 2409 3043 2467 3049
rect 2409 3009 2421 3043
rect 2455 3040 2467 3043
rect 2866 3040 2872 3052
rect 2455 3012 2872 3040
rect 2455 3009 2467 3012
rect 2409 3003 2467 3009
rect 2866 3000 2872 3012
rect 2924 3000 2930 3052
rect 6822 3000 6828 3052
rect 6880 3040 6886 3052
rect 7466 3040 7472 3052
rect 6880 3012 7472 3040
rect 6880 3000 6886 3012
rect 7466 3000 7472 3012
rect 7524 3040 7530 3052
rect 7561 3043 7619 3049
rect 7561 3040 7573 3043
rect 7524 3012 7573 3040
rect 7524 3000 7530 3012
rect 7561 3009 7573 3012
rect 7607 3009 7619 3043
rect 9674 3040 9680 3052
rect 9635 3012 9680 3040
rect 7561 3003 7619 3009
rect 9674 3000 9680 3012
rect 9732 3000 9738 3052
rect 9769 3043 9827 3049
rect 9769 3009 9781 3043
rect 9815 3040 9827 3043
rect 10410 3040 10416 3052
rect 9815 3012 10416 3040
rect 9815 3009 9827 3012
rect 9769 3003 9827 3009
rect 1486 2932 1492 2984
rect 1544 2972 1550 2984
rect 2225 2975 2283 2981
rect 2225 2972 2237 2975
rect 1544 2944 2237 2972
rect 1544 2932 1550 2944
rect 2225 2941 2237 2944
rect 2271 2972 2283 2975
rect 2682 2972 2688 2984
rect 2271 2944 2688 2972
rect 2271 2941 2283 2944
rect 2225 2935 2283 2941
rect 2682 2932 2688 2944
rect 2740 2932 2746 2984
rect 5258 2972 5264 2984
rect 5219 2944 5264 2972
rect 5258 2932 5264 2944
rect 5316 2932 5322 2984
rect 6730 2932 6736 2984
rect 6788 2972 6794 2984
rect 9784 2972 9812 3003
rect 10410 3000 10416 3012
rect 10468 3000 10474 3052
rect 11885 3043 11943 3049
rect 11885 3009 11897 3043
rect 11931 3040 11943 3043
rect 12434 3040 12440 3052
rect 11931 3012 12440 3040
rect 11931 3009 11943 3012
rect 11885 3003 11943 3009
rect 12434 3000 12440 3012
rect 12492 3040 12498 3052
rect 12989 3043 13047 3049
rect 12989 3040 13001 3043
rect 12492 3012 13001 3040
rect 12492 3000 12498 3012
rect 12989 3009 13001 3012
rect 13035 3009 13047 3043
rect 13556 3040 13584 3080
rect 12989 3003 13047 3009
rect 13372 3012 13584 3040
rect 13633 3043 13691 3049
rect 6788 2944 9812 2972
rect 12897 2975 12955 2981
rect 6788 2932 6794 2944
rect 12897 2941 12909 2975
rect 12943 2972 12955 2975
rect 13372 2972 13400 3012
rect 13633 3009 13645 3043
rect 13679 3040 13691 3043
rect 14660 3040 14688 3136
rect 15194 3108 15200 3120
rect 15155 3080 15200 3108
rect 15194 3068 15200 3080
rect 15252 3068 15258 3120
rect 13679 3012 14504 3040
rect 14660 3012 15148 3040
rect 13679 3009 13691 3012
rect 13633 3003 13691 3009
rect 13538 2972 13544 2984
rect 12943 2944 13400 2972
rect 13499 2944 13544 2972
rect 12943 2941 12955 2944
rect 12897 2935 12955 2941
rect 13538 2932 13544 2944
rect 13596 2932 13602 2984
rect 14476 2981 14504 3012
rect 13725 2975 13783 2981
rect 13725 2941 13737 2975
rect 13771 2941 13783 2975
rect 13725 2935 13783 2941
rect 14461 2975 14519 2981
rect 14461 2941 14473 2975
rect 14507 2941 14519 2975
rect 14461 2935 14519 2941
rect 6914 2864 6920 2916
rect 6972 2904 6978 2916
rect 7466 2904 7472 2916
rect 6972 2876 7472 2904
rect 6972 2864 6978 2876
rect 7466 2864 7472 2876
rect 7524 2864 7530 2916
rect 12986 2864 12992 2916
rect 13044 2904 13050 2916
rect 13740 2904 13768 2935
rect 14642 2932 14648 2984
rect 14700 2972 14706 2984
rect 14737 2975 14795 2981
rect 14737 2972 14749 2975
rect 14700 2944 14749 2972
rect 14700 2932 14706 2944
rect 14737 2941 14749 2944
rect 14783 2972 14795 2975
rect 14826 2972 14832 2984
rect 14783 2944 14832 2972
rect 14783 2941 14795 2944
rect 14737 2935 14795 2941
rect 14826 2932 14832 2944
rect 14884 2932 14890 2984
rect 14918 2932 14924 2984
rect 14976 2972 14982 2984
rect 15120 2981 15148 3012
rect 15105 2975 15163 2981
rect 14976 2944 15021 2972
rect 14976 2932 14982 2944
rect 15105 2941 15117 2975
rect 15151 2941 15163 2975
rect 15105 2935 15163 2941
rect 15381 2975 15439 2981
rect 15381 2941 15393 2975
rect 15427 2941 15439 2975
rect 15381 2935 15439 2941
rect 13044 2876 13768 2904
rect 13044 2864 13050 2876
rect 13814 2864 13820 2916
rect 13872 2904 13878 2916
rect 15010 2904 15016 2916
rect 13872 2876 15016 2904
rect 13872 2864 13878 2876
rect 15010 2864 15016 2876
rect 15068 2904 15074 2916
rect 15396 2904 15424 2935
rect 15838 2904 15844 2916
rect 15068 2876 15844 2904
rect 15068 2864 15074 2876
rect 15838 2864 15844 2876
rect 15896 2864 15902 2916
rect 1762 2836 1768 2848
rect 1723 2808 1768 2836
rect 1762 2796 1768 2808
rect 1820 2796 1826 2848
rect 2130 2836 2136 2848
rect 2091 2808 2136 2836
rect 2130 2796 2136 2808
rect 2188 2796 2194 2848
rect 7374 2836 7380 2848
rect 7335 2808 7380 2836
rect 7374 2796 7380 2808
rect 7432 2796 7438 2848
rect 9858 2796 9864 2848
rect 9916 2836 9922 2848
rect 11606 2836 11612 2848
rect 9916 2808 9961 2836
rect 11567 2808 11612 2836
rect 9916 2796 9922 2808
rect 11606 2796 11612 2808
rect 11664 2796 11670 2848
rect 11701 2839 11759 2845
rect 11701 2805 11713 2839
rect 11747 2836 11759 2839
rect 12250 2836 12256 2848
rect 11747 2808 12256 2836
rect 11747 2805 11759 2808
rect 11701 2799 11759 2805
rect 12250 2796 12256 2808
rect 12308 2796 12314 2848
rect 12802 2836 12808 2848
rect 12763 2808 12808 2836
rect 12802 2796 12808 2808
rect 12860 2796 12866 2848
rect 184 2746 18920 2768
rect 184 2694 3106 2746
rect 3158 2694 3170 2746
rect 3222 2694 3234 2746
rect 3286 2694 3298 2746
rect 3350 2694 3362 2746
rect 3414 2694 6206 2746
rect 6258 2694 6270 2746
rect 6322 2694 6334 2746
rect 6386 2694 6398 2746
rect 6450 2694 6462 2746
rect 6514 2694 9306 2746
rect 9358 2694 9370 2746
rect 9422 2694 9434 2746
rect 9486 2694 9498 2746
rect 9550 2694 9562 2746
rect 9614 2694 12406 2746
rect 12458 2694 12470 2746
rect 12522 2694 12534 2746
rect 12586 2694 12598 2746
rect 12650 2694 12662 2746
rect 12714 2694 15506 2746
rect 15558 2694 15570 2746
rect 15622 2694 15634 2746
rect 15686 2694 15698 2746
rect 15750 2694 15762 2746
rect 15814 2694 18606 2746
rect 18658 2694 18670 2746
rect 18722 2694 18734 2746
rect 18786 2694 18798 2746
rect 18850 2694 18862 2746
rect 18914 2694 18920 2746
rect 184 2672 18920 2694
rect 934 2592 940 2644
rect 992 2632 998 2644
rect 1029 2635 1087 2641
rect 1029 2632 1041 2635
rect 992 2604 1041 2632
rect 992 2592 998 2604
rect 1029 2601 1041 2604
rect 1075 2601 1087 2635
rect 1029 2595 1087 2601
rect 1397 2635 1455 2641
rect 1397 2601 1409 2635
rect 1443 2632 1455 2635
rect 1762 2632 1768 2644
rect 1443 2604 1768 2632
rect 1443 2601 1455 2604
rect 1397 2595 1455 2601
rect 1762 2592 1768 2604
rect 1820 2592 1826 2644
rect 2130 2632 2136 2644
rect 2091 2604 2136 2632
rect 2130 2592 2136 2604
rect 2188 2592 2194 2644
rect 2774 2592 2780 2644
rect 2832 2632 2838 2644
rect 2869 2635 2927 2641
rect 2869 2632 2881 2635
rect 2832 2604 2881 2632
rect 2832 2592 2838 2604
rect 2869 2601 2881 2604
rect 2915 2601 2927 2635
rect 3326 2632 3332 2644
rect 3287 2604 3332 2632
rect 2869 2595 2927 2601
rect 3326 2592 3332 2604
rect 3384 2632 3390 2644
rect 5074 2632 5080 2644
rect 3384 2604 5080 2632
rect 3384 2592 3390 2604
rect 5074 2592 5080 2604
rect 5132 2592 5138 2644
rect 5258 2592 5264 2644
rect 5316 2632 5322 2644
rect 5353 2635 5411 2641
rect 5353 2632 5365 2635
rect 5316 2604 5365 2632
rect 5316 2592 5322 2604
rect 5353 2601 5365 2604
rect 5399 2601 5411 2635
rect 8202 2632 8208 2644
rect 8163 2604 8208 2632
rect 5353 2595 5411 2601
rect 8202 2592 8208 2604
rect 8260 2592 8266 2644
rect 8573 2635 8631 2641
rect 8573 2601 8585 2635
rect 8619 2632 8631 2635
rect 9030 2632 9036 2644
rect 8619 2604 9036 2632
rect 8619 2601 8631 2604
rect 8573 2595 8631 2601
rect 9030 2592 9036 2604
rect 9088 2592 9094 2644
rect 13722 2592 13728 2644
rect 13780 2632 13786 2644
rect 15105 2635 15163 2641
rect 15105 2632 15117 2635
rect 13780 2604 15117 2632
rect 13780 2592 13786 2604
rect 15105 2601 15117 2604
rect 15151 2601 15163 2635
rect 15105 2595 15163 2601
rect 15378 2592 15384 2644
rect 15436 2632 15442 2644
rect 15473 2635 15531 2641
rect 15473 2632 15485 2635
rect 15436 2604 15485 2632
rect 15436 2592 15442 2604
rect 15473 2601 15485 2604
rect 15519 2601 15531 2635
rect 15473 2595 15531 2601
rect 1486 2564 1492 2576
rect 1447 2536 1492 2564
rect 1486 2524 1492 2536
rect 1544 2524 1550 2576
rect 3970 2564 3976 2576
rect 2332 2536 3976 2564
rect 2332 2508 2360 2536
rect 3970 2524 3976 2536
rect 4028 2524 4034 2576
rect 8386 2524 8392 2576
rect 8444 2564 8450 2576
rect 8665 2567 8723 2573
rect 8665 2564 8677 2567
rect 8444 2536 8677 2564
rect 8444 2524 8450 2536
rect 8665 2533 8677 2536
rect 8711 2533 8723 2567
rect 8665 2527 8723 2533
rect 12250 2524 12256 2576
rect 12308 2564 12314 2576
rect 12437 2567 12495 2573
rect 12437 2564 12449 2567
rect 12308 2536 12449 2564
rect 12308 2524 12314 2536
rect 12437 2533 12449 2536
rect 12483 2564 12495 2567
rect 13814 2564 13820 2576
rect 12483 2536 13820 2564
rect 12483 2533 12495 2536
rect 12437 2527 12495 2533
rect 13814 2524 13820 2536
rect 13872 2524 13878 2576
rect 14182 2564 14188 2576
rect 14143 2536 14188 2564
rect 14182 2524 14188 2536
rect 14240 2524 14246 2576
rect 17129 2567 17187 2573
rect 17129 2533 17141 2567
rect 17175 2564 17187 2567
rect 17586 2564 17592 2576
rect 17175 2536 17592 2564
rect 17175 2533 17187 2536
rect 17129 2527 17187 2533
rect 17586 2524 17592 2536
rect 17644 2524 17650 2576
rect 18322 2524 18328 2576
rect 18380 2564 18386 2576
rect 18417 2567 18475 2573
rect 18417 2564 18429 2567
rect 18380 2536 18429 2564
rect 18380 2524 18386 2536
rect 18417 2533 18429 2536
rect 18463 2533 18475 2567
rect 18417 2527 18475 2533
rect 2314 2496 2320 2508
rect 2275 2468 2320 2496
rect 2314 2456 2320 2468
rect 2372 2456 2378 2508
rect 3237 2499 3295 2505
rect 3237 2465 3249 2499
rect 3283 2496 3295 2499
rect 3602 2496 3608 2508
rect 3283 2468 3608 2496
rect 3283 2465 3295 2468
rect 3237 2459 3295 2465
rect 3602 2456 3608 2468
rect 3660 2456 3666 2508
rect 5721 2499 5779 2505
rect 5721 2465 5733 2499
rect 5767 2496 5779 2499
rect 6362 2496 6368 2508
rect 5767 2468 6368 2496
rect 5767 2465 5779 2468
rect 5721 2459 5779 2465
rect 6362 2456 6368 2468
rect 6420 2456 6426 2508
rect 16758 2456 16764 2508
rect 16816 2496 16822 2508
rect 17310 2496 17316 2508
rect 16816 2468 17316 2496
rect 16816 2456 16822 2468
rect 17310 2456 17316 2468
rect 17368 2456 17374 2508
rect 17405 2499 17463 2505
rect 17405 2465 17417 2499
rect 17451 2496 17463 2499
rect 17494 2496 17500 2508
rect 17451 2468 17500 2496
rect 17451 2465 17463 2468
rect 17405 2459 17463 2465
rect 17494 2456 17500 2468
rect 17552 2456 17558 2508
rect 17954 2496 17960 2508
rect 17915 2468 17960 2496
rect 17954 2456 17960 2468
rect 18012 2456 18018 2508
rect 1673 2431 1731 2437
rect 1673 2397 1685 2431
rect 1719 2428 1731 2431
rect 1946 2428 1952 2440
rect 1719 2400 1952 2428
rect 1719 2397 1731 2400
rect 1673 2391 1731 2397
rect 1946 2388 1952 2400
rect 2004 2428 2010 2440
rect 3421 2431 3479 2437
rect 3421 2428 3433 2431
rect 2004 2400 3433 2428
rect 2004 2388 2010 2400
rect 3421 2397 3433 2400
rect 3467 2397 3479 2431
rect 5810 2428 5816 2440
rect 5771 2400 5816 2428
rect 3421 2391 3479 2397
rect 5810 2388 5816 2400
rect 5868 2388 5874 2440
rect 5997 2431 6055 2437
rect 5997 2397 6009 2431
rect 6043 2428 6055 2431
rect 6822 2428 6828 2440
rect 6043 2400 6828 2428
rect 6043 2397 6055 2400
rect 5997 2391 6055 2397
rect 6822 2388 6828 2400
rect 6880 2388 6886 2440
rect 8849 2431 8907 2437
rect 8849 2397 8861 2431
rect 8895 2428 8907 2431
rect 9674 2428 9680 2440
rect 8895 2400 9680 2428
rect 8895 2397 8907 2400
rect 8849 2391 8907 2397
rect 9674 2388 9680 2400
rect 9732 2388 9738 2440
rect 14366 2388 14372 2440
rect 14424 2428 14430 2440
rect 14829 2431 14887 2437
rect 14829 2428 14841 2431
rect 14424 2400 14841 2428
rect 14424 2388 14430 2400
rect 14829 2397 14841 2400
rect 14875 2397 14887 2431
rect 14829 2391 14887 2397
rect 15010 2388 15016 2440
rect 15068 2428 15074 2440
rect 16482 2428 16488 2440
rect 15068 2400 16488 2428
rect 15068 2388 15074 2400
rect 16482 2388 16488 2400
rect 16540 2388 16546 2440
rect 17402 2292 17408 2304
rect 17363 2264 17408 2292
rect 17402 2252 17408 2264
rect 17460 2252 17466 2304
rect 184 2202 18860 2224
rect 184 2150 1556 2202
rect 1608 2150 1620 2202
rect 1672 2150 1684 2202
rect 1736 2150 1748 2202
rect 1800 2150 1812 2202
rect 1864 2150 4656 2202
rect 4708 2150 4720 2202
rect 4772 2150 4784 2202
rect 4836 2150 4848 2202
rect 4900 2150 4912 2202
rect 4964 2150 7756 2202
rect 7808 2150 7820 2202
rect 7872 2150 7884 2202
rect 7936 2150 7948 2202
rect 8000 2150 8012 2202
rect 8064 2150 10856 2202
rect 10908 2150 10920 2202
rect 10972 2150 10984 2202
rect 11036 2150 11048 2202
rect 11100 2150 11112 2202
rect 11164 2150 13956 2202
rect 14008 2150 14020 2202
rect 14072 2150 14084 2202
rect 14136 2150 14148 2202
rect 14200 2150 14212 2202
rect 14264 2150 17056 2202
rect 17108 2150 17120 2202
rect 17172 2150 17184 2202
rect 17236 2150 17248 2202
rect 17300 2150 17312 2202
rect 17364 2150 18860 2202
rect 184 2128 18860 2150
rect 3602 2088 3608 2100
rect 3563 2060 3608 2088
rect 3602 2048 3608 2060
rect 3660 2048 3666 2100
rect 3970 2048 3976 2100
rect 4028 2088 4034 2100
rect 6362 2088 6368 2100
rect 4028 2060 5396 2088
rect 6323 2060 6368 2088
rect 4028 2048 4034 2060
rect 4246 1980 4252 2032
rect 4304 2020 4310 2032
rect 5258 2020 5264 2032
rect 4304 1992 5264 2020
rect 4304 1980 4310 1992
rect 5258 1980 5264 1992
rect 5316 1980 5322 2032
rect 5368 2029 5396 2060
rect 6362 2048 6368 2060
rect 6420 2048 6426 2100
rect 7374 2048 7380 2100
rect 7432 2088 7438 2100
rect 7653 2091 7711 2097
rect 7653 2088 7665 2091
rect 7432 2060 7665 2088
rect 7432 2048 7438 2060
rect 7653 2057 7665 2060
rect 7699 2057 7711 2091
rect 9858 2088 9864 2100
rect 9819 2060 9864 2088
rect 7653 2051 7711 2057
rect 9858 2048 9864 2060
rect 9916 2048 9922 2100
rect 10410 2088 10416 2100
rect 10323 2060 10416 2088
rect 10410 2048 10416 2060
rect 10468 2088 10474 2100
rect 10778 2088 10784 2100
rect 10468 2060 10784 2088
rect 10468 2048 10474 2060
rect 10778 2048 10784 2060
rect 10836 2048 10842 2100
rect 11517 2091 11575 2097
rect 11517 2057 11529 2091
rect 11563 2088 11575 2091
rect 11606 2088 11612 2100
rect 11563 2060 11612 2088
rect 11563 2057 11575 2060
rect 11517 2051 11575 2057
rect 11606 2048 11612 2060
rect 11664 2048 11670 2100
rect 12802 2048 12808 2100
rect 12860 2088 12866 2100
rect 13725 2091 13783 2097
rect 13725 2088 13737 2091
rect 12860 2060 13737 2088
rect 12860 2048 12866 2060
rect 13725 2057 13737 2060
rect 13771 2057 13783 2091
rect 14826 2088 14832 2100
rect 14787 2060 14832 2088
rect 13725 2051 13783 2057
rect 14826 2048 14832 2060
rect 14884 2048 14890 2100
rect 15933 2091 15991 2097
rect 15933 2057 15945 2091
rect 15979 2088 15991 2091
rect 16206 2088 16212 2100
rect 15979 2060 16212 2088
rect 15979 2057 15991 2060
rect 15933 2051 15991 2057
rect 16206 2048 16212 2060
rect 16264 2048 16270 2100
rect 5353 2023 5411 2029
rect 5353 1989 5365 2023
rect 5399 1989 5411 2023
rect 9030 2020 9036 2032
rect 5353 1983 5411 1989
rect 8956 1992 9036 2020
rect 2866 1912 2872 1964
rect 2924 1952 2930 1964
rect 3053 1955 3111 1961
rect 3053 1952 3065 1955
rect 2924 1924 3065 1952
rect 2924 1912 2930 1924
rect 3053 1921 3065 1924
rect 3099 1952 3111 1955
rect 5534 1952 5540 1964
rect 3099 1924 5540 1952
rect 3099 1921 3111 1924
rect 3053 1915 3111 1921
rect 5534 1912 5540 1924
rect 5592 1952 5598 1964
rect 6917 1955 6975 1961
rect 6917 1952 6929 1955
rect 5592 1924 6929 1952
rect 5592 1912 5598 1924
rect 3145 1887 3203 1893
rect 3145 1853 3157 1887
rect 3191 1884 3203 1887
rect 3326 1884 3332 1896
rect 3191 1856 3332 1884
rect 3191 1853 3203 1856
rect 3145 1847 3203 1853
rect 3326 1844 3332 1856
rect 3384 1844 3390 1896
rect 3510 1844 3516 1896
rect 3568 1844 3574 1896
rect 3970 1884 3976 1896
rect 3931 1856 3976 1884
rect 3970 1844 3976 1856
rect 4028 1844 4034 1896
rect 4246 1844 4252 1896
rect 4304 1884 4310 1896
rect 4341 1887 4399 1893
rect 4341 1884 4353 1887
rect 4304 1856 4353 1884
rect 4304 1844 4310 1856
rect 4341 1853 4353 1856
rect 4387 1853 4399 1887
rect 4341 1847 4399 1853
rect 4709 1887 4767 1893
rect 4709 1853 4721 1887
rect 4755 1884 4767 1887
rect 5166 1884 5172 1896
rect 4755 1856 5172 1884
rect 4755 1853 4767 1856
rect 4709 1847 4767 1853
rect 3528 1816 3556 1844
rect 4724 1816 4752 1847
rect 5166 1844 5172 1856
rect 5224 1844 5230 1896
rect 5258 1844 5264 1896
rect 5316 1884 5322 1896
rect 5445 1887 5503 1893
rect 5445 1884 5457 1887
rect 5316 1856 5457 1884
rect 5316 1844 5322 1856
rect 5445 1853 5457 1856
rect 5491 1853 5503 1887
rect 5445 1847 5503 1853
rect 5644 1816 5672 1924
rect 6917 1921 6929 1924
rect 6963 1921 6975 1955
rect 6917 1915 6975 1921
rect 7466 1912 7472 1964
rect 7524 1952 7530 1964
rect 8956 1961 8984 1992
rect 9030 1980 9036 1992
rect 9088 1980 9094 2032
rect 15838 1980 15844 2032
rect 15896 2020 15902 2032
rect 15896 1992 17356 2020
rect 15896 1980 15902 1992
rect 8113 1955 8171 1961
rect 8113 1952 8125 1955
rect 7524 1924 8125 1952
rect 7524 1912 7530 1924
rect 8113 1921 8125 1924
rect 8159 1921 8171 1955
rect 8113 1915 8171 1921
rect 8297 1955 8355 1961
rect 8297 1921 8309 1955
rect 8343 1952 8355 1955
rect 8941 1955 8999 1961
rect 8343 1924 8892 1952
rect 8343 1921 8355 1924
rect 8297 1915 8355 1921
rect 5810 1844 5816 1896
rect 5868 1884 5874 1896
rect 6730 1884 6736 1896
rect 5868 1856 6736 1884
rect 5868 1844 5874 1856
rect 6730 1844 6736 1856
rect 6788 1884 6794 1896
rect 6825 1887 6883 1893
rect 6825 1884 6837 1887
rect 6788 1856 6837 1884
rect 6788 1844 6794 1856
rect 6825 1853 6837 1856
rect 6871 1853 6883 1887
rect 6825 1847 6883 1853
rect 3528 1788 4752 1816
rect 4816 1788 5672 1816
rect 8864 1816 8892 1924
rect 8941 1921 8953 1955
rect 8987 1921 8999 1955
rect 9766 1952 9772 1964
rect 8941 1915 8999 1921
rect 9140 1924 9772 1952
rect 9140 1893 9168 1924
rect 9766 1912 9772 1924
rect 9824 1952 9830 1964
rect 10597 1955 10655 1961
rect 10597 1952 10609 1955
rect 9824 1924 10609 1952
rect 9824 1912 9830 1924
rect 10597 1921 10609 1924
rect 10643 1921 10655 1955
rect 10597 1915 10655 1921
rect 12161 1955 12219 1961
rect 12161 1921 12173 1955
rect 12207 1952 12219 1955
rect 13173 1955 13231 1961
rect 13173 1952 13185 1955
rect 12207 1924 13185 1952
rect 12207 1921 12219 1924
rect 12161 1915 12219 1921
rect 13173 1921 13185 1924
rect 13219 1952 13231 1955
rect 14366 1952 14372 1964
rect 13219 1924 14372 1952
rect 13219 1921 13231 1924
rect 13173 1915 13231 1921
rect 14366 1912 14372 1924
rect 14424 1912 14430 1964
rect 16482 1952 16488 1964
rect 16443 1924 16488 1952
rect 16482 1912 16488 1924
rect 16540 1912 16546 1964
rect 9125 1887 9183 1893
rect 9125 1853 9137 1887
rect 9171 1853 9183 1887
rect 9125 1847 9183 1853
rect 9214 1844 9220 1896
rect 9272 1884 9278 1896
rect 9309 1887 9367 1893
rect 9309 1884 9321 1887
rect 9272 1856 9321 1884
rect 9272 1844 9278 1856
rect 9309 1853 9321 1856
rect 9355 1853 9367 1887
rect 9309 1847 9367 1853
rect 9952 1887 10010 1893
rect 9952 1853 9964 1887
rect 9998 1853 10010 1887
rect 9952 1847 10010 1853
rect 9968 1816 9996 1847
rect 10042 1844 10048 1896
rect 10100 1884 10106 1896
rect 10318 1884 10324 1896
rect 10100 1856 10145 1884
rect 10279 1856 10324 1884
rect 10100 1844 10106 1856
rect 10318 1844 10324 1856
rect 10376 1844 10382 1896
rect 11977 1887 12035 1893
rect 11977 1853 11989 1887
rect 12023 1884 12035 1887
rect 12250 1884 12256 1896
rect 12023 1856 12256 1884
rect 12023 1853 12035 1856
rect 11977 1847 12035 1853
rect 12250 1844 12256 1856
rect 12308 1844 12314 1896
rect 12621 1887 12679 1893
rect 12621 1853 12633 1887
rect 12667 1853 12679 1887
rect 12802 1884 12808 1896
rect 12763 1856 12808 1884
rect 12621 1847 12679 1853
rect 10597 1819 10655 1825
rect 10597 1816 10609 1819
rect 8864 1788 9352 1816
rect 9968 1788 10609 1816
rect 3237 1751 3295 1757
rect 3237 1717 3249 1751
rect 3283 1748 3295 1751
rect 3510 1748 3516 1760
rect 3283 1720 3516 1748
rect 3283 1717 3295 1720
rect 3237 1711 3295 1717
rect 3510 1708 3516 1720
rect 3568 1708 3574 1760
rect 4709 1751 4767 1757
rect 4709 1717 4721 1751
rect 4755 1748 4767 1751
rect 4816 1748 4844 1788
rect 4755 1720 4844 1748
rect 5445 1751 5503 1757
rect 4755 1717 4767 1720
rect 4709 1711 4767 1717
rect 5445 1717 5457 1751
rect 5491 1748 5503 1751
rect 5534 1748 5540 1760
rect 5491 1720 5540 1748
rect 5491 1717 5503 1720
rect 5445 1711 5503 1717
rect 5534 1708 5540 1720
rect 5592 1708 5598 1760
rect 6730 1748 6736 1760
rect 6691 1720 6736 1748
rect 6730 1708 6736 1720
rect 6788 1708 6794 1760
rect 8018 1748 8024 1760
rect 7979 1720 8024 1748
rect 8018 1708 8024 1720
rect 8076 1708 8082 1760
rect 9324 1757 9352 1788
rect 10597 1785 10609 1788
rect 10643 1785 10655 1819
rect 10597 1779 10655 1785
rect 11146 1776 11152 1828
rect 11204 1816 11210 1828
rect 11606 1816 11612 1828
rect 11204 1788 11612 1816
rect 11204 1776 11210 1788
rect 11606 1776 11612 1788
rect 11664 1816 11670 1828
rect 12636 1816 12664 1847
rect 12802 1844 12808 1856
rect 12860 1844 12866 1896
rect 12989 1887 13047 1893
rect 12989 1853 13001 1887
rect 13035 1884 13047 1887
rect 13722 1884 13728 1896
rect 13035 1856 13728 1884
rect 13035 1853 13047 1856
rect 12989 1847 13047 1853
rect 13722 1844 13728 1856
rect 13780 1844 13786 1896
rect 14185 1887 14243 1893
rect 14185 1853 14197 1887
rect 14231 1884 14243 1887
rect 14826 1884 14832 1896
rect 14231 1856 14832 1884
rect 14231 1853 14243 1856
rect 14185 1847 14243 1853
rect 14826 1844 14832 1856
rect 14884 1884 14890 1896
rect 17218 1884 17224 1896
rect 14884 1856 17224 1884
rect 14884 1844 14890 1856
rect 17218 1844 17224 1856
rect 17276 1844 17282 1896
rect 17328 1884 17356 1992
rect 17402 1912 17408 1964
rect 17460 1952 17466 1964
rect 17497 1955 17555 1961
rect 17497 1952 17509 1955
rect 17460 1924 17509 1952
rect 17460 1912 17466 1924
rect 17497 1921 17509 1924
rect 17543 1921 17555 1955
rect 17497 1915 17555 1921
rect 17328 1856 17448 1884
rect 13538 1816 13544 1828
rect 11664 1788 13544 1816
rect 11664 1776 11670 1788
rect 13538 1776 13544 1788
rect 13596 1776 13602 1828
rect 17420 1825 17448 1856
rect 16301 1819 16359 1825
rect 16301 1785 16313 1819
rect 16347 1816 16359 1819
rect 17405 1819 17463 1825
rect 16347 1788 16988 1816
rect 16347 1785 16359 1788
rect 16301 1779 16359 1785
rect 9309 1751 9367 1757
rect 9309 1717 9321 1751
rect 9355 1748 9367 1751
rect 9674 1748 9680 1760
rect 9355 1720 9680 1748
rect 9355 1717 9367 1720
rect 9309 1711 9367 1717
rect 9674 1708 9680 1720
rect 9732 1708 9738 1760
rect 11882 1748 11888 1760
rect 11843 1720 11888 1748
rect 11882 1708 11888 1720
rect 11940 1708 11946 1760
rect 14090 1748 14096 1760
rect 14051 1720 14096 1748
rect 14090 1708 14096 1720
rect 14148 1708 14154 1760
rect 16393 1751 16451 1757
rect 16393 1717 16405 1751
rect 16439 1748 16451 1751
rect 16758 1748 16764 1760
rect 16439 1720 16764 1748
rect 16439 1717 16451 1720
rect 16393 1711 16451 1717
rect 16758 1708 16764 1720
rect 16816 1708 16822 1760
rect 16960 1757 16988 1788
rect 17405 1785 17417 1819
rect 17451 1816 17463 1819
rect 18325 1819 18383 1825
rect 18325 1816 18337 1819
rect 17451 1788 18337 1816
rect 17451 1785 17463 1788
rect 17405 1779 17463 1785
rect 18325 1785 18337 1788
rect 18371 1785 18383 1819
rect 18325 1779 18383 1785
rect 16945 1751 17003 1757
rect 16945 1717 16957 1751
rect 16991 1717 17003 1751
rect 17310 1748 17316 1760
rect 17271 1720 17316 1748
rect 16945 1711 17003 1717
rect 17310 1708 17316 1720
rect 17368 1708 17374 1760
rect 184 1658 18920 1680
rect 184 1606 3106 1658
rect 3158 1606 3170 1658
rect 3222 1606 3234 1658
rect 3286 1606 3298 1658
rect 3350 1606 3362 1658
rect 3414 1606 6206 1658
rect 6258 1606 6270 1658
rect 6322 1606 6334 1658
rect 6386 1606 6398 1658
rect 6450 1606 6462 1658
rect 6514 1606 9306 1658
rect 9358 1606 9370 1658
rect 9422 1606 9434 1658
rect 9486 1606 9498 1658
rect 9550 1606 9562 1658
rect 9614 1606 12406 1658
rect 12458 1606 12470 1658
rect 12522 1606 12534 1658
rect 12586 1606 12598 1658
rect 12650 1606 12662 1658
rect 12714 1606 15506 1658
rect 15558 1606 15570 1658
rect 15622 1606 15634 1658
rect 15686 1606 15698 1658
rect 15750 1606 15762 1658
rect 15814 1606 18606 1658
rect 18658 1606 18670 1658
rect 18722 1606 18734 1658
rect 18786 1606 18798 1658
rect 18850 1606 18862 1658
rect 18914 1606 18920 1658
rect 184 1584 18920 1606
rect 3421 1547 3479 1553
rect 3421 1513 3433 1547
rect 3467 1544 3479 1547
rect 3510 1544 3516 1556
rect 3467 1516 3516 1544
rect 3467 1513 3479 1516
rect 3421 1507 3479 1513
rect 3510 1504 3516 1516
rect 3568 1504 3574 1556
rect 5905 1547 5963 1553
rect 5905 1513 5917 1547
rect 5951 1544 5963 1547
rect 6730 1544 6736 1556
rect 5951 1516 6736 1544
rect 5951 1513 5963 1516
rect 5905 1507 5963 1513
rect 6730 1504 6736 1516
rect 6788 1504 6794 1556
rect 7193 1547 7251 1553
rect 7193 1513 7205 1547
rect 7239 1544 7251 1547
rect 8018 1544 8024 1556
rect 7239 1516 8024 1544
rect 7239 1513 7251 1516
rect 7193 1507 7251 1513
rect 8018 1504 8024 1516
rect 8076 1504 8082 1556
rect 9214 1544 9220 1556
rect 8680 1516 9220 1544
rect 3053 1411 3111 1417
rect 3053 1377 3065 1411
rect 3099 1408 3111 1411
rect 3602 1408 3608 1420
rect 3099 1380 3608 1408
rect 3099 1377 3111 1380
rect 3053 1371 3111 1377
rect 3602 1368 3608 1380
rect 3660 1368 3666 1420
rect 5534 1408 5540 1420
rect 5495 1380 5540 1408
rect 5534 1368 5540 1380
rect 5592 1368 5598 1420
rect 5626 1368 5632 1420
rect 5684 1408 5690 1420
rect 6825 1411 6883 1417
rect 5684 1380 5729 1408
rect 5684 1368 5690 1380
rect 6825 1377 6837 1411
rect 6871 1408 6883 1411
rect 7650 1408 7656 1420
rect 6871 1380 7656 1408
rect 6871 1377 6883 1380
rect 6825 1371 6883 1377
rect 7650 1368 7656 1380
rect 7708 1408 7714 1420
rect 8680 1408 8708 1516
rect 9214 1504 9220 1516
rect 9272 1504 9278 1556
rect 9953 1547 10011 1553
rect 9953 1513 9965 1547
rect 9999 1544 10011 1547
rect 10042 1544 10048 1556
rect 9999 1516 10048 1544
rect 9999 1513 10011 1516
rect 9953 1507 10011 1513
rect 10042 1504 10048 1516
rect 10100 1504 10106 1556
rect 11701 1547 11759 1553
rect 11701 1513 11713 1547
rect 11747 1544 11759 1547
rect 11882 1544 11888 1556
rect 11747 1516 11888 1544
rect 11747 1513 11759 1516
rect 11701 1507 11759 1513
rect 11882 1504 11888 1516
rect 11940 1504 11946 1556
rect 12250 1504 12256 1556
rect 12308 1544 12314 1556
rect 12345 1547 12403 1553
rect 12345 1544 12357 1547
rect 12308 1516 12357 1544
rect 12308 1504 12314 1516
rect 12345 1513 12357 1516
rect 12391 1513 12403 1547
rect 12345 1507 12403 1513
rect 16850 1504 16856 1556
rect 16908 1544 16914 1556
rect 17129 1547 17187 1553
rect 17129 1544 17141 1547
rect 16908 1516 17141 1544
rect 16908 1504 16914 1516
rect 17129 1513 17141 1516
rect 17175 1513 17187 1547
rect 17494 1544 17500 1556
rect 17455 1516 17500 1544
rect 17129 1507 17187 1513
rect 17494 1504 17500 1516
rect 17552 1544 17558 1556
rect 18233 1547 18291 1553
rect 18233 1544 18245 1547
rect 17552 1516 18245 1544
rect 17552 1504 17558 1516
rect 18233 1513 18245 1516
rect 18279 1513 18291 1547
rect 18233 1507 18291 1513
rect 8849 1479 8907 1485
rect 8849 1445 8861 1479
rect 8895 1476 8907 1479
rect 9030 1476 9036 1488
rect 8895 1448 9036 1476
rect 8895 1445 8907 1448
rect 8849 1439 8907 1445
rect 9030 1436 9036 1448
rect 9088 1436 9094 1488
rect 9232 1476 9260 1504
rect 10229 1479 10287 1485
rect 10229 1476 10241 1479
rect 9232 1448 10241 1476
rect 10229 1445 10241 1448
rect 10275 1476 10287 1479
rect 10318 1476 10324 1488
rect 10275 1448 10324 1476
rect 10275 1445 10287 1448
rect 10229 1439 10287 1445
rect 10318 1436 10324 1448
rect 10376 1436 10382 1488
rect 11057 1479 11115 1485
rect 11057 1445 11069 1479
rect 11103 1476 11115 1479
rect 11103 1448 11468 1476
rect 11103 1445 11115 1448
rect 11057 1439 11115 1445
rect 7708 1380 8708 1408
rect 8757 1411 8815 1417
rect 7708 1368 7714 1380
rect 8757 1377 8769 1411
rect 8803 1377 8815 1411
rect 8757 1371 8815 1377
rect 3145 1343 3203 1349
rect 3145 1309 3157 1343
rect 3191 1340 3203 1343
rect 3970 1340 3976 1352
rect 3191 1312 3976 1340
rect 3191 1309 3203 1312
rect 3145 1303 3203 1309
rect 3970 1300 3976 1312
rect 4028 1300 4034 1352
rect 6733 1343 6791 1349
rect 6733 1309 6745 1343
rect 6779 1340 6791 1343
rect 8772 1340 8800 1371
rect 9766 1368 9772 1420
rect 9824 1408 9830 1420
rect 9953 1411 10011 1417
rect 9953 1408 9965 1411
rect 9824 1380 9965 1408
rect 9824 1368 9830 1380
rect 9953 1377 9965 1380
rect 9999 1377 10011 1411
rect 9953 1371 10011 1377
rect 10045 1411 10103 1417
rect 10045 1377 10057 1411
rect 10091 1408 10103 1411
rect 10410 1408 10416 1420
rect 10091 1380 10416 1408
rect 10091 1377 10103 1380
rect 10045 1371 10103 1377
rect 10060 1340 10088 1371
rect 10410 1368 10416 1380
rect 10468 1368 10474 1420
rect 10781 1411 10839 1417
rect 10781 1377 10793 1411
rect 10827 1408 10839 1411
rect 11146 1408 11152 1420
rect 10827 1380 11152 1408
rect 10827 1377 10839 1380
rect 10781 1371 10839 1377
rect 11146 1368 11152 1380
rect 11204 1368 11210 1420
rect 11330 1408 11336 1420
rect 11291 1380 11336 1408
rect 11330 1368 11336 1380
rect 11388 1368 11394 1420
rect 11440 1417 11468 1448
rect 13722 1436 13728 1488
rect 13780 1476 13786 1488
rect 14737 1479 14795 1485
rect 14737 1476 14749 1479
rect 13780 1448 14749 1476
rect 13780 1436 13786 1448
rect 14737 1445 14749 1448
rect 14783 1445 14795 1479
rect 14737 1439 14795 1445
rect 17218 1436 17224 1488
rect 17276 1476 17282 1488
rect 17586 1476 17592 1488
rect 17276 1448 17592 1476
rect 17276 1436 17282 1448
rect 17586 1436 17592 1448
rect 17644 1436 17650 1488
rect 11426 1411 11484 1417
rect 11426 1377 11438 1411
rect 11472 1377 11484 1411
rect 11426 1371 11484 1377
rect 13357 1411 13415 1417
rect 13357 1377 13369 1411
rect 13403 1408 13415 1411
rect 13538 1408 13544 1420
rect 13403 1380 13544 1408
rect 13403 1377 13415 1380
rect 13357 1371 13415 1377
rect 13538 1368 13544 1380
rect 13596 1368 13602 1420
rect 14642 1368 14648 1420
rect 14700 1408 14706 1420
rect 14829 1411 14887 1417
rect 14829 1408 14841 1411
rect 14700 1380 14841 1408
rect 14700 1368 14706 1380
rect 14829 1377 14841 1380
rect 14875 1377 14887 1411
rect 14829 1371 14887 1377
rect 16117 1411 16175 1417
rect 16117 1377 16129 1411
rect 16163 1408 16175 1411
rect 16758 1408 16764 1420
rect 16163 1380 16764 1408
rect 16163 1377 16175 1380
rect 16117 1371 16175 1377
rect 16758 1368 16764 1380
rect 16816 1368 16822 1420
rect 18141 1411 18199 1417
rect 18141 1408 18153 1411
rect 16868 1380 18153 1408
rect 6779 1312 10088 1340
rect 11057 1343 11115 1349
rect 6779 1309 6791 1312
rect 6733 1303 6791 1309
rect 11057 1309 11069 1343
rect 11103 1340 11115 1343
rect 11238 1340 11244 1352
rect 11103 1312 11244 1340
rect 11103 1309 11115 1312
rect 11057 1303 11115 1309
rect 11238 1300 11244 1312
rect 11296 1340 11302 1352
rect 12802 1340 12808 1352
rect 11296 1312 12808 1340
rect 11296 1300 11302 1312
rect 12802 1300 12808 1312
rect 12860 1300 12866 1352
rect 13449 1343 13507 1349
rect 13449 1309 13461 1343
rect 13495 1340 13507 1343
rect 13814 1340 13820 1352
rect 13495 1312 13820 1340
rect 13495 1309 13507 1312
rect 13449 1303 13507 1309
rect 13814 1300 13820 1312
rect 13872 1340 13878 1352
rect 14660 1340 14688 1368
rect 13872 1312 14688 1340
rect 16209 1343 16267 1349
rect 13872 1300 13878 1312
rect 16209 1309 16221 1343
rect 16255 1340 16267 1343
rect 16574 1340 16580 1352
rect 16255 1312 16580 1340
rect 16255 1309 16267 1312
rect 16209 1303 16267 1309
rect 16574 1300 16580 1312
rect 16632 1340 16638 1352
rect 16868 1340 16896 1380
rect 18141 1377 18153 1380
rect 18187 1377 18199 1411
rect 18141 1371 18199 1377
rect 16632 1312 16896 1340
rect 17681 1343 17739 1349
rect 16632 1300 16638 1312
rect 17681 1309 17693 1343
rect 17727 1309 17739 1343
rect 17681 1303 17739 1309
rect 13725 1275 13783 1281
rect 13725 1241 13737 1275
rect 13771 1272 13783 1275
rect 14090 1272 14096 1284
rect 13771 1244 14096 1272
rect 13771 1241 13783 1244
rect 13725 1235 13783 1241
rect 14090 1232 14096 1244
rect 14148 1232 14154 1284
rect 16485 1275 16543 1281
rect 16485 1241 16497 1275
rect 16531 1272 16543 1275
rect 17310 1272 17316 1284
rect 16531 1244 17316 1272
rect 16531 1241 16543 1244
rect 16485 1235 16543 1241
rect 17310 1232 17316 1244
rect 17368 1232 17374 1284
rect 17402 1232 17408 1284
rect 17460 1272 17466 1284
rect 17696 1272 17724 1303
rect 17460 1244 17724 1272
rect 17460 1232 17466 1244
rect 10873 1207 10931 1213
rect 10873 1173 10885 1207
rect 10919 1204 10931 1207
rect 11422 1204 11428 1216
rect 10919 1176 11428 1204
rect 10919 1173 10931 1176
rect 10873 1167 10931 1173
rect 11422 1164 11428 1176
rect 11480 1164 11486 1216
rect 184 1114 18860 1136
rect 184 1062 1556 1114
rect 1608 1062 1620 1114
rect 1672 1062 1684 1114
rect 1736 1062 1748 1114
rect 1800 1062 1812 1114
rect 1864 1062 4656 1114
rect 4708 1062 4720 1114
rect 4772 1062 4784 1114
rect 4836 1062 4848 1114
rect 4900 1062 4912 1114
rect 4964 1062 7756 1114
rect 7808 1062 7820 1114
rect 7872 1062 7884 1114
rect 7936 1062 7948 1114
rect 8000 1062 8012 1114
rect 8064 1062 10856 1114
rect 10908 1062 10920 1114
rect 10972 1062 10984 1114
rect 11036 1062 11048 1114
rect 11100 1062 11112 1114
rect 11164 1062 13956 1114
rect 14008 1062 14020 1114
rect 14072 1062 14084 1114
rect 14136 1062 14148 1114
rect 14200 1062 14212 1114
rect 14264 1062 17056 1114
rect 17108 1062 17120 1114
rect 17172 1062 17184 1114
rect 17236 1062 17248 1114
rect 17300 1062 17312 1114
rect 17364 1062 18860 1114
rect 184 1040 18860 1062
rect 3970 960 3976 1012
rect 4028 1000 4034 1012
rect 5353 1003 5411 1009
rect 5353 1000 5365 1003
rect 4028 972 5365 1000
rect 4028 960 4034 972
rect 5353 969 5365 972
rect 5399 969 5411 1003
rect 5353 963 5411 969
rect 5445 1003 5503 1009
rect 5445 969 5457 1003
rect 5491 1000 5503 1003
rect 5626 1000 5632 1012
rect 5491 972 5632 1000
rect 5491 969 5503 972
rect 5445 963 5503 969
rect 5626 960 5632 972
rect 5684 960 5690 1012
rect 11330 1000 11336 1012
rect 11291 972 11336 1000
rect 11330 960 11336 972
rect 11388 960 11394 1012
rect 17221 1003 17279 1009
rect 17221 969 17233 1003
rect 17267 1000 17279 1003
rect 17586 1000 17592 1012
rect 17267 972 17592 1000
rect 17267 969 17279 972
rect 17221 963 17279 969
rect 17586 960 17592 972
rect 17644 960 17650 1012
rect 17954 1000 17960 1012
rect 17915 972 17960 1000
rect 17954 960 17960 972
rect 18012 960 18018 1012
rect 18414 1000 18420 1012
rect 18375 972 18420 1000
rect 18414 960 18420 972
rect 18472 960 18478 1012
rect 5258 892 5264 944
rect 5316 892 5322 944
rect 11422 932 11428 944
rect 11335 904 11428 932
rect 11422 892 11428 904
rect 11480 932 11486 944
rect 13814 932 13820 944
rect 11480 904 13820 932
rect 11480 892 11486 904
rect 13814 892 13820 904
rect 13872 892 13878 944
rect 5276 864 5304 892
rect 5537 867 5595 873
rect 5537 864 5549 867
rect 5276 836 5549 864
rect 5537 833 5549 836
rect 5583 833 5595 867
rect 11606 864 11612 876
rect 11567 836 11612 864
rect 5537 827 5595 833
rect 11606 824 11612 836
rect 11664 824 11670 876
rect 5166 756 5172 808
rect 5224 796 5230 808
rect 5261 799 5319 805
rect 5261 796 5273 799
rect 5224 768 5273 796
rect 5224 756 5230 768
rect 5261 765 5273 768
rect 5307 765 5319 799
rect 5261 759 5319 765
rect 11238 756 11244 808
rect 11296 796 11302 808
rect 11333 799 11391 805
rect 11333 796 11345 799
rect 11296 768 11345 796
rect 11296 756 11302 768
rect 11333 765 11345 768
rect 11379 765 11391 799
rect 11333 759 11391 765
rect 17773 799 17831 805
rect 17773 765 17785 799
rect 17819 796 17831 799
rect 18432 796 18460 960
rect 17819 768 18460 796
rect 17819 765 17831 768
rect 17773 759 17831 765
rect 184 570 18920 592
rect 184 518 3106 570
rect 3158 518 3170 570
rect 3222 518 3234 570
rect 3286 518 3298 570
rect 3350 518 3362 570
rect 3414 518 6206 570
rect 6258 518 6270 570
rect 6322 518 6334 570
rect 6386 518 6398 570
rect 6450 518 6462 570
rect 6514 518 9306 570
rect 9358 518 9370 570
rect 9422 518 9434 570
rect 9486 518 9498 570
rect 9550 518 9562 570
rect 9614 518 12406 570
rect 12458 518 12470 570
rect 12522 518 12534 570
rect 12586 518 12598 570
rect 12650 518 12662 570
rect 12714 518 15506 570
rect 15558 518 15570 570
rect 15622 518 15634 570
rect 15686 518 15698 570
rect 15750 518 15762 570
rect 15814 518 18606 570
rect 18658 518 18670 570
rect 18722 518 18734 570
rect 18786 518 18798 570
rect 18850 518 18862 570
rect 18914 518 18920 570
rect 184 496 18920 518
<< via1 >>
rect 1556 18470 1608 18522
rect 1620 18470 1672 18522
rect 1684 18470 1736 18522
rect 1748 18470 1800 18522
rect 1812 18470 1864 18522
rect 4656 18470 4708 18522
rect 4720 18470 4772 18522
rect 4784 18470 4836 18522
rect 4848 18470 4900 18522
rect 4912 18470 4964 18522
rect 7756 18470 7808 18522
rect 7820 18470 7872 18522
rect 7884 18470 7936 18522
rect 7948 18470 8000 18522
rect 8012 18470 8064 18522
rect 10856 18470 10908 18522
rect 10920 18470 10972 18522
rect 10984 18470 11036 18522
rect 11048 18470 11100 18522
rect 11112 18470 11164 18522
rect 13956 18470 14008 18522
rect 14020 18470 14072 18522
rect 14084 18470 14136 18522
rect 14148 18470 14200 18522
rect 14212 18470 14264 18522
rect 17056 18470 17108 18522
rect 17120 18470 17172 18522
rect 17184 18470 17236 18522
rect 17248 18470 17300 18522
rect 17312 18470 17364 18522
rect 4252 18368 4304 18420
rect 18420 18411 18472 18420
rect 18420 18377 18429 18411
rect 18429 18377 18463 18411
rect 18463 18377 18472 18411
rect 18420 18368 18472 18377
rect 5816 18300 5868 18352
rect 9864 18300 9916 18352
rect 5724 18232 5776 18284
rect 8208 18275 8260 18284
rect 8208 18241 8217 18275
rect 8217 18241 8251 18275
rect 8251 18241 8260 18275
rect 8208 18232 8260 18241
rect 1400 18164 1452 18216
rect 3976 18207 4028 18216
rect 2780 18096 2832 18148
rect 2872 18096 2924 18148
rect 3976 18173 3985 18207
rect 3985 18173 4019 18207
rect 4019 18173 4028 18207
rect 3976 18164 4028 18173
rect 4160 18207 4212 18216
rect 4160 18173 4169 18207
rect 4169 18173 4203 18207
rect 4203 18173 4212 18207
rect 4160 18164 4212 18173
rect 4528 18207 4580 18216
rect 4528 18173 4537 18207
rect 4537 18173 4571 18207
rect 4571 18173 4580 18207
rect 4528 18164 4580 18173
rect 3884 18096 3936 18148
rect 6828 18164 6880 18216
rect 8760 18207 8812 18216
rect 8760 18173 8769 18207
rect 8769 18173 8803 18207
rect 8803 18173 8812 18207
rect 8760 18164 8812 18173
rect 11336 18164 11388 18216
rect 12992 18232 13044 18284
rect 12900 18207 12952 18216
rect 12900 18173 12909 18207
rect 12909 18173 12943 18207
rect 12943 18173 12952 18207
rect 12900 18164 12952 18173
rect 14372 18164 14424 18216
rect 14924 18207 14976 18216
rect 14924 18173 14933 18207
rect 14933 18173 14967 18207
rect 14967 18173 14976 18207
rect 14924 18164 14976 18173
rect 16672 18164 16724 18216
rect 18420 18164 18472 18216
rect 9220 18096 9272 18148
rect 13820 18096 13872 18148
rect 14648 18096 14700 18148
rect 14832 18139 14884 18148
rect 14832 18105 14841 18139
rect 14841 18105 14875 18139
rect 14875 18105 14884 18139
rect 14832 18096 14884 18105
rect 2504 18028 2556 18080
rect 4436 18071 4488 18080
rect 4436 18037 4445 18071
rect 4445 18037 4479 18071
rect 4479 18037 4488 18071
rect 4436 18028 4488 18037
rect 5540 18071 5592 18080
rect 5540 18037 5549 18071
rect 5549 18037 5583 18071
rect 5583 18037 5592 18071
rect 5540 18028 5592 18037
rect 5632 18071 5684 18080
rect 5632 18037 5641 18071
rect 5641 18037 5675 18071
rect 5675 18037 5684 18071
rect 7564 18071 7616 18080
rect 5632 18028 5684 18037
rect 7564 18037 7573 18071
rect 7573 18037 7607 18071
rect 7607 18037 7616 18071
rect 7564 18028 7616 18037
rect 8116 18028 8168 18080
rect 9128 18028 9180 18080
rect 9956 18071 10008 18080
rect 9956 18037 9965 18071
rect 9965 18037 9999 18071
rect 9999 18037 10008 18071
rect 9956 18028 10008 18037
rect 10324 18071 10376 18080
rect 10324 18037 10333 18071
rect 10333 18037 10367 18071
rect 10367 18037 10376 18071
rect 10324 18028 10376 18037
rect 11244 18028 11296 18080
rect 13268 18028 13320 18080
rect 15936 18071 15988 18080
rect 15936 18037 15945 18071
rect 15945 18037 15979 18071
rect 15979 18037 15988 18071
rect 15936 18028 15988 18037
rect 16580 18028 16632 18080
rect 3106 17926 3158 17978
rect 3170 17926 3222 17978
rect 3234 17926 3286 17978
rect 3298 17926 3350 17978
rect 3362 17926 3414 17978
rect 6206 17926 6258 17978
rect 6270 17926 6322 17978
rect 6334 17926 6386 17978
rect 6398 17926 6450 17978
rect 6462 17926 6514 17978
rect 9306 17926 9358 17978
rect 9370 17926 9422 17978
rect 9434 17926 9486 17978
rect 9498 17926 9550 17978
rect 9562 17926 9614 17978
rect 12406 17926 12458 17978
rect 12470 17926 12522 17978
rect 12534 17926 12586 17978
rect 12598 17926 12650 17978
rect 12662 17926 12714 17978
rect 15506 17926 15558 17978
rect 15570 17926 15622 17978
rect 15634 17926 15686 17978
rect 15698 17926 15750 17978
rect 15762 17926 15814 17978
rect 18606 17926 18658 17978
rect 18670 17926 18722 17978
rect 18734 17926 18786 17978
rect 18798 17926 18850 17978
rect 18862 17926 18914 17978
rect 3056 17824 3108 17876
rect 3976 17824 4028 17876
rect 13636 17824 13688 17876
rect 2412 17756 2464 17808
rect 4160 17756 4212 17808
rect 4436 17756 4488 17808
rect 7564 17756 7616 17808
rect 9864 17756 9916 17808
rect 2688 17688 2740 17740
rect 4252 17688 4304 17740
rect 12440 17688 12492 17740
rect 16120 17756 16172 17808
rect 12900 17731 12952 17740
rect 12900 17697 12909 17731
rect 12909 17697 12943 17731
rect 12943 17697 12952 17731
rect 12900 17688 12952 17697
rect 14832 17688 14884 17740
rect 16764 17688 16816 17740
rect 572 17663 624 17672
rect 572 17629 581 17663
rect 581 17629 615 17663
rect 615 17629 624 17663
rect 572 17620 624 17629
rect 848 17663 900 17672
rect 848 17629 857 17663
rect 857 17629 891 17663
rect 891 17629 900 17663
rect 848 17620 900 17629
rect 2780 17552 2832 17604
rect 5172 17552 5224 17604
rect 9220 17552 9272 17604
rect 11520 17552 11572 17604
rect 11980 17552 12032 17604
rect 12808 17620 12860 17672
rect 15108 17663 15160 17672
rect 15108 17629 15117 17663
rect 15117 17629 15151 17663
rect 15151 17629 15160 17663
rect 15108 17620 15160 17629
rect 2044 17484 2096 17536
rect 4436 17484 4488 17536
rect 7012 17484 7064 17536
rect 11428 17527 11480 17536
rect 11428 17493 11437 17527
rect 11437 17493 11471 17527
rect 11471 17493 11480 17527
rect 11428 17484 11480 17493
rect 11888 17484 11940 17536
rect 13084 17552 13136 17604
rect 12716 17484 12768 17536
rect 16304 17552 16356 17604
rect 16856 17484 16908 17536
rect 1556 17382 1608 17434
rect 1620 17382 1672 17434
rect 1684 17382 1736 17434
rect 1748 17382 1800 17434
rect 1812 17382 1864 17434
rect 4656 17382 4708 17434
rect 4720 17382 4772 17434
rect 4784 17382 4836 17434
rect 4848 17382 4900 17434
rect 4912 17382 4964 17434
rect 7756 17382 7808 17434
rect 7820 17382 7872 17434
rect 7884 17382 7936 17434
rect 7948 17382 8000 17434
rect 8012 17382 8064 17434
rect 10856 17382 10908 17434
rect 10920 17382 10972 17434
rect 10984 17382 11036 17434
rect 11048 17382 11100 17434
rect 11112 17382 11164 17434
rect 13956 17382 14008 17434
rect 14020 17382 14072 17434
rect 14084 17382 14136 17434
rect 14148 17382 14200 17434
rect 14212 17382 14264 17434
rect 17056 17382 17108 17434
rect 17120 17382 17172 17434
rect 17184 17382 17236 17434
rect 17248 17382 17300 17434
rect 17312 17382 17364 17434
rect 1400 17280 1452 17332
rect 2688 17323 2740 17332
rect 848 17255 900 17264
rect 848 17221 857 17255
rect 857 17221 891 17255
rect 891 17221 900 17255
rect 848 17212 900 17221
rect 2688 17289 2697 17323
rect 2697 17289 2731 17323
rect 2731 17289 2740 17323
rect 2688 17280 2740 17289
rect 5632 17280 5684 17332
rect 8760 17280 8812 17332
rect 2596 17212 2648 17264
rect 3056 17187 3108 17196
rect 3056 17153 3065 17187
rect 3065 17153 3099 17187
rect 3099 17153 3108 17187
rect 3056 17144 3108 17153
rect 5816 17144 5868 17196
rect 12992 17280 13044 17332
rect 13176 17280 13228 17332
rect 12808 17212 12860 17264
rect 12900 17212 12952 17264
rect 13452 17212 13504 17264
rect 11244 17144 11296 17196
rect 13820 17187 13872 17196
rect 1124 17119 1176 17128
rect 1124 17085 1132 17119
rect 1132 17085 1166 17119
rect 1166 17085 1176 17119
rect 1124 17076 1176 17085
rect 1216 17119 1268 17128
rect 1216 17085 1225 17119
rect 1225 17085 1259 17119
rect 1259 17085 1268 17119
rect 1216 17076 1268 17085
rect 2412 17076 2464 17128
rect 2688 17076 2740 17128
rect 4436 17076 4488 17128
rect 5908 17076 5960 17128
rect 4804 17008 4856 17060
rect 7380 17008 7432 17060
rect 9220 17008 9272 17060
rect 12440 17119 12492 17128
rect 12440 17085 12449 17119
rect 12449 17085 12483 17119
rect 12483 17085 12492 17119
rect 12716 17119 12768 17128
rect 12440 17076 12492 17085
rect 12716 17085 12725 17119
rect 12725 17085 12759 17119
rect 12759 17085 12768 17119
rect 12716 17076 12768 17085
rect 12900 17008 12952 17060
rect 2504 16983 2556 16992
rect 2504 16949 2513 16983
rect 2513 16949 2547 16983
rect 2547 16949 2556 16983
rect 2504 16940 2556 16949
rect 4344 16940 4396 16992
rect 11612 16983 11664 16992
rect 11612 16949 11621 16983
rect 11621 16949 11655 16983
rect 11655 16949 11664 16983
rect 11612 16940 11664 16949
rect 11704 16983 11756 16992
rect 11704 16949 11713 16983
rect 11713 16949 11747 16983
rect 11747 16949 11756 16983
rect 11704 16940 11756 16949
rect 13820 17153 13829 17187
rect 13829 17153 13863 17187
rect 13863 17153 13872 17187
rect 13820 17144 13872 17153
rect 13084 17076 13136 17128
rect 13360 17076 13412 17128
rect 16672 17280 16724 17332
rect 18236 17144 18288 17196
rect 16028 17076 16080 17128
rect 16212 17076 16264 17128
rect 14096 17051 14148 17060
rect 14096 17017 14105 17051
rect 14105 17017 14139 17051
rect 14139 17017 14148 17051
rect 14096 17008 14148 17017
rect 17500 17008 17552 17060
rect 13728 16940 13780 16992
rect 14004 16940 14056 16992
rect 16580 16940 16632 16992
rect 17776 16940 17828 16992
rect 3106 16838 3158 16890
rect 3170 16838 3222 16890
rect 3234 16838 3286 16890
rect 3298 16838 3350 16890
rect 3362 16838 3414 16890
rect 6206 16838 6258 16890
rect 6270 16838 6322 16890
rect 6334 16838 6386 16890
rect 6398 16838 6450 16890
rect 6462 16838 6514 16890
rect 9306 16838 9358 16890
rect 9370 16838 9422 16890
rect 9434 16838 9486 16890
rect 9498 16838 9550 16890
rect 9562 16838 9614 16890
rect 12406 16838 12458 16890
rect 12470 16838 12522 16890
rect 12534 16838 12586 16890
rect 12598 16838 12650 16890
rect 12662 16838 12714 16890
rect 15506 16838 15558 16890
rect 15570 16838 15622 16890
rect 15634 16838 15686 16890
rect 15698 16838 15750 16890
rect 15762 16838 15814 16890
rect 18606 16838 18658 16890
rect 18670 16838 18722 16890
rect 18734 16838 18786 16890
rect 18798 16838 18850 16890
rect 18862 16838 18914 16890
rect 1216 16736 1268 16788
rect 2504 16736 2556 16788
rect 11336 16736 11388 16788
rect 11612 16736 11664 16788
rect 12716 16736 12768 16788
rect 1124 16668 1176 16720
rect 2044 16643 2096 16652
rect 2044 16609 2053 16643
rect 2053 16609 2087 16643
rect 2087 16609 2096 16643
rect 2044 16600 2096 16609
rect 2136 16600 2188 16652
rect 2596 16668 2648 16720
rect 2688 16600 2740 16652
rect 2872 16643 2924 16652
rect 2872 16609 2881 16643
rect 2881 16609 2915 16643
rect 2915 16609 2924 16643
rect 2872 16600 2924 16609
rect 4068 16643 4120 16652
rect 4068 16609 4077 16643
rect 4077 16609 4111 16643
rect 4111 16609 4120 16643
rect 4068 16600 4120 16609
rect 5632 16668 5684 16720
rect 7012 16711 7064 16720
rect 7012 16677 7021 16711
rect 7021 16677 7055 16711
rect 7055 16677 7064 16711
rect 7012 16668 7064 16677
rect 7472 16668 7524 16720
rect 14004 16736 14056 16788
rect 14096 16736 14148 16788
rect 4804 16643 4856 16652
rect 4804 16609 4813 16643
rect 4813 16609 4847 16643
rect 4847 16609 4856 16643
rect 4804 16600 4856 16609
rect 4528 16532 4580 16584
rect 9128 16600 9180 16652
rect 9864 16600 9916 16652
rect 9956 16643 10008 16652
rect 9956 16609 9965 16643
rect 9965 16609 9999 16643
rect 9999 16609 10008 16643
rect 9956 16600 10008 16609
rect 11336 16532 11388 16584
rect 2596 16464 2648 16516
rect 5816 16464 5868 16516
rect 7104 16464 7156 16516
rect 10048 16464 10100 16516
rect 11520 16464 11572 16516
rect 13176 16464 13228 16516
rect 13452 16507 13504 16516
rect 13452 16473 13461 16507
rect 13461 16473 13495 16507
rect 13495 16473 13504 16507
rect 13452 16464 13504 16473
rect 13820 16668 13872 16720
rect 13636 16600 13688 16652
rect 16764 16668 16816 16720
rect 17500 16668 17552 16720
rect 17776 16643 17828 16652
rect 17776 16609 17785 16643
rect 17785 16609 17819 16643
rect 17819 16609 17828 16643
rect 17776 16600 17828 16609
rect 18420 16643 18472 16652
rect 18420 16609 18429 16643
rect 18429 16609 18463 16643
rect 18463 16609 18472 16643
rect 18420 16600 18472 16609
rect 14280 16575 14332 16584
rect 14280 16541 14289 16575
rect 14289 16541 14323 16575
rect 14323 16541 14332 16575
rect 14280 16532 14332 16541
rect 15936 16532 15988 16584
rect 2228 16439 2280 16448
rect 2228 16405 2237 16439
rect 2237 16405 2271 16439
rect 2271 16405 2280 16439
rect 2228 16396 2280 16405
rect 12716 16439 12768 16448
rect 12716 16405 12725 16439
rect 12725 16405 12759 16439
rect 12759 16405 12768 16439
rect 12716 16396 12768 16405
rect 13268 16396 13320 16448
rect 14280 16396 14332 16448
rect 16396 16396 16448 16448
rect 16764 16396 16816 16448
rect 1556 16294 1608 16346
rect 1620 16294 1672 16346
rect 1684 16294 1736 16346
rect 1748 16294 1800 16346
rect 1812 16294 1864 16346
rect 4656 16294 4708 16346
rect 4720 16294 4772 16346
rect 4784 16294 4836 16346
rect 4848 16294 4900 16346
rect 4912 16294 4964 16346
rect 7756 16294 7808 16346
rect 7820 16294 7872 16346
rect 7884 16294 7936 16346
rect 7948 16294 8000 16346
rect 8012 16294 8064 16346
rect 10856 16294 10908 16346
rect 10920 16294 10972 16346
rect 10984 16294 11036 16346
rect 11048 16294 11100 16346
rect 11112 16294 11164 16346
rect 13956 16294 14008 16346
rect 14020 16294 14072 16346
rect 14084 16294 14136 16346
rect 14148 16294 14200 16346
rect 14212 16294 14264 16346
rect 17056 16294 17108 16346
rect 17120 16294 17172 16346
rect 17184 16294 17236 16346
rect 17248 16294 17300 16346
rect 17312 16294 17364 16346
rect 5540 16192 5592 16244
rect 10324 16192 10376 16244
rect 13820 16235 13872 16244
rect 13820 16201 13829 16235
rect 13829 16201 13863 16235
rect 13863 16201 13872 16235
rect 13820 16192 13872 16201
rect 18420 16167 18472 16176
rect 18420 16133 18429 16167
rect 18429 16133 18463 16167
rect 18463 16133 18472 16167
rect 18420 16124 18472 16133
rect 5172 16056 5224 16108
rect 5632 16056 5684 16108
rect 16764 16056 16816 16108
rect 2320 15988 2372 16040
rect 2596 16031 2648 16040
rect 2596 15997 2605 16031
rect 2605 15997 2639 16031
rect 2639 15997 2648 16031
rect 2596 15988 2648 15997
rect 4344 15920 4396 15972
rect 7012 15988 7064 16040
rect 11336 15988 11388 16040
rect 16212 15988 16264 16040
rect 6552 15920 6604 15972
rect 9036 15920 9088 15972
rect 11152 15963 11204 15972
rect 11152 15929 11161 15963
rect 11161 15929 11195 15963
rect 11195 15929 11204 15963
rect 11152 15920 11204 15929
rect 11428 15920 11480 15972
rect 15016 15920 15068 15972
rect 17500 15920 17552 15972
rect 3608 15852 3660 15904
rect 8024 15852 8076 15904
rect 17868 15852 17920 15904
rect 3106 15750 3158 15802
rect 3170 15750 3222 15802
rect 3234 15750 3286 15802
rect 3298 15750 3350 15802
rect 3362 15750 3414 15802
rect 6206 15750 6258 15802
rect 6270 15750 6322 15802
rect 6334 15750 6386 15802
rect 6398 15750 6450 15802
rect 6462 15750 6514 15802
rect 9306 15750 9358 15802
rect 9370 15750 9422 15802
rect 9434 15750 9486 15802
rect 9498 15750 9550 15802
rect 9562 15750 9614 15802
rect 12406 15750 12458 15802
rect 12470 15750 12522 15802
rect 12534 15750 12586 15802
rect 12598 15750 12650 15802
rect 12662 15750 12714 15802
rect 15506 15750 15558 15802
rect 15570 15750 15622 15802
rect 15634 15750 15686 15802
rect 15698 15750 15750 15802
rect 15762 15750 15814 15802
rect 18606 15750 18658 15802
rect 18670 15750 18722 15802
rect 18734 15750 18786 15802
rect 18798 15750 18850 15802
rect 18862 15750 18914 15802
rect 4068 15648 4120 15700
rect 6828 15648 6880 15700
rect 4436 15580 4488 15632
rect 11152 15648 11204 15700
rect 11980 15691 12032 15700
rect 11980 15657 11989 15691
rect 11989 15657 12023 15691
rect 12023 15657 12032 15691
rect 11980 15648 12032 15657
rect 12808 15648 12860 15700
rect 14280 15648 14332 15700
rect 18236 15691 18288 15700
rect 18236 15657 18245 15691
rect 18245 15657 18279 15691
rect 18279 15657 18288 15691
rect 18236 15648 18288 15657
rect 8024 15580 8076 15632
rect 8300 15580 8352 15632
rect 11520 15580 11572 15632
rect 13452 15580 13504 15632
rect 14372 15580 14424 15632
rect 16304 15580 16356 15632
rect 17868 15580 17920 15632
rect 12808 15555 12860 15564
rect 12808 15521 12817 15555
rect 12817 15521 12851 15555
rect 12851 15521 12860 15555
rect 12808 15512 12860 15521
rect 13268 15512 13320 15564
rect 16488 15555 16540 15564
rect 16488 15521 16497 15555
rect 16497 15521 16531 15555
rect 16531 15521 16540 15555
rect 16488 15512 16540 15521
rect 19064 15512 19116 15564
rect 7656 15444 7708 15496
rect 10232 15487 10284 15496
rect 10232 15453 10241 15487
rect 10241 15453 10275 15487
rect 10275 15453 10284 15487
rect 10232 15444 10284 15453
rect 11520 15444 11572 15496
rect 12900 15487 12952 15496
rect 12900 15453 12909 15487
rect 12909 15453 12943 15487
rect 12943 15453 12952 15487
rect 12900 15444 12952 15453
rect 13820 15487 13872 15496
rect 13820 15453 13829 15487
rect 13829 15453 13863 15487
rect 13863 15453 13872 15487
rect 13820 15444 13872 15453
rect 9496 15351 9548 15360
rect 9496 15317 9505 15351
rect 9505 15317 9539 15351
rect 9539 15317 9548 15351
rect 9496 15308 9548 15317
rect 12348 15351 12400 15360
rect 12348 15317 12357 15351
rect 12357 15317 12391 15351
rect 12391 15317 12400 15351
rect 12348 15308 12400 15317
rect 14832 15308 14884 15360
rect 15016 15308 15068 15360
rect 1556 15206 1608 15258
rect 1620 15206 1672 15258
rect 1684 15206 1736 15258
rect 1748 15206 1800 15258
rect 1812 15206 1864 15258
rect 4656 15206 4708 15258
rect 4720 15206 4772 15258
rect 4784 15206 4836 15258
rect 4848 15206 4900 15258
rect 4912 15206 4964 15258
rect 7756 15206 7808 15258
rect 7820 15206 7872 15258
rect 7884 15206 7936 15258
rect 7948 15206 8000 15258
rect 8012 15206 8064 15258
rect 10856 15206 10908 15258
rect 10920 15206 10972 15258
rect 10984 15206 11036 15258
rect 11048 15206 11100 15258
rect 11112 15206 11164 15258
rect 13956 15206 14008 15258
rect 14020 15206 14072 15258
rect 14084 15206 14136 15258
rect 14148 15206 14200 15258
rect 14212 15206 14264 15258
rect 17056 15206 17108 15258
rect 17120 15206 17172 15258
rect 17184 15206 17236 15258
rect 17248 15206 17300 15258
rect 17312 15206 17364 15258
rect 5908 15147 5960 15156
rect 5908 15113 5917 15147
rect 5917 15113 5951 15147
rect 5951 15113 5960 15147
rect 5908 15104 5960 15113
rect 8208 15104 8260 15156
rect 9864 15104 9916 15156
rect 12992 15104 13044 15156
rect 13636 15104 13688 15156
rect 15108 15104 15160 15156
rect 2136 15011 2188 15020
rect 2136 14977 2145 15011
rect 2145 14977 2179 15011
rect 2179 14977 2188 15011
rect 2136 14968 2188 14977
rect 2228 14968 2280 15020
rect 2596 14900 2648 14952
rect 3608 14943 3660 14952
rect 2688 14832 2740 14884
rect 3608 14909 3617 14943
rect 3617 14909 3651 14943
rect 3651 14909 3660 14943
rect 3608 14900 3660 14909
rect 4068 14943 4120 14952
rect 4068 14909 4077 14943
rect 4077 14909 4111 14943
rect 4111 14909 4120 14943
rect 4068 14900 4120 14909
rect 8760 15036 8812 15088
rect 9496 15036 9548 15088
rect 11980 15036 12032 15088
rect 6644 14968 6696 15020
rect 5816 14943 5868 14952
rect 5816 14909 5825 14943
rect 5825 14909 5859 14943
rect 5859 14909 5868 14943
rect 5816 14900 5868 14909
rect 8116 14900 8168 14952
rect 11336 14943 11388 14952
rect 11336 14909 11345 14943
rect 11345 14909 11379 14943
rect 11379 14909 11388 14943
rect 11336 14900 11388 14909
rect 12348 14900 12400 14952
rect 4988 14875 5040 14884
rect 4988 14841 4997 14875
rect 4997 14841 5031 14875
rect 5031 14841 5040 14875
rect 4988 14832 5040 14841
rect 6920 14832 6972 14884
rect 848 14764 900 14816
rect 2964 14764 3016 14816
rect 3516 14807 3568 14816
rect 3516 14773 3525 14807
rect 3525 14773 3559 14807
rect 3559 14773 3568 14807
rect 3516 14764 3568 14773
rect 4804 14764 4856 14816
rect 7564 14764 7616 14816
rect 12900 14900 12952 14952
rect 12992 14943 13044 14952
rect 12992 14909 13001 14943
rect 13001 14909 13035 14943
rect 13035 14909 13044 14943
rect 12992 14900 13044 14909
rect 13912 14943 13964 14952
rect 13912 14909 13921 14943
rect 13921 14909 13955 14943
rect 13955 14909 13964 14943
rect 13912 14900 13964 14909
rect 15200 14968 15252 15020
rect 14832 14900 14884 14952
rect 13728 14832 13780 14884
rect 16856 14968 16908 15020
rect 16212 14943 16264 14952
rect 16212 14909 16221 14943
rect 16221 14909 16255 14943
rect 16255 14909 16264 14943
rect 16212 14900 16264 14909
rect 17592 14900 17644 14952
rect 16764 14832 16816 14884
rect 9036 14764 9088 14816
rect 11336 14764 11388 14816
rect 12256 14807 12308 14816
rect 12256 14773 12265 14807
rect 12265 14773 12299 14807
rect 12299 14773 12308 14807
rect 12256 14764 12308 14773
rect 12992 14764 13044 14816
rect 14280 14807 14332 14816
rect 14280 14773 14289 14807
rect 14289 14773 14323 14807
rect 14323 14773 14332 14807
rect 14280 14764 14332 14773
rect 14648 14764 14700 14816
rect 14832 14764 14884 14816
rect 16580 14764 16632 14816
rect 17960 14807 18012 14816
rect 17960 14773 17969 14807
rect 17969 14773 18003 14807
rect 18003 14773 18012 14807
rect 17960 14764 18012 14773
rect 3106 14662 3158 14714
rect 3170 14662 3222 14714
rect 3234 14662 3286 14714
rect 3298 14662 3350 14714
rect 3362 14662 3414 14714
rect 6206 14662 6258 14714
rect 6270 14662 6322 14714
rect 6334 14662 6386 14714
rect 6398 14662 6450 14714
rect 6462 14662 6514 14714
rect 9306 14662 9358 14714
rect 9370 14662 9422 14714
rect 9434 14662 9486 14714
rect 9498 14662 9550 14714
rect 9562 14662 9614 14714
rect 12406 14662 12458 14714
rect 12470 14662 12522 14714
rect 12534 14662 12586 14714
rect 12598 14662 12650 14714
rect 12662 14662 12714 14714
rect 15506 14662 15558 14714
rect 15570 14662 15622 14714
rect 15634 14662 15686 14714
rect 15698 14662 15750 14714
rect 15762 14662 15814 14714
rect 18606 14662 18658 14714
rect 18670 14662 18722 14714
rect 18734 14662 18786 14714
rect 18798 14662 18850 14714
rect 18862 14662 18914 14714
rect 2596 14560 2648 14612
rect 2688 14560 2740 14612
rect 2964 14560 3016 14612
rect 848 14535 900 14544
rect 848 14501 857 14535
rect 857 14501 891 14535
rect 891 14501 900 14535
rect 848 14492 900 14501
rect 2136 14492 2188 14544
rect 4988 14560 5040 14612
rect 7656 14603 7708 14612
rect 7656 14569 7665 14603
rect 7665 14569 7699 14603
rect 7699 14569 7708 14603
rect 7656 14560 7708 14569
rect 11520 14560 11572 14612
rect 11704 14560 11756 14612
rect 12808 14560 12860 14612
rect 14280 14560 14332 14612
rect 14372 14560 14424 14612
rect 16672 14560 16724 14612
rect 16764 14560 16816 14612
rect 572 14467 624 14476
rect 572 14433 581 14467
rect 581 14433 615 14467
rect 615 14433 624 14467
rect 572 14424 624 14433
rect 2320 14424 2372 14476
rect 2504 14424 2556 14476
rect 3148 14467 3200 14476
rect 3148 14433 3157 14467
rect 3157 14433 3191 14467
rect 3191 14433 3200 14467
rect 3148 14424 3200 14433
rect 6552 14492 6604 14544
rect 4804 14467 4856 14476
rect 4804 14433 4813 14467
rect 4813 14433 4847 14467
rect 4847 14433 4856 14467
rect 4804 14424 4856 14433
rect 5172 14467 5224 14476
rect 5172 14433 5181 14467
rect 5181 14433 5215 14467
rect 5215 14433 5224 14467
rect 5172 14424 5224 14433
rect 3516 14356 3568 14408
rect 4068 14399 4120 14408
rect 4068 14365 4077 14399
rect 4077 14365 4111 14399
rect 4111 14365 4120 14399
rect 4068 14356 4120 14365
rect 7472 14424 7524 14476
rect 6644 14356 6696 14408
rect 8116 14356 8168 14408
rect 7012 14220 7064 14272
rect 9128 14220 9180 14272
rect 11336 14467 11388 14476
rect 11336 14433 11345 14467
rect 11345 14433 11379 14467
rect 11379 14433 11388 14467
rect 11336 14424 11388 14433
rect 11888 14467 11940 14476
rect 11888 14433 11896 14467
rect 11896 14433 11930 14467
rect 11930 14433 11940 14467
rect 11888 14424 11940 14433
rect 13728 14492 13780 14544
rect 14648 14492 14700 14544
rect 17960 14492 18012 14544
rect 12900 14467 12952 14476
rect 12900 14433 12909 14467
rect 12909 14433 12943 14467
rect 12943 14433 12952 14467
rect 12900 14424 12952 14433
rect 12992 14467 13044 14476
rect 12992 14433 13002 14467
rect 13002 14433 13036 14467
rect 13036 14433 13044 14467
rect 12992 14424 13044 14433
rect 14280 14424 14332 14476
rect 12256 14356 12308 14408
rect 12900 14288 12952 14340
rect 13912 14288 13964 14340
rect 15200 14356 15252 14408
rect 15752 14424 15804 14476
rect 15936 14424 15988 14476
rect 16396 14467 16448 14476
rect 16396 14433 16405 14467
rect 16405 14433 16439 14467
rect 16439 14433 16448 14467
rect 16396 14424 16448 14433
rect 16580 14424 16632 14476
rect 16948 14424 17000 14476
rect 14648 14288 14700 14340
rect 16304 14399 16356 14408
rect 16304 14365 16313 14399
rect 16313 14365 16347 14399
rect 16347 14365 16356 14399
rect 16304 14356 16356 14365
rect 17960 14356 18012 14408
rect 17500 14288 17552 14340
rect 10048 14263 10100 14272
rect 10048 14229 10057 14263
rect 10057 14229 10091 14263
rect 10091 14229 10100 14263
rect 10048 14220 10100 14229
rect 11336 14220 11388 14272
rect 13544 14263 13596 14272
rect 13544 14229 13553 14263
rect 13553 14229 13587 14263
rect 13587 14229 13596 14263
rect 13544 14220 13596 14229
rect 15292 14220 15344 14272
rect 15752 14220 15804 14272
rect 16120 14220 16172 14272
rect 1556 14118 1608 14170
rect 1620 14118 1672 14170
rect 1684 14118 1736 14170
rect 1748 14118 1800 14170
rect 1812 14118 1864 14170
rect 4656 14118 4708 14170
rect 4720 14118 4772 14170
rect 4784 14118 4836 14170
rect 4848 14118 4900 14170
rect 4912 14118 4964 14170
rect 7756 14118 7808 14170
rect 7820 14118 7872 14170
rect 7884 14118 7936 14170
rect 7948 14118 8000 14170
rect 8012 14118 8064 14170
rect 10856 14118 10908 14170
rect 10920 14118 10972 14170
rect 10984 14118 11036 14170
rect 11048 14118 11100 14170
rect 11112 14118 11164 14170
rect 13956 14118 14008 14170
rect 14020 14118 14072 14170
rect 14084 14118 14136 14170
rect 14148 14118 14200 14170
rect 14212 14118 14264 14170
rect 17056 14118 17108 14170
rect 17120 14118 17172 14170
rect 17184 14118 17236 14170
rect 17248 14118 17300 14170
rect 17312 14118 17364 14170
rect 3884 14016 3936 14068
rect 5632 14016 5684 14068
rect 6920 14016 6972 14068
rect 3148 13948 3200 14000
rect 8208 14016 8260 14068
rect 5724 13880 5776 13932
rect 9128 13880 9180 13932
rect 10048 13880 10100 13932
rect 13820 14016 13872 14068
rect 14280 14059 14332 14068
rect 14280 14025 14289 14059
rect 14289 14025 14323 14059
rect 14323 14025 14332 14059
rect 14280 14016 14332 14025
rect 15200 14059 15252 14068
rect 15200 14025 15209 14059
rect 15209 14025 15243 14059
rect 15243 14025 15252 14059
rect 15200 14016 15252 14025
rect 17960 14059 18012 14068
rect 2228 13812 2280 13864
rect 5632 13812 5684 13864
rect 7748 13855 7800 13864
rect 7748 13821 7757 13855
rect 7757 13821 7791 13855
rect 7791 13821 7800 13855
rect 8300 13855 8352 13864
rect 7748 13812 7800 13821
rect 8300 13821 8309 13855
rect 8309 13821 8343 13855
rect 8343 13821 8352 13855
rect 8300 13812 8352 13821
rect 13544 13812 13596 13864
rect 14372 13880 14424 13932
rect 17960 14025 17969 14059
rect 17969 14025 18003 14059
rect 18003 14025 18012 14059
rect 17960 14016 18012 14025
rect 18052 13948 18104 14000
rect 18236 13880 18288 13932
rect 14740 13855 14792 13864
rect 14740 13821 14749 13855
rect 14749 13821 14783 13855
rect 14783 13821 14792 13855
rect 14740 13812 14792 13821
rect 15844 13812 15896 13864
rect 16212 13855 16264 13864
rect 16212 13821 16221 13855
rect 16221 13821 16255 13855
rect 16255 13821 16264 13855
rect 16212 13812 16264 13821
rect 17592 13812 17644 13864
rect 2964 13676 3016 13728
rect 8392 13744 8444 13796
rect 9680 13676 9732 13728
rect 11244 13719 11296 13728
rect 11244 13685 11253 13719
rect 11253 13685 11287 13719
rect 11287 13685 11296 13719
rect 11244 13676 11296 13685
rect 3106 13574 3158 13626
rect 3170 13574 3222 13626
rect 3234 13574 3286 13626
rect 3298 13574 3350 13626
rect 3362 13574 3414 13626
rect 6206 13574 6258 13626
rect 6270 13574 6322 13626
rect 6334 13574 6386 13626
rect 6398 13574 6450 13626
rect 6462 13574 6514 13626
rect 9306 13574 9358 13626
rect 9370 13574 9422 13626
rect 9434 13574 9486 13626
rect 9498 13574 9550 13626
rect 9562 13574 9614 13626
rect 12406 13574 12458 13626
rect 12470 13574 12522 13626
rect 12534 13574 12586 13626
rect 12598 13574 12650 13626
rect 12662 13574 12714 13626
rect 15506 13574 15558 13626
rect 15570 13574 15622 13626
rect 15634 13574 15686 13626
rect 15698 13574 15750 13626
rect 15762 13574 15814 13626
rect 18606 13574 18658 13626
rect 18670 13574 18722 13626
rect 18734 13574 18786 13626
rect 18798 13574 18850 13626
rect 18862 13574 18914 13626
rect 2320 13404 2372 13456
rect 572 13379 624 13388
rect 572 13345 581 13379
rect 581 13345 615 13379
rect 615 13345 624 13379
rect 572 13336 624 13345
rect 940 13311 992 13320
rect 940 13277 949 13311
rect 949 13277 983 13311
rect 983 13277 992 13311
rect 940 13268 992 13277
rect 2228 13336 2280 13388
rect 5172 13472 5224 13524
rect 5724 13472 5776 13524
rect 8392 13472 8444 13524
rect 6644 13404 6696 13456
rect 4528 13379 4580 13388
rect 4528 13345 4537 13379
rect 4537 13345 4571 13379
rect 4571 13345 4580 13379
rect 4528 13336 4580 13345
rect 5632 13336 5684 13388
rect 2780 13268 2832 13320
rect 6736 13311 6788 13320
rect 6736 13277 6745 13311
rect 6745 13277 6779 13311
rect 6779 13277 6788 13311
rect 6736 13268 6788 13277
rect 7748 13404 7800 13456
rect 9956 13336 10008 13388
rect 10232 13379 10284 13388
rect 10232 13345 10241 13379
rect 10241 13345 10275 13379
rect 10275 13345 10284 13379
rect 10232 13336 10284 13345
rect 11612 13336 11664 13388
rect 7656 13268 7708 13320
rect 8944 13268 8996 13320
rect 9312 13311 9364 13320
rect 9312 13277 9321 13311
rect 9321 13277 9355 13311
rect 9355 13277 9364 13311
rect 9312 13268 9364 13277
rect 10508 13311 10560 13320
rect 10508 13277 10517 13311
rect 10517 13277 10551 13311
rect 10551 13277 10560 13311
rect 10508 13268 10560 13277
rect 13820 13472 13872 13524
rect 14924 13472 14976 13524
rect 15016 13447 15068 13456
rect 15016 13413 15025 13447
rect 15025 13413 15059 13447
rect 15059 13413 15068 13447
rect 15016 13404 15068 13413
rect 16212 13472 16264 13524
rect 16580 13404 16632 13456
rect 14372 13379 14424 13388
rect 14372 13345 14381 13379
rect 14381 13345 14415 13379
rect 14415 13345 14424 13379
rect 14372 13336 14424 13345
rect 17684 13379 17736 13388
rect 17684 13345 17693 13379
rect 17693 13345 17727 13379
rect 17727 13345 17736 13379
rect 17684 13336 17736 13345
rect 17592 13268 17644 13320
rect 10232 13132 10284 13184
rect 12440 13132 12492 13184
rect 14740 13132 14792 13184
rect 17408 13132 17460 13184
rect 1556 13030 1608 13082
rect 1620 13030 1672 13082
rect 1684 13030 1736 13082
rect 1748 13030 1800 13082
rect 1812 13030 1864 13082
rect 4656 13030 4708 13082
rect 4720 13030 4772 13082
rect 4784 13030 4836 13082
rect 4848 13030 4900 13082
rect 4912 13030 4964 13082
rect 7756 13030 7808 13082
rect 7820 13030 7872 13082
rect 7884 13030 7936 13082
rect 7948 13030 8000 13082
rect 8012 13030 8064 13082
rect 10856 13030 10908 13082
rect 10920 13030 10972 13082
rect 10984 13030 11036 13082
rect 11048 13030 11100 13082
rect 11112 13030 11164 13082
rect 13956 13030 14008 13082
rect 14020 13030 14072 13082
rect 14084 13030 14136 13082
rect 14148 13030 14200 13082
rect 14212 13030 14264 13082
rect 17056 13030 17108 13082
rect 17120 13030 17172 13082
rect 17184 13030 17236 13082
rect 17248 13030 17300 13082
rect 17312 13030 17364 13082
rect 940 12928 992 12980
rect 11336 12928 11388 12980
rect 15936 12928 15988 12980
rect 16396 12928 16448 12980
rect 16488 12928 16540 12980
rect 16948 12928 17000 12980
rect 8944 12860 8996 12912
rect 12532 12860 12584 12912
rect 12716 12860 12768 12912
rect 18144 12860 18196 12912
rect 2136 12835 2188 12844
rect 2136 12801 2145 12835
rect 2145 12801 2179 12835
rect 2179 12801 2188 12835
rect 2136 12792 2188 12801
rect 2964 12792 3016 12844
rect 3516 12792 3568 12844
rect 7472 12792 7524 12844
rect 7656 12792 7708 12844
rect 12440 12792 12492 12844
rect 2228 12724 2280 12776
rect 5172 12724 5224 12776
rect 7012 12724 7064 12776
rect 11152 12767 11204 12776
rect 11152 12733 11161 12767
rect 11161 12733 11195 12767
rect 11195 12733 11204 12767
rect 11152 12724 11204 12733
rect 12532 12767 12584 12776
rect 12532 12733 12541 12767
rect 12541 12733 12575 12767
rect 12575 12733 12584 12767
rect 12532 12724 12584 12733
rect 12992 12792 13044 12844
rect 17408 12792 17460 12844
rect 12900 12724 12952 12776
rect 14004 12724 14056 12776
rect 14648 12767 14700 12776
rect 14648 12733 14657 12767
rect 14657 12733 14691 12767
rect 14691 12733 14700 12767
rect 14648 12724 14700 12733
rect 14832 12767 14884 12776
rect 14832 12733 14841 12767
rect 14841 12733 14875 12767
rect 14875 12733 14884 12767
rect 14832 12724 14884 12733
rect 15936 12724 15988 12776
rect 3700 12656 3752 12708
rect 4988 12656 5040 12708
rect 6736 12656 6788 12708
rect 5816 12631 5868 12640
rect 5816 12597 5825 12631
rect 5825 12597 5859 12631
rect 5859 12597 5868 12631
rect 5816 12588 5868 12597
rect 8116 12588 8168 12640
rect 10508 12656 10560 12708
rect 16120 12724 16172 12776
rect 16304 12724 16356 12776
rect 17500 12767 17552 12776
rect 17500 12733 17509 12767
rect 17509 12733 17543 12767
rect 17543 12733 17552 12767
rect 17500 12724 17552 12733
rect 12532 12588 12584 12640
rect 12808 12588 12860 12640
rect 12992 12588 13044 12640
rect 16672 12656 16724 12708
rect 18328 12656 18380 12708
rect 3106 12486 3158 12538
rect 3170 12486 3222 12538
rect 3234 12486 3286 12538
rect 3298 12486 3350 12538
rect 3362 12486 3414 12538
rect 6206 12486 6258 12538
rect 6270 12486 6322 12538
rect 6334 12486 6386 12538
rect 6398 12486 6450 12538
rect 6462 12486 6514 12538
rect 9306 12486 9358 12538
rect 9370 12486 9422 12538
rect 9434 12486 9486 12538
rect 9498 12486 9550 12538
rect 9562 12486 9614 12538
rect 12406 12486 12458 12538
rect 12470 12486 12522 12538
rect 12534 12486 12586 12538
rect 12598 12486 12650 12538
rect 12662 12486 12714 12538
rect 15506 12486 15558 12538
rect 15570 12486 15622 12538
rect 15634 12486 15686 12538
rect 15698 12486 15750 12538
rect 15762 12486 15814 12538
rect 18606 12486 18658 12538
rect 18670 12486 18722 12538
rect 18734 12486 18786 12538
rect 18798 12486 18850 12538
rect 18862 12486 18914 12538
rect 8024 12384 8076 12436
rect 9496 12384 9548 12436
rect 2780 12248 2832 12300
rect 3608 12291 3660 12300
rect 3608 12257 3642 12291
rect 3642 12257 3660 12291
rect 3608 12248 3660 12257
rect 5264 12291 5316 12300
rect 5264 12257 5273 12291
rect 5273 12257 5307 12291
rect 5307 12257 5316 12291
rect 5264 12248 5316 12257
rect 5816 12316 5868 12368
rect 12900 12384 12952 12436
rect 14188 12384 14240 12436
rect 14648 12384 14700 12436
rect 15568 12384 15620 12436
rect 18512 12384 18564 12436
rect 5540 12180 5592 12232
rect 11888 12316 11940 12368
rect 14004 12316 14056 12368
rect 15016 12316 15068 12368
rect 16304 12359 16356 12368
rect 16304 12325 16313 12359
rect 16313 12325 16347 12359
rect 16347 12325 16356 12359
rect 16304 12316 16356 12325
rect 16672 12359 16724 12368
rect 16672 12325 16681 12359
rect 16681 12325 16715 12359
rect 16715 12325 16724 12359
rect 16672 12316 16724 12325
rect 16948 12316 17000 12368
rect 17592 12359 17644 12368
rect 17592 12325 17601 12359
rect 17601 12325 17635 12359
rect 17635 12325 17644 12359
rect 17592 12316 17644 12325
rect 9128 12248 9180 12300
rect 9312 12248 9364 12300
rect 9680 12180 9732 12232
rect 12808 12248 12860 12300
rect 13728 12291 13780 12300
rect 13728 12257 13737 12291
rect 13737 12257 13771 12291
rect 13771 12257 13780 12291
rect 13728 12248 13780 12257
rect 16212 12248 16264 12300
rect 14004 12223 14056 12232
rect 14004 12189 14013 12223
rect 14013 12189 14047 12223
rect 14047 12189 14056 12223
rect 14004 12180 14056 12189
rect 11336 12112 11388 12164
rect 14188 12223 14240 12232
rect 14188 12189 14196 12223
rect 14196 12189 14230 12223
rect 14230 12189 14240 12223
rect 14188 12180 14240 12189
rect 14280 12112 14332 12164
rect 15016 12223 15068 12232
rect 15016 12189 15025 12223
rect 15025 12189 15059 12223
rect 15059 12189 15068 12223
rect 15016 12180 15068 12189
rect 15200 12223 15252 12232
rect 15200 12189 15209 12223
rect 15209 12189 15243 12223
rect 15243 12189 15252 12223
rect 15936 12223 15988 12232
rect 15200 12180 15252 12189
rect 15936 12189 15945 12223
rect 15945 12189 15979 12223
rect 15979 12189 15988 12223
rect 15936 12180 15988 12189
rect 1952 12087 2004 12096
rect 1952 12053 1961 12087
rect 1961 12053 1995 12087
rect 1995 12053 2004 12087
rect 1952 12044 2004 12053
rect 6736 12044 6788 12096
rect 8852 12044 8904 12096
rect 12900 12044 12952 12096
rect 14004 12044 14056 12096
rect 15108 12112 15160 12164
rect 14464 12044 14516 12096
rect 16396 12044 16448 12096
rect 17868 12248 17920 12300
rect 18420 12291 18472 12300
rect 18420 12257 18429 12291
rect 18429 12257 18463 12291
rect 18463 12257 18472 12291
rect 18420 12248 18472 12257
rect 18236 12155 18288 12164
rect 18236 12121 18245 12155
rect 18245 12121 18279 12155
rect 18279 12121 18288 12155
rect 18236 12112 18288 12121
rect 1556 11942 1608 11994
rect 1620 11942 1672 11994
rect 1684 11942 1736 11994
rect 1748 11942 1800 11994
rect 1812 11942 1864 11994
rect 4656 11942 4708 11994
rect 4720 11942 4772 11994
rect 4784 11942 4836 11994
rect 4848 11942 4900 11994
rect 4912 11942 4964 11994
rect 7756 11942 7808 11994
rect 7820 11942 7872 11994
rect 7884 11942 7936 11994
rect 7948 11942 8000 11994
rect 8012 11942 8064 11994
rect 10856 11942 10908 11994
rect 10920 11942 10972 11994
rect 10984 11942 11036 11994
rect 11048 11942 11100 11994
rect 11112 11942 11164 11994
rect 13956 11942 14008 11994
rect 14020 11942 14072 11994
rect 14084 11942 14136 11994
rect 14148 11942 14200 11994
rect 14212 11942 14264 11994
rect 17056 11942 17108 11994
rect 17120 11942 17172 11994
rect 17184 11942 17236 11994
rect 17248 11942 17300 11994
rect 17312 11942 17364 11994
rect 1952 11840 2004 11892
rect 7564 11840 7616 11892
rect 14280 11840 14332 11892
rect 15200 11840 15252 11892
rect 7472 11772 7524 11824
rect 2044 11636 2096 11688
rect 12900 11747 12952 11756
rect 7104 11679 7156 11688
rect 7104 11645 7113 11679
rect 7113 11645 7147 11679
rect 7147 11645 7156 11679
rect 7104 11636 7156 11645
rect 7380 11679 7432 11688
rect 2320 11568 2372 11620
rect 7380 11645 7389 11679
rect 7389 11645 7423 11679
rect 7423 11645 7432 11679
rect 7380 11636 7432 11645
rect 8024 11679 8076 11688
rect 8024 11645 8033 11679
rect 8033 11645 8067 11679
rect 8067 11645 8076 11679
rect 8024 11636 8076 11645
rect 8208 11679 8260 11688
rect 8208 11645 8217 11679
rect 8217 11645 8251 11679
rect 8251 11645 8260 11679
rect 8208 11636 8260 11645
rect 8300 11636 8352 11688
rect 7472 11568 7524 11620
rect 7656 11568 7708 11620
rect 1676 11500 1728 11552
rect 2228 11500 2280 11552
rect 4528 11543 4580 11552
rect 4528 11509 4537 11543
rect 4537 11509 4571 11543
rect 4571 11509 4580 11543
rect 4528 11500 4580 11509
rect 7012 11500 7064 11552
rect 8852 11636 8904 11688
rect 9496 11568 9548 11620
rect 12900 11713 12909 11747
rect 12909 11713 12943 11747
rect 12943 11713 12952 11747
rect 12900 11704 12952 11713
rect 16580 11747 16632 11756
rect 12808 11679 12860 11688
rect 12808 11645 12817 11679
rect 12817 11645 12851 11679
rect 12851 11645 12860 11679
rect 12808 11636 12860 11645
rect 14188 11636 14240 11688
rect 15292 11636 15344 11688
rect 15568 11679 15620 11688
rect 15568 11645 15577 11679
rect 15577 11645 15611 11679
rect 15611 11645 15620 11679
rect 15568 11636 15620 11645
rect 16580 11713 16589 11747
rect 16589 11713 16623 11747
rect 16623 11713 16632 11747
rect 16580 11704 16632 11713
rect 15384 11568 15436 11620
rect 16948 11568 17000 11620
rect 9220 11500 9272 11552
rect 9772 11500 9824 11552
rect 11796 11500 11848 11552
rect 14188 11500 14240 11552
rect 14372 11500 14424 11552
rect 14740 11500 14792 11552
rect 17776 11500 17828 11552
rect 18420 11543 18472 11552
rect 18420 11509 18429 11543
rect 18429 11509 18463 11543
rect 18463 11509 18472 11543
rect 18420 11500 18472 11509
rect 3106 11398 3158 11450
rect 3170 11398 3222 11450
rect 3234 11398 3286 11450
rect 3298 11398 3350 11450
rect 3362 11398 3414 11450
rect 6206 11398 6258 11450
rect 6270 11398 6322 11450
rect 6334 11398 6386 11450
rect 6398 11398 6450 11450
rect 6462 11398 6514 11450
rect 9306 11398 9358 11450
rect 9370 11398 9422 11450
rect 9434 11398 9486 11450
rect 9498 11398 9550 11450
rect 9562 11398 9614 11450
rect 12406 11398 12458 11450
rect 12470 11398 12522 11450
rect 12534 11398 12586 11450
rect 12598 11398 12650 11450
rect 12662 11398 12714 11450
rect 15506 11398 15558 11450
rect 15570 11398 15622 11450
rect 15634 11398 15686 11450
rect 15698 11398 15750 11450
rect 15762 11398 15814 11450
rect 18606 11398 18658 11450
rect 18670 11398 18722 11450
rect 18734 11398 18786 11450
rect 18798 11398 18850 11450
rect 18862 11398 18914 11450
rect 1676 11339 1728 11348
rect 1676 11305 1685 11339
rect 1685 11305 1719 11339
rect 1719 11305 1728 11339
rect 1676 11296 1728 11305
rect 2044 11339 2096 11348
rect 2044 11305 2053 11339
rect 2053 11305 2087 11339
rect 2087 11305 2096 11339
rect 2044 11296 2096 11305
rect 5540 11339 5592 11348
rect 5540 11305 5549 11339
rect 5549 11305 5583 11339
rect 5583 11305 5592 11339
rect 5540 11296 5592 11305
rect 8300 11339 8352 11348
rect 8300 11305 8309 11339
rect 8309 11305 8343 11339
rect 8343 11305 8352 11339
rect 8300 11296 8352 11305
rect 3792 11203 3844 11212
rect 3792 11169 3801 11203
rect 3801 11169 3835 11203
rect 3835 11169 3844 11203
rect 3792 11160 3844 11169
rect 4068 11160 4120 11212
rect 8024 11228 8076 11280
rect 9036 11228 9088 11280
rect 11612 11228 11664 11280
rect 2688 11092 2740 11144
rect 3608 11092 3660 11144
rect 5264 11203 5316 11212
rect 5264 11169 5274 11203
rect 5274 11169 5308 11203
rect 5308 11169 5316 11203
rect 5264 11160 5316 11169
rect 9772 11160 9824 11212
rect 9956 11203 10008 11212
rect 9956 11169 9965 11203
rect 9965 11169 9999 11203
rect 9999 11169 10008 11203
rect 9956 11160 10008 11169
rect 14648 11228 14700 11280
rect 16120 11228 16172 11280
rect 14464 11160 14516 11212
rect 14740 11203 14792 11212
rect 14740 11169 14749 11203
rect 14749 11169 14783 11203
rect 14783 11169 14792 11203
rect 14740 11160 14792 11169
rect 16948 11160 17000 11212
rect 17776 11203 17828 11212
rect 10232 11135 10284 11144
rect 10232 11101 10241 11135
rect 10241 11101 10275 11135
rect 10275 11101 10284 11135
rect 10232 11092 10284 11101
rect 17776 11169 17785 11203
rect 17785 11169 17819 11203
rect 17819 11169 17828 11203
rect 17776 11160 17828 11169
rect 2136 11024 2188 11076
rect 17500 11024 17552 11076
rect 3148 10956 3200 11008
rect 11520 10956 11572 11008
rect 15568 10956 15620 11008
rect 15936 10956 15988 11008
rect 17408 10956 17460 11008
rect 1556 10854 1608 10906
rect 1620 10854 1672 10906
rect 1684 10854 1736 10906
rect 1748 10854 1800 10906
rect 1812 10854 1864 10906
rect 4656 10854 4708 10906
rect 4720 10854 4772 10906
rect 4784 10854 4836 10906
rect 4848 10854 4900 10906
rect 4912 10854 4964 10906
rect 7756 10854 7808 10906
rect 7820 10854 7872 10906
rect 7884 10854 7936 10906
rect 7948 10854 8000 10906
rect 8012 10854 8064 10906
rect 10856 10854 10908 10906
rect 10920 10854 10972 10906
rect 10984 10854 11036 10906
rect 11048 10854 11100 10906
rect 11112 10854 11164 10906
rect 13956 10854 14008 10906
rect 14020 10854 14072 10906
rect 14084 10854 14136 10906
rect 14148 10854 14200 10906
rect 14212 10854 14264 10906
rect 17056 10854 17108 10906
rect 17120 10854 17172 10906
rect 17184 10854 17236 10906
rect 17248 10854 17300 10906
rect 17312 10854 17364 10906
rect 2688 10795 2740 10804
rect 2688 10761 2697 10795
rect 2697 10761 2731 10795
rect 2731 10761 2740 10795
rect 2688 10752 2740 10761
rect 6644 10752 6696 10804
rect 7656 10752 7708 10804
rect 10232 10752 10284 10804
rect 15200 10752 15252 10804
rect 16948 10795 17000 10804
rect 16948 10761 16957 10795
rect 16957 10761 16991 10795
rect 16991 10761 17000 10795
rect 16948 10752 17000 10761
rect 3700 10684 3752 10736
rect 2596 10616 2648 10668
rect 3148 10659 3200 10668
rect 3148 10625 3157 10659
rect 3157 10625 3191 10659
rect 3191 10625 3200 10659
rect 3148 10616 3200 10625
rect 2228 10548 2280 10600
rect 2688 10548 2740 10600
rect 3884 10616 3936 10668
rect 4988 10684 5040 10736
rect 6920 10616 6972 10668
rect 4252 10591 4304 10600
rect 4252 10557 4261 10591
rect 4261 10557 4295 10591
rect 4295 10557 4304 10591
rect 4252 10548 4304 10557
rect 4344 10480 4396 10532
rect 6552 10548 6604 10600
rect 6736 10591 6788 10600
rect 6736 10557 6745 10591
rect 6745 10557 6779 10591
rect 6779 10557 6788 10591
rect 11796 10659 11848 10668
rect 11796 10625 11805 10659
rect 11805 10625 11839 10659
rect 11839 10625 11848 10659
rect 11796 10616 11848 10625
rect 12808 10659 12860 10668
rect 12808 10625 12817 10659
rect 12817 10625 12851 10659
rect 12851 10625 12860 10659
rect 12808 10616 12860 10625
rect 6736 10548 6788 10557
rect 8116 10591 8168 10600
rect 8116 10557 8125 10591
rect 8125 10557 8159 10591
rect 8159 10557 8168 10591
rect 8116 10548 8168 10557
rect 11520 10591 11572 10600
rect 11520 10557 11529 10591
rect 11529 10557 11563 10591
rect 11563 10557 11572 10591
rect 11520 10548 11572 10557
rect 15568 10591 15620 10600
rect 15568 10557 15577 10591
rect 15577 10557 15611 10591
rect 15611 10557 15620 10591
rect 15568 10548 15620 10557
rect 8576 10480 8628 10532
rect 12808 10480 12860 10532
rect 4068 10455 4120 10464
rect 4068 10421 4077 10455
rect 4077 10421 4111 10455
rect 4111 10421 4120 10455
rect 4068 10412 4120 10421
rect 8116 10412 8168 10464
rect 13176 10412 13228 10464
rect 3106 10310 3158 10362
rect 3170 10310 3222 10362
rect 3234 10310 3286 10362
rect 3298 10310 3350 10362
rect 3362 10310 3414 10362
rect 6206 10310 6258 10362
rect 6270 10310 6322 10362
rect 6334 10310 6386 10362
rect 6398 10310 6450 10362
rect 6462 10310 6514 10362
rect 9306 10310 9358 10362
rect 9370 10310 9422 10362
rect 9434 10310 9486 10362
rect 9498 10310 9550 10362
rect 9562 10310 9614 10362
rect 12406 10310 12458 10362
rect 12470 10310 12522 10362
rect 12534 10310 12586 10362
rect 12598 10310 12650 10362
rect 12662 10310 12714 10362
rect 15506 10310 15558 10362
rect 15570 10310 15622 10362
rect 15634 10310 15686 10362
rect 15698 10310 15750 10362
rect 15762 10310 15814 10362
rect 18606 10310 18658 10362
rect 18670 10310 18722 10362
rect 18734 10310 18786 10362
rect 18798 10310 18850 10362
rect 18862 10310 18914 10362
rect 1400 10208 1452 10260
rect 3792 10251 3844 10260
rect 3792 10217 3801 10251
rect 3801 10217 3835 10251
rect 3835 10217 3844 10251
rect 3792 10208 3844 10217
rect 6552 10251 6604 10260
rect 6552 10217 6561 10251
rect 6561 10217 6595 10251
rect 6595 10217 6604 10251
rect 6552 10208 6604 10217
rect 7380 10208 7432 10260
rect 11888 10251 11940 10260
rect 11888 10217 11897 10251
rect 11897 10217 11931 10251
rect 11931 10217 11940 10251
rect 11888 10208 11940 10217
rect 12348 10208 12400 10260
rect 12808 10251 12860 10260
rect 12808 10217 12817 10251
rect 12817 10217 12851 10251
rect 12851 10217 12860 10251
rect 12808 10208 12860 10217
rect 8116 10183 8168 10192
rect 940 10072 992 10124
rect 3792 10115 3844 10124
rect 3792 10081 3801 10115
rect 3801 10081 3835 10115
rect 3835 10081 3844 10115
rect 3792 10072 3844 10081
rect 5356 10115 5408 10124
rect 3700 10004 3752 10056
rect 4252 10004 4304 10056
rect 5356 10081 5365 10115
rect 5365 10081 5399 10115
rect 5399 10081 5408 10115
rect 8116 10149 8125 10183
rect 8125 10149 8159 10183
rect 8159 10149 8168 10183
rect 8116 10140 8168 10149
rect 8668 10140 8720 10192
rect 17500 10183 17552 10192
rect 5356 10072 5408 10081
rect 7196 10072 7248 10124
rect 11520 10072 11572 10124
rect 12348 10115 12400 10124
rect 6552 10047 6604 10056
rect 6552 10013 6561 10047
rect 6561 10013 6595 10047
rect 6595 10013 6604 10047
rect 6552 10004 6604 10013
rect 6828 10047 6880 10056
rect 6828 10013 6837 10047
rect 6837 10013 6871 10047
rect 6871 10013 6880 10047
rect 6828 10004 6880 10013
rect 7564 10004 7616 10056
rect 12348 10081 12357 10115
rect 12357 10081 12391 10115
rect 12391 10081 12400 10115
rect 12348 10072 12400 10081
rect 17500 10149 17509 10183
rect 17509 10149 17543 10183
rect 17543 10149 17552 10183
rect 17500 10140 17552 10149
rect 13268 10115 13320 10124
rect 11980 10004 12032 10056
rect 13268 10081 13277 10115
rect 13277 10081 13311 10115
rect 13311 10081 13320 10115
rect 13268 10072 13320 10081
rect 13636 10072 13688 10124
rect 17408 10115 17460 10124
rect 17408 10081 17417 10115
rect 17417 10081 17451 10115
rect 17451 10081 17460 10115
rect 17408 10072 17460 10081
rect 17960 10072 18012 10124
rect 12900 10004 12952 10056
rect 13728 10004 13780 10056
rect 14556 10004 14608 10056
rect 7380 9936 7432 9988
rect 9128 9868 9180 9920
rect 10784 9868 10836 9920
rect 13176 9868 13228 9920
rect 16672 9868 16724 9920
rect 1556 9766 1608 9818
rect 1620 9766 1672 9818
rect 1684 9766 1736 9818
rect 1748 9766 1800 9818
rect 1812 9766 1864 9818
rect 4656 9766 4708 9818
rect 4720 9766 4772 9818
rect 4784 9766 4836 9818
rect 4848 9766 4900 9818
rect 4912 9766 4964 9818
rect 7756 9766 7808 9818
rect 7820 9766 7872 9818
rect 7884 9766 7936 9818
rect 7948 9766 8000 9818
rect 8012 9766 8064 9818
rect 10856 9766 10908 9818
rect 10920 9766 10972 9818
rect 10984 9766 11036 9818
rect 11048 9766 11100 9818
rect 11112 9766 11164 9818
rect 13956 9766 14008 9818
rect 14020 9766 14072 9818
rect 14084 9766 14136 9818
rect 14148 9766 14200 9818
rect 14212 9766 14264 9818
rect 17056 9766 17108 9818
rect 17120 9766 17172 9818
rect 17184 9766 17236 9818
rect 17248 9766 17300 9818
rect 17312 9766 17364 9818
rect 10784 9664 10836 9716
rect 4344 9596 4396 9648
rect 2136 9571 2188 9580
rect 2136 9537 2145 9571
rect 2145 9537 2179 9571
rect 2179 9537 2188 9571
rect 2136 9528 2188 9537
rect 2320 9460 2372 9512
rect 2688 9460 2740 9512
rect 4068 9528 4120 9580
rect 8208 9596 8260 9648
rect 13268 9664 13320 9716
rect 7104 9571 7156 9580
rect 7104 9537 7113 9571
rect 7113 9537 7147 9571
rect 7147 9537 7156 9571
rect 7104 9528 7156 9537
rect 17960 9639 18012 9648
rect 17960 9605 17969 9639
rect 17969 9605 18003 9639
rect 18003 9605 18012 9639
rect 17960 9596 18012 9605
rect 6828 9460 6880 9512
rect 7196 9503 7248 9512
rect 7196 9469 7205 9503
rect 7205 9469 7239 9503
rect 7239 9469 7248 9503
rect 7196 9460 7248 9469
rect 9220 9460 9272 9512
rect 10140 9503 10192 9512
rect 10140 9469 10149 9503
rect 10149 9469 10183 9503
rect 10183 9469 10192 9503
rect 10140 9460 10192 9469
rect 11980 9503 12032 9512
rect 11980 9469 11989 9503
rect 11989 9469 12023 9503
rect 12023 9469 12032 9503
rect 11980 9460 12032 9469
rect 15200 9503 15252 9512
rect 15200 9469 15209 9503
rect 15209 9469 15243 9503
rect 15243 9469 15252 9503
rect 15200 9460 15252 9469
rect 16212 9503 16264 9512
rect 16212 9469 16221 9503
rect 16221 9469 16255 9503
rect 16255 9469 16264 9503
rect 16212 9460 16264 9469
rect 16304 9460 16356 9512
rect 16856 9503 16908 9512
rect 16856 9469 16890 9503
rect 16890 9469 16908 9503
rect 16856 9460 16908 9469
rect 848 9324 900 9376
rect 2964 9367 3016 9376
rect 2964 9333 2973 9367
rect 2973 9333 3007 9367
rect 3007 9333 3016 9367
rect 2964 9324 3016 9333
rect 8576 9392 8628 9444
rect 15936 9435 15988 9444
rect 15936 9401 15945 9435
rect 15945 9401 15979 9435
rect 15979 9401 15988 9435
rect 15936 9392 15988 9401
rect 4344 9367 4396 9376
rect 4344 9333 4353 9367
rect 4353 9333 4387 9367
rect 4387 9333 4396 9367
rect 4344 9324 4396 9333
rect 7288 9324 7340 9376
rect 8668 9324 8720 9376
rect 8944 9367 8996 9376
rect 8944 9333 8953 9367
rect 8953 9333 8987 9367
rect 8987 9333 8996 9367
rect 8944 9324 8996 9333
rect 9956 9324 10008 9376
rect 12808 9324 12860 9376
rect 15108 9324 15160 9376
rect 15292 9324 15344 9376
rect 3106 9222 3158 9274
rect 3170 9222 3222 9274
rect 3234 9222 3286 9274
rect 3298 9222 3350 9274
rect 3362 9222 3414 9274
rect 6206 9222 6258 9274
rect 6270 9222 6322 9274
rect 6334 9222 6386 9274
rect 6398 9222 6450 9274
rect 6462 9222 6514 9274
rect 9306 9222 9358 9274
rect 9370 9222 9422 9274
rect 9434 9222 9486 9274
rect 9498 9222 9550 9274
rect 9562 9222 9614 9274
rect 12406 9222 12458 9274
rect 12470 9222 12522 9274
rect 12534 9222 12586 9274
rect 12598 9222 12650 9274
rect 12662 9222 12714 9274
rect 15506 9222 15558 9274
rect 15570 9222 15622 9274
rect 15634 9222 15686 9274
rect 15698 9222 15750 9274
rect 15762 9222 15814 9274
rect 18606 9222 18658 9274
rect 18670 9222 18722 9274
rect 18734 9222 18786 9274
rect 18798 9222 18850 9274
rect 18862 9222 18914 9274
rect 2320 9163 2372 9172
rect 2320 9129 2329 9163
rect 2329 9129 2363 9163
rect 2363 9129 2372 9163
rect 2320 9120 2372 9129
rect 4344 9120 4396 9172
rect 5356 9120 5408 9172
rect 7288 9120 7340 9172
rect 9220 9120 9272 9172
rect 11980 9120 12032 9172
rect 12808 9120 12860 9172
rect 18144 9120 18196 9172
rect 848 9095 900 9104
rect 848 9061 857 9095
rect 857 9061 891 9095
rect 891 9061 900 9095
rect 848 9052 900 9061
rect 2872 9052 2924 9104
rect 8668 9052 8720 9104
rect 11244 9052 11296 9104
rect 13268 9052 13320 9104
rect 13544 9052 13596 9104
rect 16120 9052 16172 9104
rect 16488 9052 16540 9104
rect 2964 8984 3016 9036
rect 3424 9027 3476 9036
rect 572 8959 624 8968
rect 572 8925 581 8959
rect 581 8925 615 8959
rect 615 8925 624 8959
rect 572 8916 624 8925
rect 3424 8993 3433 9027
rect 3433 8993 3467 9027
rect 3467 8993 3476 9027
rect 3424 8984 3476 8993
rect 7012 8984 7064 9036
rect 9956 9027 10008 9036
rect 9956 8993 9965 9027
rect 9965 8993 9999 9027
rect 9999 8993 10008 9027
rect 9956 8984 10008 8993
rect 13728 8984 13780 9036
rect 13820 8984 13872 9036
rect 15108 9027 15160 9036
rect 15108 8993 15117 9027
rect 15117 8993 15151 9027
rect 15151 8993 15160 9027
rect 15108 8984 15160 8993
rect 18420 9027 18472 9036
rect 18420 8993 18429 9027
rect 18429 8993 18463 9027
rect 18463 8993 18472 9027
rect 18420 8984 18472 8993
rect 4344 8916 4396 8968
rect 7564 8959 7616 8968
rect 4436 8848 4488 8900
rect 2872 8823 2924 8832
rect 2872 8789 2881 8823
rect 2881 8789 2915 8823
rect 2915 8789 2924 8823
rect 2872 8780 2924 8789
rect 5540 8780 5592 8832
rect 7564 8925 7573 8959
rect 7573 8925 7607 8959
rect 7607 8925 7616 8959
rect 7564 8916 7616 8925
rect 8116 8916 8168 8968
rect 10324 8959 10376 8968
rect 10324 8925 10333 8959
rect 10333 8925 10367 8959
rect 10367 8925 10376 8959
rect 10324 8916 10376 8925
rect 13084 8959 13136 8968
rect 13084 8925 13093 8959
rect 13093 8925 13127 8959
rect 13127 8925 13136 8959
rect 13084 8916 13136 8925
rect 13268 8959 13320 8968
rect 13268 8925 13277 8959
rect 13277 8925 13311 8959
rect 13311 8925 13320 8959
rect 13268 8916 13320 8925
rect 16212 8916 16264 8968
rect 13820 8848 13872 8900
rect 14740 8848 14792 8900
rect 12624 8823 12676 8832
rect 12624 8789 12633 8823
rect 12633 8789 12667 8823
rect 12667 8789 12676 8823
rect 12624 8780 12676 8789
rect 13636 8823 13688 8832
rect 13636 8789 13645 8823
rect 13645 8789 13679 8823
rect 13679 8789 13688 8823
rect 13636 8780 13688 8789
rect 1556 8678 1608 8730
rect 1620 8678 1672 8730
rect 1684 8678 1736 8730
rect 1748 8678 1800 8730
rect 1812 8678 1864 8730
rect 4656 8678 4708 8730
rect 4720 8678 4772 8730
rect 4784 8678 4836 8730
rect 4848 8678 4900 8730
rect 4912 8678 4964 8730
rect 7756 8678 7808 8730
rect 7820 8678 7872 8730
rect 7884 8678 7936 8730
rect 7948 8678 8000 8730
rect 8012 8678 8064 8730
rect 10856 8678 10908 8730
rect 10920 8678 10972 8730
rect 10984 8678 11036 8730
rect 11048 8678 11100 8730
rect 11112 8678 11164 8730
rect 13956 8678 14008 8730
rect 14020 8678 14072 8730
rect 14084 8678 14136 8730
rect 14148 8678 14200 8730
rect 14212 8678 14264 8730
rect 17056 8678 17108 8730
rect 17120 8678 17172 8730
rect 17184 8678 17236 8730
rect 17248 8678 17300 8730
rect 17312 8678 17364 8730
rect 2596 8619 2648 8628
rect 2596 8585 2605 8619
rect 2605 8585 2639 8619
rect 2639 8585 2648 8619
rect 2596 8576 2648 8585
rect 3424 8576 3476 8628
rect 6920 8619 6972 8628
rect 6920 8585 6929 8619
rect 6929 8585 6963 8619
rect 6963 8585 6972 8619
rect 6920 8576 6972 8585
rect 8116 8619 8168 8628
rect 8116 8585 8125 8619
rect 8125 8585 8159 8619
rect 8159 8585 8168 8619
rect 8116 8576 8168 8585
rect 8576 8576 8628 8628
rect 10324 8576 10376 8628
rect 13084 8576 13136 8628
rect 13820 8576 13872 8628
rect 17684 8576 17736 8628
rect 2320 8440 2372 8492
rect 8944 8508 8996 8560
rect 8208 8483 8260 8492
rect 5540 8415 5592 8424
rect 5540 8381 5549 8415
rect 5549 8381 5583 8415
rect 5583 8381 5592 8415
rect 5540 8372 5592 8381
rect 7012 8415 7064 8424
rect 7012 8381 7021 8415
rect 7021 8381 7055 8415
rect 7055 8381 7064 8415
rect 7012 8372 7064 8381
rect 7196 8372 7248 8424
rect 8208 8449 8217 8483
rect 8217 8449 8251 8483
rect 8251 8449 8260 8483
rect 8208 8440 8260 8449
rect 12624 8508 12676 8560
rect 11796 8483 11848 8492
rect 11796 8449 11805 8483
rect 11805 8449 11839 8483
rect 11839 8449 11848 8483
rect 11796 8440 11848 8449
rect 16304 8440 16356 8492
rect 8392 8372 8444 8424
rect 9128 8415 9180 8424
rect 9128 8381 9137 8415
rect 9137 8381 9171 8415
rect 9171 8381 9180 8415
rect 9128 8372 9180 8381
rect 11980 8372 12032 8424
rect 13176 8372 13228 8424
rect 13636 8372 13688 8424
rect 16580 8372 16632 8424
rect 2688 8304 2740 8356
rect 4344 8304 4396 8356
rect 5264 8347 5316 8356
rect 5264 8313 5273 8347
rect 5273 8313 5307 8347
rect 5307 8313 5316 8347
rect 5264 8304 5316 8313
rect 6552 8347 6604 8356
rect 6552 8313 6561 8347
rect 6561 8313 6595 8347
rect 6595 8313 6604 8347
rect 6552 8304 6604 8313
rect 9956 8304 10008 8356
rect 9680 8236 9732 8288
rect 10876 8236 10928 8288
rect 16488 8236 16540 8288
rect 3106 8134 3158 8186
rect 3170 8134 3222 8186
rect 3234 8134 3286 8186
rect 3298 8134 3350 8186
rect 3362 8134 3414 8186
rect 6206 8134 6258 8186
rect 6270 8134 6322 8186
rect 6334 8134 6386 8186
rect 6398 8134 6450 8186
rect 6462 8134 6514 8186
rect 9306 8134 9358 8186
rect 9370 8134 9422 8186
rect 9434 8134 9486 8186
rect 9498 8134 9550 8186
rect 9562 8134 9614 8186
rect 12406 8134 12458 8186
rect 12470 8134 12522 8186
rect 12534 8134 12586 8186
rect 12598 8134 12650 8186
rect 12662 8134 12714 8186
rect 15506 8134 15558 8186
rect 15570 8134 15622 8186
rect 15634 8134 15686 8186
rect 15698 8134 15750 8186
rect 15762 8134 15814 8186
rect 18606 8134 18658 8186
rect 18670 8134 18722 8186
rect 18734 8134 18786 8186
rect 18798 8134 18850 8186
rect 18862 8134 18914 8186
rect 2596 8032 2648 8084
rect 5448 8032 5500 8084
rect 13268 8032 13320 8084
rect 15936 8075 15988 8084
rect 2872 7964 2924 8016
rect 4528 8007 4580 8016
rect 4528 7973 4537 8007
rect 4537 7973 4571 8007
rect 4571 7973 4580 8007
rect 4528 7964 4580 7973
rect 7288 7964 7340 8016
rect 9772 7964 9824 8016
rect 11244 7964 11296 8016
rect 14372 8007 14424 8016
rect 14372 7973 14381 8007
rect 14381 7973 14415 8007
rect 14415 7973 14424 8007
rect 14372 7964 14424 7973
rect 5264 7896 5316 7948
rect 6920 7896 6972 7948
rect 572 7828 624 7880
rect 940 7871 992 7880
rect 940 7837 949 7871
rect 949 7837 983 7871
rect 983 7837 992 7871
rect 940 7828 992 7837
rect 5724 7828 5776 7880
rect 7380 7828 7432 7880
rect 8116 7871 8168 7880
rect 8116 7837 8125 7871
rect 8125 7837 8159 7871
rect 8159 7837 8168 7871
rect 8116 7828 8168 7837
rect 7472 7760 7524 7812
rect 7656 7760 7708 7812
rect 8392 7896 8444 7948
rect 8760 7896 8812 7948
rect 10876 7939 10928 7948
rect 10876 7905 10885 7939
rect 10885 7905 10919 7939
rect 10919 7905 10928 7939
rect 10876 7896 10928 7905
rect 15200 7896 15252 7948
rect 15936 8041 15945 8075
rect 15945 8041 15979 8075
rect 15979 8041 15988 8075
rect 15936 8032 15988 8041
rect 16580 8075 16632 8084
rect 16580 8041 16589 8075
rect 16589 8041 16623 8075
rect 16623 8041 16632 8075
rect 16580 8032 16632 8041
rect 17684 8032 17736 8084
rect 15844 7964 15896 8016
rect 16580 7939 16632 7948
rect 16580 7905 16589 7939
rect 16589 7905 16623 7939
rect 16623 7905 16632 7939
rect 16580 7896 16632 7905
rect 16672 7828 16724 7880
rect 17316 7871 17368 7880
rect 17316 7837 17325 7871
rect 17325 7837 17359 7871
rect 17359 7837 17368 7871
rect 17316 7828 17368 7837
rect 17776 7828 17828 7880
rect 9220 7760 9272 7812
rect 15384 7760 15436 7812
rect 6828 7692 6880 7744
rect 13820 7692 13872 7744
rect 14740 7735 14792 7744
rect 14740 7701 14749 7735
rect 14749 7701 14783 7735
rect 14783 7701 14792 7735
rect 14740 7692 14792 7701
rect 1556 7590 1608 7642
rect 1620 7590 1672 7642
rect 1684 7590 1736 7642
rect 1748 7590 1800 7642
rect 1812 7590 1864 7642
rect 4656 7590 4708 7642
rect 4720 7590 4772 7642
rect 4784 7590 4836 7642
rect 4848 7590 4900 7642
rect 4912 7590 4964 7642
rect 7756 7590 7808 7642
rect 7820 7590 7872 7642
rect 7884 7590 7936 7642
rect 7948 7590 8000 7642
rect 8012 7590 8064 7642
rect 10856 7590 10908 7642
rect 10920 7590 10972 7642
rect 10984 7590 11036 7642
rect 11048 7590 11100 7642
rect 11112 7590 11164 7642
rect 13956 7590 14008 7642
rect 14020 7590 14072 7642
rect 14084 7590 14136 7642
rect 14148 7590 14200 7642
rect 14212 7590 14264 7642
rect 17056 7590 17108 7642
rect 17120 7590 17172 7642
rect 17184 7590 17236 7642
rect 17248 7590 17300 7642
rect 17312 7590 17364 7642
rect 940 7488 992 7540
rect 4252 7488 4304 7540
rect 2136 7395 2188 7404
rect 2136 7361 2145 7395
rect 2145 7361 2179 7395
rect 2179 7361 2188 7395
rect 2136 7352 2188 7361
rect 2780 7352 2832 7404
rect 3792 7352 3844 7404
rect 8116 7488 8168 7540
rect 8944 7463 8996 7472
rect 8944 7429 8953 7463
rect 8953 7429 8987 7463
rect 8987 7429 8996 7463
rect 8944 7420 8996 7429
rect 9220 7463 9272 7472
rect 9220 7429 9229 7463
rect 9229 7429 9263 7463
rect 9263 7429 9272 7463
rect 9220 7420 9272 7429
rect 8392 7352 8444 7404
rect 10416 7488 10468 7540
rect 11244 7488 11296 7540
rect 12256 7488 12308 7540
rect 11796 7395 11848 7404
rect 11796 7361 11805 7395
rect 11805 7361 11839 7395
rect 11839 7361 11848 7395
rect 11796 7352 11848 7361
rect 13268 7352 13320 7404
rect 14740 7352 14792 7404
rect 2596 7284 2648 7336
rect 3608 7284 3660 7336
rect 4344 7327 4396 7336
rect 4344 7293 4353 7327
rect 4353 7293 4387 7327
rect 4387 7293 4396 7327
rect 4344 7284 4396 7293
rect 6828 7327 6880 7336
rect 6828 7293 6837 7327
rect 6837 7293 6871 7327
rect 6871 7293 6880 7327
rect 6828 7284 6880 7293
rect 8300 7284 8352 7336
rect 9956 7327 10008 7336
rect 9956 7293 9965 7327
rect 9965 7293 9999 7327
rect 9999 7293 10008 7327
rect 9956 7284 10008 7293
rect 10784 7327 10836 7336
rect 10784 7293 10793 7327
rect 10793 7293 10827 7327
rect 10827 7293 10836 7327
rect 10784 7284 10836 7293
rect 11888 7284 11940 7336
rect 2872 7148 2924 7200
rect 5816 7216 5868 7268
rect 5908 7148 5960 7200
rect 12900 7284 12952 7336
rect 13820 7327 13872 7336
rect 13820 7293 13829 7327
rect 13829 7293 13863 7327
rect 13863 7293 13872 7327
rect 13820 7284 13872 7293
rect 15844 7488 15896 7540
rect 16580 7488 16632 7540
rect 15844 7352 15896 7404
rect 15936 7327 15988 7336
rect 15936 7293 15945 7327
rect 15945 7293 15979 7327
rect 15979 7293 15988 7327
rect 15936 7284 15988 7293
rect 17408 7327 17460 7336
rect 17408 7293 17417 7327
rect 17417 7293 17451 7327
rect 17451 7293 17460 7327
rect 17408 7284 17460 7293
rect 16488 7216 16540 7268
rect 17684 7284 17736 7336
rect 17776 7216 17828 7268
rect 10784 7148 10836 7200
rect 11152 7191 11204 7200
rect 11152 7157 11161 7191
rect 11161 7157 11195 7191
rect 11195 7157 11204 7191
rect 11152 7148 11204 7157
rect 12808 7148 12860 7200
rect 15016 7148 15068 7200
rect 15844 7148 15896 7200
rect 16028 7191 16080 7200
rect 16028 7157 16037 7191
rect 16037 7157 16071 7191
rect 16071 7157 16080 7191
rect 16028 7148 16080 7157
rect 3106 7046 3158 7098
rect 3170 7046 3222 7098
rect 3234 7046 3286 7098
rect 3298 7046 3350 7098
rect 3362 7046 3414 7098
rect 6206 7046 6258 7098
rect 6270 7046 6322 7098
rect 6334 7046 6386 7098
rect 6398 7046 6450 7098
rect 6462 7046 6514 7098
rect 9306 7046 9358 7098
rect 9370 7046 9422 7098
rect 9434 7046 9486 7098
rect 9498 7046 9550 7098
rect 9562 7046 9614 7098
rect 12406 7046 12458 7098
rect 12470 7046 12522 7098
rect 12534 7046 12586 7098
rect 12598 7046 12650 7098
rect 12662 7046 12714 7098
rect 15506 7046 15558 7098
rect 15570 7046 15622 7098
rect 15634 7046 15686 7098
rect 15698 7046 15750 7098
rect 15762 7046 15814 7098
rect 18606 7046 18658 7098
rect 18670 7046 18722 7098
rect 18734 7046 18786 7098
rect 18798 7046 18850 7098
rect 18862 7046 18914 7098
rect 11888 6987 11940 6996
rect 11888 6953 11897 6987
rect 11897 6953 11931 6987
rect 11931 6953 11940 6987
rect 11888 6944 11940 6953
rect 15200 6944 15252 6996
rect 572 6876 624 6928
rect 4252 6876 4304 6928
rect 11428 6876 11480 6928
rect 4160 6808 4212 6860
rect 5264 6851 5316 6860
rect 5264 6817 5273 6851
rect 5273 6817 5307 6851
rect 5307 6817 5316 6851
rect 5264 6808 5316 6817
rect 5816 6808 5868 6860
rect 10140 6851 10192 6860
rect 10140 6817 10149 6851
rect 10149 6817 10183 6851
rect 10183 6817 10192 6851
rect 10140 6808 10192 6817
rect 13820 6876 13872 6928
rect 13544 6808 13596 6860
rect 5724 6672 5776 6724
rect 15936 6876 15988 6928
rect 16028 6808 16080 6860
rect 18420 6851 18472 6860
rect 18420 6817 18429 6851
rect 18429 6817 18463 6851
rect 18463 6817 18472 6851
rect 18420 6808 18472 6817
rect 1952 6647 2004 6656
rect 1952 6613 1961 6647
rect 1961 6613 1995 6647
rect 1995 6613 2004 6647
rect 1952 6604 2004 6613
rect 5632 6647 5684 6656
rect 5632 6613 5641 6647
rect 5641 6613 5675 6647
rect 5675 6613 5684 6647
rect 5632 6604 5684 6613
rect 11152 6604 11204 6656
rect 13544 6604 13596 6656
rect 14556 6740 14608 6792
rect 15016 6740 15068 6792
rect 15384 6783 15436 6792
rect 15384 6749 15393 6783
rect 15393 6749 15427 6783
rect 15427 6749 15436 6783
rect 15384 6740 15436 6749
rect 15292 6604 15344 6656
rect 1556 6502 1608 6554
rect 1620 6502 1672 6554
rect 1684 6502 1736 6554
rect 1748 6502 1800 6554
rect 1812 6502 1864 6554
rect 4656 6502 4708 6554
rect 4720 6502 4772 6554
rect 4784 6502 4836 6554
rect 4848 6502 4900 6554
rect 4912 6502 4964 6554
rect 7756 6502 7808 6554
rect 7820 6502 7872 6554
rect 7884 6502 7936 6554
rect 7948 6502 8000 6554
rect 8012 6502 8064 6554
rect 10856 6502 10908 6554
rect 10920 6502 10972 6554
rect 10984 6502 11036 6554
rect 11048 6502 11100 6554
rect 11112 6502 11164 6554
rect 13956 6502 14008 6554
rect 14020 6502 14072 6554
rect 14084 6502 14136 6554
rect 14148 6502 14200 6554
rect 14212 6502 14264 6554
rect 17056 6502 17108 6554
rect 17120 6502 17172 6554
rect 17184 6502 17236 6554
rect 17248 6502 17300 6554
rect 17312 6502 17364 6554
rect 1952 6400 2004 6452
rect 9036 6400 9088 6452
rect 12808 6400 12860 6452
rect 13728 6400 13780 6452
rect 14556 6443 14608 6452
rect 14556 6409 14565 6443
rect 14565 6409 14599 6443
rect 14599 6409 14608 6443
rect 14556 6400 14608 6409
rect 15292 6332 15344 6384
rect 2964 6264 3016 6316
rect 4252 6307 4304 6316
rect 4252 6273 4261 6307
rect 4261 6273 4295 6307
rect 4295 6273 4304 6307
rect 4252 6264 4304 6273
rect 5540 6264 5592 6316
rect 16856 6400 16908 6452
rect 16212 6264 16264 6316
rect 6736 6239 6788 6248
rect 6736 6205 6745 6239
rect 6745 6205 6779 6239
rect 6779 6205 6788 6239
rect 6736 6196 6788 6205
rect 8760 6239 8812 6248
rect 8760 6205 8769 6239
rect 8769 6205 8803 6239
rect 8803 6205 8812 6239
rect 8760 6196 8812 6205
rect 13728 6196 13780 6248
rect 14740 6196 14792 6248
rect 16304 6239 16356 6248
rect 16304 6205 16313 6239
rect 16313 6205 16347 6239
rect 16347 6205 16356 6239
rect 16304 6196 16356 6205
rect 2872 6128 2924 6180
rect 3516 6128 3568 6180
rect 4528 6171 4580 6180
rect 4528 6137 4537 6171
rect 4537 6137 4571 6171
rect 4571 6137 4580 6171
rect 4528 6128 4580 6137
rect 5908 6128 5960 6180
rect 7288 6128 7340 6180
rect 8116 6128 8168 6180
rect 8944 6128 8996 6180
rect 9128 6128 9180 6180
rect 10784 6171 10836 6180
rect 4804 6060 4856 6112
rect 10784 6137 10793 6171
rect 10793 6137 10827 6171
rect 10827 6137 10836 6171
rect 10784 6128 10836 6137
rect 16672 6128 16724 6180
rect 17776 6171 17828 6180
rect 17776 6137 17785 6171
rect 17785 6137 17819 6171
rect 17819 6137 17828 6171
rect 17776 6128 17828 6137
rect 9680 6060 9732 6112
rect 3106 5958 3158 6010
rect 3170 5958 3222 6010
rect 3234 5958 3286 6010
rect 3298 5958 3350 6010
rect 3362 5958 3414 6010
rect 6206 5958 6258 6010
rect 6270 5958 6322 6010
rect 6334 5958 6386 6010
rect 6398 5958 6450 6010
rect 6462 5958 6514 6010
rect 9306 5958 9358 6010
rect 9370 5958 9422 6010
rect 9434 5958 9486 6010
rect 9498 5958 9550 6010
rect 9562 5958 9614 6010
rect 12406 5958 12458 6010
rect 12470 5958 12522 6010
rect 12534 5958 12586 6010
rect 12598 5958 12650 6010
rect 12662 5958 12714 6010
rect 15506 5958 15558 6010
rect 15570 5958 15622 6010
rect 15634 5958 15686 6010
rect 15698 5958 15750 6010
rect 15762 5958 15814 6010
rect 18606 5958 18658 6010
rect 18670 5958 18722 6010
rect 18734 5958 18786 6010
rect 18798 5958 18850 6010
rect 18862 5958 18914 6010
rect 2320 5899 2372 5908
rect 2320 5865 2329 5899
rect 2329 5865 2363 5899
rect 2363 5865 2372 5899
rect 2320 5856 2372 5865
rect 2872 5788 2924 5840
rect 5264 5856 5316 5908
rect 5908 5856 5960 5908
rect 7288 5856 7340 5908
rect 9128 5856 9180 5908
rect 13544 5856 13596 5908
rect 13820 5856 13872 5908
rect 572 5763 624 5772
rect 572 5729 581 5763
rect 581 5729 615 5763
rect 615 5729 624 5763
rect 572 5720 624 5729
rect 3516 5720 3568 5772
rect 4804 5763 4856 5772
rect 4804 5729 4813 5763
rect 4813 5729 4847 5763
rect 4847 5729 4856 5763
rect 4804 5720 4856 5729
rect 5816 5720 5868 5772
rect 8116 5763 8168 5772
rect 8116 5729 8125 5763
rect 8125 5729 8159 5763
rect 8159 5729 8168 5763
rect 8116 5720 8168 5729
rect 8484 5720 8536 5772
rect 16212 5856 16264 5908
rect 17408 5856 17460 5908
rect 16672 5788 16724 5840
rect 16856 5720 16908 5772
rect 17500 5720 17552 5772
rect 940 5652 992 5704
rect 4252 5652 4304 5704
rect 5724 5652 5776 5704
rect 16948 5652 17000 5704
rect 8300 5627 8352 5636
rect 8300 5593 8309 5627
rect 8309 5593 8343 5627
rect 8343 5593 8352 5627
rect 8300 5584 8352 5593
rect 17592 5627 17644 5636
rect 17592 5593 17601 5627
rect 17601 5593 17635 5627
rect 17635 5593 17644 5627
rect 17592 5584 17644 5593
rect 2872 5559 2924 5568
rect 2872 5525 2881 5559
rect 2881 5525 2915 5559
rect 2915 5525 2924 5559
rect 2872 5516 2924 5525
rect 5908 5516 5960 5568
rect 1556 5414 1608 5466
rect 1620 5414 1672 5466
rect 1684 5414 1736 5466
rect 1748 5414 1800 5466
rect 1812 5414 1864 5466
rect 4656 5414 4708 5466
rect 4720 5414 4772 5466
rect 4784 5414 4836 5466
rect 4848 5414 4900 5466
rect 4912 5414 4964 5466
rect 7756 5414 7808 5466
rect 7820 5414 7872 5466
rect 7884 5414 7936 5466
rect 7948 5414 8000 5466
rect 8012 5414 8064 5466
rect 10856 5414 10908 5466
rect 10920 5414 10972 5466
rect 10984 5414 11036 5466
rect 11048 5414 11100 5466
rect 11112 5414 11164 5466
rect 13956 5414 14008 5466
rect 14020 5414 14072 5466
rect 14084 5414 14136 5466
rect 14148 5414 14200 5466
rect 14212 5414 14264 5466
rect 17056 5414 17108 5466
rect 17120 5414 17172 5466
rect 17184 5414 17236 5466
rect 17248 5414 17300 5466
rect 17312 5414 17364 5466
rect 2136 5312 2188 5364
rect 6736 5312 6788 5364
rect 7472 5312 7524 5364
rect 8668 5312 8720 5364
rect 1952 5176 2004 5228
rect 5724 5108 5776 5160
rect 7564 5244 7616 5296
rect 8760 5219 8812 5228
rect 8760 5185 8769 5219
rect 8769 5185 8803 5219
rect 8803 5185 8812 5219
rect 8760 5176 8812 5185
rect 13544 5219 13596 5228
rect 13544 5185 13553 5219
rect 13553 5185 13587 5219
rect 13587 5185 13596 5219
rect 13544 5176 13596 5185
rect 14832 5176 14884 5228
rect 16212 5176 16264 5228
rect 7196 5151 7248 5160
rect 7196 5117 7205 5151
rect 7205 5117 7239 5151
rect 7239 5117 7248 5151
rect 7196 5108 7248 5117
rect 7472 5151 7524 5160
rect 7472 5117 7481 5151
rect 7481 5117 7515 5151
rect 7515 5117 7524 5151
rect 7472 5108 7524 5117
rect 7656 5108 7708 5160
rect 7840 5108 7892 5160
rect 7104 5083 7156 5092
rect 7104 5049 7113 5083
rect 7113 5049 7147 5083
rect 7147 5049 7156 5083
rect 7104 5040 7156 5049
rect 7748 5040 7800 5092
rect 8116 5040 8168 5092
rect 12808 5108 12860 5160
rect 8760 5040 8812 5092
rect 9680 5040 9732 5092
rect 13820 5083 13872 5092
rect 2136 5015 2188 5024
rect 2136 4981 2145 5015
rect 2145 4981 2179 5015
rect 2179 4981 2188 5015
rect 2136 4972 2188 4981
rect 9772 4972 9824 5024
rect 11888 4972 11940 5024
rect 12256 4972 12308 5024
rect 13820 5049 13829 5083
rect 13829 5049 13863 5083
rect 13863 5049 13872 5083
rect 13820 5040 13872 5049
rect 16212 5083 16264 5092
rect 16212 5049 16221 5083
rect 16221 5049 16255 5083
rect 16255 5049 16264 5083
rect 16212 5040 16264 5049
rect 16672 5040 16724 5092
rect 17500 4972 17552 5024
rect 3106 4870 3158 4922
rect 3170 4870 3222 4922
rect 3234 4870 3286 4922
rect 3298 4870 3350 4922
rect 3362 4870 3414 4922
rect 6206 4870 6258 4922
rect 6270 4870 6322 4922
rect 6334 4870 6386 4922
rect 6398 4870 6450 4922
rect 6462 4870 6514 4922
rect 9306 4870 9358 4922
rect 9370 4870 9422 4922
rect 9434 4870 9486 4922
rect 9498 4870 9550 4922
rect 9562 4870 9614 4922
rect 12406 4870 12458 4922
rect 12470 4870 12522 4922
rect 12534 4870 12586 4922
rect 12598 4870 12650 4922
rect 12662 4870 12714 4922
rect 15506 4870 15558 4922
rect 15570 4870 15622 4922
rect 15634 4870 15686 4922
rect 15698 4870 15750 4922
rect 15762 4870 15814 4922
rect 18606 4870 18658 4922
rect 18670 4870 18722 4922
rect 18734 4870 18786 4922
rect 18798 4870 18850 4922
rect 18862 4870 18914 4922
rect 1952 4811 2004 4820
rect 1952 4777 1961 4811
rect 1961 4777 1995 4811
rect 1995 4777 2004 4811
rect 1952 4768 2004 4777
rect 2964 4768 3016 4820
rect 4160 4768 4212 4820
rect 4528 4811 4580 4820
rect 4528 4777 4537 4811
rect 4537 4777 4571 4811
rect 4571 4777 4580 4811
rect 4528 4768 4580 4777
rect 7196 4768 7248 4820
rect 8852 4768 8904 4820
rect 12808 4768 12860 4820
rect 13820 4768 13872 4820
rect 14740 4811 14792 4820
rect 14740 4777 14749 4811
rect 14749 4777 14783 4811
rect 14783 4777 14792 4811
rect 14740 4768 14792 4777
rect 15016 4768 15068 4820
rect 15476 4768 15528 4820
rect 1952 4632 2004 4684
rect 2780 4675 2832 4684
rect 2780 4641 2789 4675
rect 2789 4641 2823 4675
rect 2823 4641 2832 4675
rect 3332 4675 3384 4684
rect 2780 4632 2832 4641
rect 3332 4641 3341 4675
rect 3341 4641 3375 4675
rect 3375 4641 3384 4675
rect 3332 4632 3384 4641
rect 3884 4675 3936 4684
rect 3884 4641 3892 4675
rect 3892 4641 3926 4675
rect 3926 4641 3936 4675
rect 3884 4632 3936 4641
rect 5172 4632 5224 4684
rect 7564 4675 7616 4684
rect 7564 4641 7573 4675
rect 7573 4641 7607 4675
rect 7607 4641 7616 4675
rect 7564 4632 7616 4641
rect 7840 4632 7892 4684
rect 8484 4675 8536 4684
rect 8484 4641 8493 4675
rect 8493 4641 8527 4675
rect 8527 4641 8536 4675
rect 8484 4632 8536 4641
rect 8668 4632 8720 4684
rect 12256 4700 12308 4752
rect 9956 4632 10008 4684
rect 10140 4632 10192 4684
rect 13268 4700 13320 4752
rect 14280 4700 14332 4752
rect 12716 4632 12768 4684
rect 13728 4675 13780 4684
rect 13728 4641 13737 4675
rect 13737 4641 13771 4675
rect 13771 4641 13780 4675
rect 13728 4632 13780 4641
rect 4528 4607 4580 4616
rect 2044 4428 2096 4480
rect 4528 4573 4537 4607
rect 4537 4573 4571 4607
rect 4571 4573 4580 4607
rect 4528 4564 4580 4573
rect 5724 4564 5776 4616
rect 8116 4564 8168 4616
rect 4160 4496 4212 4548
rect 5540 4496 5592 4548
rect 11244 4564 11296 4616
rect 11888 4564 11940 4616
rect 13544 4564 13596 4616
rect 14280 4564 14332 4616
rect 9772 4496 9824 4548
rect 14464 4496 14516 4548
rect 15384 4496 15436 4548
rect 5724 4428 5776 4480
rect 8760 4471 8812 4480
rect 8760 4437 8769 4471
rect 8769 4437 8803 4471
rect 8803 4437 8812 4471
rect 8760 4428 8812 4437
rect 12440 4428 12492 4480
rect 1556 4326 1608 4378
rect 1620 4326 1672 4378
rect 1684 4326 1736 4378
rect 1748 4326 1800 4378
rect 1812 4326 1864 4378
rect 4656 4326 4708 4378
rect 4720 4326 4772 4378
rect 4784 4326 4836 4378
rect 4848 4326 4900 4378
rect 4912 4326 4964 4378
rect 7756 4326 7808 4378
rect 7820 4326 7872 4378
rect 7884 4326 7936 4378
rect 7948 4326 8000 4378
rect 8012 4326 8064 4378
rect 10856 4326 10908 4378
rect 10920 4326 10972 4378
rect 10984 4326 11036 4378
rect 11048 4326 11100 4378
rect 11112 4326 11164 4378
rect 13956 4326 14008 4378
rect 14020 4326 14072 4378
rect 14084 4326 14136 4378
rect 14148 4326 14200 4378
rect 14212 4326 14264 4378
rect 17056 4326 17108 4378
rect 17120 4326 17172 4378
rect 17184 4326 17236 4378
rect 17248 4326 17300 4378
rect 17312 4326 17364 4378
rect 1952 4156 2004 4208
rect 3332 4224 3384 4276
rect 5724 4267 5776 4276
rect 5724 4233 5733 4267
rect 5733 4233 5767 4267
rect 5767 4233 5776 4267
rect 5724 4224 5776 4233
rect 8852 4224 8904 4276
rect 756 4063 808 4072
rect 756 4029 765 4063
rect 765 4029 799 4063
rect 799 4029 808 4063
rect 756 4020 808 4029
rect 940 3952 992 4004
rect 1952 4063 2004 4072
rect 1952 4029 1961 4063
rect 1961 4029 1995 4063
rect 1995 4029 2004 4063
rect 3884 4088 3936 4140
rect 1952 4020 2004 4029
rect 3516 4063 3568 4072
rect 3516 4029 3525 4063
rect 3525 4029 3559 4063
rect 3559 4029 3568 4063
rect 3516 4020 3568 4029
rect 2320 3952 2372 4004
rect 2688 3952 2740 4004
rect 5448 4088 5500 4140
rect 4344 4063 4396 4072
rect 4344 4029 4353 4063
rect 4353 4029 4387 4063
rect 4387 4029 4396 4063
rect 5080 4063 5132 4072
rect 4344 4020 4396 4029
rect 5080 4029 5089 4063
rect 5089 4029 5123 4063
rect 5123 4029 5132 4063
rect 5080 4020 5132 4029
rect 5264 4063 5316 4072
rect 5264 4029 5273 4063
rect 5273 4029 5307 4063
rect 5307 4029 5316 4063
rect 5264 4020 5316 4029
rect 5540 4020 5592 4072
rect 6552 4156 6604 4208
rect 12440 4224 12492 4276
rect 12992 4224 13044 4276
rect 14280 4267 14332 4276
rect 14280 4233 14289 4267
rect 14289 4233 14323 4267
rect 14323 4233 14332 4267
rect 14280 4224 14332 4233
rect 14740 4224 14792 4276
rect 12808 4156 12860 4208
rect 7564 4088 7616 4140
rect 7472 4020 7524 4072
rect 5356 3952 5408 4004
rect 11244 4088 11296 4140
rect 11520 4131 11572 4140
rect 11520 4097 11529 4131
rect 11529 4097 11563 4131
rect 11563 4097 11572 4131
rect 14464 4156 14516 4208
rect 16948 4224 17000 4276
rect 17592 4156 17644 4208
rect 11520 4088 11572 4097
rect 9036 4063 9088 4072
rect 9036 4029 9045 4063
rect 9045 4029 9079 4063
rect 9079 4029 9088 4063
rect 9036 4020 9088 4029
rect 11612 4063 11664 4072
rect 11612 4029 11621 4063
rect 11621 4029 11655 4063
rect 11655 4029 11664 4063
rect 14740 4088 14792 4140
rect 15292 4088 15344 4140
rect 16856 4088 16908 4140
rect 17408 4088 17460 4140
rect 11612 4020 11664 4029
rect 12900 3952 12952 4004
rect 13268 4020 13320 4072
rect 15476 4063 15528 4072
rect 15476 4029 15485 4063
rect 15485 4029 15519 4063
rect 15519 4029 15528 4063
rect 15476 4020 15528 4029
rect 17776 4088 17828 4140
rect 17316 3995 17368 4004
rect 17316 3961 17325 3995
rect 17325 3961 17359 3995
rect 17359 3961 17368 3995
rect 17316 3952 17368 3961
rect 8944 3884 8996 3936
rect 12716 3927 12768 3936
rect 12716 3893 12725 3927
rect 12725 3893 12759 3927
rect 12759 3893 12768 3927
rect 12716 3884 12768 3893
rect 17684 4063 17736 4072
rect 17684 4029 17694 4063
rect 17694 4029 17728 4063
rect 17728 4029 17736 4063
rect 17684 4020 17736 4029
rect 3106 3782 3158 3834
rect 3170 3782 3222 3834
rect 3234 3782 3286 3834
rect 3298 3782 3350 3834
rect 3362 3782 3414 3834
rect 6206 3782 6258 3834
rect 6270 3782 6322 3834
rect 6334 3782 6386 3834
rect 6398 3782 6450 3834
rect 6462 3782 6514 3834
rect 9306 3782 9358 3834
rect 9370 3782 9422 3834
rect 9434 3782 9486 3834
rect 9498 3782 9550 3834
rect 9562 3782 9614 3834
rect 12406 3782 12458 3834
rect 12470 3782 12522 3834
rect 12534 3782 12586 3834
rect 12598 3782 12650 3834
rect 12662 3782 12714 3834
rect 15506 3782 15558 3834
rect 15570 3782 15622 3834
rect 15634 3782 15686 3834
rect 15698 3782 15750 3834
rect 15762 3782 15814 3834
rect 18606 3782 18658 3834
rect 18670 3782 18722 3834
rect 18734 3782 18786 3834
rect 18798 3782 18850 3834
rect 18862 3782 18914 3834
rect 756 3680 808 3732
rect 3884 3680 3936 3732
rect 4528 3723 4580 3732
rect 4528 3689 4537 3723
rect 4537 3689 4571 3723
rect 4571 3689 4580 3723
rect 4528 3680 4580 3689
rect 5448 3723 5500 3732
rect 5448 3689 5457 3723
rect 5457 3689 5491 3723
rect 5491 3689 5500 3723
rect 5448 3680 5500 3689
rect 5632 3680 5684 3732
rect 7564 3723 7616 3732
rect 7564 3689 7573 3723
rect 7573 3689 7607 3723
rect 7607 3689 7616 3723
rect 7564 3680 7616 3689
rect 9956 3723 10008 3732
rect 9956 3689 9965 3723
rect 9965 3689 9999 3723
rect 9999 3689 10008 3723
rect 9956 3680 10008 3689
rect 11612 3680 11664 3732
rect 14740 3723 14792 3732
rect 14740 3689 14749 3723
rect 14749 3689 14783 3723
rect 14783 3689 14792 3723
rect 14740 3680 14792 3689
rect 14924 3680 14976 3732
rect 15292 3680 15344 3732
rect 16304 3680 16356 3732
rect 17684 3680 17736 3732
rect 18052 3680 18104 3732
rect 940 3587 992 3596
rect 940 3553 949 3587
rect 949 3553 983 3587
rect 983 3553 992 3587
rect 940 3544 992 3553
rect 4142 3587 4194 3596
rect 4142 3553 4151 3587
rect 4151 3553 4185 3587
rect 4185 3553 4194 3587
rect 4142 3544 4194 3553
rect 5540 3587 5592 3596
rect 5540 3553 5549 3587
rect 5549 3553 5583 3587
rect 5583 3553 5592 3587
rect 5540 3544 5592 3553
rect 4344 3476 4396 3528
rect 5264 3476 5316 3528
rect 5356 3476 5408 3528
rect 8208 3544 8260 3596
rect 10232 3544 10284 3596
rect 11520 3612 11572 3664
rect 15016 3612 15068 3664
rect 16580 3612 16632 3664
rect 12440 3544 12492 3596
rect 12900 3544 12952 3596
rect 15384 3544 15436 3596
rect 16856 3544 16908 3596
rect 16948 3544 17000 3596
rect 17592 3587 17644 3596
rect 17592 3553 17601 3587
rect 17601 3553 17635 3587
rect 17635 3553 17644 3587
rect 17592 3544 17644 3553
rect 19064 3544 19116 3596
rect 5080 3340 5132 3392
rect 5264 3383 5316 3392
rect 5264 3349 5273 3383
rect 5273 3349 5307 3383
rect 5307 3349 5316 3383
rect 5264 3340 5316 3349
rect 5448 3408 5500 3460
rect 8116 3519 8168 3528
rect 8116 3485 8125 3519
rect 8125 3485 8159 3519
rect 8159 3485 8168 3519
rect 10416 3519 10468 3528
rect 8116 3476 8168 3485
rect 10416 3485 10425 3519
rect 10425 3485 10459 3519
rect 10459 3485 10468 3519
rect 10416 3476 10468 3485
rect 8392 3408 8444 3460
rect 8668 3408 8720 3460
rect 11336 3408 11388 3460
rect 17408 3476 17460 3528
rect 6736 3340 6788 3392
rect 16580 3340 16632 3392
rect 17316 3340 17368 3392
rect 1556 3238 1608 3290
rect 1620 3238 1672 3290
rect 1684 3238 1736 3290
rect 1748 3238 1800 3290
rect 1812 3238 1864 3290
rect 4656 3238 4708 3290
rect 4720 3238 4772 3290
rect 4784 3238 4836 3290
rect 4848 3238 4900 3290
rect 4912 3238 4964 3290
rect 7756 3238 7808 3290
rect 7820 3238 7872 3290
rect 7884 3238 7936 3290
rect 7948 3238 8000 3290
rect 8012 3238 8064 3290
rect 10856 3238 10908 3290
rect 10920 3238 10972 3290
rect 10984 3238 11036 3290
rect 11048 3238 11100 3290
rect 11112 3238 11164 3290
rect 13956 3238 14008 3290
rect 14020 3238 14072 3290
rect 14084 3238 14136 3290
rect 14148 3238 14200 3290
rect 14212 3238 14264 3290
rect 17056 3238 17108 3290
rect 17120 3238 17172 3290
rect 17184 3238 17236 3290
rect 17248 3238 17300 3290
rect 17312 3238 17364 3290
rect 5172 3179 5224 3188
rect 5172 3145 5181 3179
rect 5181 3145 5215 3179
rect 5215 3145 5224 3179
rect 5172 3136 5224 3145
rect 5264 3136 5316 3188
rect 6920 3136 6972 3188
rect 7104 3136 7156 3188
rect 10232 3179 10284 3188
rect 10232 3145 10241 3179
rect 10241 3145 10275 3179
rect 10275 3145 10284 3179
rect 10232 3136 10284 3145
rect 11336 3136 11388 3188
rect 12808 3136 12860 3188
rect 14188 3136 14240 3188
rect 14648 3136 14700 3188
rect 2872 3000 2924 3052
rect 6828 3000 6880 3052
rect 7472 3000 7524 3052
rect 9680 3043 9732 3052
rect 9680 3009 9689 3043
rect 9689 3009 9723 3043
rect 9723 3009 9732 3043
rect 9680 3000 9732 3009
rect 1492 2932 1544 2984
rect 2688 2932 2740 2984
rect 5264 2975 5316 2984
rect 5264 2941 5273 2975
rect 5273 2941 5307 2975
rect 5307 2941 5316 2975
rect 5264 2932 5316 2941
rect 6736 2932 6788 2984
rect 10416 3000 10468 3052
rect 12440 3000 12492 3052
rect 15200 3111 15252 3120
rect 15200 3077 15209 3111
rect 15209 3077 15243 3111
rect 15243 3077 15252 3111
rect 15200 3068 15252 3077
rect 13544 2975 13596 2984
rect 13544 2941 13553 2975
rect 13553 2941 13587 2975
rect 13587 2941 13596 2975
rect 13544 2932 13596 2941
rect 6920 2864 6972 2916
rect 7472 2907 7524 2916
rect 7472 2873 7481 2907
rect 7481 2873 7515 2907
rect 7515 2873 7524 2907
rect 7472 2864 7524 2873
rect 12992 2864 13044 2916
rect 14648 2932 14700 2984
rect 14832 2932 14884 2984
rect 14924 2975 14976 2984
rect 14924 2941 14933 2975
rect 14933 2941 14967 2975
rect 14967 2941 14976 2975
rect 14924 2932 14976 2941
rect 13820 2864 13872 2916
rect 15016 2864 15068 2916
rect 15844 2864 15896 2916
rect 1768 2839 1820 2848
rect 1768 2805 1777 2839
rect 1777 2805 1811 2839
rect 1811 2805 1820 2839
rect 1768 2796 1820 2805
rect 2136 2839 2188 2848
rect 2136 2805 2145 2839
rect 2145 2805 2179 2839
rect 2179 2805 2188 2839
rect 2136 2796 2188 2805
rect 7380 2839 7432 2848
rect 7380 2805 7389 2839
rect 7389 2805 7423 2839
rect 7423 2805 7432 2839
rect 7380 2796 7432 2805
rect 9864 2839 9916 2848
rect 9864 2805 9873 2839
rect 9873 2805 9907 2839
rect 9907 2805 9916 2839
rect 11612 2839 11664 2848
rect 9864 2796 9916 2805
rect 11612 2805 11621 2839
rect 11621 2805 11655 2839
rect 11655 2805 11664 2839
rect 11612 2796 11664 2805
rect 12256 2796 12308 2848
rect 12808 2839 12860 2848
rect 12808 2805 12817 2839
rect 12817 2805 12851 2839
rect 12851 2805 12860 2839
rect 12808 2796 12860 2805
rect 3106 2694 3158 2746
rect 3170 2694 3222 2746
rect 3234 2694 3286 2746
rect 3298 2694 3350 2746
rect 3362 2694 3414 2746
rect 6206 2694 6258 2746
rect 6270 2694 6322 2746
rect 6334 2694 6386 2746
rect 6398 2694 6450 2746
rect 6462 2694 6514 2746
rect 9306 2694 9358 2746
rect 9370 2694 9422 2746
rect 9434 2694 9486 2746
rect 9498 2694 9550 2746
rect 9562 2694 9614 2746
rect 12406 2694 12458 2746
rect 12470 2694 12522 2746
rect 12534 2694 12586 2746
rect 12598 2694 12650 2746
rect 12662 2694 12714 2746
rect 15506 2694 15558 2746
rect 15570 2694 15622 2746
rect 15634 2694 15686 2746
rect 15698 2694 15750 2746
rect 15762 2694 15814 2746
rect 18606 2694 18658 2746
rect 18670 2694 18722 2746
rect 18734 2694 18786 2746
rect 18798 2694 18850 2746
rect 18862 2694 18914 2746
rect 940 2592 992 2644
rect 1768 2592 1820 2644
rect 2136 2635 2188 2644
rect 2136 2601 2145 2635
rect 2145 2601 2179 2635
rect 2179 2601 2188 2635
rect 2136 2592 2188 2601
rect 2780 2592 2832 2644
rect 3332 2635 3384 2644
rect 3332 2601 3341 2635
rect 3341 2601 3375 2635
rect 3375 2601 3384 2635
rect 3332 2592 3384 2601
rect 5080 2592 5132 2644
rect 5264 2592 5316 2644
rect 8208 2635 8260 2644
rect 8208 2601 8217 2635
rect 8217 2601 8251 2635
rect 8251 2601 8260 2635
rect 8208 2592 8260 2601
rect 9036 2592 9088 2644
rect 13728 2592 13780 2644
rect 15384 2592 15436 2644
rect 1492 2567 1544 2576
rect 1492 2533 1501 2567
rect 1501 2533 1535 2567
rect 1535 2533 1544 2567
rect 1492 2524 1544 2533
rect 3976 2524 4028 2576
rect 8392 2524 8444 2576
rect 12256 2524 12308 2576
rect 13820 2524 13872 2576
rect 14188 2567 14240 2576
rect 14188 2533 14197 2567
rect 14197 2533 14231 2567
rect 14231 2533 14240 2567
rect 14188 2524 14240 2533
rect 17592 2524 17644 2576
rect 18328 2524 18380 2576
rect 2320 2499 2372 2508
rect 2320 2465 2329 2499
rect 2329 2465 2363 2499
rect 2363 2465 2372 2499
rect 2320 2456 2372 2465
rect 3608 2456 3660 2508
rect 6368 2456 6420 2508
rect 16764 2456 16816 2508
rect 17316 2499 17368 2508
rect 17316 2465 17325 2499
rect 17325 2465 17359 2499
rect 17359 2465 17368 2499
rect 17316 2456 17368 2465
rect 17500 2456 17552 2508
rect 17960 2499 18012 2508
rect 17960 2465 17969 2499
rect 17969 2465 18003 2499
rect 18003 2465 18012 2499
rect 17960 2456 18012 2465
rect 1952 2388 2004 2440
rect 5816 2431 5868 2440
rect 5816 2397 5825 2431
rect 5825 2397 5859 2431
rect 5859 2397 5868 2431
rect 5816 2388 5868 2397
rect 6828 2388 6880 2440
rect 9680 2388 9732 2440
rect 14372 2388 14424 2440
rect 15016 2431 15068 2440
rect 15016 2397 15025 2431
rect 15025 2397 15059 2431
rect 15059 2397 15068 2431
rect 15016 2388 15068 2397
rect 16488 2388 16540 2440
rect 17408 2295 17460 2304
rect 17408 2261 17417 2295
rect 17417 2261 17451 2295
rect 17451 2261 17460 2295
rect 17408 2252 17460 2261
rect 1556 2150 1608 2202
rect 1620 2150 1672 2202
rect 1684 2150 1736 2202
rect 1748 2150 1800 2202
rect 1812 2150 1864 2202
rect 4656 2150 4708 2202
rect 4720 2150 4772 2202
rect 4784 2150 4836 2202
rect 4848 2150 4900 2202
rect 4912 2150 4964 2202
rect 7756 2150 7808 2202
rect 7820 2150 7872 2202
rect 7884 2150 7936 2202
rect 7948 2150 8000 2202
rect 8012 2150 8064 2202
rect 10856 2150 10908 2202
rect 10920 2150 10972 2202
rect 10984 2150 11036 2202
rect 11048 2150 11100 2202
rect 11112 2150 11164 2202
rect 13956 2150 14008 2202
rect 14020 2150 14072 2202
rect 14084 2150 14136 2202
rect 14148 2150 14200 2202
rect 14212 2150 14264 2202
rect 17056 2150 17108 2202
rect 17120 2150 17172 2202
rect 17184 2150 17236 2202
rect 17248 2150 17300 2202
rect 17312 2150 17364 2202
rect 3608 2091 3660 2100
rect 3608 2057 3617 2091
rect 3617 2057 3651 2091
rect 3651 2057 3660 2091
rect 3608 2048 3660 2057
rect 3976 2048 4028 2100
rect 6368 2091 6420 2100
rect 4252 1980 4304 2032
rect 5264 1980 5316 2032
rect 6368 2057 6377 2091
rect 6377 2057 6411 2091
rect 6411 2057 6420 2091
rect 6368 2048 6420 2057
rect 7380 2048 7432 2100
rect 9864 2091 9916 2100
rect 9864 2057 9873 2091
rect 9873 2057 9907 2091
rect 9907 2057 9916 2091
rect 9864 2048 9916 2057
rect 10416 2091 10468 2100
rect 10416 2057 10425 2091
rect 10425 2057 10459 2091
rect 10459 2057 10468 2091
rect 10416 2048 10468 2057
rect 10784 2048 10836 2100
rect 11612 2048 11664 2100
rect 12808 2048 12860 2100
rect 14832 2091 14884 2100
rect 14832 2057 14841 2091
rect 14841 2057 14875 2091
rect 14875 2057 14884 2091
rect 14832 2048 14884 2057
rect 16212 2048 16264 2100
rect 2872 1912 2924 1964
rect 5540 1912 5592 1964
rect 3332 1844 3384 1896
rect 3516 1844 3568 1896
rect 3976 1887 4028 1896
rect 3976 1853 3985 1887
rect 3985 1853 4019 1887
rect 4019 1853 4028 1887
rect 3976 1844 4028 1853
rect 4252 1844 4304 1896
rect 5172 1887 5224 1896
rect 5172 1853 5181 1887
rect 5181 1853 5215 1887
rect 5215 1853 5224 1887
rect 5172 1844 5224 1853
rect 5264 1844 5316 1896
rect 7472 1912 7524 1964
rect 9036 1980 9088 2032
rect 15844 1980 15896 2032
rect 5816 1844 5868 1896
rect 6736 1844 6788 1896
rect 9772 1912 9824 1964
rect 14372 1955 14424 1964
rect 14372 1921 14381 1955
rect 14381 1921 14415 1955
rect 14415 1921 14424 1955
rect 14372 1912 14424 1921
rect 16488 1955 16540 1964
rect 16488 1921 16497 1955
rect 16497 1921 16531 1955
rect 16531 1921 16540 1955
rect 16488 1912 16540 1921
rect 9220 1844 9272 1896
rect 10048 1887 10100 1896
rect 10048 1853 10057 1887
rect 10057 1853 10091 1887
rect 10091 1853 10100 1887
rect 10324 1887 10376 1896
rect 10048 1844 10100 1853
rect 10324 1853 10333 1887
rect 10333 1853 10367 1887
rect 10367 1853 10376 1887
rect 10324 1844 10376 1853
rect 12256 1844 12308 1896
rect 12808 1887 12860 1896
rect 3516 1708 3568 1760
rect 5540 1708 5592 1760
rect 6736 1751 6788 1760
rect 6736 1717 6745 1751
rect 6745 1717 6779 1751
rect 6779 1717 6788 1751
rect 6736 1708 6788 1717
rect 8024 1751 8076 1760
rect 8024 1717 8033 1751
rect 8033 1717 8067 1751
rect 8067 1717 8076 1751
rect 8024 1708 8076 1717
rect 11152 1776 11204 1828
rect 11612 1776 11664 1828
rect 12808 1853 12817 1887
rect 12817 1853 12851 1887
rect 12851 1853 12860 1887
rect 12808 1844 12860 1853
rect 13728 1844 13780 1896
rect 14832 1844 14884 1896
rect 17224 1844 17276 1896
rect 17408 1912 17460 1964
rect 13544 1776 13596 1828
rect 9680 1708 9732 1760
rect 11888 1751 11940 1760
rect 11888 1717 11897 1751
rect 11897 1717 11931 1751
rect 11931 1717 11940 1751
rect 11888 1708 11940 1717
rect 14096 1751 14148 1760
rect 14096 1717 14105 1751
rect 14105 1717 14139 1751
rect 14139 1717 14148 1751
rect 14096 1708 14148 1717
rect 16764 1708 16816 1760
rect 17316 1751 17368 1760
rect 17316 1717 17325 1751
rect 17325 1717 17359 1751
rect 17359 1717 17368 1751
rect 17316 1708 17368 1717
rect 3106 1606 3158 1658
rect 3170 1606 3222 1658
rect 3234 1606 3286 1658
rect 3298 1606 3350 1658
rect 3362 1606 3414 1658
rect 6206 1606 6258 1658
rect 6270 1606 6322 1658
rect 6334 1606 6386 1658
rect 6398 1606 6450 1658
rect 6462 1606 6514 1658
rect 9306 1606 9358 1658
rect 9370 1606 9422 1658
rect 9434 1606 9486 1658
rect 9498 1606 9550 1658
rect 9562 1606 9614 1658
rect 12406 1606 12458 1658
rect 12470 1606 12522 1658
rect 12534 1606 12586 1658
rect 12598 1606 12650 1658
rect 12662 1606 12714 1658
rect 15506 1606 15558 1658
rect 15570 1606 15622 1658
rect 15634 1606 15686 1658
rect 15698 1606 15750 1658
rect 15762 1606 15814 1658
rect 18606 1606 18658 1658
rect 18670 1606 18722 1658
rect 18734 1606 18786 1658
rect 18798 1606 18850 1658
rect 18862 1606 18914 1658
rect 3516 1504 3568 1556
rect 6736 1504 6788 1556
rect 8024 1504 8076 1556
rect 3608 1368 3660 1420
rect 5540 1411 5592 1420
rect 5540 1377 5549 1411
rect 5549 1377 5583 1411
rect 5583 1377 5592 1411
rect 5540 1368 5592 1377
rect 5632 1411 5684 1420
rect 5632 1377 5642 1411
rect 5642 1377 5676 1411
rect 5676 1377 5684 1411
rect 5632 1368 5684 1377
rect 7656 1368 7708 1420
rect 9220 1504 9272 1556
rect 10048 1504 10100 1556
rect 11888 1504 11940 1556
rect 12256 1504 12308 1556
rect 16856 1504 16908 1556
rect 17500 1547 17552 1556
rect 17500 1513 17509 1547
rect 17509 1513 17543 1547
rect 17543 1513 17552 1547
rect 17500 1504 17552 1513
rect 9036 1436 9088 1488
rect 10324 1436 10376 1488
rect 3976 1300 4028 1352
rect 9772 1368 9824 1420
rect 10416 1368 10468 1420
rect 11152 1368 11204 1420
rect 11336 1411 11388 1420
rect 11336 1377 11345 1411
rect 11345 1377 11379 1411
rect 11379 1377 11388 1411
rect 11336 1368 11388 1377
rect 13728 1436 13780 1488
rect 17224 1436 17276 1488
rect 17592 1479 17644 1488
rect 17592 1445 17601 1479
rect 17601 1445 17635 1479
rect 17635 1445 17644 1479
rect 17592 1436 17644 1445
rect 13544 1368 13596 1420
rect 14648 1368 14700 1420
rect 16764 1368 16816 1420
rect 11244 1300 11296 1352
rect 12808 1300 12860 1352
rect 13820 1300 13872 1352
rect 16580 1300 16632 1352
rect 14096 1232 14148 1284
rect 17316 1232 17368 1284
rect 17408 1232 17460 1284
rect 11428 1164 11480 1216
rect 1556 1062 1608 1114
rect 1620 1062 1672 1114
rect 1684 1062 1736 1114
rect 1748 1062 1800 1114
rect 1812 1062 1864 1114
rect 4656 1062 4708 1114
rect 4720 1062 4772 1114
rect 4784 1062 4836 1114
rect 4848 1062 4900 1114
rect 4912 1062 4964 1114
rect 7756 1062 7808 1114
rect 7820 1062 7872 1114
rect 7884 1062 7936 1114
rect 7948 1062 8000 1114
rect 8012 1062 8064 1114
rect 10856 1062 10908 1114
rect 10920 1062 10972 1114
rect 10984 1062 11036 1114
rect 11048 1062 11100 1114
rect 11112 1062 11164 1114
rect 13956 1062 14008 1114
rect 14020 1062 14072 1114
rect 14084 1062 14136 1114
rect 14148 1062 14200 1114
rect 14212 1062 14264 1114
rect 17056 1062 17108 1114
rect 17120 1062 17172 1114
rect 17184 1062 17236 1114
rect 17248 1062 17300 1114
rect 17312 1062 17364 1114
rect 3976 960 4028 1012
rect 5632 960 5684 1012
rect 11336 1003 11388 1012
rect 11336 969 11345 1003
rect 11345 969 11379 1003
rect 11379 969 11388 1003
rect 11336 960 11388 969
rect 17592 960 17644 1012
rect 17960 1003 18012 1012
rect 17960 969 17969 1003
rect 17969 969 18003 1003
rect 18003 969 18012 1003
rect 17960 960 18012 969
rect 18420 1003 18472 1012
rect 18420 969 18429 1003
rect 18429 969 18463 1003
rect 18463 969 18472 1003
rect 18420 960 18472 969
rect 5264 892 5316 944
rect 11428 935 11480 944
rect 11428 901 11437 935
rect 11437 901 11471 935
rect 11471 901 11480 935
rect 11428 892 11480 901
rect 13820 892 13872 944
rect 11612 867 11664 876
rect 11612 833 11621 867
rect 11621 833 11655 867
rect 11655 833 11664 867
rect 11612 824 11664 833
rect 5172 756 5224 808
rect 11244 756 11296 808
rect 3106 518 3158 570
rect 3170 518 3222 570
rect 3234 518 3286 570
rect 3298 518 3350 570
rect 3362 518 3414 570
rect 6206 518 6258 570
rect 6270 518 6322 570
rect 6334 518 6386 570
rect 6398 518 6450 570
rect 6462 518 6514 570
rect 9306 518 9358 570
rect 9370 518 9422 570
rect 9434 518 9486 570
rect 9498 518 9550 570
rect 9562 518 9614 570
rect 12406 518 12458 570
rect 12470 518 12522 570
rect 12534 518 12586 570
rect 12598 518 12650 570
rect 12662 518 12714 570
rect 15506 518 15558 570
rect 15570 518 15622 570
rect 15634 518 15686 570
rect 15698 518 15750 570
rect 15762 518 15814 570
rect 18606 518 18658 570
rect 18670 518 18722 570
rect 18734 518 18786 570
rect 18798 518 18850 570
rect 18862 518 18914 570
<< metal2 >>
rect 1398 19200 1454 20000
rect 4250 19200 4306 20000
rect 7102 19200 7158 20000
rect 9954 19200 10010 20000
rect 12806 19200 12862 20000
rect 15396 19230 15608 19258
rect 1412 18222 1440 19200
rect 1556 18524 1864 18533
rect 1556 18522 1562 18524
rect 1618 18522 1642 18524
rect 1698 18522 1722 18524
rect 1778 18522 1802 18524
rect 1858 18522 1864 18524
rect 1618 18470 1620 18522
rect 1800 18470 1802 18522
rect 1556 18468 1562 18470
rect 1618 18468 1642 18470
rect 1698 18468 1722 18470
rect 1778 18468 1802 18470
rect 1858 18468 1864 18470
rect 1556 18459 1864 18468
rect 4264 18426 4292 19200
rect 4656 18524 4964 18533
rect 4656 18522 4662 18524
rect 4718 18522 4742 18524
rect 4798 18522 4822 18524
rect 4878 18522 4902 18524
rect 4958 18522 4964 18524
rect 4718 18470 4720 18522
rect 4900 18470 4902 18522
rect 4656 18468 4662 18470
rect 4718 18468 4742 18470
rect 4798 18468 4822 18470
rect 4878 18468 4902 18470
rect 4958 18468 4964 18470
rect 4656 18459 4964 18468
rect 4252 18420 4304 18426
rect 4252 18362 4304 18368
rect 1400 18216 1452 18222
rect 1400 18158 1452 18164
rect 3976 18216 4028 18222
rect 3976 18158 4028 18164
rect 4160 18216 4212 18222
rect 4160 18158 4212 18164
rect 2780 18148 2832 18154
rect 2780 18090 2832 18096
rect 2872 18148 2924 18154
rect 2872 18090 2924 18096
rect 3884 18148 3936 18154
rect 3884 18090 3936 18096
rect 2504 18080 2556 18086
rect 2504 18022 2556 18028
rect 2412 17808 2464 17814
rect 2412 17750 2464 17756
rect 572 17672 624 17678
rect 572 17614 624 17620
rect 848 17672 900 17678
rect 848 17614 900 17620
rect 584 14482 612 17614
rect 860 17270 888 17614
rect 2044 17536 2096 17542
rect 2044 17478 2096 17484
rect 1556 17436 1864 17445
rect 1556 17434 1562 17436
rect 1618 17434 1642 17436
rect 1698 17434 1722 17436
rect 1778 17434 1802 17436
rect 1858 17434 1864 17436
rect 1618 17382 1620 17434
rect 1800 17382 1802 17434
rect 1556 17380 1562 17382
rect 1618 17380 1642 17382
rect 1698 17380 1722 17382
rect 1778 17380 1802 17382
rect 1858 17380 1864 17382
rect 1556 17371 1864 17380
rect 1400 17332 1452 17338
rect 1400 17274 1452 17280
rect 848 17264 900 17270
rect 848 17206 900 17212
rect 1124 17128 1176 17134
rect 1124 17070 1176 17076
rect 1216 17128 1268 17134
rect 1216 17070 1268 17076
rect 1136 16726 1164 17070
rect 1228 16794 1256 17070
rect 1216 16788 1268 16794
rect 1216 16730 1268 16736
rect 1124 16720 1176 16726
rect 1124 16662 1176 16668
rect 848 14816 900 14822
rect 848 14758 900 14764
rect 860 14550 888 14758
rect 848 14544 900 14550
rect 848 14486 900 14492
rect 572 14476 624 14482
rect 572 14418 624 14424
rect 584 13394 612 14418
rect 572 13388 624 13394
rect 572 13330 624 13336
rect 940 13320 992 13326
rect 940 13262 992 13268
rect 952 12986 980 13262
rect 940 12980 992 12986
rect 940 12922 992 12928
rect 1412 10266 1440 17274
rect 2056 16810 2084 17478
rect 2424 17134 2452 17750
rect 2412 17128 2464 17134
rect 2412 17070 2464 17076
rect 2056 16782 2360 16810
rect 2056 16658 2084 16782
rect 2044 16652 2096 16658
rect 2044 16594 2096 16600
rect 2136 16652 2188 16658
rect 2136 16594 2188 16600
rect 1556 16348 1864 16357
rect 1556 16346 1562 16348
rect 1618 16346 1642 16348
rect 1698 16346 1722 16348
rect 1778 16346 1802 16348
rect 1858 16346 1864 16348
rect 1618 16294 1620 16346
rect 1800 16294 1802 16346
rect 1556 16292 1562 16294
rect 1618 16292 1642 16294
rect 1698 16292 1722 16294
rect 1778 16292 1802 16294
rect 1858 16292 1864 16294
rect 1556 16283 1864 16292
rect 1556 15260 1864 15269
rect 1556 15258 1562 15260
rect 1618 15258 1642 15260
rect 1698 15258 1722 15260
rect 1778 15258 1802 15260
rect 1858 15258 1864 15260
rect 1618 15206 1620 15258
rect 1800 15206 1802 15258
rect 1556 15204 1562 15206
rect 1618 15204 1642 15206
rect 1698 15204 1722 15206
rect 1778 15204 1802 15206
rect 1858 15204 1864 15206
rect 1556 15195 1864 15204
rect 2148 15026 2176 16594
rect 2228 16448 2280 16454
rect 2228 16390 2280 16396
rect 2240 15026 2268 16390
rect 2332 16046 2360 16782
rect 2424 16674 2452 17070
rect 2516 16998 2544 18022
rect 2688 17740 2740 17746
rect 2688 17682 2740 17688
rect 2700 17338 2728 17682
rect 2792 17610 2820 18090
rect 2780 17604 2832 17610
rect 2780 17546 2832 17552
rect 2688 17332 2740 17338
rect 2688 17274 2740 17280
rect 2596 17264 2648 17270
rect 2596 17206 2648 17212
rect 2504 16992 2556 16998
rect 2504 16934 2556 16940
rect 2516 16794 2544 16934
rect 2504 16788 2556 16794
rect 2504 16730 2556 16736
rect 2608 16726 2636 17206
rect 2688 17128 2740 17134
rect 2688 17070 2740 17076
rect 2596 16720 2648 16726
rect 2424 16646 2544 16674
rect 2596 16662 2648 16668
rect 2700 16658 2728 17070
rect 2884 16658 2912 18090
rect 3106 17980 3414 17989
rect 3106 17978 3112 17980
rect 3168 17978 3192 17980
rect 3248 17978 3272 17980
rect 3328 17978 3352 17980
rect 3408 17978 3414 17980
rect 3168 17926 3170 17978
rect 3350 17926 3352 17978
rect 3106 17924 3112 17926
rect 3168 17924 3192 17926
rect 3248 17924 3272 17926
rect 3328 17924 3352 17926
rect 3408 17924 3414 17926
rect 3106 17915 3414 17924
rect 3056 17876 3108 17882
rect 3056 17818 3108 17824
rect 3068 17202 3096 17818
rect 3056 17196 3108 17202
rect 3056 17138 3108 17144
rect 3106 16892 3414 16901
rect 3106 16890 3112 16892
rect 3168 16890 3192 16892
rect 3248 16890 3272 16892
rect 3328 16890 3352 16892
rect 3408 16890 3414 16892
rect 3168 16838 3170 16890
rect 3350 16838 3352 16890
rect 3106 16836 3112 16838
rect 3168 16836 3192 16838
rect 3248 16836 3272 16838
rect 3328 16836 3352 16838
rect 3408 16836 3414 16838
rect 3106 16827 3414 16836
rect 2320 16040 2372 16046
rect 2320 15982 2372 15988
rect 2136 15020 2188 15026
rect 2136 14962 2188 14968
rect 2228 15020 2280 15026
rect 2228 14962 2280 14968
rect 2148 14550 2176 14962
rect 2136 14544 2188 14550
rect 2136 14486 2188 14492
rect 1556 14172 1864 14181
rect 1556 14170 1562 14172
rect 1618 14170 1642 14172
rect 1698 14170 1722 14172
rect 1778 14170 1802 14172
rect 1858 14170 1864 14172
rect 1618 14118 1620 14170
rect 1800 14118 1802 14170
rect 1556 14116 1562 14118
rect 1618 14116 1642 14118
rect 1698 14116 1722 14118
rect 1778 14116 1802 14118
rect 1858 14116 1864 14118
rect 1556 14107 1864 14116
rect 1556 13084 1864 13093
rect 1556 13082 1562 13084
rect 1618 13082 1642 13084
rect 1698 13082 1722 13084
rect 1778 13082 1802 13084
rect 1858 13082 1864 13084
rect 1618 13030 1620 13082
rect 1800 13030 1802 13082
rect 1556 13028 1562 13030
rect 1618 13028 1642 13030
rect 1698 13028 1722 13030
rect 1778 13028 1802 13030
rect 1858 13028 1864 13030
rect 1556 13019 1864 13028
rect 2148 12850 2176 14486
rect 2240 13870 2268 14962
rect 2516 14482 2544 16646
rect 2688 16652 2740 16658
rect 2688 16594 2740 16600
rect 2872 16652 2924 16658
rect 2872 16594 2924 16600
rect 2596 16516 2648 16522
rect 2596 16458 2648 16464
rect 2608 16046 2636 16458
rect 2596 16040 2648 16046
rect 2596 15982 2648 15988
rect 2608 14958 2636 15982
rect 2596 14952 2648 14958
rect 2596 14894 2648 14900
rect 2608 14618 2636 14894
rect 2688 14884 2740 14890
rect 2688 14826 2740 14832
rect 2700 14618 2728 14826
rect 2596 14612 2648 14618
rect 2596 14554 2648 14560
rect 2688 14612 2740 14618
rect 2688 14554 2740 14560
rect 2320 14476 2372 14482
rect 2320 14418 2372 14424
rect 2504 14476 2556 14482
rect 2504 14418 2556 14424
rect 2228 13864 2280 13870
rect 2228 13806 2280 13812
rect 2240 13394 2268 13806
rect 2332 13462 2360 14418
rect 2320 13456 2372 13462
rect 2320 13398 2372 13404
rect 2228 13388 2280 13394
rect 2228 13330 2280 13336
rect 2136 12844 2188 12850
rect 2136 12786 2188 12792
rect 2240 12782 2268 13330
rect 2228 12776 2280 12782
rect 2228 12718 2280 12724
rect 1952 12096 2004 12102
rect 1952 12038 2004 12044
rect 1556 11996 1864 12005
rect 1556 11994 1562 11996
rect 1618 11994 1642 11996
rect 1698 11994 1722 11996
rect 1778 11994 1802 11996
rect 1858 11994 1864 11996
rect 1618 11942 1620 11994
rect 1800 11942 1802 11994
rect 1556 11940 1562 11942
rect 1618 11940 1642 11942
rect 1698 11940 1722 11942
rect 1778 11940 1802 11942
rect 1858 11940 1864 11942
rect 1556 11931 1864 11940
rect 1964 11898 1992 12038
rect 1952 11892 2004 11898
rect 1952 11834 2004 11840
rect 2044 11688 2096 11694
rect 2044 11630 2096 11636
rect 1676 11552 1728 11558
rect 1676 11494 1728 11500
rect 1688 11354 1716 11494
rect 2056 11354 2084 11630
rect 2332 11626 2360 13398
rect 2780 13320 2832 13326
rect 2780 13262 2832 13268
rect 2792 12306 2820 13262
rect 2780 12300 2832 12306
rect 2780 12242 2832 12248
rect 2320 11620 2372 11626
rect 2320 11562 2372 11568
rect 2228 11552 2280 11558
rect 2228 11494 2280 11500
rect 1676 11348 1728 11354
rect 1676 11290 1728 11296
rect 2044 11348 2096 11354
rect 2044 11290 2096 11296
rect 2136 11076 2188 11082
rect 2136 11018 2188 11024
rect 1556 10908 1864 10917
rect 1556 10906 1562 10908
rect 1618 10906 1642 10908
rect 1698 10906 1722 10908
rect 1778 10906 1802 10908
rect 1858 10906 1864 10908
rect 1618 10854 1620 10906
rect 1800 10854 1802 10906
rect 1556 10852 1562 10854
rect 1618 10852 1642 10854
rect 1698 10852 1722 10854
rect 1778 10852 1802 10854
rect 1858 10852 1864 10854
rect 1556 10843 1864 10852
rect 1400 10260 1452 10266
rect 1400 10202 1452 10208
rect 940 10124 992 10130
rect 940 10066 992 10072
rect 952 10033 980 10066
rect 938 10024 994 10033
rect 938 9959 994 9968
rect 1556 9820 1864 9829
rect 1556 9818 1562 9820
rect 1618 9818 1642 9820
rect 1698 9818 1722 9820
rect 1778 9818 1802 9820
rect 1858 9818 1864 9820
rect 1618 9766 1620 9818
rect 1800 9766 1802 9818
rect 1556 9764 1562 9766
rect 1618 9764 1642 9766
rect 1698 9764 1722 9766
rect 1778 9764 1802 9766
rect 1858 9764 1864 9766
rect 1556 9755 1864 9764
rect 2148 9586 2176 11018
rect 2240 10606 2268 11494
rect 2688 11144 2740 11150
rect 2688 11086 2740 11092
rect 2700 10810 2728 11086
rect 2688 10804 2740 10810
rect 2688 10746 2740 10752
rect 2596 10668 2648 10674
rect 2596 10610 2648 10616
rect 2228 10600 2280 10606
rect 2228 10542 2280 10548
rect 2136 9580 2188 9586
rect 2136 9522 2188 9528
rect 848 9376 900 9382
rect 848 9318 900 9324
rect 860 9110 888 9318
rect 848 9104 900 9110
rect 848 9046 900 9052
rect 572 8968 624 8974
rect 572 8910 624 8916
rect 584 7886 612 8910
rect 1556 8732 1864 8741
rect 1556 8730 1562 8732
rect 1618 8730 1642 8732
rect 1698 8730 1722 8732
rect 1778 8730 1802 8732
rect 1858 8730 1864 8732
rect 1618 8678 1620 8730
rect 1800 8678 1802 8730
rect 1556 8676 1562 8678
rect 1618 8676 1642 8678
rect 1698 8676 1722 8678
rect 1778 8676 1802 8678
rect 1858 8676 1864 8678
rect 1556 8667 1864 8676
rect 572 7880 624 7886
rect 572 7822 624 7828
rect 940 7880 992 7886
rect 940 7822 992 7828
rect 584 6934 612 7822
rect 952 7546 980 7822
rect 1556 7644 1864 7653
rect 1556 7642 1562 7644
rect 1618 7642 1642 7644
rect 1698 7642 1722 7644
rect 1778 7642 1802 7644
rect 1858 7642 1864 7644
rect 1618 7590 1620 7642
rect 1800 7590 1802 7642
rect 1556 7588 1562 7590
rect 1618 7588 1642 7590
rect 1698 7588 1722 7590
rect 1778 7588 1802 7590
rect 1858 7588 1864 7590
rect 1556 7579 1864 7588
rect 940 7540 992 7546
rect 940 7482 992 7488
rect 2148 7410 2176 9522
rect 2320 9512 2372 9518
rect 2320 9454 2372 9460
rect 2332 9178 2360 9454
rect 2320 9172 2372 9178
rect 2320 9114 2372 9120
rect 2332 8498 2360 9114
rect 2608 8634 2636 10610
rect 2688 10600 2740 10606
rect 2688 10542 2740 10548
rect 2700 9518 2728 10542
rect 2688 9512 2740 9518
rect 2688 9454 2740 9460
rect 2596 8628 2648 8634
rect 2596 8570 2648 8576
rect 2320 8492 2372 8498
rect 2320 8434 2372 8440
rect 2608 8090 2636 8570
rect 2700 8362 2728 9454
rect 2884 9110 2912 16594
rect 3608 15904 3660 15910
rect 3608 15846 3660 15852
rect 3106 15804 3414 15813
rect 3106 15802 3112 15804
rect 3168 15802 3192 15804
rect 3248 15802 3272 15804
rect 3328 15802 3352 15804
rect 3408 15802 3414 15804
rect 3168 15750 3170 15802
rect 3350 15750 3352 15802
rect 3106 15748 3112 15750
rect 3168 15748 3192 15750
rect 3248 15748 3272 15750
rect 3328 15748 3352 15750
rect 3408 15748 3414 15750
rect 3106 15739 3414 15748
rect 3620 14958 3648 15846
rect 3608 14952 3660 14958
rect 3608 14894 3660 14900
rect 2964 14816 3016 14822
rect 2964 14758 3016 14764
rect 3516 14816 3568 14822
rect 3516 14758 3568 14764
rect 2976 14618 3004 14758
rect 3106 14716 3414 14725
rect 3106 14714 3112 14716
rect 3168 14714 3192 14716
rect 3248 14714 3272 14716
rect 3328 14714 3352 14716
rect 3408 14714 3414 14716
rect 3168 14662 3170 14714
rect 3350 14662 3352 14714
rect 3106 14660 3112 14662
rect 3168 14660 3192 14662
rect 3248 14660 3272 14662
rect 3328 14660 3352 14662
rect 3408 14660 3414 14662
rect 3106 14651 3414 14660
rect 2964 14612 3016 14618
rect 2964 14554 3016 14560
rect 3148 14476 3200 14482
rect 3148 14418 3200 14424
rect 3160 14006 3188 14418
rect 3528 14414 3556 14758
rect 3516 14408 3568 14414
rect 3516 14350 3568 14356
rect 3148 14000 3200 14006
rect 3148 13942 3200 13948
rect 2964 13728 3016 13734
rect 2964 13670 3016 13676
rect 2976 12850 3004 13670
rect 3106 13628 3414 13637
rect 3106 13626 3112 13628
rect 3168 13626 3192 13628
rect 3248 13626 3272 13628
rect 3328 13626 3352 13628
rect 3408 13626 3414 13628
rect 3168 13574 3170 13626
rect 3350 13574 3352 13626
rect 3106 13572 3112 13574
rect 3168 13572 3192 13574
rect 3248 13572 3272 13574
rect 3328 13572 3352 13574
rect 3408 13572 3414 13574
rect 3106 13563 3414 13572
rect 3528 12850 3556 14350
rect 3896 14074 3924 18090
rect 3988 17882 4016 18158
rect 3976 17876 4028 17882
rect 3976 17818 4028 17824
rect 4172 17814 4200 18158
rect 4160 17808 4212 17814
rect 4160 17750 4212 17756
rect 4264 17746 4292 18362
rect 5816 18352 5868 18358
rect 5816 18294 5868 18300
rect 5724 18284 5776 18290
rect 5724 18226 5776 18232
rect 4528 18216 4580 18222
rect 4528 18158 4580 18164
rect 4436 18080 4488 18086
rect 4436 18022 4488 18028
rect 4448 17814 4476 18022
rect 4436 17808 4488 17814
rect 4436 17750 4488 17756
rect 4252 17740 4304 17746
rect 4252 17682 4304 17688
rect 4436 17536 4488 17542
rect 4436 17478 4488 17484
rect 4448 17134 4476 17478
rect 4436 17128 4488 17134
rect 4436 17070 4488 17076
rect 4344 16992 4396 16998
rect 4344 16934 4396 16940
rect 4068 16652 4120 16658
rect 4068 16594 4120 16600
rect 4080 15706 4108 16594
rect 4356 15978 4384 16934
rect 4344 15972 4396 15978
rect 4344 15914 4396 15920
rect 4068 15700 4120 15706
rect 4068 15642 4120 15648
rect 4448 15638 4476 17070
rect 4540 16590 4568 18158
rect 5540 18080 5592 18086
rect 5540 18022 5592 18028
rect 5632 18080 5684 18086
rect 5632 18022 5684 18028
rect 5172 17604 5224 17610
rect 5172 17546 5224 17552
rect 4656 17436 4964 17445
rect 4656 17434 4662 17436
rect 4718 17434 4742 17436
rect 4798 17434 4822 17436
rect 4878 17434 4902 17436
rect 4958 17434 4964 17436
rect 4718 17382 4720 17434
rect 4900 17382 4902 17434
rect 4656 17380 4662 17382
rect 4718 17380 4742 17382
rect 4798 17380 4822 17382
rect 4878 17380 4902 17382
rect 4958 17380 4964 17382
rect 4656 17371 4964 17380
rect 4804 17060 4856 17066
rect 4804 17002 4856 17008
rect 4816 16658 4844 17002
rect 4804 16652 4856 16658
rect 4804 16594 4856 16600
rect 4528 16584 4580 16590
rect 4528 16526 4580 16532
rect 4656 16348 4964 16357
rect 4656 16346 4662 16348
rect 4718 16346 4742 16348
rect 4798 16346 4822 16348
rect 4878 16346 4902 16348
rect 4958 16346 4964 16348
rect 4718 16294 4720 16346
rect 4900 16294 4902 16346
rect 4656 16292 4662 16294
rect 4718 16292 4742 16294
rect 4798 16292 4822 16294
rect 4878 16292 4902 16294
rect 4958 16292 4964 16294
rect 4656 16283 4964 16292
rect 5184 16114 5212 17546
rect 5552 16250 5580 18022
rect 5644 17338 5672 18022
rect 5632 17332 5684 17338
rect 5632 17274 5684 17280
rect 5632 16720 5684 16726
rect 5632 16662 5684 16668
rect 5540 16244 5592 16250
rect 5540 16186 5592 16192
rect 5644 16114 5672 16662
rect 5172 16108 5224 16114
rect 5172 16050 5224 16056
rect 5632 16108 5684 16114
rect 5632 16050 5684 16056
rect 4436 15632 4488 15638
rect 4436 15574 4488 15580
rect 4656 15260 4964 15269
rect 4656 15258 4662 15260
rect 4718 15258 4742 15260
rect 4798 15258 4822 15260
rect 4878 15258 4902 15260
rect 4958 15258 4964 15260
rect 4718 15206 4720 15258
rect 4900 15206 4902 15258
rect 4656 15204 4662 15206
rect 4718 15204 4742 15206
rect 4798 15204 4822 15206
rect 4878 15204 4902 15206
rect 4958 15204 4964 15206
rect 4656 15195 4964 15204
rect 4068 14952 4120 14958
rect 4068 14894 4120 14900
rect 4080 14414 4108 14894
rect 4988 14884 5040 14890
rect 4988 14826 5040 14832
rect 4804 14816 4856 14822
rect 4804 14758 4856 14764
rect 4816 14482 4844 14758
rect 5000 14618 5028 14826
rect 4988 14612 5040 14618
rect 4988 14554 5040 14560
rect 4804 14476 4856 14482
rect 4804 14418 4856 14424
rect 4068 14408 4120 14414
rect 4068 14350 4120 14356
rect 4656 14172 4964 14181
rect 4656 14170 4662 14172
rect 4718 14170 4742 14172
rect 4798 14170 4822 14172
rect 4878 14170 4902 14172
rect 4958 14170 4964 14172
rect 4718 14118 4720 14170
rect 4900 14118 4902 14170
rect 4656 14116 4662 14118
rect 4718 14116 4742 14118
rect 4798 14116 4822 14118
rect 4878 14116 4902 14118
rect 4958 14116 4964 14118
rect 4656 14107 4964 14116
rect 3884 14068 3936 14074
rect 3884 14010 3936 14016
rect 4528 13388 4580 13394
rect 4528 13330 4580 13336
rect 2964 12844 3016 12850
rect 2964 12786 3016 12792
rect 3516 12844 3568 12850
rect 3516 12786 3568 12792
rect 3700 12708 3752 12714
rect 3700 12650 3752 12656
rect 3106 12540 3414 12549
rect 3106 12538 3112 12540
rect 3168 12538 3192 12540
rect 3248 12538 3272 12540
rect 3328 12538 3352 12540
rect 3408 12538 3414 12540
rect 3168 12486 3170 12538
rect 3350 12486 3352 12538
rect 3106 12484 3112 12486
rect 3168 12484 3192 12486
rect 3248 12484 3272 12486
rect 3328 12484 3352 12486
rect 3408 12484 3414 12486
rect 3106 12475 3414 12484
rect 3608 12300 3660 12306
rect 3608 12242 3660 12248
rect 3106 11452 3414 11461
rect 3106 11450 3112 11452
rect 3168 11450 3192 11452
rect 3248 11450 3272 11452
rect 3328 11450 3352 11452
rect 3408 11450 3414 11452
rect 3168 11398 3170 11450
rect 3350 11398 3352 11450
rect 3106 11396 3112 11398
rect 3168 11396 3192 11398
rect 3248 11396 3272 11398
rect 3328 11396 3352 11398
rect 3408 11396 3414 11398
rect 3106 11387 3414 11396
rect 3620 11150 3648 12242
rect 3608 11144 3660 11150
rect 3608 11086 3660 11092
rect 3148 11008 3200 11014
rect 3148 10950 3200 10956
rect 3160 10674 3188 10950
rect 3148 10668 3200 10674
rect 3148 10610 3200 10616
rect 3106 10364 3414 10373
rect 3106 10362 3112 10364
rect 3168 10362 3192 10364
rect 3248 10362 3272 10364
rect 3328 10362 3352 10364
rect 3408 10362 3414 10364
rect 3168 10310 3170 10362
rect 3350 10310 3352 10362
rect 3106 10308 3112 10310
rect 3168 10308 3192 10310
rect 3248 10308 3272 10310
rect 3328 10308 3352 10310
rect 3408 10308 3414 10310
rect 3106 10299 3414 10308
rect 2964 9376 3016 9382
rect 2964 9318 3016 9324
rect 2872 9104 2924 9110
rect 2872 9046 2924 9052
rect 2884 8838 2912 9046
rect 2976 9042 3004 9318
rect 3106 9276 3414 9285
rect 3106 9274 3112 9276
rect 3168 9274 3192 9276
rect 3248 9274 3272 9276
rect 3328 9274 3352 9276
rect 3408 9274 3414 9276
rect 3168 9222 3170 9274
rect 3350 9222 3352 9274
rect 3106 9220 3112 9222
rect 3168 9220 3192 9222
rect 3248 9220 3272 9222
rect 3328 9220 3352 9222
rect 3408 9220 3414 9222
rect 3106 9211 3414 9220
rect 2964 9036 3016 9042
rect 2964 8978 3016 8984
rect 3424 9036 3476 9042
rect 3424 8978 3476 8984
rect 2872 8832 2924 8838
rect 2872 8774 2924 8780
rect 2688 8356 2740 8362
rect 2688 8298 2740 8304
rect 2596 8084 2648 8090
rect 2596 8026 2648 8032
rect 2136 7404 2188 7410
rect 2136 7346 2188 7352
rect 572 6928 624 6934
rect 572 6870 624 6876
rect 584 5778 612 6870
rect 1952 6656 2004 6662
rect 1952 6598 2004 6604
rect 1556 6556 1864 6565
rect 1556 6554 1562 6556
rect 1618 6554 1642 6556
rect 1698 6554 1722 6556
rect 1778 6554 1802 6556
rect 1858 6554 1864 6556
rect 1618 6502 1620 6554
rect 1800 6502 1802 6554
rect 1556 6500 1562 6502
rect 1618 6500 1642 6502
rect 1698 6500 1722 6502
rect 1778 6500 1802 6502
rect 1858 6500 1864 6502
rect 1556 6491 1864 6500
rect 1964 6458 1992 6598
rect 1952 6452 2004 6458
rect 1952 6394 2004 6400
rect 572 5772 624 5778
rect 572 5714 624 5720
rect 940 5704 992 5710
rect 940 5646 992 5652
rect 756 4072 808 4078
rect 756 4014 808 4020
rect 768 3738 796 4014
rect 952 4010 980 5646
rect 1556 5468 1864 5477
rect 1556 5466 1562 5468
rect 1618 5466 1642 5468
rect 1698 5466 1722 5468
rect 1778 5466 1802 5468
rect 1858 5466 1864 5468
rect 1618 5414 1620 5466
rect 1800 5414 1802 5466
rect 1556 5412 1562 5414
rect 1618 5412 1642 5414
rect 1698 5412 1722 5414
rect 1778 5412 1802 5414
rect 1858 5412 1864 5414
rect 1556 5403 1864 5412
rect 2148 5370 2176 7346
rect 2608 7342 2636 8026
rect 2884 8022 2912 8774
rect 3436 8634 3464 8978
rect 3424 8628 3476 8634
rect 3424 8570 3476 8576
rect 3106 8188 3414 8197
rect 3106 8186 3112 8188
rect 3168 8186 3192 8188
rect 3248 8186 3272 8188
rect 3328 8186 3352 8188
rect 3408 8186 3414 8188
rect 3168 8134 3170 8186
rect 3350 8134 3352 8186
rect 3106 8132 3112 8134
rect 3168 8132 3192 8134
rect 3248 8132 3272 8134
rect 3328 8132 3352 8134
rect 3408 8132 3414 8134
rect 3106 8123 3414 8132
rect 2872 8016 2924 8022
rect 2872 7958 2924 7964
rect 2780 7404 2832 7410
rect 2780 7346 2832 7352
rect 2596 7336 2648 7342
rect 2596 7278 2648 7284
rect 2792 6914 2820 7346
rect 2884 7206 2912 7958
rect 3620 7342 3648 11086
rect 3712 10742 3740 12650
rect 4540 11558 4568 13330
rect 4656 13084 4964 13093
rect 4656 13082 4662 13084
rect 4718 13082 4742 13084
rect 4798 13082 4822 13084
rect 4878 13082 4902 13084
rect 4958 13082 4964 13084
rect 4718 13030 4720 13082
rect 4900 13030 4902 13082
rect 4656 13028 4662 13030
rect 4718 13028 4742 13030
rect 4798 13028 4822 13030
rect 4878 13028 4902 13030
rect 4958 13028 4964 13030
rect 4656 13019 4964 13028
rect 5000 12714 5028 14554
rect 5184 14482 5212 16050
rect 5172 14476 5224 14482
rect 5172 14418 5224 14424
rect 5184 13530 5212 14418
rect 5632 14068 5684 14074
rect 5632 14010 5684 14016
rect 5644 13870 5672 14010
rect 5736 13938 5764 18226
rect 5828 17202 5856 18294
rect 6828 18216 6880 18222
rect 6828 18158 6880 18164
rect 6206 17980 6514 17989
rect 6206 17978 6212 17980
rect 6268 17978 6292 17980
rect 6348 17978 6372 17980
rect 6428 17978 6452 17980
rect 6508 17978 6514 17980
rect 6268 17926 6270 17978
rect 6450 17926 6452 17978
rect 6206 17924 6212 17926
rect 6268 17924 6292 17926
rect 6348 17924 6372 17926
rect 6428 17924 6452 17926
rect 6508 17924 6514 17926
rect 6206 17915 6514 17924
rect 5816 17196 5868 17202
rect 5816 17138 5868 17144
rect 5908 17128 5960 17134
rect 5908 17070 5960 17076
rect 5816 16516 5868 16522
rect 5816 16458 5868 16464
rect 5828 14958 5856 16458
rect 5920 15162 5948 17070
rect 6206 16892 6514 16901
rect 6206 16890 6212 16892
rect 6268 16890 6292 16892
rect 6348 16890 6372 16892
rect 6428 16890 6452 16892
rect 6508 16890 6514 16892
rect 6268 16838 6270 16890
rect 6450 16838 6452 16890
rect 6206 16836 6212 16838
rect 6268 16836 6292 16838
rect 6348 16836 6372 16838
rect 6428 16836 6452 16838
rect 6508 16836 6514 16838
rect 6206 16827 6514 16836
rect 6552 15972 6604 15978
rect 6552 15914 6604 15920
rect 6206 15804 6514 15813
rect 6206 15802 6212 15804
rect 6268 15802 6292 15804
rect 6348 15802 6372 15804
rect 6428 15802 6452 15804
rect 6508 15802 6514 15804
rect 6268 15750 6270 15802
rect 6450 15750 6452 15802
rect 6206 15748 6212 15750
rect 6268 15748 6292 15750
rect 6348 15748 6372 15750
rect 6428 15748 6452 15750
rect 6508 15748 6514 15750
rect 6206 15739 6514 15748
rect 5908 15156 5960 15162
rect 5908 15098 5960 15104
rect 5816 14952 5868 14958
rect 5816 14894 5868 14900
rect 6206 14716 6514 14725
rect 6206 14714 6212 14716
rect 6268 14714 6292 14716
rect 6348 14714 6372 14716
rect 6428 14714 6452 14716
rect 6508 14714 6514 14716
rect 6268 14662 6270 14714
rect 6450 14662 6452 14714
rect 6206 14660 6212 14662
rect 6268 14660 6292 14662
rect 6348 14660 6372 14662
rect 6428 14660 6452 14662
rect 6508 14660 6514 14662
rect 6206 14651 6514 14660
rect 6564 14550 6592 15914
rect 6840 15706 6868 18158
rect 7012 17536 7064 17542
rect 7012 17478 7064 17484
rect 7024 16726 7052 17478
rect 7012 16720 7064 16726
rect 7012 16662 7064 16668
rect 7024 16046 7052 16662
rect 7116 16522 7144 19200
rect 7756 18524 8064 18533
rect 7756 18522 7762 18524
rect 7818 18522 7842 18524
rect 7898 18522 7922 18524
rect 7978 18522 8002 18524
rect 8058 18522 8064 18524
rect 7818 18470 7820 18522
rect 8000 18470 8002 18522
rect 7756 18468 7762 18470
rect 7818 18468 7842 18470
rect 7898 18468 7922 18470
rect 7978 18468 8002 18470
rect 8058 18468 8064 18470
rect 7756 18459 8064 18468
rect 9864 18352 9916 18358
rect 9864 18294 9916 18300
rect 8208 18284 8260 18290
rect 8208 18226 8260 18232
rect 7564 18080 7616 18086
rect 7564 18022 7616 18028
rect 8116 18080 8168 18086
rect 8116 18022 8168 18028
rect 7576 17814 7604 18022
rect 7564 17808 7616 17814
rect 7564 17750 7616 17756
rect 7756 17436 8064 17445
rect 7756 17434 7762 17436
rect 7818 17434 7842 17436
rect 7898 17434 7922 17436
rect 7978 17434 8002 17436
rect 8058 17434 8064 17436
rect 7818 17382 7820 17434
rect 8000 17382 8002 17434
rect 7756 17380 7762 17382
rect 7818 17380 7842 17382
rect 7898 17380 7922 17382
rect 7978 17380 8002 17382
rect 8058 17380 8064 17382
rect 7756 17371 8064 17380
rect 7380 17060 7432 17066
rect 7380 17002 7432 17008
rect 7392 16708 7420 17002
rect 7472 16720 7524 16726
rect 7392 16680 7472 16708
rect 7472 16662 7524 16668
rect 7104 16516 7156 16522
rect 7104 16458 7156 16464
rect 7012 16040 7064 16046
rect 7012 15982 7064 15988
rect 6828 15700 6880 15706
rect 6828 15642 6880 15648
rect 6644 15020 6696 15026
rect 6644 14962 6696 14968
rect 6552 14544 6604 14550
rect 6552 14486 6604 14492
rect 6656 14414 6684 14962
rect 6920 14884 6972 14890
rect 6920 14826 6972 14832
rect 6644 14408 6696 14414
rect 6644 14350 6696 14356
rect 5724 13932 5776 13938
rect 5724 13874 5776 13880
rect 5632 13864 5684 13870
rect 5632 13806 5684 13812
rect 5172 13524 5224 13530
rect 5172 13466 5224 13472
rect 5184 12782 5212 13466
rect 5644 13394 5672 13806
rect 5736 13530 5764 13874
rect 6206 13628 6514 13637
rect 6206 13626 6212 13628
rect 6268 13626 6292 13628
rect 6348 13626 6372 13628
rect 6428 13626 6452 13628
rect 6508 13626 6514 13628
rect 6268 13574 6270 13626
rect 6450 13574 6452 13626
rect 6206 13572 6212 13574
rect 6268 13572 6292 13574
rect 6348 13572 6372 13574
rect 6428 13572 6452 13574
rect 6508 13572 6514 13574
rect 6206 13563 6514 13572
rect 5724 13524 5776 13530
rect 5724 13466 5776 13472
rect 6656 13462 6684 14350
rect 6932 14074 6960 14826
rect 7484 14482 7512 16662
rect 7756 16348 8064 16357
rect 7756 16346 7762 16348
rect 7818 16346 7842 16348
rect 7898 16346 7922 16348
rect 7978 16346 8002 16348
rect 8058 16346 8064 16348
rect 7818 16294 7820 16346
rect 8000 16294 8002 16346
rect 7756 16292 7762 16294
rect 7818 16292 7842 16294
rect 7898 16292 7922 16294
rect 7978 16292 8002 16294
rect 8058 16292 8064 16294
rect 7756 16283 8064 16292
rect 8128 16130 8156 18022
rect 8220 16810 8248 18226
rect 8760 18216 8812 18222
rect 8760 18158 8812 18164
rect 8772 17338 8800 18158
rect 9220 18148 9272 18154
rect 9220 18090 9272 18096
rect 9128 18080 9180 18086
rect 9128 18022 9180 18028
rect 8760 17332 8812 17338
rect 8760 17274 8812 17280
rect 8220 16782 8340 16810
rect 8312 16538 8340 16782
rect 9140 16658 9168 18022
rect 9232 17610 9260 18090
rect 9306 17980 9614 17989
rect 9306 17978 9312 17980
rect 9368 17978 9392 17980
rect 9448 17978 9472 17980
rect 9528 17978 9552 17980
rect 9608 17978 9614 17980
rect 9368 17926 9370 17978
rect 9550 17926 9552 17978
rect 9306 17924 9312 17926
rect 9368 17924 9392 17926
rect 9448 17924 9472 17926
rect 9528 17924 9552 17926
rect 9608 17924 9614 17926
rect 9306 17915 9614 17924
rect 9876 17814 9904 18294
rect 9968 18170 9996 19200
rect 10856 18524 11164 18533
rect 10856 18522 10862 18524
rect 10918 18522 10942 18524
rect 10998 18522 11022 18524
rect 11078 18522 11102 18524
rect 11158 18522 11164 18524
rect 10918 18470 10920 18522
rect 11100 18470 11102 18522
rect 10856 18468 10862 18470
rect 10918 18468 10942 18470
rect 10998 18468 11022 18470
rect 11078 18468 11102 18470
rect 11158 18468 11164 18470
rect 10856 18459 11164 18468
rect 11336 18216 11388 18222
rect 9968 18142 10088 18170
rect 11336 18158 11388 18164
rect 9956 18080 10008 18086
rect 9956 18022 10008 18028
rect 9864 17808 9916 17814
rect 9864 17750 9916 17756
rect 9220 17604 9272 17610
rect 9220 17546 9272 17552
rect 9232 17066 9260 17546
rect 9220 17060 9272 17066
rect 9220 17002 9272 17008
rect 9306 16892 9614 16901
rect 9306 16890 9312 16892
rect 9368 16890 9392 16892
rect 9448 16890 9472 16892
rect 9528 16890 9552 16892
rect 9608 16890 9614 16892
rect 9368 16838 9370 16890
rect 9550 16838 9552 16890
rect 9306 16836 9312 16838
rect 9368 16836 9392 16838
rect 9448 16836 9472 16838
rect 9528 16836 9552 16838
rect 9608 16836 9614 16838
rect 9306 16827 9614 16836
rect 9968 16658 9996 18022
rect 9128 16652 9180 16658
rect 9128 16594 9180 16600
rect 9864 16652 9916 16658
rect 9864 16594 9916 16600
rect 9956 16652 10008 16658
rect 9956 16594 10008 16600
rect 8036 16102 8156 16130
rect 8220 16510 8340 16538
rect 8036 15910 8064 16102
rect 8024 15904 8076 15910
rect 8024 15846 8076 15852
rect 8036 15638 8064 15846
rect 8024 15632 8076 15638
rect 8024 15574 8076 15580
rect 7656 15496 7708 15502
rect 7656 15438 7708 15444
rect 7564 14816 7616 14822
rect 7564 14758 7616 14764
rect 7472 14476 7524 14482
rect 7472 14418 7524 14424
rect 7012 14272 7064 14278
rect 7012 14214 7064 14220
rect 6920 14068 6972 14074
rect 6920 14010 6972 14016
rect 6644 13456 6696 13462
rect 6644 13398 6696 13404
rect 5632 13388 5684 13394
rect 5632 13330 5684 13336
rect 6736 13320 6788 13326
rect 6736 13262 6788 13268
rect 5172 12776 5224 12782
rect 5172 12718 5224 12724
rect 6748 12714 6776 13262
rect 7024 12782 7052 14214
rect 7472 12844 7524 12850
rect 7472 12786 7524 12792
rect 7012 12776 7064 12782
rect 7012 12718 7064 12724
rect 4988 12708 5040 12714
rect 4988 12650 5040 12656
rect 6736 12708 6788 12714
rect 6736 12650 6788 12656
rect 4656 11996 4964 12005
rect 4656 11994 4662 11996
rect 4718 11994 4742 11996
rect 4798 11994 4822 11996
rect 4878 11994 4902 11996
rect 4958 11994 4964 11996
rect 4718 11942 4720 11994
rect 4900 11942 4902 11994
rect 4656 11940 4662 11942
rect 4718 11940 4742 11942
rect 4798 11940 4822 11942
rect 4878 11940 4902 11942
rect 4958 11940 4964 11942
rect 4656 11931 4964 11940
rect 4528 11552 4580 11558
rect 4528 11494 4580 11500
rect 3792 11212 3844 11218
rect 3792 11154 3844 11160
rect 4068 11212 4120 11218
rect 4068 11154 4120 11160
rect 3700 10736 3752 10742
rect 3700 10678 3752 10684
rect 3712 10062 3740 10678
rect 3804 10266 3832 11154
rect 3884 10668 3936 10674
rect 3884 10610 3936 10616
rect 3792 10260 3844 10266
rect 3792 10202 3844 10208
rect 3896 10146 3924 10610
rect 4080 10470 4108 11154
rect 4252 10600 4304 10606
rect 4252 10542 4304 10548
rect 4068 10464 4120 10470
rect 4068 10406 4120 10412
rect 3804 10130 3924 10146
rect 3792 10124 3924 10130
rect 3844 10118 3924 10124
rect 3792 10066 3844 10072
rect 3700 10056 3752 10062
rect 3700 9998 3752 10004
rect 3804 7410 3832 10066
rect 4080 9586 4108 10406
rect 4264 10062 4292 10542
rect 4344 10532 4396 10538
rect 4344 10474 4396 10480
rect 4252 10056 4304 10062
rect 4252 9998 4304 10004
rect 4356 9654 4384 10474
rect 4344 9648 4396 9654
rect 4344 9590 4396 9596
rect 4068 9580 4120 9586
rect 4068 9522 4120 9528
rect 4356 9466 4384 9590
rect 4264 9438 4384 9466
rect 4264 7546 4292 9438
rect 4344 9376 4396 9382
rect 4344 9318 4396 9324
rect 4356 9178 4384 9318
rect 4344 9172 4396 9178
rect 4344 9114 4396 9120
rect 4344 8968 4396 8974
rect 4344 8910 4396 8916
rect 4356 8362 4384 8910
rect 4436 8900 4488 8906
rect 4436 8842 4488 8848
rect 4344 8356 4396 8362
rect 4344 8298 4396 8304
rect 4252 7540 4304 7546
rect 4252 7482 4304 7488
rect 3792 7404 3844 7410
rect 3792 7346 3844 7352
rect 4356 7342 4384 8298
rect 3608 7336 3660 7342
rect 3608 7278 3660 7284
rect 4344 7336 4396 7342
rect 4344 7278 4396 7284
rect 2872 7200 2924 7206
rect 2872 7142 2924 7148
rect 2700 6886 2820 6914
rect 2320 5908 2372 5914
rect 2320 5850 2372 5856
rect 2136 5364 2188 5370
rect 2136 5306 2188 5312
rect 1952 5228 2004 5234
rect 1952 5170 2004 5176
rect 1964 4826 1992 5170
rect 2136 5024 2188 5030
rect 2056 4984 2136 5012
rect 1952 4820 2004 4826
rect 1952 4762 2004 4768
rect 1952 4684 2004 4690
rect 1952 4626 2004 4632
rect 1556 4380 1864 4389
rect 1556 4378 1562 4380
rect 1618 4378 1642 4380
rect 1698 4378 1722 4380
rect 1778 4378 1802 4380
rect 1858 4378 1864 4380
rect 1618 4326 1620 4378
rect 1800 4326 1802 4378
rect 1556 4324 1562 4326
rect 1618 4324 1642 4326
rect 1698 4324 1722 4326
rect 1778 4324 1802 4326
rect 1858 4324 1864 4326
rect 1556 4315 1864 4324
rect 1964 4214 1992 4626
rect 2056 4486 2084 4984
rect 2136 4966 2188 4972
rect 2044 4480 2096 4486
rect 2044 4422 2096 4428
rect 1952 4208 2004 4214
rect 1952 4150 2004 4156
rect 1952 4072 2004 4078
rect 2056 4060 2084 4422
rect 2004 4032 2084 4060
rect 1952 4014 2004 4020
rect 940 4004 992 4010
rect 940 3946 992 3952
rect 756 3732 808 3738
rect 756 3674 808 3680
rect 940 3596 992 3602
rect 940 3538 992 3544
rect 952 2650 980 3538
rect 1556 3292 1864 3301
rect 1556 3290 1562 3292
rect 1618 3290 1642 3292
rect 1698 3290 1722 3292
rect 1778 3290 1802 3292
rect 1858 3290 1864 3292
rect 1618 3238 1620 3290
rect 1800 3238 1802 3290
rect 1556 3236 1562 3238
rect 1618 3236 1642 3238
rect 1698 3236 1722 3238
rect 1778 3236 1802 3238
rect 1858 3236 1864 3238
rect 1556 3227 1864 3236
rect 1492 2984 1544 2990
rect 1492 2926 1544 2932
rect 940 2644 992 2650
rect 940 2586 992 2592
rect 1504 2582 1532 2926
rect 1768 2848 1820 2854
rect 1768 2790 1820 2796
rect 1780 2650 1808 2790
rect 1768 2644 1820 2650
rect 1768 2586 1820 2592
rect 1492 2576 1544 2582
rect 1492 2518 1544 2524
rect 1964 2446 1992 4014
rect 2332 4010 2360 5850
rect 2700 4010 2728 6886
rect 2884 6186 2912 7142
rect 3106 7100 3414 7109
rect 3106 7098 3112 7100
rect 3168 7098 3192 7100
rect 3248 7098 3272 7100
rect 3328 7098 3352 7100
rect 3408 7098 3414 7100
rect 3168 7046 3170 7098
rect 3350 7046 3352 7098
rect 3106 7044 3112 7046
rect 3168 7044 3192 7046
rect 3248 7044 3272 7046
rect 3328 7044 3352 7046
rect 3408 7044 3414 7046
rect 3106 7035 3414 7044
rect 4252 6928 4304 6934
rect 4252 6870 4304 6876
rect 4160 6860 4212 6866
rect 4160 6802 4212 6808
rect 2964 6316 3016 6322
rect 2964 6258 3016 6264
rect 2872 6180 2924 6186
rect 2872 6122 2924 6128
rect 2884 5846 2912 6122
rect 2872 5840 2924 5846
rect 2872 5782 2924 5788
rect 2884 5574 2912 5782
rect 2872 5568 2924 5574
rect 2872 5510 2924 5516
rect 2976 4826 3004 6258
rect 3516 6180 3568 6186
rect 3516 6122 3568 6128
rect 3106 6012 3414 6021
rect 3106 6010 3112 6012
rect 3168 6010 3192 6012
rect 3248 6010 3272 6012
rect 3328 6010 3352 6012
rect 3408 6010 3414 6012
rect 3168 5958 3170 6010
rect 3350 5958 3352 6010
rect 3106 5956 3112 5958
rect 3168 5956 3192 5958
rect 3248 5956 3272 5958
rect 3328 5956 3352 5958
rect 3408 5956 3414 5958
rect 3106 5947 3414 5956
rect 3528 5778 3556 6122
rect 3516 5772 3568 5778
rect 3516 5714 3568 5720
rect 3106 4924 3414 4933
rect 3106 4922 3112 4924
rect 3168 4922 3192 4924
rect 3248 4922 3272 4924
rect 3328 4922 3352 4924
rect 3408 4922 3414 4924
rect 3168 4870 3170 4922
rect 3350 4870 3352 4922
rect 3106 4868 3112 4870
rect 3168 4868 3192 4870
rect 3248 4868 3272 4870
rect 3328 4868 3352 4870
rect 3408 4868 3414 4870
rect 3106 4859 3414 4868
rect 2964 4820 3016 4826
rect 2964 4762 3016 4768
rect 2780 4684 2832 4690
rect 2780 4626 2832 4632
rect 3332 4684 3384 4690
rect 3332 4626 3384 4632
rect 2320 4004 2372 4010
rect 2320 3946 2372 3952
rect 2688 4004 2740 4010
rect 2688 3946 2740 3952
rect 2136 2848 2188 2854
rect 2136 2790 2188 2796
rect 2148 2650 2176 2790
rect 2136 2644 2188 2650
rect 2136 2586 2188 2592
rect 2332 2514 2360 3946
rect 2700 2990 2728 3946
rect 2688 2984 2740 2990
rect 2688 2926 2740 2932
rect 2792 2650 2820 4626
rect 3344 4282 3372 4626
rect 3332 4276 3384 4282
rect 3332 4218 3384 4224
rect 3528 4078 3556 5714
rect 4172 4826 4200 6802
rect 4264 6322 4292 6870
rect 4252 6316 4304 6322
rect 4252 6258 4304 6264
rect 4252 5704 4304 5710
rect 4252 5646 4304 5652
rect 4160 4820 4212 4826
rect 4160 4762 4212 4768
rect 3884 4684 3936 4690
rect 3884 4626 3936 4632
rect 3896 4146 3924 4626
rect 4160 4548 4212 4554
rect 4160 4490 4212 4496
rect 3884 4140 3936 4146
rect 3884 4082 3936 4088
rect 3516 4072 3568 4078
rect 3516 4014 3568 4020
rect 3106 3836 3414 3845
rect 3106 3834 3112 3836
rect 3168 3834 3192 3836
rect 3248 3834 3272 3836
rect 3328 3834 3352 3836
rect 3408 3834 3414 3836
rect 3168 3782 3170 3834
rect 3350 3782 3352 3834
rect 3106 3780 3112 3782
rect 3168 3780 3192 3782
rect 3248 3780 3272 3782
rect 3328 3780 3352 3782
rect 3408 3780 3414 3782
rect 3106 3771 3414 3780
rect 2872 3052 2924 3058
rect 2872 2994 2924 3000
rect 2780 2644 2832 2650
rect 2780 2586 2832 2592
rect 2320 2508 2372 2514
rect 2320 2450 2372 2456
rect 1952 2440 2004 2446
rect 1952 2382 2004 2388
rect 1556 2204 1864 2213
rect 1556 2202 1562 2204
rect 1618 2202 1642 2204
rect 1698 2202 1722 2204
rect 1778 2202 1802 2204
rect 1858 2202 1864 2204
rect 1618 2150 1620 2202
rect 1800 2150 1802 2202
rect 1556 2148 1562 2150
rect 1618 2148 1642 2150
rect 1698 2148 1722 2150
rect 1778 2148 1802 2150
rect 1858 2148 1864 2150
rect 1556 2139 1864 2148
rect 2884 1970 2912 2994
rect 3106 2748 3414 2757
rect 3106 2746 3112 2748
rect 3168 2746 3192 2748
rect 3248 2746 3272 2748
rect 3328 2746 3352 2748
rect 3408 2746 3414 2748
rect 3168 2694 3170 2746
rect 3350 2694 3352 2746
rect 3106 2692 3112 2694
rect 3168 2692 3192 2694
rect 3248 2692 3272 2694
rect 3328 2692 3352 2694
rect 3408 2692 3414 2694
rect 3106 2683 3414 2692
rect 3332 2644 3384 2650
rect 3332 2586 3384 2592
rect 2872 1964 2924 1970
rect 2872 1906 2924 1912
rect 3344 1902 3372 2586
rect 3528 1902 3556 4014
rect 3896 3738 3924 4082
rect 3884 3732 3936 3738
rect 3884 3674 3936 3680
rect 4172 3602 4200 4490
rect 4142 3596 4200 3602
rect 4194 3556 4200 3596
rect 4142 3538 4194 3544
rect 4264 3516 4292 5646
rect 4448 5522 4476 8842
rect 4540 8022 4568 11494
rect 4656 10908 4964 10917
rect 4656 10906 4662 10908
rect 4718 10906 4742 10908
rect 4798 10906 4822 10908
rect 4878 10906 4902 10908
rect 4958 10906 4964 10908
rect 4718 10854 4720 10906
rect 4900 10854 4902 10906
rect 4656 10852 4662 10854
rect 4718 10852 4742 10854
rect 4798 10852 4822 10854
rect 4878 10852 4902 10854
rect 4958 10852 4964 10854
rect 4656 10843 4964 10852
rect 5000 10742 5028 12650
rect 5816 12640 5868 12646
rect 5816 12582 5868 12588
rect 5828 12374 5856 12582
rect 6206 12540 6514 12549
rect 6206 12538 6212 12540
rect 6268 12538 6292 12540
rect 6348 12538 6372 12540
rect 6428 12538 6452 12540
rect 6508 12538 6514 12540
rect 6268 12486 6270 12538
rect 6450 12486 6452 12538
rect 6206 12484 6212 12486
rect 6268 12484 6292 12486
rect 6348 12484 6372 12486
rect 6428 12484 6452 12486
rect 6508 12484 6514 12486
rect 6206 12475 6514 12484
rect 5816 12368 5868 12374
rect 5816 12310 5868 12316
rect 5264 12300 5316 12306
rect 5264 12242 5316 12248
rect 5276 11218 5304 12242
rect 5540 12232 5592 12238
rect 5540 12174 5592 12180
rect 5552 11354 5580 12174
rect 6736 12096 6788 12102
rect 6736 12038 6788 12044
rect 6206 11452 6514 11461
rect 6206 11450 6212 11452
rect 6268 11450 6292 11452
rect 6348 11450 6372 11452
rect 6428 11450 6452 11452
rect 6508 11450 6514 11452
rect 6268 11398 6270 11450
rect 6450 11398 6452 11450
rect 6206 11396 6212 11398
rect 6268 11396 6292 11398
rect 6348 11396 6372 11398
rect 6428 11396 6452 11398
rect 6508 11396 6514 11398
rect 6206 11387 6514 11396
rect 5540 11348 5592 11354
rect 5540 11290 5592 11296
rect 5264 11212 5316 11218
rect 5264 11154 5316 11160
rect 6644 10804 6696 10810
rect 6644 10746 6696 10752
rect 4988 10736 5040 10742
rect 4988 10678 5040 10684
rect 6552 10600 6604 10606
rect 6552 10542 6604 10548
rect 6206 10364 6514 10373
rect 6206 10362 6212 10364
rect 6268 10362 6292 10364
rect 6348 10362 6372 10364
rect 6428 10362 6452 10364
rect 6508 10362 6514 10364
rect 6268 10310 6270 10362
rect 6450 10310 6452 10362
rect 6206 10308 6212 10310
rect 6268 10308 6292 10310
rect 6348 10308 6372 10310
rect 6428 10308 6452 10310
rect 6508 10308 6514 10310
rect 6206 10299 6514 10308
rect 6564 10266 6592 10542
rect 6552 10260 6604 10266
rect 6552 10202 6604 10208
rect 6656 10146 6684 10746
rect 6748 10606 6776 12038
rect 7484 11830 7512 12786
rect 7576 11898 7604 14758
rect 7668 14618 7696 15438
rect 7756 15260 8064 15269
rect 7756 15258 7762 15260
rect 7818 15258 7842 15260
rect 7898 15258 7922 15260
rect 7978 15258 8002 15260
rect 8058 15258 8064 15260
rect 7818 15206 7820 15258
rect 8000 15206 8002 15258
rect 7756 15204 7762 15206
rect 7818 15204 7842 15206
rect 7898 15204 7922 15206
rect 7978 15204 8002 15206
rect 8058 15204 8064 15206
rect 7756 15195 8064 15204
rect 8220 15162 8248 16510
rect 9036 15972 9088 15978
rect 9036 15914 9088 15920
rect 8300 15632 8352 15638
rect 8300 15574 8352 15580
rect 8208 15156 8260 15162
rect 8208 15098 8260 15104
rect 8116 14952 8168 14958
rect 8116 14894 8168 14900
rect 7656 14612 7708 14618
rect 7656 14554 7708 14560
rect 8128 14414 8156 14894
rect 8116 14408 8168 14414
rect 8116 14350 8168 14356
rect 7756 14172 8064 14181
rect 7756 14170 7762 14172
rect 7818 14170 7842 14172
rect 7898 14170 7922 14172
rect 7978 14170 8002 14172
rect 8058 14170 8064 14172
rect 7818 14118 7820 14170
rect 8000 14118 8002 14170
rect 7756 14116 7762 14118
rect 7818 14116 7842 14118
rect 7898 14116 7922 14118
rect 7978 14116 8002 14118
rect 8058 14116 8064 14118
rect 7756 14107 8064 14116
rect 7748 13864 7800 13870
rect 7748 13806 7800 13812
rect 7760 13462 7788 13806
rect 7748 13456 7800 13462
rect 7748 13398 7800 13404
rect 7656 13320 7708 13326
rect 7656 13262 7708 13268
rect 7668 12850 7696 13262
rect 7756 13084 8064 13093
rect 7756 13082 7762 13084
rect 7818 13082 7842 13084
rect 7898 13082 7922 13084
rect 7978 13082 8002 13084
rect 8058 13082 8064 13084
rect 7818 13030 7820 13082
rect 8000 13030 8002 13082
rect 7756 13028 7762 13030
rect 7818 13028 7842 13030
rect 7898 13028 7922 13030
rect 7978 13028 8002 13030
rect 8058 13028 8064 13030
rect 7756 13019 8064 13028
rect 8128 12900 8156 14350
rect 8208 14068 8260 14074
rect 8208 14010 8260 14016
rect 8036 12872 8156 12900
rect 7656 12844 7708 12850
rect 7656 12786 7708 12792
rect 8036 12442 8064 12872
rect 8116 12640 8168 12646
rect 8116 12582 8168 12588
rect 8024 12436 8076 12442
rect 8024 12378 8076 12384
rect 7756 11996 8064 12005
rect 7756 11994 7762 11996
rect 7818 11994 7842 11996
rect 7898 11994 7922 11996
rect 7978 11994 8002 11996
rect 8058 11994 8064 11996
rect 7818 11942 7820 11994
rect 8000 11942 8002 11994
rect 7756 11940 7762 11942
rect 7818 11940 7842 11942
rect 7898 11940 7922 11942
rect 7978 11940 8002 11942
rect 8058 11940 8064 11942
rect 7756 11931 8064 11940
rect 7564 11892 7616 11898
rect 7564 11834 7616 11840
rect 7472 11824 7524 11830
rect 7472 11766 7524 11772
rect 7104 11688 7156 11694
rect 7104 11630 7156 11636
rect 7380 11688 7432 11694
rect 7380 11630 7432 11636
rect 8024 11688 8076 11694
rect 8024 11630 8076 11636
rect 7012 11552 7064 11558
rect 7012 11494 7064 11500
rect 6920 10668 6972 10674
rect 6920 10610 6972 10616
rect 6736 10600 6788 10606
rect 6736 10542 6788 10548
rect 5356 10124 5408 10130
rect 5356 10066 5408 10072
rect 6564 10118 6684 10146
rect 4656 9820 4964 9829
rect 4656 9818 4662 9820
rect 4718 9818 4742 9820
rect 4798 9818 4822 9820
rect 4878 9818 4902 9820
rect 4958 9818 4964 9820
rect 4718 9766 4720 9818
rect 4900 9766 4902 9818
rect 4656 9764 4662 9766
rect 4718 9764 4742 9766
rect 4798 9764 4822 9766
rect 4878 9764 4902 9766
rect 4958 9764 4964 9766
rect 4656 9755 4964 9764
rect 5368 9178 5396 10066
rect 6564 10062 6592 10118
rect 6552 10056 6604 10062
rect 6552 9998 6604 10004
rect 6828 10056 6880 10062
rect 6828 9998 6880 10004
rect 6206 9276 6514 9285
rect 6206 9274 6212 9276
rect 6268 9274 6292 9276
rect 6348 9274 6372 9276
rect 6428 9274 6452 9276
rect 6508 9274 6514 9276
rect 6268 9222 6270 9274
rect 6450 9222 6452 9274
rect 6206 9220 6212 9222
rect 6268 9220 6292 9222
rect 6348 9220 6372 9222
rect 6428 9220 6452 9222
rect 6508 9220 6514 9222
rect 6206 9211 6514 9220
rect 5356 9172 5408 9178
rect 5356 9114 5408 9120
rect 5540 8832 5592 8838
rect 5540 8774 5592 8780
rect 4656 8732 4964 8741
rect 4656 8730 4662 8732
rect 4718 8730 4742 8732
rect 4798 8730 4822 8732
rect 4878 8730 4902 8732
rect 4958 8730 4964 8732
rect 4718 8678 4720 8730
rect 4900 8678 4902 8730
rect 4656 8676 4662 8678
rect 4718 8676 4742 8678
rect 4798 8676 4822 8678
rect 4878 8676 4902 8678
rect 4958 8676 4964 8678
rect 4656 8667 4964 8676
rect 5552 8430 5580 8774
rect 5540 8424 5592 8430
rect 5540 8366 5592 8372
rect 5264 8356 5316 8362
rect 5264 8298 5316 8304
rect 4528 8016 4580 8022
rect 4528 7958 4580 7964
rect 5276 7954 5304 8298
rect 5448 8084 5500 8090
rect 5552 8072 5580 8366
rect 6564 8362 6592 9998
rect 6840 9518 6868 9998
rect 6828 9512 6880 9518
rect 6828 9454 6880 9460
rect 6552 8356 6604 8362
rect 6552 8298 6604 8304
rect 6206 8188 6514 8197
rect 6206 8186 6212 8188
rect 6268 8186 6292 8188
rect 6348 8186 6372 8188
rect 6428 8186 6452 8188
rect 6508 8186 6514 8188
rect 6268 8134 6270 8186
rect 6450 8134 6452 8186
rect 6206 8132 6212 8134
rect 6268 8132 6292 8134
rect 6348 8132 6372 8134
rect 6428 8132 6452 8134
rect 6508 8132 6514 8134
rect 6206 8123 6514 8132
rect 5500 8044 5580 8072
rect 5448 8026 5500 8032
rect 5264 7948 5316 7954
rect 5264 7890 5316 7896
rect 4656 7644 4964 7653
rect 4656 7642 4662 7644
rect 4718 7642 4742 7644
rect 4798 7642 4822 7644
rect 4878 7642 4902 7644
rect 4958 7642 4964 7644
rect 4718 7590 4720 7642
rect 4900 7590 4902 7642
rect 4656 7588 4662 7590
rect 4718 7588 4742 7590
rect 4798 7588 4822 7590
rect 4878 7588 4902 7590
rect 4958 7588 4964 7590
rect 4656 7579 4964 7588
rect 5264 6860 5316 6866
rect 5264 6802 5316 6808
rect 4656 6556 4964 6565
rect 4656 6554 4662 6556
rect 4718 6554 4742 6556
rect 4798 6554 4822 6556
rect 4878 6554 4902 6556
rect 4958 6554 4964 6556
rect 4718 6502 4720 6554
rect 4900 6502 4902 6554
rect 4656 6500 4662 6502
rect 4718 6500 4742 6502
rect 4798 6500 4822 6502
rect 4878 6500 4902 6502
rect 4958 6500 4964 6502
rect 4656 6491 4964 6500
rect 4528 6180 4580 6186
rect 4528 6122 4580 6128
rect 4356 5494 4476 5522
rect 4356 4078 4384 5494
rect 4540 4826 4568 6122
rect 4804 6112 4856 6118
rect 4804 6054 4856 6060
rect 4816 5778 4844 6054
rect 5276 5914 5304 6802
rect 5552 6322 5580 8044
rect 5724 7880 5776 7886
rect 5724 7822 5776 7828
rect 5736 6730 5764 7822
rect 5816 7268 5868 7274
rect 5816 7210 5868 7216
rect 5828 6866 5856 7210
rect 5908 7200 5960 7206
rect 5908 7142 5960 7148
rect 5816 6860 5868 6866
rect 5816 6802 5868 6808
rect 5724 6724 5776 6730
rect 5724 6666 5776 6672
rect 5632 6656 5684 6662
rect 5632 6598 5684 6604
rect 5540 6316 5592 6322
rect 5540 6258 5592 6264
rect 5264 5908 5316 5914
rect 5264 5850 5316 5856
rect 4804 5772 4856 5778
rect 4804 5714 4856 5720
rect 4656 5468 4964 5477
rect 4656 5466 4662 5468
rect 4718 5466 4742 5468
rect 4798 5466 4822 5468
rect 4878 5466 4902 5468
rect 4958 5466 4964 5468
rect 4718 5414 4720 5466
rect 4900 5414 4902 5466
rect 4656 5412 4662 5414
rect 4718 5412 4742 5414
rect 4798 5412 4822 5414
rect 4878 5412 4902 5414
rect 4958 5412 4964 5414
rect 4656 5403 4964 5412
rect 4528 4820 4580 4826
rect 4528 4762 4580 4768
rect 5172 4684 5224 4690
rect 5172 4626 5224 4632
rect 4528 4616 4580 4622
rect 4528 4558 4580 4564
rect 4344 4072 4396 4078
rect 4344 4014 4396 4020
rect 4540 3738 4568 4558
rect 4656 4380 4964 4389
rect 4656 4378 4662 4380
rect 4718 4378 4742 4380
rect 4798 4378 4822 4380
rect 4878 4378 4902 4380
rect 4958 4378 4964 4380
rect 4718 4326 4720 4378
rect 4900 4326 4902 4378
rect 4656 4324 4662 4326
rect 4718 4324 4742 4326
rect 4798 4324 4822 4326
rect 4878 4324 4902 4326
rect 4958 4324 4964 4326
rect 4656 4315 4964 4324
rect 5080 4072 5132 4078
rect 5080 4014 5132 4020
rect 4528 3732 4580 3738
rect 4528 3674 4580 3680
rect 4344 3528 4396 3534
rect 4264 3488 4344 3516
rect 3976 2576 4028 2582
rect 3976 2518 4028 2524
rect 3608 2508 3660 2514
rect 3608 2450 3660 2456
rect 3620 2106 3648 2450
rect 3988 2106 4016 2518
rect 3608 2100 3660 2106
rect 3608 2042 3660 2048
rect 3976 2100 4028 2106
rect 3976 2042 4028 2048
rect 3988 1902 4016 2042
rect 4264 2038 4292 3488
rect 4344 3470 4396 3476
rect 5092 3398 5120 4014
rect 5080 3392 5132 3398
rect 5080 3334 5132 3340
rect 4656 3292 4964 3301
rect 4656 3290 4662 3292
rect 4718 3290 4742 3292
rect 4798 3290 4822 3292
rect 4878 3290 4902 3292
rect 4958 3290 4964 3292
rect 4718 3238 4720 3290
rect 4900 3238 4902 3290
rect 4656 3236 4662 3238
rect 4718 3236 4742 3238
rect 4798 3236 4822 3238
rect 4878 3236 4902 3238
rect 4958 3236 4964 3238
rect 4656 3227 4964 3236
rect 5092 2650 5120 3334
rect 5184 3194 5212 4626
rect 5540 4548 5592 4554
rect 5540 4490 5592 4496
rect 5448 4140 5500 4146
rect 5448 4082 5500 4088
rect 5264 4072 5316 4078
rect 5264 4014 5316 4020
rect 5276 3534 5304 4014
rect 5356 4004 5408 4010
rect 5356 3946 5408 3952
rect 5368 3534 5396 3946
rect 5460 3738 5488 4082
rect 5552 4078 5580 4490
rect 5540 4072 5592 4078
rect 5540 4014 5592 4020
rect 5644 3738 5672 6598
rect 5828 5778 5856 6802
rect 5920 6186 5948 7142
rect 6206 7100 6514 7109
rect 6206 7098 6212 7100
rect 6268 7098 6292 7100
rect 6348 7098 6372 7100
rect 6428 7098 6452 7100
rect 6508 7098 6514 7100
rect 6268 7046 6270 7098
rect 6450 7046 6452 7098
rect 6206 7044 6212 7046
rect 6268 7044 6292 7046
rect 6348 7044 6372 7046
rect 6428 7044 6452 7046
rect 6508 7044 6514 7046
rect 6206 7035 6514 7044
rect 5908 6180 5960 6186
rect 5908 6122 5960 6128
rect 5920 5914 5948 6122
rect 6206 6012 6514 6021
rect 6206 6010 6212 6012
rect 6268 6010 6292 6012
rect 6348 6010 6372 6012
rect 6428 6010 6452 6012
rect 6508 6010 6514 6012
rect 6268 5958 6270 6010
rect 6450 5958 6452 6010
rect 6206 5956 6212 5958
rect 6268 5956 6292 5958
rect 6348 5956 6372 5958
rect 6428 5956 6452 5958
rect 6508 5956 6514 5958
rect 6206 5947 6514 5956
rect 5908 5908 5960 5914
rect 5908 5850 5960 5856
rect 5816 5772 5868 5778
rect 5816 5714 5868 5720
rect 5724 5704 5776 5710
rect 5724 5646 5776 5652
rect 5736 5166 5764 5646
rect 5920 5574 5948 5850
rect 5908 5568 5960 5574
rect 5908 5510 5960 5516
rect 5724 5160 5776 5166
rect 5724 5102 5776 5108
rect 5736 4622 5764 5102
rect 6206 4924 6514 4933
rect 6206 4922 6212 4924
rect 6268 4922 6292 4924
rect 6348 4922 6372 4924
rect 6428 4922 6452 4924
rect 6508 4922 6514 4924
rect 6268 4870 6270 4922
rect 6450 4870 6452 4922
rect 6206 4868 6212 4870
rect 6268 4868 6292 4870
rect 6348 4868 6372 4870
rect 6428 4868 6452 4870
rect 6508 4868 6514 4870
rect 6206 4859 6514 4868
rect 5724 4616 5776 4622
rect 5724 4558 5776 4564
rect 5724 4480 5776 4486
rect 5724 4422 5776 4428
rect 5736 4282 5764 4422
rect 5724 4276 5776 4282
rect 5724 4218 5776 4224
rect 6564 4214 6592 8298
rect 6840 7750 6868 9454
rect 6932 8634 6960 10610
rect 7024 9042 7052 11494
rect 7116 9586 7144 11630
rect 7392 10266 7420 11630
rect 7472 11620 7524 11626
rect 7472 11562 7524 11568
rect 7656 11620 7708 11626
rect 7656 11562 7708 11568
rect 7380 10260 7432 10266
rect 7380 10202 7432 10208
rect 7196 10124 7248 10130
rect 7196 10066 7248 10072
rect 7104 9580 7156 9586
rect 7104 9522 7156 9528
rect 7208 9518 7236 10066
rect 7380 9988 7432 9994
rect 7380 9930 7432 9936
rect 7196 9512 7248 9518
rect 7196 9454 7248 9460
rect 7012 9036 7064 9042
rect 7012 8978 7064 8984
rect 6920 8628 6972 8634
rect 6920 8570 6972 8576
rect 6932 7954 6960 8570
rect 7024 8430 7052 8978
rect 7208 8430 7236 9454
rect 7288 9376 7340 9382
rect 7288 9318 7340 9324
rect 7300 9178 7328 9318
rect 7288 9172 7340 9178
rect 7288 9114 7340 9120
rect 7012 8424 7064 8430
rect 7012 8366 7064 8372
rect 7196 8424 7248 8430
rect 7196 8366 7248 8372
rect 7300 8022 7328 9114
rect 7288 8016 7340 8022
rect 7288 7958 7340 7964
rect 6920 7948 6972 7954
rect 6920 7890 6972 7896
rect 6828 7744 6880 7750
rect 6828 7686 6880 7692
rect 6840 7342 6868 7686
rect 6828 7336 6880 7342
rect 6828 7278 6880 7284
rect 6736 6248 6788 6254
rect 6736 6190 6788 6196
rect 6748 5370 6776 6190
rect 6736 5364 6788 5370
rect 6736 5306 6788 5312
rect 6552 4208 6604 4214
rect 6552 4150 6604 4156
rect 6206 3836 6514 3845
rect 6206 3834 6212 3836
rect 6268 3834 6292 3836
rect 6348 3834 6372 3836
rect 6428 3834 6452 3836
rect 6508 3834 6514 3836
rect 6268 3782 6270 3834
rect 6450 3782 6452 3834
rect 6206 3780 6212 3782
rect 6268 3780 6292 3782
rect 6348 3780 6372 3782
rect 6428 3780 6452 3782
rect 6508 3780 6514 3782
rect 6206 3771 6514 3780
rect 5448 3732 5500 3738
rect 5448 3674 5500 3680
rect 5632 3732 5684 3738
rect 5632 3674 5684 3680
rect 5264 3528 5316 3534
rect 5264 3470 5316 3476
rect 5356 3528 5408 3534
rect 5356 3470 5408 3476
rect 5460 3466 5488 3674
rect 5540 3596 5592 3602
rect 5540 3538 5592 3544
rect 5448 3460 5500 3466
rect 5448 3402 5500 3408
rect 5264 3392 5316 3398
rect 5264 3334 5316 3340
rect 5276 3194 5304 3334
rect 5172 3188 5224 3194
rect 5172 3130 5224 3136
rect 5264 3188 5316 3194
rect 5264 3130 5316 3136
rect 5264 2984 5316 2990
rect 5264 2926 5316 2932
rect 5276 2650 5304 2926
rect 5080 2644 5132 2650
rect 5080 2586 5132 2592
rect 5264 2644 5316 2650
rect 5264 2586 5316 2592
rect 4656 2204 4964 2213
rect 4656 2202 4662 2204
rect 4718 2202 4742 2204
rect 4798 2202 4822 2204
rect 4878 2202 4902 2204
rect 4958 2202 4964 2204
rect 4718 2150 4720 2202
rect 4900 2150 4902 2202
rect 4656 2148 4662 2150
rect 4718 2148 4742 2150
rect 4798 2148 4822 2150
rect 4878 2148 4902 2150
rect 4958 2148 4964 2150
rect 4656 2139 4964 2148
rect 4252 2032 4304 2038
rect 4252 1974 4304 1980
rect 5264 2032 5316 2038
rect 5264 1974 5316 1980
rect 4264 1902 4292 1974
rect 5276 1902 5304 1974
rect 5552 1970 5580 3538
rect 6736 3392 6788 3398
rect 6736 3334 6788 3340
rect 6748 2990 6776 3334
rect 6932 3194 6960 7890
rect 7300 6186 7328 7958
rect 7392 7886 7420 9930
rect 7380 7880 7432 7886
rect 7380 7822 7432 7828
rect 7484 7818 7512 11562
rect 7668 10810 7696 11562
rect 8036 11286 8064 11630
rect 8024 11280 8076 11286
rect 8024 11222 8076 11228
rect 7756 10908 8064 10917
rect 7756 10906 7762 10908
rect 7818 10906 7842 10908
rect 7898 10906 7922 10908
rect 7978 10906 8002 10908
rect 8058 10906 8064 10908
rect 7818 10854 7820 10906
rect 8000 10854 8002 10906
rect 7756 10852 7762 10854
rect 7818 10852 7842 10854
rect 7898 10852 7922 10854
rect 7978 10852 8002 10854
rect 8058 10852 8064 10854
rect 7756 10843 8064 10852
rect 7656 10804 7708 10810
rect 7656 10746 7708 10752
rect 8128 10606 8156 12582
rect 8220 11694 8248 14010
rect 8312 13870 8340 15574
rect 8760 15088 8812 15094
rect 8760 15030 8812 15036
rect 8300 13864 8352 13870
rect 8300 13806 8352 13812
rect 8392 13796 8444 13802
rect 8392 13738 8444 13744
rect 8404 13530 8432 13738
rect 8392 13524 8444 13530
rect 8392 13466 8444 13472
rect 8208 11688 8260 11694
rect 8208 11630 8260 11636
rect 8300 11688 8352 11694
rect 8300 11630 8352 11636
rect 8312 11354 8340 11630
rect 8300 11348 8352 11354
rect 8300 11290 8352 11296
rect 8116 10600 8168 10606
rect 8116 10542 8168 10548
rect 8576 10532 8628 10538
rect 8576 10474 8628 10480
rect 8116 10464 8168 10470
rect 8116 10406 8168 10412
rect 8128 10198 8156 10406
rect 8116 10192 8168 10198
rect 8116 10134 8168 10140
rect 7564 10056 7616 10062
rect 7564 9998 7616 10004
rect 7576 8974 7604 9998
rect 7756 9820 8064 9829
rect 7756 9818 7762 9820
rect 7818 9818 7842 9820
rect 7898 9818 7922 9820
rect 7978 9818 8002 9820
rect 8058 9818 8064 9820
rect 7818 9766 7820 9818
rect 8000 9766 8002 9818
rect 7756 9764 7762 9766
rect 7818 9764 7842 9766
rect 7898 9764 7922 9766
rect 7978 9764 8002 9766
rect 8058 9764 8064 9766
rect 7756 9755 8064 9764
rect 8208 9648 8260 9654
rect 8208 9590 8260 9596
rect 7564 8968 7616 8974
rect 7564 8910 7616 8916
rect 8116 8968 8168 8974
rect 8116 8910 8168 8916
rect 7756 8732 8064 8741
rect 7756 8730 7762 8732
rect 7818 8730 7842 8732
rect 7898 8730 7922 8732
rect 7978 8730 8002 8732
rect 8058 8730 8064 8732
rect 7818 8678 7820 8730
rect 8000 8678 8002 8730
rect 7756 8676 7762 8678
rect 7818 8676 7842 8678
rect 7898 8676 7922 8678
rect 7978 8676 8002 8678
rect 8058 8676 8064 8678
rect 7756 8667 8064 8676
rect 8128 8634 8156 8910
rect 8116 8628 8168 8634
rect 8116 8570 8168 8576
rect 8220 8498 8248 9590
rect 8588 9450 8616 10474
rect 8668 10192 8720 10198
rect 8668 10134 8720 10140
rect 8576 9444 8628 9450
rect 8576 9386 8628 9392
rect 8588 8634 8616 9386
rect 8680 9382 8708 10134
rect 8668 9376 8720 9382
rect 8668 9318 8720 9324
rect 8680 9110 8708 9318
rect 8668 9104 8720 9110
rect 8668 9046 8720 9052
rect 8576 8628 8628 8634
rect 8628 8588 8708 8616
rect 8576 8570 8628 8576
rect 8208 8492 8260 8498
rect 8208 8434 8260 8440
rect 8392 8424 8444 8430
rect 8392 8366 8444 8372
rect 8404 7954 8432 8366
rect 8392 7948 8444 7954
rect 8392 7890 8444 7896
rect 8116 7880 8168 7886
rect 8116 7822 8168 7828
rect 7472 7812 7524 7818
rect 7472 7754 7524 7760
rect 7656 7812 7708 7818
rect 7656 7754 7708 7760
rect 7288 6180 7340 6186
rect 7288 6122 7340 6128
rect 7300 5914 7328 6122
rect 7288 5908 7340 5914
rect 7288 5850 7340 5856
rect 7472 5364 7524 5370
rect 7472 5306 7524 5312
rect 7484 5166 7512 5306
rect 7564 5296 7616 5302
rect 7564 5238 7616 5244
rect 7196 5160 7248 5166
rect 7196 5102 7248 5108
rect 7472 5160 7524 5166
rect 7472 5102 7524 5108
rect 7104 5092 7156 5098
rect 7104 5034 7156 5040
rect 7116 3194 7144 5034
rect 7208 4826 7236 5102
rect 7196 4820 7248 4826
rect 7196 4762 7248 4768
rect 7484 4078 7512 5102
rect 7576 4690 7604 5238
rect 7668 5166 7696 7754
rect 7756 7644 8064 7653
rect 7756 7642 7762 7644
rect 7818 7642 7842 7644
rect 7898 7642 7922 7644
rect 7978 7642 8002 7644
rect 8058 7642 8064 7644
rect 7818 7590 7820 7642
rect 8000 7590 8002 7642
rect 7756 7588 7762 7590
rect 7818 7588 7842 7590
rect 7898 7588 7922 7590
rect 7978 7588 8002 7590
rect 8058 7588 8064 7590
rect 7756 7579 8064 7588
rect 8128 7546 8156 7822
rect 8116 7540 8168 7546
rect 8116 7482 8168 7488
rect 8404 7410 8432 7890
rect 8392 7404 8444 7410
rect 8392 7346 8444 7352
rect 8300 7336 8352 7342
rect 8300 7278 8352 7284
rect 7756 6556 8064 6565
rect 7756 6554 7762 6556
rect 7818 6554 7842 6556
rect 7898 6554 7922 6556
rect 7978 6554 8002 6556
rect 8058 6554 8064 6556
rect 7818 6502 7820 6554
rect 8000 6502 8002 6554
rect 7756 6500 7762 6502
rect 7818 6500 7842 6502
rect 7898 6500 7922 6502
rect 7978 6500 8002 6502
rect 8058 6500 8064 6502
rect 7756 6491 8064 6500
rect 8116 6180 8168 6186
rect 8116 6122 8168 6128
rect 8128 5778 8156 6122
rect 8116 5772 8168 5778
rect 8116 5714 8168 5720
rect 7756 5468 8064 5477
rect 7756 5466 7762 5468
rect 7818 5466 7842 5468
rect 7898 5466 7922 5468
rect 7978 5466 8002 5468
rect 8058 5466 8064 5468
rect 7818 5414 7820 5466
rect 8000 5414 8002 5466
rect 7756 5412 7762 5414
rect 7818 5412 7842 5414
rect 7898 5412 7922 5414
rect 7978 5412 8002 5414
rect 8058 5412 8064 5414
rect 7756 5403 8064 5412
rect 7656 5160 7708 5166
rect 7656 5102 7708 5108
rect 7840 5160 7892 5166
rect 7840 5102 7892 5108
rect 7748 5092 7800 5098
rect 7748 5034 7800 5040
rect 7760 4978 7788 5034
rect 7668 4950 7788 4978
rect 7564 4684 7616 4690
rect 7564 4626 7616 4632
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 7472 4072 7524 4078
rect 7472 4014 7524 4020
rect 6920 3188 6972 3194
rect 6920 3130 6972 3136
rect 7104 3188 7156 3194
rect 7104 3130 7156 3136
rect 6828 3052 6880 3058
rect 6828 2994 6880 3000
rect 6736 2984 6788 2990
rect 6736 2926 6788 2932
rect 6206 2748 6514 2757
rect 6206 2746 6212 2748
rect 6268 2746 6292 2748
rect 6348 2746 6372 2748
rect 6428 2746 6452 2748
rect 6508 2746 6514 2748
rect 6268 2694 6270 2746
rect 6450 2694 6452 2746
rect 6206 2692 6212 2694
rect 6268 2692 6292 2694
rect 6348 2692 6372 2694
rect 6428 2692 6452 2694
rect 6508 2692 6514 2694
rect 6206 2683 6514 2692
rect 6368 2508 6420 2514
rect 6368 2450 6420 2456
rect 5816 2440 5868 2446
rect 5816 2382 5868 2388
rect 5540 1964 5592 1970
rect 5540 1906 5592 1912
rect 5828 1902 5856 2382
rect 6380 2106 6408 2450
rect 6368 2100 6420 2106
rect 6368 2042 6420 2048
rect 6748 1902 6776 2926
rect 6840 2446 6868 2994
rect 6932 2922 6960 3130
rect 7484 3058 7512 4014
rect 7576 3738 7604 4082
rect 7564 3732 7616 3738
rect 7564 3674 7616 3680
rect 7472 3052 7524 3058
rect 7472 2994 7524 3000
rect 6920 2916 6972 2922
rect 6920 2858 6972 2864
rect 7472 2916 7524 2922
rect 7472 2858 7524 2864
rect 7380 2848 7432 2854
rect 7380 2790 7432 2796
rect 6828 2440 6880 2446
rect 6828 2382 6880 2388
rect 7392 2106 7420 2790
rect 7380 2100 7432 2106
rect 7380 2042 7432 2048
rect 7484 1970 7512 2858
rect 7472 1964 7524 1970
rect 7472 1906 7524 1912
rect 3332 1896 3384 1902
rect 3332 1838 3384 1844
rect 3516 1896 3568 1902
rect 3976 1896 4028 1902
rect 3568 1844 3648 1850
rect 3516 1838 3648 1844
rect 3976 1838 4028 1844
rect 4252 1896 4304 1902
rect 4252 1838 4304 1844
rect 5172 1896 5224 1902
rect 5172 1838 5224 1844
rect 5264 1896 5316 1902
rect 5264 1838 5316 1844
rect 5816 1896 5868 1902
rect 5816 1838 5868 1844
rect 6736 1896 6788 1902
rect 6736 1838 6788 1844
rect 3528 1822 3648 1838
rect 3516 1760 3568 1766
rect 3516 1702 3568 1708
rect 3106 1660 3414 1669
rect 3106 1658 3112 1660
rect 3168 1658 3192 1660
rect 3248 1658 3272 1660
rect 3328 1658 3352 1660
rect 3408 1658 3414 1660
rect 3168 1606 3170 1658
rect 3350 1606 3352 1658
rect 3106 1604 3112 1606
rect 3168 1604 3192 1606
rect 3248 1604 3272 1606
rect 3328 1604 3352 1606
rect 3408 1604 3414 1606
rect 3106 1595 3414 1604
rect 3528 1562 3556 1702
rect 3516 1556 3568 1562
rect 3516 1498 3568 1504
rect 3620 1426 3648 1822
rect 3608 1420 3660 1426
rect 3608 1362 3660 1368
rect 3988 1358 4016 1838
rect 3976 1352 4028 1358
rect 3976 1294 4028 1300
rect 1556 1116 1864 1125
rect 1556 1114 1562 1116
rect 1618 1114 1642 1116
rect 1698 1114 1722 1116
rect 1778 1114 1802 1116
rect 1858 1114 1864 1116
rect 1618 1062 1620 1114
rect 1800 1062 1802 1114
rect 1556 1060 1562 1062
rect 1618 1060 1642 1062
rect 1698 1060 1722 1062
rect 1778 1060 1802 1062
rect 1858 1060 1864 1062
rect 1556 1051 1864 1060
rect 3988 1018 4016 1294
rect 4656 1116 4964 1125
rect 4656 1114 4662 1116
rect 4718 1114 4742 1116
rect 4798 1114 4822 1116
rect 4878 1114 4902 1116
rect 4958 1114 4964 1116
rect 4718 1062 4720 1114
rect 4900 1062 4902 1114
rect 4656 1060 4662 1062
rect 4718 1060 4742 1062
rect 4798 1060 4822 1062
rect 4878 1060 4902 1062
rect 4958 1060 4964 1062
rect 4656 1051 4964 1060
rect 3976 1012 4028 1018
rect 3976 954 4028 960
rect 5184 814 5212 1838
rect 5276 950 5304 1838
rect 5540 1760 5592 1766
rect 5540 1702 5592 1708
rect 6736 1760 6788 1766
rect 6736 1702 6788 1708
rect 5552 1426 5580 1702
rect 6206 1660 6514 1669
rect 6206 1658 6212 1660
rect 6268 1658 6292 1660
rect 6348 1658 6372 1660
rect 6428 1658 6452 1660
rect 6508 1658 6514 1660
rect 6268 1606 6270 1658
rect 6450 1606 6452 1658
rect 6206 1604 6212 1606
rect 6268 1604 6292 1606
rect 6348 1604 6372 1606
rect 6428 1604 6452 1606
rect 6508 1604 6514 1606
rect 6206 1595 6514 1604
rect 6748 1562 6776 1702
rect 6736 1556 6788 1562
rect 6736 1498 6788 1504
rect 7668 1426 7696 4950
rect 7852 4690 7880 5102
rect 8128 5098 8156 5714
rect 8312 5642 8340 7278
rect 8300 5636 8352 5642
rect 8300 5578 8352 5584
rect 8116 5092 8168 5098
rect 8116 5034 8168 5040
rect 7840 4684 7892 4690
rect 7840 4626 7892 4632
rect 8116 4616 8168 4622
rect 8116 4558 8168 4564
rect 7756 4380 8064 4389
rect 7756 4378 7762 4380
rect 7818 4378 7842 4380
rect 7898 4378 7922 4380
rect 7978 4378 8002 4380
rect 8058 4378 8064 4380
rect 7818 4326 7820 4378
rect 8000 4326 8002 4378
rect 7756 4324 7762 4326
rect 7818 4324 7842 4326
rect 7898 4324 7922 4326
rect 7978 4324 8002 4326
rect 8058 4324 8064 4326
rect 7756 4315 8064 4324
rect 8128 3534 8156 4558
rect 8208 3596 8260 3602
rect 8208 3538 8260 3544
rect 8116 3528 8168 3534
rect 8116 3470 8168 3476
rect 7756 3292 8064 3301
rect 7756 3290 7762 3292
rect 7818 3290 7842 3292
rect 7898 3290 7922 3292
rect 7978 3290 8002 3292
rect 8058 3290 8064 3292
rect 7818 3238 7820 3290
rect 8000 3238 8002 3290
rect 7756 3236 7762 3238
rect 7818 3236 7842 3238
rect 7898 3236 7922 3238
rect 7978 3236 8002 3238
rect 8058 3236 8064 3238
rect 7756 3227 8064 3236
rect 8220 2650 8248 3538
rect 8404 3466 8432 7346
rect 8484 5772 8536 5778
rect 8484 5714 8536 5720
rect 8496 4690 8524 5714
rect 8680 5370 8708 8588
rect 8772 7954 8800 15030
rect 9048 14822 9076 15914
rect 9306 15804 9614 15813
rect 9306 15802 9312 15804
rect 9368 15802 9392 15804
rect 9448 15802 9472 15804
rect 9528 15802 9552 15804
rect 9608 15802 9614 15804
rect 9368 15750 9370 15802
rect 9550 15750 9552 15802
rect 9306 15748 9312 15750
rect 9368 15748 9392 15750
rect 9448 15748 9472 15750
rect 9528 15748 9552 15750
rect 9608 15748 9614 15750
rect 9306 15739 9614 15748
rect 9496 15360 9548 15366
rect 9496 15302 9548 15308
rect 9508 15094 9536 15302
rect 9876 15162 9904 16594
rect 10060 16522 10088 18142
rect 10324 18080 10376 18086
rect 10324 18022 10376 18028
rect 11244 18080 11296 18086
rect 11244 18022 11296 18028
rect 10048 16516 10100 16522
rect 10048 16458 10100 16464
rect 10336 16250 10364 18022
rect 10856 17436 11164 17445
rect 10856 17434 10862 17436
rect 10918 17434 10942 17436
rect 10998 17434 11022 17436
rect 11078 17434 11102 17436
rect 11158 17434 11164 17436
rect 10918 17382 10920 17434
rect 11100 17382 11102 17434
rect 10856 17380 10862 17382
rect 10918 17380 10942 17382
rect 10998 17380 11022 17382
rect 11078 17380 11102 17382
rect 11158 17380 11164 17382
rect 10856 17371 11164 17380
rect 11256 17202 11284 18022
rect 11244 17196 11296 17202
rect 11244 17138 11296 17144
rect 11348 16794 11376 18158
rect 12406 17980 12714 17989
rect 12406 17978 12412 17980
rect 12468 17978 12492 17980
rect 12548 17978 12572 17980
rect 12628 17978 12652 17980
rect 12708 17978 12714 17980
rect 12468 17926 12470 17978
rect 12650 17926 12652 17978
rect 12406 17924 12412 17926
rect 12468 17924 12492 17926
rect 12548 17924 12572 17926
rect 12628 17924 12652 17926
rect 12708 17924 12714 17926
rect 12406 17915 12714 17924
rect 12440 17740 12492 17746
rect 12440 17682 12492 17688
rect 11520 17604 11572 17610
rect 11520 17546 11572 17552
rect 11980 17604 12032 17610
rect 11980 17546 12032 17552
rect 11428 17536 11480 17542
rect 11428 17478 11480 17484
rect 11336 16788 11388 16794
rect 11336 16730 11388 16736
rect 11336 16584 11388 16590
rect 11336 16526 11388 16532
rect 10856 16348 11164 16357
rect 10856 16346 10862 16348
rect 10918 16346 10942 16348
rect 10998 16346 11022 16348
rect 11078 16346 11102 16348
rect 11158 16346 11164 16348
rect 10918 16294 10920 16346
rect 11100 16294 11102 16346
rect 10856 16292 10862 16294
rect 10918 16292 10942 16294
rect 10998 16292 11022 16294
rect 11078 16292 11102 16294
rect 11158 16292 11164 16294
rect 10856 16283 11164 16292
rect 10324 16244 10376 16250
rect 10324 16186 10376 16192
rect 11348 16046 11376 16526
rect 11336 16040 11388 16046
rect 11336 15982 11388 15988
rect 11152 15972 11204 15978
rect 11152 15914 11204 15920
rect 11164 15706 11192 15914
rect 11152 15700 11204 15706
rect 11152 15642 11204 15648
rect 10232 15496 10284 15502
rect 10232 15438 10284 15444
rect 9864 15156 9916 15162
rect 9864 15098 9916 15104
rect 9496 15088 9548 15094
rect 9496 15030 9548 15036
rect 9036 14816 9088 14822
rect 9036 14758 9088 14764
rect 8944 13320 8996 13326
rect 8944 13262 8996 13268
rect 8956 12918 8984 13262
rect 8944 12912 8996 12918
rect 8944 12854 8996 12860
rect 8852 12096 8904 12102
rect 8852 12038 8904 12044
rect 8864 11694 8892 12038
rect 8852 11688 8904 11694
rect 8852 11630 8904 11636
rect 9048 11286 9076 14758
rect 9306 14716 9614 14725
rect 9306 14714 9312 14716
rect 9368 14714 9392 14716
rect 9448 14714 9472 14716
rect 9528 14714 9552 14716
rect 9608 14714 9614 14716
rect 9368 14662 9370 14714
rect 9550 14662 9552 14714
rect 9306 14660 9312 14662
rect 9368 14660 9392 14662
rect 9448 14660 9472 14662
rect 9528 14660 9552 14662
rect 9608 14660 9614 14662
rect 9306 14651 9614 14660
rect 9128 14272 9180 14278
rect 9128 14214 9180 14220
rect 10048 14272 10100 14278
rect 10048 14214 10100 14220
rect 9140 13938 9168 14214
rect 10060 13938 10088 14214
rect 9128 13932 9180 13938
rect 9128 13874 9180 13880
rect 10048 13932 10100 13938
rect 10048 13874 10100 13880
rect 9140 13274 9168 13874
rect 9680 13728 9732 13734
rect 9680 13670 9732 13676
rect 9306 13628 9614 13637
rect 9306 13626 9312 13628
rect 9368 13626 9392 13628
rect 9448 13626 9472 13628
rect 9528 13626 9552 13628
rect 9608 13626 9614 13628
rect 9368 13574 9370 13626
rect 9550 13574 9552 13626
rect 9306 13572 9312 13574
rect 9368 13572 9392 13574
rect 9448 13572 9472 13574
rect 9528 13572 9552 13574
rect 9608 13572 9614 13574
rect 9306 13563 9614 13572
rect 9312 13320 9364 13326
rect 9140 13268 9312 13274
rect 9140 13262 9364 13268
rect 9140 13246 9352 13262
rect 9128 12300 9180 12306
rect 9128 12242 9180 12248
rect 9232 12288 9260 13246
rect 9306 12540 9614 12549
rect 9306 12538 9312 12540
rect 9368 12538 9392 12540
rect 9448 12538 9472 12540
rect 9528 12538 9552 12540
rect 9608 12538 9614 12540
rect 9368 12486 9370 12538
rect 9550 12486 9552 12538
rect 9306 12484 9312 12486
rect 9368 12484 9392 12486
rect 9448 12484 9472 12486
rect 9528 12484 9552 12486
rect 9608 12484 9614 12486
rect 9306 12475 9614 12484
rect 9496 12436 9548 12442
rect 9496 12378 9548 12384
rect 9312 12300 9364 12306
rect 9232 12260 9312 12288
rect 9036 11280 9088 11286
rect 9036 11222 9088 11228
rect 9140 10010 9168 12242
rect 9232 11558 9260 12260
rect 9312 12242 9364 12248
rect 9508 11626 9536 12378
rect 9692 12238 9720 13670
rect 10244 13394 10272 15438
rect 10856 15260 11164 15269
rect 10856 15258 10862 15260
rect 10918 15258 10942 15260
rect 10998 15258 11022 15260
rect 11078 15258 11102 15260
rect 11158 15258 11164 15260
rect 10918 15206 10920 15258
rect 11100 15206 11102 15258
rect 10856 15204 10862 15206
rect 10918 15204 10942 15206
rect 10998 15204 11022 15206
rect 11078 15204 11102 15206
rect 11158 15204 11164 15206
rect 10856 15195 11164 15204
rect 11348 14958 11376 15982
rect 11440 15978 11468 17478
rect 11532 16522 11560 17546
rect 11888 17536 11940 17542
rect 11888 17478 11940 17484
rect 11612 16992 11664 16998
rect 11612 16934 11664 16940
rect 11704 16992 11756 16998
rect 11704 16934 11756 16940
rect 11624 16794 11652 16934
rect 11612 16788 11664 16794
rect 11612 16730 11664 16736
rect 11520 16516 11572 16522
rect 11520 16458 11572 16464
rect 11428 15972 11480 15978
rect 11428 15914 11480 15920
rect 11532 15638 11560 16458
rect 11520 15632 11572 15638
rect 11572 15580 11652 15586
rect 11520 15574 11652 15580
rect 11532 15558 11652 15574
rect 11520 15496 11572 15502
rect 11520 15438 11572 15444
rect 11336 14952 11388 14958
rect 11336 14894 11388 14900
rect 11336 14816 11388 14822
rect 11336 14758 11388 14764
rect 11348 14482 11376 14758
rect 11532 14618 11560 15438
rect 11520 14612 11572 14618
rect 11520 14554 11572 14560
rect 11336 14476 11388 14482
rect 11336 14418 11388 14424
rect 11336 14272 11388 14278
rect 11336 14214 11388 14220
rect 10856 14172 11164 14181
rect 10856 14170 10862 14172
rect 10918 14170 10942 14172
rect 10998 14170 11022 14172
rect 11078 14170 11102 14172
rect 11158 14170 11164 14172
rect 10918 14118 10920 14170
rect 11100 14118 11102 14170
rect 10856 14116 10862 14118
rect 10918 14116 10942 14118
rect 10998 14116 11022 14118
rect 11078 14116 11102 14118
rect 11158 14116 11164 14118
rect 10856 14107 11164 14116
rect 11244 13728 11296 13734
rect 11244 13670 11296 13676
rect 9956 13388 10008 13394
rect 9956 13330 10008 13336
rect 10232 13388 10284 13394
rect 10232 13330 10284 13336
rect 9680 12232 9732 12238
rect 9680 12174 9732 12180
rect 9496 11620 9548 11626
rect 9496 11562 9548 11568
rect 9220 11552 9272 11558
rect 9220 11494 9272 11500
rect 9306 11452 9614 11461
rect 9306 11450 9312 11452
rect 9368 11450 9392 11452
rect 9448 11450 9472 11452
rect 9528 11450 9552 11452
rect 9608 11450 9614 11452
rect 9368 11398 9370 11450
rect 9550 11398 9552 11450
rect 9306 11396 9312 11398
rect 9368 11396 9392 11398
rect 9448 11396 9472 11398
rect 9528 11396 9552 11398
rect 9608 11396 9614 11398
rect 9306 11387 9614 11396
rect 9306 10364 9614 10373
rect 9306 10362 9312 10364
rect 9368 10362 9392 10364
rect 9448 10362 9472 10364
rect 9528 10362 9552 10364
rect 9608 10362 9614 10364
rect 9368 10310 9370 10362
rect 9550 10310 9552 10362
rect 9306 10308 9312 10310
rect 9368 10308 9392 10310
rect 9448 10308 9472 10310
rect 9528 10308 9552 10310
rect 9608 10308 9614 10310
rect 9306 10299 9614 10308
rect 9048 9982 9168 10010
rect 8944 9376 8996 9382
rect 8944 9318 8996 9324
rect 8956 8566 8984 9318
rect 8944 8560 8996 8566
rect 8944 8502 8996 8508
rect 8760 7948 8812 7954
rect 8760 7890 8812 7896
rect 8956 7478 8984 8502
rect 8944 7472 8996 7478
rect 8944 7414 8996 7420
rect 9048 6458 9076 9982
rect 9128 9920 9180 9926
rect 9128 9862 9180 9868
rect 9140 8430 9168 9862
rect 9220 9512 9272 9518
rect 9220 9454 9272 9460
rect 9232 9178 9260 9454
rect 9306 9276 9614 9285
rect 9306 9274 9312 9276
rect 9368 9274 9392 9276
rect 9448 9274 9472 9276
rect 9528 9274 9552 9276
rect 9608 9274 9614 9276
rect 9368 9222 9370 9274
rect 9550 9222 9552 9274
rect 9306 9220 9312 9222
rect 9368 9220 9392 9222
rect 9448 9220 9472 9222
rect 9528 9220 9552 9222
rect 9608 9220 9614 9222
rect 9306 9211 9614 9220
rect 9220 9172 9272 9178
rect 9220 9114 9272 9120
rect 9128 8424 9180 8430
rect 9128 8366 9180 8372
rect 9692 8294 9720 12174
rect 9772 11552 9824 11558
rect 9772 11494 9824 11500
rect 9784 11218 9812 11494
rect 9968 11218 9996 13330
rect 10244 13190 10272 13330
rect 10508 13320 10560 13326
rect 10508 13262 10560 13268
rect 10232 13184 10284 13190
rect 10232 13126 10284 13132
rect 10520 12714 10548 13262
rect 10856 13084 11164 13093
rect 10856 13082 10862 13084
rect 10918 13082 10942 13084
rect 10998 13082 11022 13084
rect 11078 13082 11102 13084
rect 11158 13082 11164 13084
rect 10918 13030 10920 13082
rect 11100 13030 11102 13082
rect 10856 13028 10862 13030
rect 10918 13028 10942 13030
rect 10998 13028 11022 13030
rect 11078 13028 11102 13030
rect 11158 13028 11164 13030
rect 10856 13019 11164 13028
rect 11152 12776 11204 12782
rect 11256 12764 11284 13670
rect 11348 12986 11376 14214
rect 11624 13394 11652 15558
rect 11716 14618 11744 16934
rect 11704 14612 11756 14618
rect 11704 14554 11756 14560
rect 11900 14482 11928 17478
rect 11992 15706 12020 17546
rect 12452 17134 12480 17682
rect 12820 17678 12848 19200
rect 13956 18524 14264 18533
rect 13956 18522 13962 18524
rect 14018 18522 14042 18524
rect 14098 18522 14122 18524
rect 14178 18522 14202 18524
rect 14258 18522 14264 18524
rect 14018 18470 14020 18522
rect 14200 18470 14202 18522
rect 13956 18468 13962 18470
rect 14018 18468 14042 18470
rect 14098 18468 14122 18470
rect 14178 18468 14202 18470
rect 14258 18468 14264 18470
rect 13956 18459 14264 18468
rect 12992 18284 13044 18290
rect 12992 18226 13044 18232
rect 12900 18216 12952 18222
rect 12900 18158 12952 18164
rect 12912 17746 12940 18158
rect 12900 17740 12952 17746
rect 12900 17682 12952 17688
rect 12808 17672 12860 17678
rect 12808 17614 12860 17620
rect 12716 17536 12768 17542
rect 12716 17478 12768 17484
rect 12728 17134 12756 17478
rect 13004 17338 13032 18226
rect 14372 18216 14424 18222
rect 14372 18158 14424 18164
rect 14924 18216 14976 18222
rect 14924 18158 14976 18164
rect 13820 18148 13872 18154
rect 13820 18090 13872 18096
rect 13268 18080 13320 18086
rect 13268 18022 13320 18028
rect 13084 17604 13136 17610
rect 13084 17546 13136 17552
rect 12992 17332 13044 17338
rect 12992 17274 13044 17280
rect 12808 17264 12860 17270
rect 12808 17206 12860 17212
rect 12900 17264 12952 17270
rect 12900 17206 12952 17212
rect 12440 17128 12492 17134
rect 12440 17070 12492 17076
rect 12716 17128 12768 17134
rect 12716 17070 12768 17076
rect 12406 16892 12714 16901
rect 12406 16890 12412 16892
rect 12468 16890 12492 16892
rect 12548 16890 12572 16892
rect 12628 16890 12652 16892
rect 12708 16890 12714 16892
rect 12468 16838 12470 16890
rect 12650 16838 12652 16890
rect 12406 16836 12412 16838
rect 12468 16836 12492 16838
rect 12548 16836 12572 16838
rect 12628 16836 12652 16838
rect 12708 16836 12714 16838
rect 12406 16827 12714 16836
rect 12716 16788 12768 16794
rect 12716 16730 12768 16736
rect 12728 16454 12756 16730
rect 12716 16448 12768 16454
rect 12716 16390 12768 16396
rect 12406 15804 12714 15813
rect 12406 15802 12412 15804
rect 12468 15802 12492 15804
rect 12548 15802 12572 15804
rect 12628 15802 12652 15804
rect 12708 15802 12714 15804
rect 12468 15750 12470 15802
rect 12650 15750 12652 15802
rect 12406 15748 12412 15750
rect 12468 15748 12492 15750
rect 12548 15748 12572 15750
rect 12628 15748 12652 15750
rect 12708 15748 12714 15750
rect 12406 15739 12714 15748
rect 12820 15706 12848 17206
rect 12912 17066 12940 17206
rect 13096 17134 13124 17546
rect 13176 17332 13228 17338
rect 13176 17274 13228 17280
rect 13084 17128 13136 17134
rect 13084 17070 13136 17076
rect 12900 17060 12952 17066
rect 12900 17002 12952 17008
rect 13188 16522 13216 17274
rect 13176 16516 13228 16522
rect 13176 16458 13228 16464
rect 13280 16454 13308 18022
rect 13636 17876 13688 17882
rect 13636 17818 13688 17824
rect 13452 17264 13504 17270
rect 13452 17206 13504 17212
rect 13360 17128 13412 17134
rect 13360 17070 13412 17076
rect 13372 16697 13400 17070
rect 13358 16688 13414 16697
rect 13358 16623 13414 16632
rect 13464 16522 13492 17206
rect 13648 16658 13676 17818
rect 13832 17202 13860 18090
rect 13956 17436 14264 17445
rect 13956 17434 13962 17436
rect 14018 17434 14042 17436
rect 14098 17434 14122 17436
rect 14178 17434 14202 17436
rect 14258 17434 14264 17436
rect 14018 17382 14020 17434
rect 14200 17382 14202 17434
rect 13956 17380 13962 17382
rect 14018 17380 14042 17382
rect 14098 17380 14122 17382
rect 14178 17380 14202 17382
rect 14258 17380 14264 17382
rect 13956 17371 14264 17380
rect 13820 17196 13872 17202
rect 13820 17138 13872 17144
rect 13728 16992 13780 16998
rect 13728 16934 13780 16940
rect 13636 16652 13688 16658
rect 13636 16594 13688 16600
rect 13452 16516 13504 16522
rect 13452 16458 13504 16464
rect 13268 16448 13320 16454
rect 13268 16390 13320 16396
rect 11980 15700 12032 15706
rect 11980 15642 12032 15648
rect 12808 15700 12860 15706
rect 12808 15642 12860 15648
rect 11992 15094 12020 15642
rect 13280 15570 13308 16390
rect 13452 15632 13504 15638
rect 13452 15574 13504 15580
rect 12808 15564 12860 15570
rect 12808 15506 12860 15512
rect 13268 15564 13320 15570
rect 13268 15506 13320 15512
rect 12348 15360 12400 15366
rect 12348 15302 12400 15308
rect 11980 15088 12032 15094
rect 11980 15030 12032 15036
rect 12360 14958 12388 15302
rect 12348 14952 12400 14958
rect 12348 14894 12400 14900
rect 12256 14816 12308 14822
rect 12256 14758 12308 14764
rect 11888 14476 11940 14482
rect 11888 14418 11940 14424
rect 12268 14414 12296 14758
rect 12406 14716 12714 14725
rect 12406 14714 12412 14716
rect 12468 14714 12492 14716
rect 12548 14714 12572 14716
rect 12628 14714 12652 14716
rect 12708 14714 12714 14716
rect 12468 14662 12470 14714
rect 12650 14662 12652 14714
rect 12406 14660 12412 14662
rect 12468 14660 12492 14662
rect 12548 14660 12572 14662
rect 12628 14660 12652 14662
rect 12708 14660 12714 14662
rect 12406 14651 12714 14660
rect 12820 14618 12848 15506
rect 12900 15496 12952 15502
rect 12900 15438 12952 15444
rect 12912 14958 12940 15438
rect 12992 15156 13044 15162
rect 12992 15098 13044 15104
rect 13004 14958 13032 15098
rect 12900 14952 12952 14958
rect 12900 14894 12952 14900
rect 12992 14952 13044 14958
rect 12992 14894 13044 14900
rect 12808 14612 12860 14618
rect 12808 14554 12860 14560
rect 12912 14482 12940 14894
rect 12992 14816 13044 14822
rect 12992 14758 13044 14764
rect 13004 14482 13032 14758
rect 12900 14476 12952 14482
rect 12900 14418 12952 14424
rect 12992 14476 13044 14482
rect 12992 14418 13044 14424
rect 12256 14408 12308 14414
rect 12256 14350 12308 14356
rect 12912 14346 12940 14418
rect 12900 14340 12952 14346
rect 12900 14282 12952 14288
rect 12406 13628 12714 13637
rect 12406 13626 12412 13628
rect 12468 13626 12492 13628
rect 12548 13626 12572 13628
rect 12628 13626 12652 13628
rect 12708 13626 12714 13628
rect 12468 13574 12470 13626
rect 12650 13574 12652 13626
rect 12406 13572 12412 13574
rect 12468 13572 12492 13574
rect 12548 13572 12572 13574
rect 12628 13572 12652 13574
rect 12708 13572 12714 13574
rect 12406 13563 12714 13572
rect 11612 13388 11664 13394
rect 11612 13330 11664 13336
rect 11336 12980 11388 12986
rect 11336 12922 11388 12928
rect 11204 12736 11284 12764
rect 11152 12718 11204 12724
rect 10508 12708 10560 12714
rect 10508 12650 10560 12656
rect 11348 12170 11376 12922
rect 11336 12164 11388 12170
rect 11336 12106 11388 12112
rect 10856 11996 11164 12005
rect 10856 11994 10862 11996
rect 10918 11994 10942 11996
rect 10998 11994 11022 11996
rect 11078 11994 11102 11996
rect 11158 11994 11164 11996
rect 10918 11942 10920 11994
rect 11100 11942 11102 11994
rect 10856 11940 10862 11942
rect 10918 11940 10942 11942
rect 10998 11940 11022 11942
rect 11078 11940 11102 11942
rect 11158 11940 11164 11942
rect 10856 11931 11164 11940
rect 11624 11286 11652 13330
rect 12440 13184 12492 13190
rect 12440 13126 12492 13132
rect 12452 12850 12480 13126
rect 12532 12912 12584 12918
rect 12716 12912 12768 12918
rect 12584 12860 12716 12866
rect 12532 12854 12768 12860
rect 12440 12844 12492 12850
rect 12544 12838 12756 12854
rect 12440 12786 12492 12792
rect 12912 12782 12940 14282
rect 13004 12850 13032 14418
rect 12992 12844 13044 12850
rect 12992 12786 13044 12792
rect 12532 12776 12584 12782
rect 12532 12718 12584 12724
rect 12900 12776 12952 12782
rect 12900 12718 12952 12724
rect 12544 12646 12572 12718
rect 12532 12640 12584 12646
rect 12532 12582 12584 12588
rect 12808 12640 12860 12646
rect 12808 12582 12860 12588
rect 12406 12540 12714 12549
rect 12406 12538 12412 12540
rect 12468 12538 12492 12540
rect 12548 12538 12572 12540
rect 12628 12538 12652 12540
rect 12708 12538 12714 12540
rect 12468 12486 12470 12538
rect 12650 12486 12652 12538
rect 12406 12484 12412 12486
rect 12468 12484 12492 12486
rect 12548 12484 12572 12486
rect 12628 12484 12652 12486
rect 12708 12484 12714 12486
rect 12406 12475 12714 12484
rect 11888 12368 11940 12374
rect 11888 12310 11940 12316
rect 11796 11552 11848 11558
rect 11796 11494 11848 11500
rect 11612 11280 11664 11286
rect 11612 11222 11664 11228
rect 9772 11212 9824 11218
rect 9772 11154 9824 11160
rect 9956 11212 10008 11218
rect 9956 11154 10008 11160
rect 9680 8288 9732 8294
rect 9680 8230 9732 8236
rect 9306 8188 9614 8197
rect 9306 8186 9312 8188
rect 9368 8186 9392 8188
rect 9448 8186 9472 8188
rect 9528 8186 9552 8188
rect 9608 8186 9614 8188
rect 9368 8134 9370 8186
rect 9550 8134 9552 8186
rect 9306 8132 9312 8134
rect 9368 8132 9392 8134
rect 9448 8132 9472 8134
rect 9528 8132 9552 8134
rect 9608 8132 9614 8134
rect 9306 8123 9614 8132
rect 9784 8022 9812 11154
rect 10232 11144 10284 11150
rect 10232 11086 10284 11092
rect 10244 10810 10272 11086
rect 11520 11008 11572 11014
rect 11520 10950 11572 10956
rect 10856 10908 11164 10917
rect 10856 10906 10862 10908
rect 10918 10906 10942 10908
rect 10998 10906 11022 10908
rect 11078 10906 11102 10908
rect 11158 10906 11164 10908
rect 10918 10854 10920 10906
rect 11100 10854 11102 10906
rect 10856 10852 10862 10854
rect 10918 10852 10942 10854
rect 10998 10852 11022 10854
rect 11078 10852 11102 10854
rect 11158 10852 11164 10854
rect 10856 10843 11164 10852
rect 10232 10804 10284 10810
rect 10232 10746 10284 10752
rect 11532 10606 11560 10950
rect 11808 10674 11836 11494
rect 11796 10668 11848 10674
rect 11796 10610 11848 10616
rect 11520 10600 11572 10606
rect 11520 10542 11572 10548
rect 11532 10130 11560 10542
rect 11520 10124 11572 10130
rect 11520 10066 11572 10072
rect 10784 9920 10836 9926
rect 10784 9862 10836 9868
rect 10796 9722 10824 9862
rect 10856 9820 11164 9829
rect 10856 9818 10862 9820
rect 10918 9818 10942 9820
rect 10998 9818 11022 9820
rect 11078 9818 11102 9820
rect 11158 9818 11164 9820
rect 10918 9766 10920 9818
rect 11100 9766 11102 9818
rect 10856 9764 10862 9766
rect 10918 9764 10942 9766
rect 10998 9764 11022 9766
rect 11078 9764 11102 9766
rect 11158 9764 11164 9766
rect 10856 9755 11164 9764
rect 10784 9716 10836 9722
rect 10784 9658 10836 9664
rect 10140 9512 10192 9518
rect 10140 9454 10192 9460
rect 9956 9376 10008 9382
rect 9956 9318 10008 9324
rect 9968 9042 9996 9318
rect 9956 9036 10008 9042
rect 9956 8978 10008 8984
rect 9956 8356 10008 8362
rect 9956 8298 10008 8304
rect 9772 8016 9824 8022
rect 9772 7958 9824 7964
rect 9220 7812 9272 7818
rect 9220 7754 9272 7760
rect 9232 7478 9260 7754
rect 9220 7472 9272 7478
rect 9220 7414 9272 7420
rect 9968 7342 9996 8298
rect 9956 7336 10008 7342
rect 9956 7278 10008 7284
rect 9306 7100 9614 7109
rect 9306 7098 9312 7100
rect 9368 7098 9392 7100
rect 9448 7098 9472 7100
rect 9528 7098 9552 7100
rect 9608 7098 9614 7100
rect 9368 7046 9370 7098
rect 9550 7046 9552 7098
rect 9306 7044 9312 7046
rect 9368 7044 9392 7046
rect 9448 7044 9472 7046
rect 9528 7044 9552 7046
rect 9608 7044 9614 7046
rect 9306 7035 9614 7044
rect 10152 6866 10180 9454
rect 10324 8968 10376 8974
rect 10324 8910 10376 8916
rect 10336 8634 10364 8910
rect 10324 8628 10376 8634
rect 10324 8570 10376 8576
rect 10416 7540 10468 7546
rect 10416 7482 10468 7488
rect 10140 6860 10192 6866
rect 10140 6802 10192 6808
rect 9036 6452 9088 6458
rect 9036 6394 9088 6400
rect 8760 6248 8812 6254
rect 8760 6190 8812 6196
rect 8668 5364 8720 5370
rect 8668 5306 8720 5312
rect 8680 4690 8708 5306
rect 8772 5234 8800 6190
rect 8944 6180 8996 6186
rect 8944 6122 8996 6128
rect 9128 6180 9180 6186
rect 9128 6122 9180 6128
rect 8760 5228 8812 5234
rect 8760 5170 8812 5176
rect 8760 5092 8812 5098
rect 8760 5034 8812 5040
rect 8484 4684 8536 4690
rect 8484 4626 8536 4632
rect 8668 4684 8720 4690
rect 8668 4626 8720 4632
rect 8680 3466 8708 4626
rect 8772 4486 8800 5034
rect 8852 4820 8904 4826
rect 8852 4762 8904 4768
rect 8760 4480 8812 4486
rect 8760 4422 8812 4428
rect 8864 4282 8892 4762
rect 8852 4276 8904 4282
rect 8852 4218 8904 4224
rect 8956 3942 8984 6122
rect 9140 5914 9168 6122
rect 9680 6112 9732 6118
rect 9680 6054 9732 6060
rect 9306 6012 9614 6021
rect 9306 6010 9312 6012
rect 9368 6010 9392 6012
rect 9448 6010 9472 6012
rect 9528 6010 9552 6012
rect 9608 6010 9614 6012
rect 9368 5958 9370 6010
rect 9550 5958 9552 6010
rect 9306 5956 9312 5958
rect 9368 5956 9392 5958
rect 9448 5956 9472 5958
rect 9528 5956 9552 5958
rect 9608 5956 9614 5958
rect 9306 5947 9614 5956
rect 9128 5908 9180 5914
rect 9128 5850 9180 5856
rect 9692 5098 9720 6054
rect 9680 5092 9732 5098
rect 9680 5034 9732 5040
rect 9772 5024 9824 5030
rect 9772 4966 9824 4972
rect 9306 4924 9614 4933
rect 9306 4922 9312 4924
rect 9368 4922 9392 4924
rect 9448 4922 9472 4924
rect 9528 4922 9552 4924
rect 9608 4922 9614 4924
rect 9368 4870 9370 4922
rect 9550 4870 9552 4922
rect 9306 4868 9312 4870
rect 9368 4868 9392 4870
rect 9448 4868 9472 4870
rect 9528 4868 9552 4870
rect 9608 4868 9614 4870
rect 9306 4859 9614 4868
rect 9784 4554 9812 4966
rect 10152 4690 10180 6802
rect 9956 4684 10008 4690
rect 9956 4626 10008 4632
rect 10140 4684 10192 4690
rect 10140 4626 10192 4632
rect 9772 4548 9824 4554
rect 9772 4490 9824 4496
rect 9036 4072 9088 4078
rect 9036 4014 9088 4020
rect 8944 3936 8996 3942
rect 8944 3878 8996 3884
rect 8392 3460 8444 3466
rect 8392 3402 8444 3408
rect 8668 3460 8720 3466
rect 8668 3402 8720 3408
rect 8208 2644 8260 2650
rect 8208 2586 8260 2592
rect 8404 2582 8432 3402
rect 9048 2650 9076 4014
rect 9306 3836 9614 3845
rect 9306 3834 9312 3836
rect 9368 3834 9392 3836
rect 9448 3834 9472 3836
rect 9528 3834 9552 3836
rect 9608 3834 9614 3836
rect 9368 3782 9370 3834
rect 9550 3782 9552 3834
rect 9306 3780 9312 3782
rect 9368 3780 9392 3782
rect 9448 3780 9472 3782
rect 9528 3780 9552 3782
rect 9608 3780 9614 3782
rect 9306 3771 9614 3780
rect 9680 3052 9732 3058
rect 9680 2994 9732 3000
rect 9306 2748 9614 2757
rect 9306 2746 9312 2748
rect 9368 2746 9392 2748
rect 9448 2746 9472 2748
rect 9528 2746 9552 2748
rect 9608 2746 9614 2748
rect 9368 2694 9370 2746
rect 9550 2694 9552 2746
rect 9306 2692 9312 2694
rect 9368 2692 9392 2694
rect 9448 2692 9472 2694
rect 9528 2692 9552 2694
rect 9608 2692 9614 2694
rect 9306 2683 9614 2692
rect 9036 2644 9088 2650
rect 9036 2586 9088 2592
rect 8392 2576 8444 2582
rect 8392 2518 8444 2524
rect 7756 2204 8064 2213
rect 7756 2202 7762 2204
rect 7818 2202 7842 2204
rect 7898 2202 7922 2204
rect 7978 2202 8002 2204
rect 8058 2202 8064 2204
rect 7818 2150 7820 2202
rect 8000 2150 8002 2202
rect 7756 2148 7762 2150
rect 7818 2148 7842 2150
rect 7898 2148 7922 2150
rect 7978 2148 8002 2150
rect 8058 2148 8064 2150
rect 7756 2139 8064 2148
rect 9048 2038 9076 2586
rect 9692 2446 9720 2994
rect 9680 2440 9732 2446
rect 9680 2382 9732 2388
rect 9036 2032 9088 2038
rect 9036 1974 9088 1980
rect 8024 1760 8076 1766
rect 8024 1702 8076 1708
rect 8036 1562 8064 1702
rect 8024 1556 8076 1562
rect 8024 1498 8076 1504
rect 9048 1494 9076 1974
rect 9220 1896 9272 1902
rect 9220 1838 9272 1844
rect 9232 1562 9260 1838
rect 9692 1766 9720 2382
rect 9784 1970 9812 4490
rect 9968 3738 9996 4626
rect 9956 3732 10008 3738
rect 9956 3674 10008 3680
rect 10232 3596 10284 3602
rect 10232 3538 10284 3544
rect 10244 3194 10272 3538
rect 10428 3534 10456 7482
rect 10796 7342 10824 9658
rect 11244 9104 11296 9110
rect 11244 9046 11296 9052
rect 10856 8732 11164 8741
rect 10856 8730 10862 8732
rect 10918 8730 10942 8732
rect 10998 8730 11022 8732
rect 11078 8730 11102 8732
rect 11158 8730 11164 8732
rect 10918 8678 10920 8730
rect 11100 8678 11102 8730
rect 10856 8676 10862 8678
rect 10918 8676 10942 8678
rect 10998 8676 11022 8678
rect 11078 8676 11102 8678
rect 11158 8676 11164 8678
rect 10856 8667 11164 8676
rect 10876 8288 10928 8294
rect 10876 8230 10928 8236
rect 10888 7954 10916 8230
rect 11256 8022 11284 9046
rect 11808 8498 11836 10610
rect 11900 10266 11928 12310
rect 12820 12306 12848 12582
rect 12912 12442 12940 12718
rect 13004 12646 13032 12786
rect 12992 12640 13044 12646
rect 12992 12582 13044 12588
rect 12900 12436 12952 12442
rect 12900 12378 12952 12384
rect 12808 12300 12860 12306
rect 12808 12242 12860 12248
rect 12912 12186 12940 12378
rect 12820 12158 12940 12186
rect 12820 11694 12848 12158
rect 12900 12096 12952 12102
rect 12900 12038 12952 12044
rect 12912 11762 12940 12038
rect 12900 11756 12952 11762
rect 12900 11698 12952 11704
rect 12808 11688 12860 11694
rect 12808 11630 12860 11636
rect 12406 11452 12714 11461
rect 12406 11450 12412 11452
rect 12468 11450 12492 11452
rect 12548 11450 12572 11452
rect 12628 11450 12652 11452
rect 12708 11450 12714 11452
rect 12468 11398 12470 11450
rect 12650 11398 12652 11450
rect 12406 11396 12412 11398
rect 12468 11396 12492 11398
rect 12548 11396 12572 11398
rect 12628 11396 12652 11398
rect 12708 11396 12714 11398
rect 12406 11387 12714 11396
rect 12820 10674 12848 11630
rect 12808 10668 12860 10674
rect 12808 10610 12860 10616
rect 12808 10532 12860 10538
rect 12808 10474 12860 10480
rect 12406 10364 12714 10373
rect 12406 10362 12412 10364
rect 12468 10362 12492 10364
rect 12548 10362 12572 10364
rect 12628 10362 12652 10364
rect 12708 10362 12714 10364
rect 12468 10310 12470 10362
rect 12650 10310 12652 10362
rect 12406 10308 12412 10310
rect 12468 10308 12492 10310
rect 12548 10308 12572 10310
rect 12628 10308 12652 10310
rect 12708 10308 12714 10310
rect 12406 10299 12714 10308
rect 12820 10266 12848 10474
rect 13176 10464 13228 10470
rect 13176 10406 13228 10412
rect 11888 10260 11940 10266
rect 11888 10202 11940 10208
rect 12348 10260 12400 10266
rect 12348 10202 12400 10208
rect 12808 10260 12860 10266
rect 12808 10202 12860 10208
rect 12360 10130 12388 10202
rect 12348 10124 12400 10130
rect 12348 10066 12400 10072
rect 11980 10056 12032 10062
rect 11980 9998 12032 10004
rect 12900 10056 12952 10062
rect 12900 9998 12952 10004
rect 11992 9518 12020 9998
rect 11980 9512 12032 9518
rect 11980 9454 12032 9460
rect 11992 9178 12020 9454
rect 12808 9376 12860 9382
rect 12808 9318 12860 9324
rect 12406 9276 12714 9285
rect 12406 9274 12412 9276
rect 12468 9274 12492 9276
rect 12548 9274 12572 9276
rect 12628 9274 12652 9276
rect 12708 9274 12714 9276
rect 12468 9222 12470 9274
rect 12650 9222 12652 9274
rect 12406 9220 12412 9222
rect 12468 9220 12492 9222
rect 12548 9220 12572 9222
rect 12628 9220 12652 9222
rect 12708 9220 12714 9222
rect 12406 9211 12714 9220
rect 12820 9178 12848 9318
rect 11980 9172 12032 9178
rect 11980 9114 12032 9120
rect 12808 9172 12860 9178
rect 12808 9114 12860 9120
rect 11796 8492 11848 8498
rect 11796 8434 11848 8440
rect 11244 8016 11296 8022
rect 11244 7958 11296 7964
rect 10876 7948 10928 7954
rect 10876 7890 10928 7896
rect 10856 7644 11164 7653
rect 10856 7642 10862 7644
rect 10918 7642 10942 7644
rect 10998 7642 11022 7644
rect 11078 7642 11102 7644
rect 11158 7642 11164 7644
rect 10918 7590 10920 7642
rect 11100 7590 11102 7642
rect 10856 7588 10862 7590
rect 10918 7588 10942 7590
rect 10998 7588 11022 7590
rect 11078 7588 11102 7590
rect 11158 7588 11164 7590
rect 10856 7579 11164 7588
rect 11256 7546 11284 7958
rect 11244 7540 11296 7546
rect 11244 7482 11296 7488
rect 10784 7336 10836 7342
rect 10784 7278 10836 7284
rect 10784 7200 10836 7206
rect 10784 7142 10836 7148
rect 11152 7200 11204 7206
rect 11152 7142 11204 7148
rect 10796 6186 10824 7142
rect 11164 6662 11192 7142
rect 11256 7018 11284 7482
rect 11808 7410 11836 8434
rect 11992 8430 12020 9114
rect 12624 8832 12676 8838
rect 12624 8774 12676 8780
rect 12636 8566 12664 8774
rect 12624 8560 12676 8566
rect 12624 8502 12676 8508
rect 11980 8424 12032 8430
rect 11980 8366 12032 8372
rect 12406 8188 12714 8197
rect 12406 8186 12412 8188
rect 12468 8186 12492 8188
rect 12548 8186 12572 8188
rect 12628 8186 12652 8188
rect 12708 8186 12714 8188
rect 12468 8134 12470 8186
rect 12650 8134 12652 8186
rect 12406 8132 12412 8134
rect 12468 8132 12492 8134
rect 12548 8132 12572 8134
rect 12628 8132 12652 8134
rect 12708 8132 12714 8134
rect 12406 8123 12714 8132
rect 12256 7540 12308 7546
rect 12256 7482 12308 7488
rect 11796 7404 11848 7410
rect 11796 7346 11848 7352
rect 11888 7336 11940 7342
rect 11888 7278 11940 7284
rect 11256 6990 11468 7018
rect 11900 7002 11928 7278
rect 11440 6934 11468 6990
rect 11888 6996 11940 7002
rect 11888 6938 11940 6944
rect 11428 6928 11480 6934
rect 11428 6870 11480 6876
rect 11152 6656 11204 6662
rect 11152 6598 11204 6604
rect 10856 6556 11164 6565
rect 10856 6554 10862 6556
rect 10918 6554 10942 6556
rect 10998 6554 11022 6556
rect 11078 6554 11102 6556
rect 11158 6554 11164 6556
rect 10918 6502 10920 6554
rect 11100 6502 11102 6554
rect 10856 6500 10862 6502
rect 10918 6500 10942 6502
rect 10998 6500 11022 6502
rect 11078 6500 11102 6502
rect 11158 6500 11164 6502
rect 10856 6491 11164 6500
rect 10784 6180 10836 6186
rect 10784 6122 10836 6128
rect 10416 3528 10468 3534
rect 10416 3470 10468 3476
rect 10232 3188 10284 3194
rect 10232 3130 10284 3136
rect 10428 3058 10456 3470
rect 10416 3052 10468 3058
rect 10416 2994 10468 3000
rect 9864 2848 9916 2854
rect 9864 2790 9916 2796
rect 9876 2106 9904 2790
rect 10796 2106 10824 6122
rect 10856 5468 11164 5477
rect 10856 5466 10862 5468
rect 10918 5466 10942 5468
rect 10998 5466 11022 5468
rect 11078 5466 11102 5468
rect 11158 5466 11164 5468
rect 10918 5414 10920 5466
rect 11100 5414 11102 5466
rect 10856 5412 10862 5414
rect 10918 5412 10942 5414
rect 10998 5412 11022 5414
rect 11078 5412 11102 5414
rect 11158 5412 11164 5414
rect 10856 5403 11164 5412
rect 12268 5030 12296 7482
rect 12912 7342 12940 9998
rect 13188 9926 13216 10406
rect 13280 10130 13308 15506
rect 13464 12866 13492 15574
rect 13648 15162 13676 16594
rect 13740 16130 13768 16934
rect 13832 16726 13860 17138
rect 14096 17060 14148 17066
rect 14096 17002 14148 17008
rect 14004 16992 14056 16998
rect 14004 16934 14056 16940
rect 14016 16794 14044 16934
rect 14108 16794 14136 17002
rect 14004 16788 14056 16794
rect 14004 16730 14056 16736
rect 14096 16788 14148 16794
rect 14096 16730 14148 16736
rect 13820 16720 13872 16726
rect 13820 16662 13872 16668
rect 14278 16688 14334 16697
rect 13832 16250 13860 16662
rect 14278 16623 14334 16632
rect 14292 16590 14320 16623
rect 14280 16584 14332 16590
rect 14280 16526 14332 16532
rect 14280 16448 14332 16454
rect 14280 16390 14332 16396
rect 13956 16348 14264 16357
rect 13956 16346 13962 16348
rect 14018 16346 14042 16348
rect 14098 16346 14122 16348
rect 14178 16346 14202 16348
rect 14258 16346 14264 16348
rect 14018 16294 14020 16346
rect 14200 16294 14202 16346
rect 13956 16292 13962 16294
rect 14018 16292 14042 16294
rect 14098 16292 14122 16294
rect 14178 16292 14202 16294
rect 14258 16292 14264 16294
rect 13956 16283 14264 16292
rect 13820 16244 13872 16250
rect 13820 16186 13872 16192
rect 13740 16102 13860 16130
rect 13832 15502 13860 16102
rect 14292 15706 14320 16390
rect 14280 15700 14332 15706
rect 14280 15642 14332 15648
rect 14384 15638 14412 18158
rect 14648 18148 14700 18154
rect 14648 18090 14700 18096
rect 14832 18148 14884 18154
rect 14832 18090 14884 18096
rect 14372 15632 14424 15638
rect 14372 15574 14424 15580
rect 13820 15496 13872 15502
rect 13820 15438 13872 15444
rect 13636 15156 13688 15162
rect 13636 15098 13688 15104
rect 13728 14884 13780 14890
rect 13728 14826 13780 14832
rect 13740 14550 13768 14826
rect 13728 14544 13780 14550
rect 13728 14486 13780 14492
rect 13544 14272 13596 14278
rect 13544 14214 13596 14220
rect 13556 13870 13584 14214
rect 13832 14074 13860 15438
rect 13956 15260 14264 15269
rect 13956 15258 13962 15260
rect 14018 15258 14042 15260
rect 14098 15258 14122 15260
rect 14178 15258 14202 15260
rect 14258 15258 14264 15260
rect 14018 15206 14020 15258
rect 14200 15206 14202 15258
rect 13956 15204 13962 15206
rect 14018 15204 14042 15206
rect 14098 15204 14122 15206
rect 14178 15204 14202 15206
rect 14258 15204 14264 15206
rect 13956 15195 14264 15204
rect 13912 14952 13964 14958
rect 13912 14894 13964 14900
rect 13924 14346 13952 14894
rect 14660 14822 14688 18090
rect 14844 17746 14872 18090
rect 14832 17740 14884 17746
rect 14832 17682 14884 17688
rect 14738 16688 14794 16697
rect 14738 16623 14794 16632
rect 14280 14816 14332 14822
rect 14280 14758 14332 14764
rect 14648 14816 14700 14822
rect 14648 14758 14700 14764
rect 14292 14618 14320 14758
rect 14280 14612 14332 14618
rect 14280 14554 14332 14560
rect 14372 14612 14424 14618
rect 14372 14554 14424 14560
rect 14280 14476 14332 14482
rect 14280 14418 14332 14424
rect 13912 14340 13964 14346
rect 13912 14282 13964 14288
rect 13956 14172 14264 14181
rect 13956 14170 13962 14172
rect 14018 14170 14042 14172
rect 14098 14170 14122 14172
rect 14178 14170 14202 14172
rect 14258 14170 14264 14172
rect 14018 14118 14020 14170
rect 14200 14118 14202 14170
rect 13956 14116 13962 14118
rect 14018 14116 14042 14118
rect 14098 14116 14122 14118
rect 14178 14116 14202 14118
rect 14258 14116 14264 14118
rect 13956 14107 14264 14116
rect 14292 14074 14320 14418
rect 13820 14068 13872 14074
rect 13820 14010 13872 14016
rect 14280 14068 14332 14074
rect 14280 14010 14332 14016
rect 13544 13864 13596 13870
rect 13544 13806 13596 13812
rect 13832 13682 13860 14010
rect 14384 13938 14412 14554
rect 14648 14544 14700 14550
rect 14648 14486 14700 14492
rect 14660 14346 14688 14486
rect 14648 14340 14700 14346
rect 14648 14282 14700 14288
rect 14372 13932 14424 13938
rect 14372 13874 14424 13880
rect 13740 13654 13860 13682
rect 13464 12838 13676 12866
rect 13648 10130 13676 12838
rect 13740 12306 13768 13654
rect 13820 13524 13872 13530
rect 13820 13466 13872 13472
rect 13728 12300 13780 12306
rect 13728 12242 13780 12248
rect 13268 10124 13320 10130
rect 13268 10066 13320 10072
rect 13636 10124 13688 10130
rect 13636 10066 13688 10072
rect 13176 9920 13228 9926
rect 13176 9862 13228 9868
rect 13084 8968 13136 8974
rect 13084 8910 13136 8916
rect 13096 8634 13124 8910
rect 13084 8628 13136 8634
rect 13084 8570 13136 8576
rect 13188 8430 13216 9862
rect 13280 9722 13308 10066
rect 13728 10056 13780 10062
rect 13728 9998 13780 10004
rect 13268 9716 13320 9722
rect 13268 9658 13320 9664
rect 13280 9110 13308 9658
rect 13268 9104 13320 9110
rect 13268 9046 13320 9052
rect 13544 9104 13596 9110
rect 13544 9046 13596 9052
rect 13268 8968 13320 8974
rect 13268 8910 13320 8916
rect 13176 8424 13228 8430
rect 13176 8366 13228 8372
rect 13280 8090 13308 8910
rect 13268 8084 13320 8090
rect 13268 8026 13320 8032
rect 13280 7410 13308 8026
rect 13268 7404 13320 7410
rect 13268 7346 13320 7352
rect 12900 7336 12952 7342
rect 12900 7278 12952 7284
rect 12808 7200 12860 7206
rect 12808 7142 12860 7148
rect 12406 7100 12714 7109
rect 12406 7098 12412 7100
rect 12468 7098 12492 7100
rect 12548 7098 12572 7100
rect 12628 7098 12652 7100
rect 12708 7098 12714 7100
rect 12468 7046 12470 7098
rect 12650 7046 12652 7098
rect 12406 7044 12412 7046
rect 12468 7044 12492 7046
rect 12548 7044 12572 7046
rect 12628 7044 12652 7046
rect 12708 7044 12714 7046
rect 12406 7035 12714 7044
rect 12820 6458 12848 7142
rect 12808 6452 12860 6458
rect 12808 6394 12860 6400
rect 12406 6012 12714 6021
rect 12406 6010 12412 6012
rect 12468 6010 12492 6012
rect 12548 6010 12572 6012
rect 12628 6010 12652 6012
rect 12708 6010 12714 6012
rect 12468 5958 12470 6010
rect 12650 5958 12652 6010
rect 12406 5956 12412 5958
rect 12468 5956 12492 5958
rect 12548 5956 12572 5958
rect 12628 5956 12652 5958
rect 12708 5956 12714 5958
rect 12406 5947 12714 5956
rect 12808 5160 12860 5166
rect 12808 5102 12860 5108
rect 11888 5024 11940 5030
rect 11888 4966 11940 4972
rect 12256 5024 12308 5030
rect 12256 4966 12308 4972
rect 11900 4622 11928 4966
rect 12268 4758 12296 4966
rect 12406 4924 12714 4933
rect 12406 4922 12412 4924
rect 12468 4922 12492 4924
rect 12548 4922 12572 4924
rect 12628 4922 12652 4924
rect 12708 4922 12714 4924
rect 12468 4870 12470 4922
rect 12650 4870 12652 4922
rect 12406 4868 12412 4870
rect 12468 4868 12492 4870
rect 12548 4868 12572 4870
rect 12628 4868 12652 4870
rect 12708 4868 12714 4870
rect 12406 4859 12714 4868
rect 12820 4826 12848 5102
rect 12808 4820 12860 4826
rect 12808 4762 12860 4768
rect 13280 4758 13308 7346
rect 13556 6866 13584 9046
rect 13740 9042 13768 9998
rect 13832 9042 13860 13466
rect 14372 13388 14424 13394
rect 14372 13330 14424 13336
rect 13956 13084 14264 13093
rect 13956 13082 13962 13084
rect 14018 13082 14042 13084
rect 14098 13082 14122 13084
rect 14178 13082 14202 13084
rect 14258 13082 14264 13084
rect 14018 13030 14020 13082
rect 14200 13030 14202 13082
rect 13956 13028 13962 13030
rect 14018 13028 14042 13030
rect 14098 13028 14122 13030
rect 14178 13028 14202 13030
rect 14258 13028 14264 13030
rect 13956 13019 14264 13028
rect 14004 12776 14056 12782
rect 14004 12718 14056 12724
rect 14016 12374 14044 12718
rect 14188 12436 14240 12442
rect 14188 12378 14240 12384
rect 14004 12368 14056 12374
rect 14004 12310 14056 12316
rect 14200 12238 14228 12378
rect 14004 12232 14056 12238
rect 14004 12174 14056 12180
rect 14188 12232 14240 12238
rect 14188 12174 14240 12180
rect 14016 12102 14044 12174
rect 14280 12164 14332 12170
rect 14280 12106 14332 12112
rect 14004 12096 14056 12102
rect 14004 12038 14056 12044
rect 13956 11996 14264 12005
rect 13956 11994 13962 11996
rect 14018 11994 14042 11996
rect 14098 11994 14122 11996
rect 14178 11994 14202 11996
rect 14258 11994 14264 11996
rect 14018 11942 14020 11994
rect 14200 11942 14202 11994
rect 13956 11940 13962 11942
rect 14018 11940 14042 11942
rect 14098 11940 14122 11942
rect 14178 11940 14202 11942
rect 14258 11940 14264 11942
rect 13956 11931 14264 11940
rect 14292 11898 14320 12106
rect 14280 11892 14332 11898
rect 14280 11834 14332 11840
rect 14188 11688 14240 11694
rect 14188 11630 14240 11636
rect 14200 11558 14228 11630
rect 14384 11558 14412 13330
rect 14660 12782 14688 14282
rect 14752 13870 14780 16623
rect 14832 15360 14884 15366
rect 14832 15302 14884 15308
rect 14844 14958 14872 15302
rect 14832 14952 14884 14958
rect 14832 14894 14884 14900
rect 14832 14816 14884 14822
rect 14832 14758 14884 14764
rect 14740 13864 14792 13870
rect 14740 13806 14792 13812
rect 14752 13190 14780 13806
rect 14740 13184 14792 13190
rect 14740 13126 14792 13132
rect 14844 12782 14872 14758
rect 14936 13530 14964 18158
rect 15108 17672 15160 17678
rect 15108 17614 15160 17620
rect 15016 15972 15068 15978
rect 15016 15914 15068 15920
rect 15028 15366 15056 15914
rect 15016 15360 15068 15366
rect 15016 15302 15068 15308
rect 14924 13524 14976 13530
rect 14924 13466 14976 13472
rect 15028 13462 15056 15302
rect 15120 15162 15148 17614
rect 15108 15156 15160 15162
rect 15108 15098 15160 15104
rect 15200 15020 15252 15026
rect 15200 14962 15252 14968
rect 15212 14414 15240 14962
rect 15200 14408 15252 14414
rect 15200 14350 15252 14356
rect 15212 14074 15240 14350
rect 15292 14272 15344 14278
rect 15292 14214 15344 14220
rect 15200 14068 15252 14074
rect 15200 14010 15252 14016
rect 15016 13456 15068 13462
rect 15016 13398 15068 13404
rect 14648 12776 14700 12782
rect 14568 12724 14648 12730
rect 14568 12718 14700 12724
rect 14832 12776 14884 12782
rect 14832 12718 14884 12724
rect 14568 12702 14688 12718
rect 14464 12096 14516 12102
rect 14464 12038 14516 12044
rect 14188 11552 14240 11558
rect 14188 11494 14240 11500
rect 14372 11552 14424 11558
rect 14372 11494 14424 11500
rect 14200 11098 14228 11494
rect 14200 11070 14320 11098
rect 13956 10908 14264 10917
rect 13956 10906 13962 10908
rect 14018 10906 14042 10908
rect 14098 10906 14122 10908
rect 14178 10906 14202 10908
rect 14258 10906 14264 10908
rect 14018 10854 14020 10906
rect 14200 10854 14202 10906
rect 13956 10852 13962 10854
rect 14018 10852 14042 10854
rect 14098 10852 14122 10854
rect 14178 10852 14202 10854
rect 14258 10852 14264 10854
rect 13956 10843 14264 10852
rect 13956 9820 14264 9829
rect 13956 9818 13962 9820
rect 14018 9818 14042 9820
rect 14098 9818 14122 9820
rect 14178 9818 14202 9820
rect 14258 9818 14264 9820
rect 14018 9766 14020 9818
rect 14200 9766 14202 9818
rect 13956 9764 13962 9766
rect 14018 9764 14042 9766
rect 14098 9764 14122 9766
rect 14178 9764 14202 9766
rect 14258 9764 14264 9766
rect 13956 9755 14264 9764
rect 13728 9036 13780 9042
rect 13728 8978 13780 8984
rect 13820 9036 13872 9042
rect 13820 8978 13872 8984
rect 13820 8900 13872 8906
rect 13820 8842 13872 8848
rect 13636 8832 13688 8838
rect 13636 8774 13688 8780
rect 13648 8430 13676 8774
rect 13832 8634 13860 8842
rect 13956 8732 14264 8741
rect 13956 8730 13962 8732
rect 14018 8730 14042 8732
rect 14098 8730 14122 8732
rect 14178 8730 14202 8732
rect 14258 8730 14264 8732
rect 14018 8678 14020 8730
rect 14200 8678 14202 8730
rect 13956 8676 13962 8678
rect 14018 8676 14042 8678
rect 14098 8676 14122 8678
rect 14178 8676 14202 8678
rect 14258 8676 14264 8678
rect 13956 8667 14264 8676
rect 13820 8628 13872 8634
rect 13820 8570 13872 8576
rect 13636 8424 13688 8430
rect 13832 8378 13860 8570
rect 13636 8366 13688 8372
rect 13740 8350 13860 8378
rect 13544 6860 13596 6866
rect 13544 6802 13596 6808
rect 13556 6662 13584 6802
rect 13544 6656 13596 6662
rect 13544 6598 13596 6604
rect 13740 6458 13768 8350
rect 13820 7744 13872 7750
rect 13820 7686 13872 7692
rect 13832 7342 13860 7686
rect 13956 7644 14264 7653
rect 13956 7642 13962 7644
rect 14018 7642 14042 7644
rect 14098 7642 14122 7644
rect 14178 7642 14202 7644
rect 14258 7642 14264 7644
rect 14018 7590 14020 7642
rect 14200 7590 14202 7642
rect 13956 7588 13962 7590
rect 14018 7588 14042 7590
rect 14098 7588 14122 7590
rect 14178 7588 14202 7590
rect 14258 7588 14264 7590
rect 13956 7579 14264 7588
rect 13820 7336 13872 7342
rect 13820 7278 13872 7284
rect 13832 6934 13860 7278
rect 13820 6928 13872 6934
rect 13820 6870 13872 6876
rect 13728 6452 13780 6458
rect 13728 6394 13780 6400
rect 13740 6254 13768 6394
rect 13728 6248 13780 6254
rect 13728 6190 13780 6196
rect 13832 5914 13860 6870
rect 13956 6556 14264 6565
rect 13956 6554 13962 6556
rect 14018 6554 14042 6556
rect 14098 6554 14122 6556
rect 14178 6554 14202 6556
rect 14258 6554 14264 6556
rect 14018 6502 14020 6554
rect 14200 6502 14202 6554
rect 13956 6500 13962 6502
rect 14018 6500 14042 6502
rect 14098 6500 14122 6502
rect 14178 6500 14202 6502
rect 14258 6500 14264 6502
rect 13956 6491 14264 6500
rect 13544 5908 13596 5914
rect 13544 5850 13596 5856
rect 13820 5908 13872 5914
rect 13820 5850 13872 5856
rect 13556 5234 13584 5850
rect 13956 5468 14264 5477
rect 13956 5466 13962 5468
rect 14018 5466 14042 5468
rect 14098 5466 14122 5468
rect 14178 5466 14202 5468
rect 14258 5466 14264 5468
rect 14018 5414 14020 5466
rect 14200 5414 14202 5466
rect 13956 5412 13962 5414
rect 14018 5412 14042 5414
rect 14098 5412 14122 5414
rect 14178 5412 14202 5414
rect 14258 5412 14264 5414
rect 13956 5403 14264 5412
rect 13544 5228 13596 5234
rect 13544 5170 13596 5176
rect 13820 5092 13872 5098
rect 13820 5034 13872 5040
rect 13832 4826 13860 5034
rect 13820 4820 13872 4826
rect 13820 4762 13872 4768
rect 14292 4758 14320 11070
rect 14384 8022 14412 11494
rect 14476 11218 14504 12038
rect 14464 11212 14516 11218
rect 14464 11154 14516 11160
rect 14568 10062 14596 12702
rect 14648 12436 14700 12442
rect 14648 12378 14700 12384
rect 14660 11286 14688 12378
rect 14740 11552 14792 11558
rect 14740 11494 14792 11500
rect 14648 11280 14700 11286
rect 14648 11222 14700 11228
rect 14752 11218 14780 11494
rect 14740 11212 14792 11218
rect 14740 11154 14792 11160
rect 14556 10056 14608 10062
rect 14556 9998 14608 10004
rect 14844 8922 14872 12718
rect 15016 12368 15068 12374
rect 15016 12310 15068 12316
rect 15028 12238 15056 12310
rect 15016 12232 15068 12238
rect 15016 12174 15068 12180
rect 15200 12232 15252 12238
rect 15200 12174 15252 12180
rect 15108 12164 15160 12170
rect 15108 12106 15160 12112
rect 15120 9674 15148 12106
rect 15212 11898 15240 12174
rect 15200 11892 15252 11898
rect 15200 11834 15252 11840
rect 15212 10810 15240 11834
rect 15304 11694 15332 14214
rect 15292 11688 15344 11694
rect 15292 11630 15344 11636
rect 15396 11626 15424 19230
rect 15580 19122 15608 19230
rect 15658 19200 15714 20000
rect 18510 19200 18566 20000
rect 15672 19122 15700 19200
rect 15580 19094 15700 19122
rect 18418 18592 18474 18601
rect 17056 18524 17364 18533
rect 18418 18527 18474 18536
rect 17056 18522 17062 18524
rect 17118 18522 17142 18524
rect 17198 18522 17222 18524
rect 17278 18522 17302 18524
rect 17358 18522 17364 18524
rect 17118 18470 17120 18522
rect 17300 18470 17302 18522
rect 17056 18468 17062 18470
rect 17118 18468 17142 18470
rect 17198 18468 17222 18470
rect 17278 18468 17302 18470
rect 17358 18468 17364 18470
rect 17056 18459 17364 18468
rect 18432 18426 18460 18527
rect 18420 18420 18472 18426
rect 18420 18362 18472 18368
rect 18432 18222 18460 18362
rect 16672 18216 16724 18222
rect 16672 18158 16724 18164
rect 18420 18216 18472 18222
rect 18420 18158 18472 18164
rect 15936 18080 15988 18086
rect 15936 18022 15988 18028
rect 16580 18080 16632 18086
rect 16580 18022 16632 18028
rect 15506 17980 15814 17989
rect 15506 17978 15512 17980
rect 15568 17978 15592 17980
rect 15648 17978 15672 17980
rect 15728 17978 15752 17980
rect 15808 17978 15814 17980
rect 15568 17926 15570 17978
rect 15750 17926 15752 17978
rect 15506 17924 15512 17926
rect 15568 17924 15592 17926
rect 15648 17924 15672 17926
rect 15728 17924 15752 17926
rect 15808 17924 15814 17926
rect 15506 17915 15814 17924
rect 15506 16892 15814 16901
rect 15506 16890 15512 16892
rect 15568 16890 15592 16892
rect 15648 16890 15672 16892
rect 15728 16890 15752 16892
rect 15808 16890 15814 16892
rect 15568 16838 15570 16890
rect 15750 16838 15752 16890
rect 15506 16836 15512 16838
rect 15568 16836 15592 16838
rect 15648 16836 15672 16838
rect 15728 16836 15752 16838
rect 15808 16836 15814 16838
rect 15506 16827 15814 16836
rect 15948 16590 15976 18022
rect 16120 17808 16172 17814
rect 16120 17750 16172 17756
rect 16132 17218 16160 17750
rect 16304 17604 16356 17610
rect 16304 17546 16356 17552
rect 16040 17190 16160 17218
rect 16040 17134 16068 17190
rect 16028 17128 16080 17134
rect 16028 17070 16080 17076
rect 16212 17128 16264 17134
rect 16212 17070 16264 17076
rect 15936 16584 15988 16590
rect 15936 16526 15988 16532
rect 16224 16046 16252 17070
rect 16316 16697 16344 17546
rect 16592 16998 16620 18022
rect 16684 17338 16712 18158
rect 16764 17740 16816 17746
rect 16764 17682 16816 17688
rect 16672 17332 16724 17338
rect 16672 17274 16724 17280
rect 16580 16992 16632 16998
rect 16580 16934 16632 16940
rect 16776 16726 16804 17682
rect 16856 17536 16908 17542
rect 16856 17478 16908 17484
rect 16764 16720 16816 16726
rect 16302 16688 16358 16697
rect 16764 16662 16816 16668
rect 16302 16623 16358 16632
rect 16396 16448 16448 16454
rect 16396 16390 16448 16396
rect 16764 16448 16816 16454
rect 16764 16390 16816 16396
rect 16212 16040 16264 16046
rect 16212 15982 16264 15988
rect 15506 15804 15814 15813
rect 15506 15802 15512 15804
rect 15568 15802 15592 15804
rect 15648 15802 15672 15804
rect 15728 15802 15752 15804
rect 15808 15802 15814 15804
rect 15568 15750 15570 15802
rect 15750 15750 15752 15802
rect 15506 15748 15512 15750
rect 15568 15748 15592 15750
rect 15648 15748 15672 15750
rect 15728 15748 15752 15750
rect 15808 15748 15814 15750
rect 15506 15739 15814 15748
rect 16224 14958 16252 15982
rect 16304 15632 16356 15638
rect 16304 15574 16356 15580
rect 16212 14952 16264 14958
rect 16212 14894 16264 14900
rect 15506 14716 15814 14725
rect 15506 14714 15512 14716
rect 15568 14714 15592 14716
rect 15648 14714 15672 14716
rect 15728 14714 15752 14716
rect 15808 14714 15814 14716
rect 15568 14662 15570 14714
rect 15750 14662 15752 14714
rect 15506 14660 15512 14662
rect 15568 14660 15592 14662
rect 15648 14660 15672 14662
rect 15728 14660 15752 14662
rect 15808 14660 15814 14662
rect 15506 14651 15814 14660
rect 15752 14476 15804 14482
rect 15752 14418 15804 14424
rect 15936 14476 15988 14482
rect 15936 14418 15988 14424
rect 15764 14278 15792 14418
rect 15752 14272 15804 14278
rect 15752 14214 15804 14220
rect 15844 13864 15896 13870
rect 15844 13806 15896 13812
rect 15506 13628 15814 13637
rect 15506 13626 15512 13628
rect 15568 13626 15592 13628
rect 15648 13626 15672 13628
rect 15728 13626 15752 13628
rect 15808 13626 15814 13628
rect 15568 13574 15570 13626
rect 15750 13574 15752 13626
rect 15506 13572 15512 13574
rect 15568 13572 15592 13574
rect 15648 13572 15672 13574
rect 15728 13572 15752 13574
rect 15808 13572 15814 13574
rect 15506 13563 15814 13572
rect 15506 12540 15814 12549
rect 15506 12538 15512 12540
rect 15568 12538 15592 12540
rect 15648 12538 15672 12540
rect 15728 12538 15752 12540
rect 15808 12538 15814 12540
rect 15568 12486 15570 12538
rect 15750 12486 15752 12538
rect 15506 12484 15512 12486
rect 15568 12484 15592 12486
rect 15648 12484 15672 12486
rect 15728 12484 15752 12486
rect 15808 12484 15814 12486
rect 15506 12475 15814 12484
rect 15568 12436 15620 12442
rect 15568 12378 15620 12384
rect 15580 11694 15608 12378
rect 15568 11688 15620 11694
rect 15568 11630 15620 11636
rect 15384 11620 15436 11626
rect 15384 11562 15436 11568
rect 15506 11452 15814 11461
rect 15506 11450 15512 11452
rect 15568 11450 15592 11452
rect 15648 11450 15672 11452
rect 15728 11450 15752 11452
rect 15808 11450 15814 11452
rect 15568 11398 15570 11450
rect 15750 11398 15752 11450
rect 15506 11396 15512 11398
rect 15568 11396 15592 11398
rect 15648 11396 15672 11398
rect 15728 11396 15752 11398
rect 15808 11396 15814 11398
rect 15506 11387 15814 11396
rect 15568 11008 15620 11014
rect 15568 10950 15620 10956
rect 15200 10804 15252 10810
rect 15200 10746 15252 10752
rect 15580 10606 15608 10950
rect 15568 10600 15620 10606
rect 15568 10542 15620 10548
rect 15506 10364 15814 10373
rect 15506 10362 15512 10364
rect 15568 10362 15592 10364
rect 15648 10362 15672 10364
rect 15728 10362 15752 10364
rect 15808 10362 15814 10364
rect 15568 10310 15570 10362
rect 15750 10310 15752 10362
rect 15506 10308 15512 10310
rect 15568 10308 15592 10310
rect 15648 10308 15672 10310
rect 15728 10308 15752 10310
rect 15808 10308 15814 10310
rect 15506 10299 15814 10308
rect 15120 9646 15424 9674
rect 15200 9512 15252 9518
rect 15252 9472 15332 9500
rect 15200 9454 15252 9460
rect 15304 9382 15332 9472
rect 15108 9376 15160 9382
rect 15108 9318 15160 9324
rect 15292 9376 15344 9382
rect 15292 9318 15344 9324
rect 15120 9042 15148 9318
rect 15108 9036 15160 9042
rect 15108 8978 15160 8984
rect 14752 8906 14872 8922
rect 14740 8900 14872 8906
rect 14792 8894 14872 8900
rect 14740 8842 14792 8848
rect 14372 8016 14424 8022
rect 14372 7958 14424 7964
rect 15200 7948 15252 7954
rect 15200 7890 15252 7896
rect 14740 7744 14792 7750
rect 14740 7686 14792 7692
rect 14752 7410 14780 7686
rect 14740 7404 14792 7410
rect 14740 7346 14792 7352
rect 15016 7200 15068 7206
rect 15016 7142 15068 7148
rect 15028 6798 15056 7142
rect 15212 7002 15240 7890
rect 15200 6996 15252 7002
rect 15200 6938 15252 6944
rect 15304 6882 15332 9318
rect 15396 7818 15424 9646
rect 15506 9276 15814 9285
rect 15506 9274 15512 9276
rect 15568 9274 15592 9276
rect 15648 9274 15672 9276
rect 15728 9274 15752 9276
rect 15808 9274 15814 9276
rect 15568 9222 15570 9274
rect 15750 9222 15752 9274
rect 15506 9220 15512 9222
rect 15568 9220 15592 9222
rect 15648 9220 15672 9222
rect 15728 9220 15752 9222
rect 15808 9220 15814 9222
rect 15506 9211 15814 9220
rect 15506 8188 15814 8197
rect 15506 8186 15512 8188
rect 15568 8186 15592 8188
rect 15648 8186 15672 8188
rect 15728 8186 15752 8188
rect 15808 8186 15814 8188
rect 15568 8134 15570 8186
rect 15750 8134 15752 8186
rect 15506 8132 15512 8134
rect 15568 8132 15592 8134
rect 15648 8132 15672 8134
rect 15728 8132 15752 8134
rect 15808 8132 15814 8134
rect 15506 8123 15814 8132
rect 15856 8022 15884 13806
rect 15948 12986 15976 14418
rect 16120 14272 16172 14278
rect 16120 14214 16172 14220
rect 15936 12980 15988 12986
rect 15936 12922 15988 12928
rect 15948 12782 15976 12922
rect 16132 12782 16160 14214
rect 16224 13870 16252 14894
rect 16316 14414 16344 15574
rect 16408 14482 16436 16390
rect 16776 16114 16804 16390
rect 16764 16108 16816 16114
rect 16764 16050 16816 16056
rect 16488 15564 16540 15570
rect 16488 15506 16540 15512
rect 16396 14476 16448 14482
rect 16396 14418 16448 14424
rect 16304 14408 16356 14414
rect 16304 14350 16356 14356
rect 16212 13864 16264 13870
rect 16212 13806 16264 13812
rect 16224 13530 16252 13806
rect 16212 13524 16264 13530
rect 16212 13466 16264 13472
rect 16500 12986 16528 15506
rect 16868 15026 16896 17478
rect 17056 17436 17364 17445
rect 17056 17434 17062 17436
rect 17118 17434 17142 17436
rect 17198 17434 17222 17436
rect 17278 17434 17302 17436
rect 17358 17434 17364 17436
rect 17118 17382 17120 17434
rect 17300 17382 17302 17434
rect 17056 17380 17062 17382
rect 17118 17380 17142 17382
rect 17198 17380 17222 17382
rect 17278 17380 17302 17382
rect 17358 17380 17364 17382
rect 17056 17371 17364 17380
rect 18236 17196 18288 17202
rect 18236 17138 18288 17144
rect 17500 17060 17552 17066
rect 17500 17002 17552 17008
rect 17512 16726 17540 17002
rect 17776 16992 17828 16998
rect 17776 16934 17828 16940
rect 17500 16720 17552 16726
rect 17500 16662 17552 16668
rect 17056 16348 17364 16357
rect 17056 16346 17062 16348
rect 17118 16346 17142 16348
rect 17198 16346 17222 16348
rect 17278 16346 17302 16348
rect 17358 16346 17364 16348
rect 17118 16294 17120 16346
rect 17300 16294 17302 16346
rect 17056 16292 17062 16294
rect 17118 16292 17142 16294
rect 17198 16292 17222 16294
rect 17278 16292 17302 16294
rect 17358 16292 17364 16294
rect 17056 16283 17364 16292
rect 17512 15978 17540 16662
rect 17788 16658 17816 16934
rect 17776 16652 17828 16658
rect 17776 16594 17828 16600
rect 17500 15972 17552 15978
rect 17500 15914 17552 15920
rect 17056 15260 17364 15269
rect 17056 15258 17062 15260
rect 17118 15258 17142 15260
rect 17198 15258 17222 15260
rect 17278 15258 17302 15260
rect 17358 15258 17364 15260
rect 17118 15206 17120 15258
rect 17300 15206 17302 15258
rect 17056 15204 17062 15206
rect 17118 15204 17142 15206
rect 17198 15204 17222 15206
rect 17278 15204 17302 15206
rect 17358 15204 17364 15206
rect 17056 15195 17364 15204
rect 16856 15020 16908 15026
rect 16856 14962 16908 14968
rect 17512 14940 17540 15914
rect 17868 15904 17920 15910
rect 17868 15846 17920 15852
rect 17880 15638 17908 15846
rect 18248 15706 18276 17138
rect 18420 16652 18472 16658
rect 18420 16594 18472 16600
rect 18432 16182 18460 16594
rect 18420 16176 18472 16182
rect 18418 16144 18420 16153
rect 18472 16144 18474 16153
rect 18418 16079 18474 16088
rect 18236 15700 18288 15706
rect 18236 15642 18288 15648
rect 17868 15632 17920 15638
rect 17868 15574 17920 15580
rect 17592 14952 17644 14958
rect 17512 14912 17592 14940
rect 17592 14894 17644 14900
rect 16764 14884 16816 14890
rect 16764 14826 16816 14832
rect 16580 14816 16632 14822
rect 16580 14758 16632 14764
rect 16592 14482 16620 14758
rect 16776 14618 16804 14826
rect 16672 14612 16724 14618
rect 16672 14554 16724 14560
rect 16764 14612 16816 14618
rect 16764 14554 16816 14560
rect 16580 14476 16632 14482
rect 16580 14418 16632 14424
rect 16684 14396 16712 14554
rect 16948 14476 17000 14482
rect 16948 14418 17000 14424
rect 16684 14368 16896 14396
rect 16580 13456 16632 13462
rect 16580 13398 16632 13404
rect 16396 12980 16448 12986
rect 16396 12922 16448 12928
rect 16488 12980 16540 12986
rect 16488 12922 16540 12928
rect 15936 12776 15988 12782
rect 15936 12718 15988 12724
rect 16120 12776 16172 12782
rect 16120 12718 16172 12724
rect 16304 12776 16356 12782
rect 16304 12718 16356 12724
rect 16316 12374 16344 12718
rect 16304 12368 16356 12374
rect 16304 12310 16356 12316
rect 16212 12300 16264 12306
rect 16212 12242 16264 12248
rect 15936 12232 15988 12238
rect 15936 12174 15988 12180
rect 15948 11014 15976 12174
rect 16120 11280 16172 11286
rect 16120 11222 16172 11228
rect 15936 11008 15988 11014
rect 15936 10950 15988 10956
rect 15936 9444 15988 9450
rect 15936 9386 15988 9392
rect 15948 8090 15976 9386
rect 16132 9110 16160 11222
rect 16224 9518 16252 12242
rect 16408 12102 16436 12922
rect 16396 12096 16448 12102
rect 16396 12038 16448 12044
rect 16592 11762 16620 13398
rect 16672 12708 16724 12714
rect 16672 12650 16724 12656
rect 16684 12374 16712 12650
rect 16672 12368 16724 12374
rect 16672 12310 16724 12316
rect 16580 11756 16632 11762
rect 16580 11698 16632 11704
rect 16672 9920 16724 9926
rect 16672 9862 16724 9868
rect 16212 9512 16264 9518
rect 16212 9454 16264 9460
rect 16304 9512 16356 9518
rect 16304 9454 16356 9460
rect 16120 9104 16172 9110
rect 16120 9046 16172 9052
rect 16224 8974 16252 9454
rect 16212 8968 16264 8974
rect 16212 8910 16264 8916
rect 16316 8498 16344 9454
rect 16488 9104 16540 9110
rect 16488 9046 16540 9052
rect 16304 8492 16356 8498
rect 16304 8434 16356 8440
rect 15936 8084 15988 8090
rect 15936 8026 15988 8032
rect 15844 8016 15896 8022
rect 15844 7958 15896 7964
rect 15384 7812 15436 7818
rect 15384 7754 15436 7760
rect 15212 6854 15332 6882
rect 14556 6792 14608 6798
rect 14556 6734 14608 6740
rect 15016 6792 15068 6798
rect 15016 6734 15068 6740
rect 14568 6458 14596 6734
rect 14556 6452 14608 6458
rect 14556 6394 14608 6400
rect 14740 6248 14792 6254
rect 14740 6190 14792 6196
rect 14752 4826 14780 6190
rect 14832 5228 14884 5234
rect 14832 5170 14884 5176
rect 14740 4820 14792 4826
rect 14740 4762 14792 4768
rect 12256 4752 12308 4758
rect 12256 4694 12308 4700
rect 13268 4752 13320 4758
rect 13268 4694 13320 4700
rect 14280 4752 14332 4758
rect 14280 4694 14332 4700
rect 12716 4684 12768 4690
rect 12716 4626 12768 4632
rect 11244 4616 11296 4622
rect 11244 4558 11296 4564
rect 11888 4616 11940 4622
rect 11888 4558 11940 4564
rect 10856 4380 11164 4389
rect 10856 4378 10862 4380
rect 10918 4378 10942 4380
rect 10998 4378 11022 4380
rect 11078 4378 11102 4380
rect 11158 4378 11164 4380
rect 10918 4326 10920 4378
rect 11100 4326 11102 4378
rect 10856 4324 10862 4326
rect 10918 4324 10942 4326
rect 10998 4324 11022 4326
rect 11078 4324 11102 4326
rect 11158 4324 11164 4326
rect 10856 4315 11164 4324
rect 11256 4146 11284 4558
rect 12440 4480 12492 4486
rect 12440 4422 12492 4428
rect 12452 4282 12480 4422
rect 12440 4276 12492 4282
rect 12440 4218 12492 4224
rect 11244 4140 11296 4146
rect 11244 4082 11296 4088
rect 11520 4140 11572 4146
rect 11520 4082 11572 4088
rect 11532 3670 11560 4082
rect 11612 4072 11664 4078
rect 11612 4014 11664 4020
rect 11624 3738 11652 4014
rect 12728 3942 12756 4626
rect 12992 4276 13044 4282
rect 12992 4218 13044 4224
rect 12808 4208 12860 4214
rect 12808 4150 12860 4156
rect 12716 3936 12768 3942
rect 12716 3878 12768 3884
rect 12406 3836 12714 3845
rect 12406 3834 12412 3836
rect 12468 3834 12492 3836
rect 12548 3834 12572 3836
rect 12628 3834 12652 3836
rect 12708 3834 12714 3836
rect 12468 3782 12470 3834
rect 12650 3782 12652 3834
rect 12406 3780 12412 3782
rect 12468 3780 12492 3782
rect 12548 3780 12572 3782
rect 12628 3780 12652 3782
rect 12708 3780 12714 3782
rect 12406 3771 12714 3780
rect 11612 3732 11664 3738
rect 11612 3674 11664 3680
rect 11520 3664 11572 3670
rect 11520 3606 11572 3612
rect 12440 3596 12492 3602
rect 12440 3538 12492 3544
rect 11336 3460 11388 3466
rect 11336 3402 11388 3408
rect 10856 3292 11164 3301
rect 10856 3290 10862 3292
rect 10918 3290 10942 3292
rect 10998 3290 11022 3292
rect 11078 3290 11102 3292
rect 11158 3290 11164 3292
rect 10918 3238 10920 3290
rect 11100 3238 11102 3290
rect 10856 3236 10862 3238
rect 10918 3236 10942 3238
rect 10998 3236 11022 3238
rect 11078 3236 11102 3238
rect 11158 3236 11164 3238
rect 10856 3227 11164 3236
rect 11348 3194 11376 3402
rect 11336 3188 11388 3194
rect 11336 3130 11388 3136
rect 12452 3058 12480 3538
rect 12820 3194 12848 4150
rect 12900 4004 12952 4010
rect 12900 3946 12952 3952
rect 12912 3602 12940 3946
rect 12900 3596 12952 3602
rect 12900 3538 12952 3544
rect 12808 3188 12860 3194
rect 12808 3130 12860 3136
rect 12440 3052 12492 3058
rect 12440 2994 12492 3000
rect 13004 2922 13032 4218
rect 13280 4078 13308 4694
rect 13728 4684 13780 4690
rect 13728 4626 13780 4632
rect 13544 4616 13596 4622
rect 13544 4558 13596 4564
rect 13268 4072 13320 4078
rect 13268 4014 13320 4020
rect 13556 2990 13584 4558
rect 13544 2984 13596 2990
rect 13544 2926 13596 2932
rect 12992 2916 13044 2922
rect 12992 2858 13044 2864
rect 11612 2848 11664 2854
rect 11612 2790 11664 2796
rect 12256 2848 12308 2854
rect 12256 2790 12308 2796
rect 12808 2848 12860 2854
rect 12808 2790 12860 2796
rect 10856 2204 11164 2213
rect 10856 2202 10862 2204
rect 10918 2202 10942 2204
rect 10998 2202 11022 2204
rect 11078 2202 11102 2204
rect 11158 2202 11164 2204
rect 10918 2150 10920 2202
rect 11100 2150 11102 2202
rect 10856 2148 10862 2150
rect 10918 2148 10942 2150
rect 10998 2148 11022 2150
rect 11078 2148 11102 2150
rect 11158 2148 11164 2150
rect 10856 2139 11164 2148
rect 11624 2106 11652 2790
rect 12268 2582 12296 2790
rect 12406 2748 12714 2757
rect 12406 2746 12412 2748
rect 12468 2746 12492 2748
rect 12548 2746 12572 2748
rect 12628 2746 12652 2748
rect 12708 2746 12714 2748
rect 12468 2694 12470 2746
rect 12650 2694 12652 2746
rect 12406 2692 12412 2694
rect 12468 2692 12492 2694
rect 12548 2692 12572 2694
rect 12628 2692 12652 2694
rect 12708 2692 12714 2694
rect 12406 2683 12714 2692
rect 12256 2576 12308 2582
rect 12256 2518 12308 2524
rect 9864 2100 9916 2106
rect 9864 2042 9916 2048
rect 10416 2100 10468 2106
rect 10416 2042 10468 2048
rect 10784 2100 10836 2106
rect 10784 2042 10836 2048
rect 11612 2100 11664 2106
rect 11612 2042 11664 2048
rect 9772 1964 9824 1970
rect 9772 1906 9824 1912
rect 9680 1760 9732 1766
rect 9680 1702 9732 1708
rect 9306 1660 9614 1669
rect 9306 1658 9312 1660
rect 9368 1658 9392 1660
rect 9448 1658 9472 1660
rect 9528 1658 9552 1660
rect 9608 1658 9614 1660
rect 9368 1606 9370 1658
rect 9550 1606 9552 1658
rect 9306 1604 9312 1606
rect 9368 1604 9392 1606
rect 9448 1604 9472 1606
rect 9528 1604 9552 1606
rect 9608 1604 9614 1606
rect 9306 1595 9614 1604
rect 9220 1556 9272 1562
rect 9220 1498 9272 1504
rect 9036 1488 9088 1494
rect 9036 1430 9088 1436
rect 9784 1426 9812 1906
rect 10048 1896 10100 1902
rect 10048 1838 10100 1844
rect 10324 1896 10376 1902
rect 10324 1838 10376 1844
rect 10060 1562 10088 1838
rect 10048 1556 10100 1562
rect 10048 1498 10100 1504
rect 10336 1494 10364 1838
rect 10324 1488 10376 1494
rect 10324 1430 10376 1436
rect 10428 1426 10456 2042
rect 12268 1902 12296 2518
rect 12820 2106 12848 2790
rect 12808 2100 12860 2106
rect 12808 2042 12860 2048
rect 12256 1896 12308 1902
rect 12256 1838 12308 1844
rect 12808 1896 12860 1902
rect 13004 1884 13032 2858
rect 12860 1856 13032 1884
rect 12808 1838 12860 1844
rect 11152 1828 11204 1834
rect 11152 1770 11204 1776
rect 11612 1828 11664 1834
rect 11612 1770 11664 1776
rect 11164 1426 11192 1770
rect 5540 1420 5592 1426
rect 5540 1362 5592 1368
rect 5632 1420 5684 1426
rect 5632 1362 5684 1368
rect 7656 1420 7708 1426
rect 7656 1362 7708 1368
rect 9772 1420 9824 1426
rect 9772 1362 9824 1368
rect 10416 1420 10468 1426
rect 10416 1362 10468 1368
rect 11152 1420 11204 1426
rect 11152 1362 11204 1368
rect 11336 1420 11388 1426
rect 11336 1362 11388 1368
rect 5644 1018 5672 1362
rect 11244 1352 11296 1358
rect 11244 1294 11296 1300
rect 7756 1116 8064 1125
rect 7756 1114 7762 1116
rect 7818 1114 7842 1116
rect 7898 1114 7922 1116
rect 7978 1114 8002 1116
rect 8058 1114 8064 1116
rect 7818 1062 7820 1114
rect 8000 1062 8002 1114
rect 7756 1060 7762 1062
rect 7818 1060 7842 1062
rect 7898 1060 7922 1062
rect 7978 1060 8002 1062
rect 8058 1060 8064 1062
rect 7756 1051 8064 1060
rect 10856 1116 11164 1125
rect 10856 1114 10862 1116
rect 10918 1114 10942 1116
rect 10998 1114 11022 1116
rect 11078 1114 11102 1116
rect 11158 1114 11164 1116
rect 10918 1062 10920 1114
rect 11100 1062 11102 1114
rect 10856 1060 10862 1062
rect 10918 1060 10942 1062
rect 10998 1060 11022 1062
rect 11078 1060 11102 1062
rect 11158 1060 11164 1062
rect 10856 1051 11164 1060
rect 5632 1012 5684 1018
rect 5632 954 5684 960
rect 5264 944 5316 950
rect 5264 886 5316 892
rect 11256 814 11284 1294
rect 11348 1018 11376 1362
rect 11428 1216 11480 1222
rect 11428 1158 11480 1164
rect 11336 1012 11388 1018
rect 11336 954 11388 960
rect 11440 950 11468 1158
rect 11428 944 11480 950
rect 11428 886 11480 892
rect 11624 882 11652 1770
rect 11888 1760 11940 1766
rect 11888 1702 11940 1708
rect 11900 1562 11928 1702
rect 12268 1562 12296 1838
rect 12406 1660 12714 1669
rect 12406 1658 12412 1660
rect 12468 1658 12492 1660
rect 12548 1658 12572 1660
rect 12628 1658 12652 1660
rect 12708 1658 12714 1660
rect 12468 1606 12470 1658
rect 12650 1606 12652 1658
rect 12406 1604 12412 1606
rect 12468 1604 12492 1606
rect 12548 1604 12572 1606
rect 12628 1604 12652 1606
rect 12708 1604 12714 1606
rect 12406 1595 12714 1604
rect 11888 1556 11940 1562
rect 11888 1498 11940 1504
rect 12256 1556 12308 1562
rect 12256 1498 12308 1504
rect 12820 1358 12848 1838
rect 13556 1834 13584 2926
rect 13740 2650 13768 4626
rect 14280 4616 14332 4622
rect 14280 4558 14332 4564
rect 13956 4380 14264 4389
rect 13956 4378 13962 4380
rect 14018 4378 14042 4380
rect 14098 4378 14122 4380
rect 14178 4378 14202 4380
rect 14258 4378 14264 4380
rect 14018 4326 14020 4378
rect 14200 4326 14202 4378
rect 13956 4324 13962 4326
rect 14018 4324 14042 4326
rect 14098 4324 14122 4326
rect 14178 4324 14202 4326
rect 14258 4324 14264 4326
rect 13956 4315 14264 4324
rect 14292 4282 14320 4558
rect 14464 4548 14516 4554
rect 14464 4490 14516 4496
rect 14280 4276 14332 4282
rect 14280 4218 14332 4224
rect 14476 4214 14504 4490
rect 14752 4298 14780 4762
rect 14660 4282 14780 4298
rect 14660 4276 14792 4282
rect 14660 4270 14740 4276
rect 14464 4208 14516 4214
rect 14464 4150 14516 4156
rect 13956 3292 14264 3301
rect 13956 3290 13962 3292
rect 14018 3290 14042 3292
rect 14098 3290 14122 3292
rect 14178 3290 14202 3292
rect 14258 3290 14264 3292
rect 14018 3238 14020 3290
rect 14200 3238 14202 3290
rect 13956 3236 13962 3238
rect 14018 3236 14042 3238
rect 14098 3236 14122 3238
rect 14178 3236 14202 3238
rect 14258 3236 14264 3238
rect 13956 3227 14264 3236
rect 14660 3194 14688 4270
rect 14740 4218 14792 4224
rect 14740 4140 14792 4146
rect 14740 4082 14792 4088
rect 14752 3738 14780 4082
rect 14740 3732 14792 3738
rect 14740 3674 14792 3680
rect 14188 3188 14240 3194
rect 14188 3130 14240 3136
rect 14648 3188 14700 3194
rect 14648 3130 14700 3136
rect 13820 2916 13872 2922
rect 13820 2858 13872 2864
rect 13728 2644 13780 2650
rect 13728 2586 13780 2592
rect 13740 1902 13768 2586
rect 13832 2582 13860 2858
rect 14200 2582 14228 3130
rect 14660 3074 14688 3130
rect 14660 3046 14780 3074
rect 14648 2984 14700 2990
rect 14648 2926 14700 2932
rect 13820 2576 13872 2582
rect 13820 2518 13872 2524
rect 14188 2576 14240 2582
rect 14188 2518 14240 2524
rect 14372 2440 14424 2446
rect 14372 2382 14424 2388
rect 13956 2204 14264 2213
rect 13956 2202 13962 2204
rect 14018 2202 14042 2204
rect 14098 2202 14122 2204
rect 14178 2202 14202 2204
rect 14258 2202 14264 2204
rect 14018 2150 14020 2202
rect 14200 2150 14202 2202
rect 13956 2148 13962 2150
rect 14018 2148 14042 2150
rect 14098 2148 14122 2150
rect 14178 2148 14202 2150
rect 14258 2148 14264 2150
rect 13956 2139 14264 2148
rect 14384 1970 14412 2382
rect 14372 1964 14424 1970
rect 14372 1906 14424 1912
rect 13728 1896 13780 1902
rect 13728 1838 13780 1844
rect 13544 1828 13596 1834
rect 13544 1770 13596 1776
rect 13556 1426 13584 1770
rect 13740 1494 13768 1838
rect 14096 1760 14148 1766
rect 14096 1702 14148 1708
rect 13728 1488 13780 1494
rect 13728 1430 13780 1436
rect 13544 1420 13596 1426
rect 13544 1362 13596 1368
rect 12808 1352 12860 1358
rect 12808 1294 12860 1300
rect 13820 1352 13872 1358
rect 13820 1294 13872 1300
rect 13832 950 13860 1294
rect 14108 1290 14136 1702
rect 14660 1426 14688 2926
rect 14752 2774 14780 3046
rect 14844 2990 14872 5170
rect 15028 4826 15056 6734
rect 15016 4820 15068 4826
rect 15016 4762 15068 4768
rect 14924 3732 14976 3738
rect 14924 3674 14976 3680
rect 14936 2990 14964 3674
rect 15028 3670 15056 4762
rect 15016 3664 15068 3670
rect 15016 3606 15068 3612
rect 14832 2984 14884 2990
rect 14832 2926 14884 2932
rect 14924 2984 14976 2990
rect 14924 2926 14976 2932
rect 14936 2774 14964 2926
rect 15028 2922 15056 3606
rect 15212 3126 15240 6854
rect 15396 6798 15424 7754
rect 15856 7546 15884 7958
rect 15844 7540 15896 7546
rect 15844 7482 15896 7488
rect 15844 7404 15896 7410
rect 15844 7346 15896 7352
rect 15856 7206 15884 7346
rect 15936 7336 15988 7342
rect 15936 7278 15988 7284
rect 15844 7200 15896 7206
rect 15844 7142 15896 7148
rect 15506 7100 15814 7109
rect 15506 7098 15512 7100
rect 15568 7098 15592 7100
rect 15648 7098 15672 7100
rect 15728 7098 15752 7100
rect 15808 7098 15814 7100
rect 15568 7046 15570 7098
rect 15750 7046 15752 7098
rect 15506 7044 15512 7046
rect 15568 7044 15592 7046
rect 15648 7044 15672 7046
rect 15728 7044 15752 7046
rect 15808 7044 15814 7046
rect 15506 7035 15814 7044
rect 15948 6934 15976 7278
rect 16028 7200 16080 7206
rect 16028 7142 16080 7148
rect 15936 6928 15988 6934
rect 15936 6870 15988 6876
rect 16040 6866 16068 7142
rect 16028 6860 16080 6866
rect 16028 6802 16080 6808
rect 15384 6792 15436 6798
rect 15384 6734 15436 6740
rect 15292 6656 15344 6662
rect 15292 6598 15344 6604
rect 15304 6390 15332 6598
rect 15292 6384 15344 6390
rect 15292 6326 15344 6332
rect 15396 4554 15424 6734
rect 16316 6338 16344 8434
rect 16500 8294 16528 9046
rect 16580 8424 16632 8430
rect 16580 8366 16632 8372
rect 16488 8288 16540 8294
rect 16488 8230 16540 8236
rect 16500 7274 16528 8230
rect 16592 8090 16620 8366
rect 16580 8084 16632 8090
rect 16580 8026 16632 8032
rect 16580 7948 16632 7954
rect 16580 7890 16632 7896
rect 16592 7546 16620 7890
rect 16684 7886 16712 9862
rect 16868 9518 16896 14368
rect 16960 12986 16988 14418
rect 17500 14340 17552 14346
rect 17500 14282 17552 14288
rect 17056 14172 17364 14181
rect 17056 14170 17062 14172
rect 17118 14170 17142 14172
rect 17198 14170 17222 14172
rect 17278 14170 17302 14172
rect 17358 14170 17364 14172
rect 17118 14118 17120 14170
rect 17300 14118 17302 14170
rect 17056 14116 17062 14118
rect 17118 14116 17142 14118
rect 17198 14116 17222 14118
rect 17278 14116 17302 14118
rect 17358 14116 17364 14118
rect 17056 14107 17364 14116
rect 17408 13184 17460 13190
rect 17408 13126 17460 13132
rect 17056 13084 17364 13093
rect 17056 13082 17062 13084
rect 17118 13082 17142 13084
rect 17198 13082 17222 13084
rect 17278 13082 17302 13084
rect 17358 13082 17364 13084
rect 17118 13030 17120 13082
rect 17300 13030 17302 13082
rect 17056 13028 17062 13030
rect 17118 13028 17142 13030
rect 17198 13028 17222 13030
rect 17278 13028 17302 13030
rect 17358 13028 17364 13030
rect 17056 13019 17364 13028
rect 16948 12980 17000 12986
rect 16948 12922 17000 12928
rect 16960 12374 16988 12922
rect 17420 12850 17448 13126
rect 17408 12844 17460 12850
rect 17408 12786 17460 12792
rect 17512 12782 17540 14282
rect 17604 13870 17632 14894
rect 17592 13864 17644 13870
rect 17592 13806 17644 13812
rect 17684 13388 17736 13394
rect 17684 13330 17736 13336
rect 17592 13320 17644 13326
rect 17592 13262 17644 13268
rect 17500 12776 17552 12782
rect 17500 12718 17552 12724
rect 17604 12374 17632 13262
rect 16948 12368 17000 12374
rect 16948 12310 17000 12316
rect 17592 12368 17644 12374
rect 17592 12310 17644 12316
rect 16960 11626 16988 12310
rect 17056 11996 17364 12005
rect 17056 11994 17062 11996
rect 17118 11994 17142 11996
rect 17198 11994 17222 11996
rect 17278 11994 17302 11996
rect 17358 11994 17364 11996
rect 17118 11942 17120 11994
rect 17300 11942 17302 11994
rect 17056 11940 17062 11942
rect 17118 11940 17142 11942
rect 17198 11940 17222 11942
rect 17278 11940 17302 11942
rect 17358 11940 17364 11942
rect 17056 11931 17364 11940
rect 16948 11620 17000 11626
rect 16948 11562 17000 11568
rect 16960 11218 16988 11562
rect 16948 11212 17000 11218
rect 16948 11154 17000 11160
rect 16960 10810 16988 11154
rect 17500 11076 17552 11082
rect 17500 11018 17552 11024
rect 17408 11008 17460 11014
rect 17408 10950 17460 10956
rect 17056 10908 17364 10917
rect 17056 10906 17062 10908
rect 17118 10906 17142 10908
rect 17198 10906 17222 10908
rect 17278 10906 17302 10908
rect 17358 10906 17364 10908
rect 17118 10854 17120 10906
rect 17300 10854 17302 10906
rect 17056 10852 17062 10854
rect 17118 10852 17142 10854
rect 17198 10852 17222 10854
rect 17278 10852 17302 10854
rect 17358 10852 17364 10854
rect 17056 10843 17364 10852
rect 16948 10804 17000 10810
rect 16948 10746 17000 10752
rect 17420 10130 17448 10950
rect 17512 10198 17540 11018
rect 17500 10192 17552 10198
rect 17500 10134 17552 10140
rect 17408 10124 17460 10130
rect 17408 10066 17460 10072
rect 17056 9820 17364 9829
rect 17056 9818 17062 9820
rect 17118 9818 17142 9820
rect 17198 9818 17222 9820
rect 17278 9818 17302 9820
rect 17358 9818 17364 9820
rect 17118 9766 17120 9818
rect 17300 9766 17302 9818
rect 17056 9764 17062 9766
rect 17118 9764 17142 9766
rect 17198 9764 17222 9766
rect 17278 9764 17302 9766
rect 17358 9764 17364 9766
rect 17056 9755 17364 9764
rect 16856 9512 16908 9518
rect 16856 9454 16908 9460
rect 16672 7880 16724 7886
rect 16672 7822 16724 7828
rect 16580 7540 16632 7546
rect 16580 7482 16632 7488
rect 16488 7268 16540 7274
rect 16488 7210 16540 7216
rect 16500 6882 16528 7210
rect 16500 6854 16712 6882
rect 16224 6322 16344 6338
rect 16212 6316 16344 6322
rect 16264 6310 16344 6316
rect 16212 6258 16264 6264
rect 15506 6012 15814 6021
rect 15506 6010 15512 6012
rect 15568 6010 15592 6012
rect 15648 6010 15672 6012
rect 15728 6010 15752 6012
rect 15808 6010 15814 6012
rect 15568 5958 15570 6010
rect 15750 5958 15752 6010
rect 15506 5956 15512 5958
rect 15568 5956 15592 5958
rect 15648 5956 15672 5958
rect 15728 5956 15752 5958
rect 15808 5956 15814 5958
rect 15506 5947 15814 5956
rect 16224 5914 16252 6258
rect 16304 6248 16356 6254
rect 16304 6190 16356 6196
rect 16212 5908 16264 5914
rect 16212 5850 16264 5856
rect 16224 5234 16252 5850
rect 16212 5228 16264 5234
rect 16212 5170 16264 5176
rect 16212 5092 16264 5098
rect 16212 5034 16264 5040
rect 15506 4924 15814 4933
rect 15506 4922 15512 4924
rect 15568 4922 15592 4924
rect 15648 4922 15672 4924
rect 15728 4922 15752 4924
rect 15808 4922 15814 4924
rect 15568 4870 15570 4922
rect 15750 4870 15752 4922
rect 15506 4868 15512 4870
rect 15568 4868 15592 4870
rect 15648 4868 15672 4870
rect 15728 4868 15752 4870
rect 15808 4868 15814 4870
rect 15506 4859 15814 4868
rect 15476 4820 15528 4826
rect 15476 4762 15528 4768
rect 15384 4548 15436 4554
rect 15384 4490 15436 4496
rect 15292 4140 15344 4146
rect 15292 4082 15344 4088
rect 15304 3738 15332 4082
rect 15488 4078 15516 4762
rect 15476 4072 15528 4078
rect 15476 4014 15528 4020
rect 15506 3836 15814 3845
rect 15506 3834 15512 3836
rect 15568 3834 15592 3836
rect 15648 3834 15672 3836
rect 15728 3834 15752 3836
rect 15808 3834 15814 3836
rect 15568 3782 15570 3834
rect 15750 3782 15752 3834
rect 15506 3780 15512 3782
rect 15568 3780 15592 3782
rect 15648 3780 15672 3782
rect 15728 3780 15752 3782
rect 15808 3780 15814 3782
rect 15506 3771 15814 3780
rect 15292 3732 15344 3738
rect 15292 3674 15344 3680
rect 15384 3596 15436 3602
rect 15384 3538 15436 3544
rect 15200 3120 15252 3126
rect 15200 3062 15252 3068
rect 15016 2916 15068 2922
rect 15016 2858 15068 2864
rect 14752 2746 14872 2774
rect 14936 2746 15056 2774
rect 14844 2106 14872 2746
rect 15028 2446 15056 2746
rect 15396 2650 15424 3538
rect 15844 2916 15896 2922
rect 15844 2858 15896 2864
rect 15506 2748 15814 2757
rect 15506 2746 15512 2748
rect 15568 2746 15592 2748
rect 15648 2746 15672 2748
rect 15728 2746 15752 2748
rect 15808 2746 15814 2748
rect 15568 2694 15570 2746
rect 15750 2694 15752 2746
rect 15506 2692 15512 2694
rect 15568 2692 15592 2694
rect 15648 2692 15672 2694
rect 15728 2692 15752 2694
rect 15808 2692 15814 2694
rect 15506 2683 15814 2692
rect 15384 2644 15436 2650
rect 15384 2586 15436 2592
rect 15016 2440 15068 2446
rect 15016 2382 15068 2388
rect 14832 2100 14884 2106
rect 14832 2042 14884 2048
rect 14844 1902 14872 2042
rect 15856 2038 15884 2858
rect 16224 2106 16252 5034
rect 16316 3738 16344 6190
rect 16684 6186 16712 6854
rect 16868 6458 16896 9454
rect 17056 8732 17364 8741
rect 17056 8730 17062 8732
rect 17118 8730 17142 8732
rect 17198 8730 17222 8732
rect 17278 8730 17302 8732
rect 17358 8730 17364 8732
rect 17118 8678 17120 8730
rect 17300 8678 17302 8730
rect 17056 8676 17062 8678
rect 17118 8676 17142 8678
rect 17198 8676 17222 8678
rect 17278 8676 17302 8678
rect 17358 8676 17364 8678
rect 17056 8667 17364 8676
rect 17696 8634 17724 13330
rect 17880 12306 17908 15574
rect 17960 14816 18012 14822
rect 17960 14758 18012 14764
rect 17972 14550 18000 14758
rect 17960 14544 18012 14550
rect 17960 14486 18012 14492
rect 17960 14408 18012 14414
rect 17960 14350 18012 14356
rect 17972 14074 18000 14350
rect 17960 14068 18012 14074
rect 17960 14010 18012 14016
rect 18052 14000 18104 14006
rect 18052 13942 18104 13948
rect 17868 12300 17920 12306
rect 17868 12242 17920 12248
rect 17776 11552 17828 11558
rect 17776 11494 17828 11500
rect 17788 11218 17816 11494
rect 17776 11212 17828 11218
rect 17776 11154 17828 11160
rect 17960 10124 18012 10130
rect 17960 10066 18012 10072
rect 17972 9654 18000 10066
rect 17960 9648 18012 9654
rect 17960 9590 18012 9596
rect 17684 8628 17736 8634
rect 17684 8570 17736 8576
rect 17696 8090 17724 8570
rect 17684 8084 17736 8090
rect 17684 8026 17736 8032
rect 17316 7880 17368 7886
rect 17368 7828 17448 7834
rect 17316 7822 17448 7828
rect 17328 7806 17448 7822
rect 17056 7644 17364 7653
rect 17056 7642 17062 7644
rect 17118 7642 17142 7644
rect 17198 7642 17222 7644
rect 17278 7642 17302 7644
rect 17358 7642 17364 7644
rect 17118 7590 17120 7642
rect 17300 7590 17302 7642
rect 17056 7588 17062 7590
rect 17118 7588 17142 7590
rect 17198 7588 17222 7590
rect 17278 7588 17302 7590
rect 17358 7588 17364 7590
rect 17056 7579 17364 7588
rect 17420 7342 17448 7806
rect 17696 7342 17724 8026
rect 17776 7880 17828 7886
rect 17776 7822 17828 7828
rect 17408 7336 17460 7342
rect 17408 7278 17460 7284
rect 17684 7336 17736 7342
rect 17684 7278 17736 7284
rect 17056 6556 17364 6565
rect 17056 6554 17062 6556
rect 17118 6554 17142 6556
rect 17198 6554 17222 6556
rect 17278 6554 17302 6556
rect 17358 6554 17364 6556
rect 17118 6502 17120 6554
rect 17300 6502 17302 6554
rect 17056 6500 17062 6502
rect 17118 6500 17142 6502
rect 17198 6500 17222 6502
rect 17278 6500 17302 6502
rect 17358 6500 17364 6502
rect 17056 6491 17364 6500
rect 16856 6452 16908 6458
rect 16856 6394 16908 6400
rect 16672 6180 16724 6186
rect 16672 6122 16724 6128
rect 16684 5846 16712 6122
rect 16672 5840 16724 5846
rect 16672 5782 16724 5788
rect 16684 5098 16712 5782
rect 16868 5778 16896 6394
rect 17420 5914 17448 7278
rect 17788 7274 17816 7822
rect 17776 7268 17828 7274
rect 17776 7210 17828 7216
rect 17788 6186 17816 7210
rect 17776 6180 17828 6186
rect 17776 6122 17828 6128
rect 17408 5908 17460 5914
rect 17408 5850 17460 5856
rect 16856 5772 16908 5778
rect 16856 5714 16908 5720
rect 17500 5772 17552 5778
rect 17500 5714 17552 5720
rect 16672 5092 16724 5098
rect 16672 5034 16724 5040
rect 16868 4146 16896 5714
rect 16948 5704 17000 5710
rect 16948 5646 17000 5652
rect 16960 4282 16988 5646
rect 17056 5468 17364 5477
rect 17056 5466 17062 5468
rect 17118 5466 17142 5468
rect 17198 5466 17222 5468
rect 17278 5466 17302 5468
rect 17358 5466 17364 5468
rect 17118 5414 17120 5466
rect 17300 5414 17302 5466
rect 17056 5412 17062 5414
rect 17118 5412 17142 5414
rect 17198 5412 17222 5414
rect 17278 5412 17302 5414
rect 17358 5412 17364 5414
rect 17056 5403 17364 5412
rect 17512 5030 17540 5714
rect 17592 5636 17644 5642
rect 17592 5578 17644 5584
rect 17500 5024 17552 5030
rect 17420 4984 17500 5012
rect 17056 4380 17364 4389
rect 17056 4378 17062 4380
rect 17118 4378 17142 4380
rect 17198 4378 17222 4380
rect 17278 4378 17302 4380
rect 17358 4378 17364 4380
rect 17118 4326 17120 4378
rect 17300 4326 17302 4378
rect 17056 4324 17062 4326
rect 17118 4324 17142 4326
rect 17198 4324 17222 4326
rect 17278 4324 17302 4326
rect 17358 4324 17364 4326
rect 17056 4315 17364 4324
rect 16948 4276 17000 4282
rect 16948 4218 17000 4224
rect 17420 4146 17448 4984
rect 17500 4966 17552 4972
rect 17604 4214 17632 5578
rect 17592 4208 17644 4214
rect 17592 4150 17644 4156
rect 16856 4140 16908 4146
rect 16856 4082 16908 4088
rect 17408 4140 17460 4146
rect 17408 4082 17460 4088
rect 16868 3754 16896 4082
rect 17316 4004 17368 4010
rect 17316 3946 17368 3952
rect 16304 3732 16356 3738
rect 16868 3726 16988 3754
rect 16304 3674 16356 3680
rect 16580 3664 16632 3670
rect 16580 3606 16632 3612
rect 16592 3398 16620 3606
rect 16960 3602 16988 3726
rect 16856 3596 16908 3602
rect 16856 3538 16908 3544
rect 16948 3596 17000 3602
rect 16948 3538 17000 3544
rect 16580 3392 16632 3398
rect 16580 3334 16632 3340
rect 16488 2440 16540 2446
rect 16488 2382 16540 2388
rect 16212 2100 16264 2106
rect 16212 2042 16264 2048
rect 15844 2032 15896 2038
rect 15844 1974 15896 1980
rect 16500 1970 16528 2382
rect 16488 1964 16540 1970
rect 16488 1906 16540 1912
rect 14832 1896 14884 1902
rect 14832 1838 14884 1844
rect 15506 1660 15814 1669
rect 15506 1658 15512 1660
rect 15568 1658 15592 1660
rect 15648 1658 15672 1660
rect 15728 1658 15752 1660
rect 15808 1658 15814 1660
rect 15568 1606 15570 1658
rect 15750 1606 15752 1658
rect 15506 1604 15512 1606
rect 15568 1604 15592 1606
rect 15648 1604 15672 1606
rect 15728 1604 15752 1606
rect 15808 1604 15814 1606
rect 15506 1595 15814 1604
rect 14648 1420 14700 1426
rect 14648 1362 14700 1368
rect 16592 1358 16620 3334
rect 16764 2508 16816 2514
rect 16764 2450 16816 2456
rect 16776 1766 16804 2450
rect 16764 1760 16816 1766
rect 16764 1702 16816 1708
rect 16776 1426 16804 1702
rect 16868 1562 16896 3538
rect 17328 3398 17356 3946
rect 17420 3534 17448 4082
rect 17604 3602 17632 4150
rect 17788 4146 17816 6122
rect 17776 4140 17828 4146
rect 17776 4082 17828 4088
rect 17684 4072 17736 4078
rect 17684 4014 17736 4020
rect 17696 3738 17724 4014
rect 18064 3738 18092 13942
rect 18236 13932 18288 13938
rect 18236 13874 18288 13880
rect 18144 12912 18196 12918
rect 18144 12854 18196 12860
rect 18156 9178 18184 12854
rect 18248 12170 18276 13874
rect 18328 12708 18380 12714
rect 18328 12650 18380 12656
rect 18236 12164 18288 12170
rect 18236 12106 18288 12112
rect 18144 9172 18196 9178
rect 18144 9114 18196 9120
rect 17684 3732 17736 3738
rect 17684 3674 17736 3680
rect 18052 3732 18104 3738
rect 18052 3674 18104 3680
rect 17592 3596 17644 3602
rect 17592 3538 17644 3544
rect 17408 3528 17460 3534
rect 17408 3470 17460 3476
rect 17316 3392 17368 3398
rect 17316 3334 17368 3340
rect 17056 3292 17364 3301
rect 17056 3290 17062 3292
rect 17118 3290 17142 3292
rect 17198 3290 17222 3292
rect 17278 3290 17302 3292
rect 17358 3290 17364 3292
rect 17118 3238 17120 3290
rect 17300 3238 17302 3290
rect 17056 3236 17062 3238
rect 17118 3236 17142 3238
rect 17198 3236 17222 3238
rect 17278 3236 17302 3238
rect 17358 3236 17364 3238
rect 17056 3227 17364 3236
rect 17420 2530 17448 3470
rect 17604 2582 17632 3538
rect 18340 2582 18368 12650
rect 18524 12442 18552 19200
rect 18606 17980 18914 17989
rect 18606 17978 18612 17980
rect 18668 17978 18692 17980
rect 18748 17978 18772 17980
rect 18828 17978 18852 17980
rect 18908 17978 18914 17980
rect 18668 17926 18670 17978
rect 18850 17926 18852 17978
rect 18606 17924 18612 17926
rect 18668 17924 18692 17926
rect 18748 17924 18772 17926
rect 18828 17924 18852 17926
rect 18908 17924 18914 17926
rect 18606 17915 18914 17924
rect 18606 16892 18914 16901
rect 18606 16890 18612 16892
rect 18668 16890 18692 16892
rect 18748 16890 18772 16892
rect 18828 16890 18852 16892
rect 18908 16890 18914 16892
rect 18668 16838 18670 16890
rect 18850 16838 18852 16890
rect 18606 16836 18612 16838
rect 18668 16836 18692 16838
rect 18748 16836 18772 16838
rect 18828 16836 18852 16838
rect 18908 16836 18914 16838
rect 18606 16827 18914 16836
rect 18606 15804 18914 15813
rect 18606 15802 18612 15804
rect 18668 15802 18692 15804
rect 18748 15802 18772 15804
rect 18828 15802 18852 15804
rect 18908 15802 18914 15804
rect 18668 15750 18670 15802
rect 18850 15750 18852 15802
rect 18606 15748 18612 15750
rect 18668 15748 18692 15750
rect 18748 15748 18772 15750
rect 18828 15748 18852 15750
rect 18908 15748 18914 15750
rect 18606 15739 18914 15748
rect 19064 15564 19116 15570
rect 19064 15506 19116 15512
rect 18606 14716 18914 14725
rect 18606 14714 18612 14716
rect 18668 14714 18692 14716
rect 18748 14714 18772 14716
rect 18828 14714 18852 14716
rect 18908 14714 18914 14716
rect 18668 14662 18670 14714
rect 18850 14662 18852 14714
rect 18606 14660 18612 14662
rect 18668 14660 18692 14662
rect 18748 14660 18772 14662
rect 18828 14660 18852 14662
rect 18908 14660 18914 14662
rect 18606 14651 18914 14660
rect 19076 13705 19104 15506
rect 19062 13696 19118 13705
rect 18606 13628 18914 13637
rect 19062 13631 19118 13640
rect 18606 13626 18612 13628
rect 18668 13626 18692 13628
rect 18748 13626 18772 13628
rect 18828 13626 18852 13628
rect 18908 13626 18914 13628
rect 18668 13574 18670 13626
rect 18850 13574 18852 13626
rect 18606 13572 18612 13574
rect 18668 13572 18692 13574
rect 18748 13572 18772 13574
rect 18828 13572 18852 13574
rect 18908 13572 18914 13574
rect 18606 13563 18914 13572
rect 18606 12540 18914 12549
rect 18606 12538 18612 12540
rect 18668 12538 18692 12540
rect 18748 12538 18772 12540
rect 18828 12538 18852 12540
rect 18908 12538 18914 12540
rect 18668 12486 18670 12538
rect 18850 12486 18852 12538
rect 18606 12484 18612 12486
rect 18668 12484 18692 12486
rect 18748 12484 18772 12486
rect 18828 12484 18852 12486
rect 18908 12484 18914 12486
rect 18606 12475 18914 12484
rect 18512 12436 18564 12442
rect 18512 12378 18564 12384
rect 18420 12300 18472 12306
rect 18420 12242 18472 12248
rect 18432 11558 18460 12242
rect 18420 11552 18472 11558
rect 18420 11494 18472 11500
rect 18432 11257 18460 11494
rect 18606 11452 18914 11461
rect 18606 11450 18612 11452
rect 18668 11450 18692 11452
rect 18748 11450 18772 11452
rect 18828 11450 18852 11452
rect 18908 11450 18914 11452
rect 18668 11398 18670 11450
rect 18850 11398 18852 11450
rect 18606 11396 18612 11398
rect 18668 11396 18692 11398
rect 18748 11396 18772 11398
rect 18828 11396 18852 11398
rect 18908 11396 18914 11398
rect 18606 11387 18914 11396
rect 18418 11248 18474 11257
rect 18418 11183 18474 11192
rect 18606 10364 18914 10373
rect 18606 10362 18612 10364
rect 18668 10362 18692 10364
rect 18748 10362 18772 10364
rect 18828 10362 18852 10364
rect 18908 10362 18914 10364
rect 18668 10310 18670 10362
rect 18850 10310 18852 10362
rect 18606 10308 18612 10310
rect 18668 10308 18692 10310
rect 18748 10308 18772 10310
rect 18828 10308 18852 10310
rect 18908 10308 18914 10310
rect 18606 10299 18914 10308
rect 18606 9276 18914 9285
rect 18606 9274 18612 9276
rect 18668 9274 18692 9276
rect 18748 9274 18772 9276
rect 18828 9274 18852 9276
rect 18908 9274 18914 9276
rect 18668 9222 18670 9274
rect 18850 9222 18852 9274
rect 18606 9220 18612 9222
rect 18668 9220 18692 9222
rect 18748 9220 18772 9222
rect 18828 9220 18852 9222
rect 18908 9220 18914 9222
rect 18606 9211 18914 9220
rect 18420 9036 18472 9042
rect 18420 8978 18472 8984
rect 18432 8809 18460 8978
rect 18418 8800 18474 8809
rect 18418 8735 18474 8744
rect 18606 8188 18914 8197
rect 18606 8186 18612 8188
rect 18668 8186 18692 8188
rect 18748 8186 18772 8188
rect 18828 8186 18852 8188
rect 18908 8186 18914 8188
rect 18668 8134 18670 8186
rect 18850 8134 18852 8186
rect 18606 8132 18612 8134
rect 18668 8132 18692 8134
rect 18748 8132 18772 8134
rect 18828 8132 18852 8134
rect 18908 8132 18914 8134
rect 18606 8123 18914 8132
rect 18606 7100 18914 7109
rect 18606 7098 18612 7100
rect 18668 7098 18692 7100
rect 18748 7098 18772 7100
rect 18828 7098 18852 7100
rect 18908 7098 18914 7100
rect 18668 7046 18670 7098
rect 18850 7046 18852 7098
rect 18606 7044 18612 7046
rect 18668 7044 18692 7046
rect 18748 7044 18772 7046
rect 18828 7044 18852 7046
rect 18908 7044 18914 7046
rect 18606 7035 18914 7044
rect 18420 6860 18472 6866
rect 18420 6802 18472 6808
rect 18432 6361 18460 6802
rect 18418 6352 18474 6361
rect 18418 6287 18474 6296
rect 18606 6012 18914 6021
rect 18606 6010 18612 6012
rect 18668 6010 18692 6012
rect 18748 6010 18772 6012
rect 18828 6010 18852 6012
rect 18908 6010 18914 6012
rect 18668 5958 18670 6010
rect 18850 5958 18852 6010
rect 18606 5956 18612 5958
rect 18668 5956 18692 5958
rect 18748 5956 18772 5958
rect 18828 5956 18852 5958
rect 18908 5956 18914 5958
rect 18606 5947 18914 5956
rect 18606 4924 18914 4933
rect 18606 4922 18612 4924
rect 18668 4922 18692 4924
rect 18748 4922 18772 4924
rect 18828 4922 18852 4924
rect 18908 4922 18914 4924
rect 18668 4870 18670 4922
rect 18850 4870 18852 4922
rect 18606 4868 18612 4870
rect 18668 4868 18692 4870
rect 18748 4868 18772 4870
rect 18828 4868 18852 4870
rect 18908 4868 18914 4870
rect 18606 4859 18914 4868
rect 19062 3904 19118 3913
rect 18606 3836 18914 3845
rect 19062 3839 19118 3848
rect 18606 3834 18612 3836
rect 18668 3834 18692 3836
rect 18748 3834 18772 3836
rect 18828 3834 18852 3836
rect 18908 3834 18914 3836
rect 18668 3782 18670 3834
rect 18850 3782 18852 3834
rect 18606 3780 18612 3782
rect 18668 3780 18692 3782
rect 18748 3780 18772 3782
rect 18828 3780 18852 3782
rect 18908 3780 18914 3782
rect 18606 3771 18914 3780
rect 19076 3602 19104 3839
rect 19064 3596 19116 3602
rect 19064 3538 19116 3544
rect 18606 2748 18914 2757
rect 18606 2746 18612 2748
rect 18668 2746 18692 2748
rect 18748 2746 18772 2748
rect 18828 2746 18852 2748
rect 18908 2746 18914 2748
rect 18668 2694 18670 2746
rect 18850 2694 18852 2746
rect 18606 2692 18612 2694
rect 18668 2692 18692 2694
rect 18748 2692 18772 2694
rect 18828 2692 18852 2694
rect 18908 2692 18914 2694
rect 18606 2683 18914 2692
rect 17328 2514 17448 2530
rect 17592 2576 17644 2582
rect 17592 2518 17644 2524
rect 18328 2576 18380 2582
rect 18328 2518 18380 2524
rect 17316 2508 17448 2514
rect 17368 2502 17448 2508
rect 17500 2508 17552 2514
rect 17316 2450 17368 2456
rect 17500 2450 17552 2456
rect 17960 2508 18012 2514
rect 17960 2450 18012 2456
rect 17408 2304 17460 2310
rect 17408 2246 17460 2252
rect 17056 2204 17364 2213
rect 17056 2202 17062 2204
rect 17118 2202 17142 2204
rect 17198 2202 17222 2204
rect 17278 2202 17302 2204
rect 17358 2202 17364 2204
rect 17118 2150 17120 2202
rect 17300 2150 17302 2202
rect 17056 2148 17062 2150
rect 17118 2148 17142 2150
rect 17198 2148 17222 2150
rect 17278 2148 17302 2150
rect 17358 2148 17364 2150
rect 17056 2139 17364 2148
rect 17420 1970 17448 2246
rect 17408 1964 17460 1970
rect 17408 1906 17460 1912
rect 17224 1896 17276 1902
rect 17224 1838 17276 1844
rect 16856 1556 16908 1562
rect 16856 1498 16908 1504
rect 17236 1494 17264 1838
rect 17316 1760 17368 1766
rect 17316 1702 17368 1708
rect 17224 1488 17276 1494
rect 17224 1430 17276 1436
rect 16764 1420 16816 1426
rect 16764 1362 16816 1368
rect 16580 1352 16632 1358
rect 16580 1294 16632 1300
rect 17328 1290 17356 1702
rect 17420 1290 17448 1906
rect 17512 1562 17540 2450
rect 17500 1556 17552 1562
rect 17500 1498 17552 1504
rect 17592 1488 17644 1494
rect 17592 1430 17644 1436
rect 14096 1284 14148 1290
rect 14096 1226 14148 1232
rect 17316 1284 17368 1290
rect 17316 1226 17368 1232
rect 17408 1284 17460 1290
rect 17408 1226 17460 1232
rect 13956 1116 14264 1125
rect 13956 1114 13962 1116
rect 14018 1114 14042 1116
rect 14098 1114 14122 1116
rect 14178 1114 14202 1116
rect 14258 1114 14264 1116
rect 14018 1062 14020 1114
rect 14200 1062 14202 1114
rect 13956 1060 13962 1062
rect 14018 1060 14042 1062
rect 14098 1060 14122 1062
rect 14178 1060 14202 1062
rect 14258 1060 14264 1062
rect 13956 1051 14264 1060
rect 17056 1116 17364 1125
rect 17056 1114 17062 1116
rect 17118 1114 17142 1116
rect 17198 1114 17222 1116
rect 17278 1114 17302 1116
rect 17358 1114 17364 1116
rect 17118 1062 17120 1114
rect 17300 1062 17302 1114
rect 17056 1060 17062 1062
rect 17118 1060 17142 1062
rect 17198 1060 17222 1062
rect 17278 1060 17302 1062
rect 17358 1060 17364 1062
rect 17056 1051 17364 1060
rect 17604 1018 17632 1430
rect 17972 1018 18000 2450
rect 18606 1660 18914 1669
rect 18606 1658 18612 1660
rect 18668 1658 18692 1660
rect 18748 1658 18772 1660
rect 18828 1658 18852 1660
rect 18908 1658 18914 1660
rect 18668 1606 18670 1658
rect 18850 1606 18852 1658
rect 18606 1604 18612 1606
rect 18668 1604 18692 1606
rect 18748 1604 18772 1606
rect 18828 1604 18852 1606
rect 18908 1604 18914 1606
rect 18606 1595 18914 1604
rect 18418 1456 18474 1465
rect 18418 1391 18474 1400
rect 18432 1018 18460 1391
rect 17592 1012 17644 1018
rect 17592 954 17644 960
rect 17960 1012 18012 1018
rect 17960 954 18012 960
rect 18420 1012 18472 1018
rect 18420 954 18472 960
rect 13820 944 13872 950
rect 13820 886 13872 892
rect 11612 876 11664 882
rect 11612 818 11664 824
rect 5172 808 5224 814
rect 5172 750 5224 756
rect 11244 808 11296 814
rect 11244 750 11296 756
rect 3106 572 3414 581
rect 3106 570 3112 572
rect 3168 570 3192 572
rect 3248 570 3272 572
rect 3328 570 3352 572
rect 3408 570 3414 572
rect 3168 518 3170 570
rect 3350 518 3352 570
rect 3106 516 3112 518
rect 3168 516 3192 518
rect 3248 516 3272 518
rect 3328 516 3352 518
rect 3408 516 3414 518
rect 3106 507 3414 516
rect 6206 572 6514 581
rect 6206 570 6212 572
rect 6268 570 6292 572
rect 6348 570 6372 572
rect 6428 570 6452 572
rect 6508 570 6514 572
rect 6268 518 6270 570
rect 6450 518 6452 570
rect 6206 516 6212 518
rect 6268 516 6292 518
rect 6348 516 6372 518
rect 6428 516 6452 518
rect 6508 516 6514 518
rect 6206 507 6514 516
rect 9306 572 9614 581
rect 9306 570 9312 572
rect 9368 570 9392 572
rect 9448 570 9472 572
rect 9528 570 9552 572
rect 9608 570 9614 572
rect 9368 518 9370 570
rect 9550 518 9552 570
rect 9306 516 9312 518
rect 9368 516 9392 518
rect 9448 516 9472 518
rect 9528 516 9552 518
rect 9608 516 9614 518
rect 9306 507 9614 516
rect 12406 572 12714 581
rect 12406 570 12412 572
rect 12468 570 12492 572
rect 12548 570 12572 572
rect 12628 570 12652 572
rect 12708 570 12714 572
rect 12468 518 12470 570
rect 12650 518 12652 570
rect 12406 516 12412 518
rect 12468 516 12492 518
rect 12548 516 12572 518
rect 12628 516 12652 518
rect 12708 516 12714 518
rect 12406 507 12714 516
rect 15506 572 15814 581
rect 15506 570 15512 572
rect 15568 570 15592 572
rect 15648 570 15672 572
rect 15728 570 15752 572
rect 15808 570 15814 572
rect 15568 518 15570 570
rect 15750 518 15752 570
rect 15506 516 15512 518
rect 15568 516 15592 518
rect 15648 516 15672 518
rect 15728 516 15752 518
rect 15808 516 15814 518
rect 15506 507 15814 516
rect 18606 572 18914 581
rect 18606 570 18612 572
rect 18668 570 18692 572
rect 18748 570 18772 572
rect 18828 570 18852 572
rect 18908 570 18914 572
rect 18668 518 18670 570
rect 18850 518 18852 570
rect 18606 516 18612 518
rect 18668 516 18692 518
rect 18748 516 18772 518
rect 18828 516 18852 518
rect 18908 516 18914 518
rect 18606 507 18914 516
<< via2 >>
rect 1562 18522 1618 18524
rect 1642 18522 1698 18524
rect 1722 18522 1778 18524
rect 1802 18522 1858 18524
rect 1562 18470 1608 18522
rect 1608 18470 1618 18522
rect 1642 18470 1672 18522
rect 1672 18470 1684 18522
rect 1684 18470 1698 18522
rect 1722 18470 1736 18522
rect 1736 18470 1748 18522
rect 1748 18470 1778 18522
rect 1802 18470 1812 18522
rect 1812 18470 1858 18522
rect 1562 18468 1618 18470
rect 1642 18468 1698 18470
rect 1722 18468 1778 18470
rect 1802 18468 1858 18470
rect 4662 18522 4718 18524
rect 4742 18522 4798 18524
rect 4822 18522 4878 18524
rect 4902 18522 4958 18524
rect 4662 18470 4708 18522
rect 4708 18470 4718 18522
rect 4742 18470 4772 18522
rect 4772 18470 4784 18522
rect 4784 18470 4798 18522
rect 4822 18470 4836 18522
rect 4836 18470 4848 18522
rect 4848 18470 4878 18522
rect 4902 18470 4912 18522
rect 4912 18470 4958 18522
rect 4662 18468 4718 18470
rect 4742 18468 4798 18470
rect 4822 18468 4878 18470
rect 4902 18468 4958 18470
rect 1562 17434 1618 17436
rect 1642 17434 1698 17436
rect 1722 17434 1778 17436
rect 1802 17434 1858 17436
rect 1562 17382 1608 17434
rect 1608 17382 1618 17434
rect 1642 17382 1672 17434
rect 1672 17382 1684 17434
rect 1684 17382 1698 17434
rect 1722 17382 1736 17434
rect 1736 17382 1748 17434
rect 1748 17382 1778 17434
rect 1802 17382 1812 17434
rect 1812 17382 1858 17434
rect 1562 17380 1618 17382
rect 1642 17380 1698 17382
rect 1722 17380 1778 17382
rect 1802 17380 1858 17382
rect 1562 16346 1618 16348
rect 1642 16346 1698 16348
rect 1722 16346 1778 16348
rect 1802 16346 1858 16348
rect 1562 16294 1608 16346
rect 1608 16294 1618 16346
rect 1642 16294 1672 16346
rect 1672 16294 1684 16346
rect 1684 16294 1698 16346
rect 1722 16294 1736 16346
rect 1736 16294 1748 16346
rect 1748 16294 1778 16346
rect 1802 16294 1812 16346
rect 1812 16294 1858 16346
rect 1562 16292 1618 16294
rect 1642 16292 1698 16294
rect 1722 16292 1778 16294
rect 1802 16292 1858 16294
rect 1562 15258 1618 15260
rect 1642 15258 1698 15260
rect 1722 15258 1778 15260
rect 1802 15258 1858 15260
rect 1562 15206 1608 15258
rect 1608 15206 1618 15258
rect 1642 15206 1672 15258
rect 1672 15206 1684 15258
rect 1684 15206 1698 15258
rect 1722 15206 1736 15258
rect 1736 15206 1748 15258
rect 1748 15206 1778 15258
rect 1802 15206 1812 15258
rect 1812 15206 1858 15258
rect 1562 15204 1618 15206
rect 1642 15204 1698 15206
rect 1722 15204 1778 15206
rect 1802 15204 1858 15206
rect 3112 17978 3168 17980
rect 3192 17978 3248 17980
rect 3272 17978 3328 17980
rect 3352 17978 3408 17980
rect 3112 17926 3158 17978
rect 3158 17926 3168 17978
rect 3192 17926 3222 17978
rect 3222 17926 3234 17978
rect 3234 17926 3248 17978
rect 3272 17926 3286 17978
rect 3286 17926 3298 17978
rect 3298 17926 3328 17978
rect 3352 17926 3362 17978
rect 3362 17926 3408 17978
rect 3112 17924 3168 17926
rect 3192 17924 3248 17926
rect 3272 17924 3328 17926
rect 3352 17924 3408 17926
rect 3112 16890 3168 16892
rect 3192 16890 3248 16892
rect 3272 16890 3328 16892
rect 3352 16890 3408 16892
rect 3112 16838 3158 16890
rect 3158 16838 3168 16890
rect 3192 16838 3222 16890
rect 3222 16838 3234 16890
rect 3234 16838 3248 16890
rect 3272 16838 3286 16890
rect 3286 16838 3298 16890
rect 3298 16838 3328 16890
rect 3352 16838 3362 16890
rect 3362 16838 3408 16890
rect 3112 16836 3168 16838
rect 3192 16836 3248 16838
rect 3272 16836 3328 16838
rect 3352 16836 3408 16838
rect 1562 14170 1618 14172
rect 1642 14170 1698 14172
rect 1722 14170 1778 14172
rect 1802 14170 1858 14172
rect 1562 14118 1608 14170
rect 1608 14118 1618 14170
rect 1642 14118 1672 14170
rect 1672 14118 1684 14170
rect 1684 14118 1698 14170
rect 1722 14118 1736 14170
rect 1736 14118 1748 14170
rect 1748 14118 1778 14170
rect 1802 14118 1812 14170
rect 1812 14118 1858 14170
rect 1562 14116 1618 14118
rect 1642 14116 1698 14118
rect 1722 14116 1778 14118
rect 1802 14116 1858 14118
rect 1562 13082 1618 13084
rect 1642 13082 1698 13084
rect 1722 13082 1778 13084
rect 1802 13082 1858 13084
rect 1562 13030 1608 13082
rect 1608 13030 1618 13082
rect 1642 13030 1672 13082
rect 1672 13030 1684 13082
rect 1684 13030 1698 13082
rect 1722 13030 1736 13082
rect 1736 13030 1748 13082
rect 1748 13030 1778 13082
rect 1802 13030 1812 13082
rect 1812 13030 1858 13082
rect 1562 13028 1618 13030
rect 1642 13028 1698 13030
rect 1722 13028 1778 13030
rect 1802 13028 1858 13030
rect 1562 11994 1618 11996
rect 1642 11994 1698 11996
rect 1722 11994 1778 11996
rect 1802 11994 1858 11996
rect 1562 11942 1608 11994
rect 1608 11942 1618 11994
rect 1642 11942 1672 11994
rect 1672 11942 1684 11994
rect 1684 11942 1698 11994
rect 1722 11942 1736 11994
rect 1736 11942 1748 11994
rect 1748 11942 1778 11994
rect 1802 11942 1812 11994
rect 1812 11942 1858 11994
rect 1562 11940 1618 11942
rect 1642 11940 1698 11942
rect 1722 11940 1778 11942
rect 1802 11940 1858 11942
rect 1562 10906 1618 10908
rect 1642 10906 1698 10908
rect 1722 10906 1778 10908
rect 1802 10906 1858 10908
rect 1562 10854 1608 10906
rect 1608 10854 1618 10906
rect 1642 10854 1672 10906
rect 1672 10854 1684 10906
rect 1684 10854 1698 10906
rect 1722 10854 1736 10906
rect 1736 10854 1748 10906
rect 1748 10854 1778 10906
rect 1802 10854 1812 10906
rect 1812 10854 1858 10906
rect 1562 10852 1618 10854
rect 1642 10852 1698 10854
rect 1722 10852 1778 10854
rect 1802 10852 1858 10854
rect 938 9968 994 10024
rect 1562 9818 1618 9820
rect 1642 9818 1698 9820
rect 1722 9818 1778 9820
rect 1802 9818 1858 9820
rect 1562 9766 1608 9818
rect 1608 9766 1618 9818
rect 1642 9766 1672 9818
rect 1672 9766 1684 9818
rect 1684 9766 1698 9818
rect 1722 9766 1736 9818
rect 1736 9766 1748 9818
rect 1748 9766 1778 9818
rect 1802 9766 1812 9818
rect 1812 9766 1858 9818
rect 1562 9764 1618 9766
rect 1642 9764 1698 9766
rect 1722 9764 1778 9766
rect 1802 9764 1858 9766
rect 1562 8730 1618 8732
rect 1642 8730 1698 8732
rect 1722 8730 1778 8732
rect 1802 8730 1858 8732
rect 1562 8678 1608 8730
rect 1608 8678 1618 8730
rect 1642 8678 1672 8730
rect 1672 8678 1684 8730
rect 1684 8678 1698 8730
rect 1722 8678 1736 8730
rect 1736 8678 1748 8730
rect 1748 8678 1778 8730
rect 1802 8678 1812 8730
rect 1812 8678 1858 8730
rect 1562 8676 1618 8678
rect 1642 8676 1698 8678
rect 1722 8676 1778 8678
rect 1802 8676 1858 8678
rect 1562 7642 1618 7644
rect 1642 7642 1698 7644
rect 1722 7642 1778 7644
rect 1802 7642 1858 7644
rect 1562 7590 1608 7642
rect 1608 7590 1618 7642
rect 1642 7590 1672 7642
rect 1672 7590 1684 7642
rect 1684 7590 1698 7642
rect 1722 7590 1736 7642
rect 1736 7590 1748 7642
rect 1748 7590 1778 7642
rect 1802 7590 1812 7642
rect 1812 7590 1858 7642
rect 1562 7588 1618 7590
rect 1642 7588 1698 7590
rect 1722 7588 1778 7590
rect 1802 7588 1858 7590
rect 3112 15802 3168 15804
rect 3192 15802 3248 15804
rect 3272 15802 3328 15804
rect 3352 15802 3408 15804
rect 3112 15750 3158 15802
rect 3158 15750 3168 15802
rect 3192 15750 3222 15802
rect 3222 15750 3234 15802
rect 3234 15750 3248 15802
rect 3272 15750 3286 15802
rect 3286 15750 3298 15802
rect 3298 15750 3328 15802
rect 3352 15750 3362 15802
rect 3362 15750 3408 15802
rect 3112 15748 3168 15750
rect 3192 15748 3248 15750
rect 3272 15748 3328 15750
rect 3352 15748 3408 15750
rect 3112 14714 3168 14716
rect 3192 14714 3248 14716
rect 3272 14714 3328 14716
rect 3352 14714 3408 14716
rect 3112 14662 3158 14714
rect 3158 14662 3168 14714
rect 3192 14662 3222 14714
rect 3222 14662 3234 14714
rect 3234 14662 3248 14714
rect 3272 14662 3286 14714
rect 3286 14662 3298 14714
rect 3298 14662 3328 14714
rect 3352 14662 3362 14714
rect 3362 14662 3408 14714
rect 3112 14660 3168 14662
rect 3192 14660 3248 14662
rect 3272 14660 3328 14662
rect 3352 14660 3408 14662
rect 3112 13626 3168 13628
rect 3192 13626 3248 13628
rect 3272 13626 3328 13628
rect 3352 13626 3408 13628
rect 3112 13574 3158 13626
rect 3158 13574 3168 13626
rect 3192 13574 3222 13626
rect 3222 13574 3234 13626
rect 3234 13574 3248 13626
rect 3272 13574 3286 13626
rect 3286 13574 3298 13626
rect 3298 13574 3328 13626
rect 3352 13574 3362 13626
rect 3362 13574 3408 13626
rect 3112 13572 3168 13574
rect 3192 13572 3248 13574
rect 3272 13572 3328 13574
rect 3352 13572 3408 13574
rect 4662 17434 4718 17436
rect 4742 17434 4798 17436
rect 4822 17434 4878 17436
rect 4902 17434 4958 17436
rect 4662 17382 4708 17434
rect 4708 17382 4718 17434
rect 4742 17382 4772 17434
rect 4772 17382 4784 17434
rect 4784 17382 4798 17434
rect 4822 17382 4836 17434
rect 4836 17382 4848 17434
rect 4848 17382 4878 17434
rect 4902 17382 4912 17434
rect 4912 17382 4958 17434
rect 4662 17380 4718 17382
rect 4742 17380 4798 17382
rect 4822 17380 4878 17382
rect 4902 17380 4958 17382
rect 4662 16346 4718 16348
rect 4742 16346 4798 16348
rect 4822 16346 4878 16348
rect 4902 16346 4958 16348
rect 4662 16294 4708 16346
rect 4708 16294 4718 16346
rect 4742 16294 4772 16346
rect 4772 16294 4784 16346
rect 4784 16294 4798 16346
rect 4822 16294 4836 16346
rect 4836 16294 4848 16346
rect 4848 16294 4878 16346
rect 4902 16294 4912 16346
rect 4912 16294 4958 16346
rect 4662 16292 4718 16294
rect 4742 16292 4798 16294
rect 4822 16292 4878 16294
rect 4902 16292 4958 16294
rect 4662 15258 4718 15260
rect 4742 15258 4798 15260
rect 4822 15258 4878 15260
rect 4902 15258 4958 15260
rect 4662 15206 4708 15258
rect 4708 15206 4718 15258
rect 4742 15206 4772 15258
rect 4772 15206 4784 15258
rect 4784 15206 4798 15258
rect 4822 15206 4836 15258
rect 4836 15206 4848 15258
rect 4848 15206 4878 15258
rect 4902 15206 4912 15258
rect 4912 15206 4958 15258
rect 4662 15204 4718 15206
rect 4742 15204 4798 15206
rect 4822 15204 4878 15206
rect 4902 15204 4958 15206
rect 4662 14170 4718 14172
rect 4742 14170 4798 14172
rect 4822 14170 4878 14172
rect 4902 14170 4958 14172
rect 4662 14118 4708 14170
rect 4708 14118 4718 14170
rect 4742 14118 4772 14170
rect 4772 14118 4784 14170
rect 4784 14118 4798 14170
rect 4822 14118 4836 14170
rect 4836 14118 4848 14170
rect 4848 14118 4878 14170
rect 4902 14118 4912 14170
rect 4912 14118 4958 14170
rect 4662 14116 4718 14118
rect 4742 14116 4798 14118
rect 4822 14116 4878 14118
rect 4902 14116 4958 14118
rect 3112 12538 3168 12540
rect 3192 12538 3248 12540
rect 3272 12538 3328 12540
rect 3352 12538 3408 12540
rect 3112 12486 3158 12538
rect 3158 12486 3168 12538
rect 3192 12486 3222 12538
rect 3222 12486 3234 12538
rect 3234 12486 3248 12538
rect 3272 12486 3286 12538
rect 3286 12486 3298 12538
rect 3298 12486 3328 12538
rect 3352 12486 3362 12538
rect 3362 12486 3408 12538
rect 3112 12484 3168 12486
rect 3192 12484 3248 12486
rect 3272 12484 3328 12486
rect 3352 12484 3408 12486
rect 3112 11450 3168 11452
rect 3192 11450 3248 11452
rect 3272 11450 3328 11452
rect 3352 11450 3408 11452
rect 3112 11398 3158 11450
rect 3158 11398 3168 11450
rect 3192 11398 3222 11450
rect 3222 11398 3234 11450
rect 3234 11398 3248 11450
rect 3272 11398 3286 11450
rect 3286 11398 3298 11450
rect 3298 11398 3328 11450
rect 3352 11398 3362 11450
rect 3362 11398 3408 11450
rect 3112 11396 3168 11398
rect 3192 11396 3248 11398
rect 3272 11396 3328 11398
rect 3352 11396 3408 11398
rect 3112 10362 3168 10364
rect 3192 10362 3248 10364
rect 3272 10362 3328 10364
rect 3352 10362 3408 10364
rect 3112 10310 3158 10362
rect 3158 10310 3168 10362
rect 3192 10310 3222 10362
rect 3222 10310 3234 10362
rect 3234 10310 3248 10362
rect 3272 10310 3286 10362
rect 3286 10310 3298 10362
rect 3298 10310 3328 10362
rect 3352 10310 3362 10362
rect 3362 10310 3408 10362
rect 3112 10308 3168 10310
rect 3192 10308 3248 10310
rect 3272 10308 3328 10310
rect 3352 10308 3408 10310
rect 3112 9274 3168 9276
rect 3192 9274 3248 9276
rect 3272 9274 3328 9276
rect 3352 9274 3408 9276
rect 3112 9222 3158 9274
rect 3158 9222 3168 9274
rect 3192 9222 3222 9274
rect 3222 9222 3234 9274
rect 3234 9222 3248 9274
rect 3272 9222 3286 9274
rect 3286 9222 3298 9274
rect 3298 9222 3328 9274
rect 3352 9222 3362 9274
rect 3362 9222 3408 9274
rect 3112 9220 3168 9222
rect 3192 9220 3248 9222
rect 3272 9220 3328 9222
rect 3352 9220 3408 9222
rect 1562 6554 1618 6556
rect 1642 6554 1698 6556
rect 1722 6554 1778 6556
rect 1802 6554 1858 6556
rect 1562 6502 1608 6554
rect 1608 6502 1618 6554
rect 1642 6502 1672 6554
rect 1672 6502 1684 6554
rect 1684 6502 1698 6554
rect 1722 6502 1736 6554
rect 1736 6502 1748 6554
rect 1748 6502 1778 6554
rect 1802 6502 1812 6554
rect 1812 6502 1858 6554
rect 1562 6500 1618 6502
rect 1642 6500 1698 6502
rect 1722 6500 1778 6502
rect 1802 6500 1858 6502
rect 1562 5466 1618 5468
rect 1642 5466 1698 5468
rect 1722 5466 1778 5468
rect 1802 5466 1858 5468
rect 1562 5414 1608 5466
rect 1608 5414 1618 5466
rect 1642 5414 1672 5466
rect 1672 5414 1684 5466
rect 1684 5414 1698 5466
rect 1722 5414 1736 5466
rect 1736 5414 1748 5466
rect 1748 5414 1778 5466
rect 1802 5414 1812 5466
rect 1812 5414 1858 5466
rect 1562 5412 1618 5414
rect 1642 5412 1698 5414
rect 1722 5412 1778 5414
rect 1802 5412 1858 5414
rect 3112 8186 3168 8188
rect 3192 8186 3248 8188
rect 3272 8186 3328 8188
rect 3352 8186 3408 8188
rect 3112 8134 3158 8186
rect 3158 8134 3168 8186
rect 3192 8134 3222 8186
rect 3222 8134 3234 8186
rect 3234 8134 3248 8186
rect 3272 8134 3286 8186
rect 3286 8134 3298 8186
rect 3298 8134 3328 8186
rect 3352 8134 3362 8186
rect 3362 8134 3408 8186
rect 3112 8132 3168 8134
rect 3192 8132 3248 8134
rect 3272 8132 3328 8134
rect 3352 8132 3408 8134
rect 4662 13082 4718 13084
rect 4742 13082 4798 13084
rect 4822 13082 4878 13084
rect 4902 13082 4958 13084
rect 4662 13030 4708 13082
rect 4708 13030 4718 13082
rect 4742 13030 4772 13082
rect 4772 13030 4784 13082
rect 4784 13030 4798 13082
rect 4822 13030 4836 13082
rect 4836 13030 4848 13082
rect 4848 13030 4878 13082
rect 4902 13030 4912 13082
rect 4912 13030 4958 13082
rect 4662 13028 4718 13030
rect 4742 13028 4798 13030
rect 4822 13028 4878 13030
rect 4902 13028 4958 13030
rect 6212 17978 6268 17980
rect 6292 17978 6348 17980
rect 6372 17978 6428 17980
rect 6452 17978 6508 17980
rect 6212 17926 6258 17978
rect 6258 17926 6268 17978
rect 6292 17926 6322 17978
rect 6322 17926 6334 17978
rect 6334 17926 6348 17978
rect 6372 17926 6386 17978
rect 6386 17926 6398 17978
rect 6398 17926 6428 17978
rect 6452 17926 6462 17978
rect 6462 17926 6508 17978
rect 6212 17924 6268 17926
rect 6292 17924 6348 17926
rect 6372 17924 6428 17926
rect 6452 17924 6508 17926
rect 6212 16890 6268 16892
rect 6292 16890 6348 16892
rect 6372 16890 6428 16892
rect 6452 16890 6508 16892
rect 6212 16838 6258 16890
rect 6258 16838 6268 16890
rect 6292 16838 6322 16890
rect 6322 16838 6334 16890
rect 6334 16838 6348 16890
rect 6372 16838 6386 16890
rect 6386 16838 6398 16890
rect 6398 16838 6428 16890
rect 6452 16838 6462 16890
rect 6462 16838 6508 16890
rect 6212 16836 6268 16838
rect 6292 16836 6348 16838
rect 6372 16836 6428 16838
rect 6452 16836 6508 16838
rect 6212 15802 6268 15804
rect 6292 15802 6348 15804
rect 6372 15802 6428 15804
rect 6452 15802 6508 15804
rect 6212 15750 6258 15802
rect 6258 15750 6268 15802
rect 6292 15750 6322 15802
rect 6322 15750 6334 15802
rect 6334 15750 6348 15802
rect 6372 15750 6386 15802
rect 6386 15750 6398 15802
rect 6398 15750 6428 15802
rect 6452 15750 6462 15802
rect 6462 15750 6508 15802
rect 6212 15748 6268 15750
rect 6292 15748 6348 15750
rect 6372 15748 6428 15750
rect 6452 15748 6508 15750
rect 6212 14714 6268 14716
rect 6292 14714 6348 14716
rect 6372 14714 6428 14716
rect 6452 14714 6508 14716
rect 6212 14662 6258 14714
rect 6258 14662 6268 14714
rect 6292 14662 6322 14714
rect 6322 14662 6334 14714
rect 6334 14662 6348 14714
rect 6372 14662 6386 14714
rect 6386 14662 6398 14714
rect 6398 14662 6428 14714
rect 6452 14662 6462 14714
rect 6462 14662 6508 14714
rect 6212 14660 6268 14662
rect 6292 14660 6348 14662
rect 6372 14660 6428 14662
rect 6452 14660 6508 14662
rect 7762 18522 7818 18524
rect 7842 18522 7898 18524
rect 7922 18522 7978 18524
rect 8002 18522 8058 18524
rect 7762 18470 7808 18522
rect 7808 18470 7818 18522
rect 7842 18470 7872 18522
rect 7872 18470 7884 18522
rect 7884 18470 7898 18522
rect 7922 18470 7936 18522
rect 7936 18470 7948 18522
rect 7948 18470 7978 18522
rect 8002 18470 8012 18522
rect 8012 18470 8058 18522
rect 7762 18468 7818 18470
rect 7842 18468 7898 18470
rect 7922 18468 7978 18470
rect 8002 18468 8058 18470
rect 7762 17434 7818 17436
rect 7842 17434 7898 17436
rect 7922 17434 7978 17436
rect 8002 17434 8058 17436
rect 7762 17382 7808 17434
rect 7808 17382 7818 17434
rect 7842 17382 7872 17434
rect 7872 17382 7884 17434
rect 7884 17382 7898 17434
rect 7922 17382 7936 17434
rect 7936 17382 7948 17434
rect 7948 17382 7978 17434
rect 8002 17382 8012 17434
rect 8012 17382 8058 17434
rect 7762 17380 7818 17382
rect 7842 17380 7898 17382
rect 7922 17380 7978 17382
rect 8002 17380 8058 17382
rect 6212 13626 6268 13628
rect 6292 13626 6348 13628
rect 6372 13626 6428 13628
rect 6452 13626 6508 13628
rect 6212 13574 6258 13626
rect 6258 13574 6268 13626
rect 6292 13574 6322 13626
rect 6322 13574 6334 13626
rect 6334 13574 6348 13626
rect 6372 13574 6386 13626
rect 6386 13574 6398 13626
rect 6398 13574 6428 13626
rect 6452 13574 6462 13626
rect 6462 13574 6508 13626
rect 6212 13572 6268 13574
rect 6292 13572 6348 13574
rect 6372 13572 6428 13574
rect 6452 13572 6508 13574
rect 7762 16346 7818 16348
rect 7842 16346 7898 16348
rect 7922 16346 7978 16348
rect 8002 16346 8058 16348
rect 7762 16294 7808 16346
rect 7808 16294 7818 16346
rect 7842 16294 7872 16346
rect 7872 16294 7884 16346
rect 7884 16294 7898 16346
rect 7922 16294 7936 16346
rect 7936 16294 7948 16346
rect 7948 16294 7978 16346
rect 8002 16294 8012 16346
rect 8012 16294 8058 16346
rect 7762 16292 7818 16294
rect 7842 16292 7898 16294
rect 7922 16292 7978 16294
rect 8002 16292 8058 16294
rect 9312 17978 9368 17980
rect 9392 17978 9448 17980
rect 9472 17978 9528 17980
rect 9552 17978 9608 17980
rect 9312 17926 9358 17978
rect 9358 17926 9368 17978
rect 9392 17926 9422 17978
rect 9422 17926 9434 17978
rect 9434 17926 9448 17978
rect 9472 17926 9486 17978
rect 9486 17926 9498 17978
rect 9498 17926 9528 17978
rect 9552 17926 9562 17978
rect 9562 17926 9608 17978
rect 9312 17924 9368 17926
rect 9392 17924 9448 17926
rect 9472 17924 9528 17926
rect 9552 17924 9608 17926
rect 10862 18522 10918 18524
rect 10942 18522 10998 18524
rect 11022 18522 11078 18524
rect 11102 18522 11158 18524
rect 10862 18470 10908 18522
rect 10908 18470 10918 18522
rect 10942 18470 10972 18522
rect 10972 18470 10984 18522
rect 10984 18470 10998 18522
rect 11022 18470 11036 18522
rect 11036 18470 11048 18522
rect 11048 18470 11078 18522
rect 11102 18470 11112 18522
rect 11112 18470 11158 18522
rect 10862 18468 10918 18470
rect 10942 18468 10998 18470
rect 11022 18468 11078 18470
rect 11102 18468 11158 18470
rect 9312 16890 9368 16892
rect 9392 16890 9448 16892
rect 9472 16890 9528 16892
rect 9552 16890 9608 16892
rect 9312 16838 9358 16890
rect 9358 16838 9368 16890
rect 9392 16838 9422 16890
rect 9422 16838 9434 16890
rect 9434 16838 9448 16890
rect 9472 16838 9486 16890
rect 9486 16838 9498 16890
rect 9498 16838 9528 16890
rect 9552 16838 9562 16890
rect 9562 16838 9608 16890
rect 9312 16836 9368 16838
rect 9392 16836 9448 16838
rect 9472 16836 9528 16838
rect 9552 16836 9608 16838
rect 4662 11994 4718 11996
rect 4742 11994 4798 11996
rect 4822 11994 4878 11996
rect 4902 11994 4958 11996
rect 4662 11942 4708 11994
rect 4708 11942 4718 11994
rect 4742 11942 4772 11994
rect 4772 11942 4784 11994
rect 4784 11942 4798 11994
rect 4822 11942 4836 11994
rect 4836 11942 4848 11994
rect 4848 11942 4878 11994
rect 4902 11942 4912 11994
rect 4912 11942 4958 11994
rect 4662 11940 4718 11942
rect 4742 11940 4798 11942
rect 4822 11940 4878 11942
rect 4902 11940 4958 11942
rect 1562 4378 1618 4380
rect 1642 4378 1698 4380
rect 1722 4378 1778 4380
rect 1802 4378 1858 4380
rect 1562 4326 1608 4378
rect 1608 4326 1618 4378
rect 1642 4326 1672 4378
rect 1672 4326 1684 4378
rect 1684 4326 1698 4378
rect 1722 4326 1736 4378
rect 1736 4326 1748 4378
rect 1748 4326 1778 4378
rect 1802 4326 1812 4378
rect 1812 4326 1858 4378
rect 1562 4324 1618 4326
rect 1642 4324 1698 4326
rect 1722 4324 1778 4326
rect 1802 4324 1858 4326
rect 1562 3290 1618 3292
rect 1642 3290 1698 3292
rect 1722 3290 1778 3292
rect 1802 3290 1858 3292
rect 1562 3238 1608 3290
rect 1608 3238 1618 3290
rect 1642 3238 1672 3290
rect 1672 3238 1684 3290
rect 1684 3238 1698 3290
rect 1722 3238 1736 3290
rect 1736 3238 1748 3290
rect 1748 3238 1778 3290
rect 1802 3238 1812 3290
rect 1812 3238 1858 3290
rect 1562 3236 1618 3238
rect 1642 3236 1698 3238
rect 1722 3236 1778 3238
rect 1802 3236 1858 3238
rect 3112 7098 3168 7100
rect 3192 7098 3248 7100
rect 3272 7098 3328 7100
rect 3352 7098 3408 7100
rect 3112 7046 3158 7098
rect 3158 7046 3168 7098
rect 3192 7046 3222 7098
rect 3222 7046 3234 7098
rect 3234 7046 3248 7098
rect 3272 7046 3286 7098
rect 3286 7046 3298 7098
rect 3298 7046 3328 7098
rect 3352 7046 3362 7098
rect 3362 7046 3408 7098
rect 3112 7044 3168 7046
rect 3192 7044 3248 7046
rect 3272 7044 3328 7046
rect 3352 7044 3408 7046
rect 3112 6010 3168 6012
rect 3192 6010 3248 6012
rect 3272 6010 3328 6012
rect 3352 6010 3408 6012
rect 3112 5958 3158 6010
rect 3158 5958 3168 6010
rect 3192 5958 3222 6010
rect 3222 5958 3234 6010
rect 3234 5958 3248 6010
rect 3272 5958 3286 6010
rect 3286 5958 3298 6010
rect 3298 5958 3328 6010
rect 3352 5958 3362 6010
rect 3362 5958 3408 6010
rect 3112 5956 3168 5958
rect 3192 5956 3248 5958
rect 3272 5956 3328 5958
rect 3352 5956 3408 5958
rect 3112 4922 3168 4924
rect 3192 4922 3248 4924
rect 3272 4922 3328 4924
rect 3352 4922 3408 4924
rect 3112 4870 3158 4922
rect 3158 4870 3168 4922
rect 3192 4870 3222 4922
rect 3222 4870 3234 4922
rect 3234 4870 3248 4922
rect 3272 4870 3286 4922
rect 3286 4870 3298 4922
rect 3298 4870 3328 4922
rect 3352 4870 3362 4922
rect 3362 4870 3408 4922
rect 3112 4868 3168 4870
rect 3192 4868 3248 4870
rect 3272 4868 3328 4870
rect 3352 4868 3408 4870
rect 3112 3834 3168 3836
rect 3192 3834 3248 3836
rect 3272 3834 3328 3836
rect 3352 3834 3408 3836
rect 3112 3782 3158 3834
rect 3158 3782 3168 3834
rect 3192 3782 3222 3834
rect 3222 3782 3234 3834
rect 3234 3782 3248 3834
rect 3272 3782 3286 3834
rect 3286 3782 3298 3834
rect 3298 3782 3328 3834
rect 3352 3782 3362 3834
rect 3362 3782 3408 3834
rect 3112 3780 3168 3782
rect 3192 3780 3248 3782
rect 3272 3780 3328 3782
rect 3352 3780 3408 3782
rect 1562 2202 1618 2204
rect 1642 2202 1698 2204
rect 1722 2202 1778 2204
rect 1802 2202 1858 2204
rect 1562 2150 1608 2202
rect 1608 2150 1618 2202
rect 1642 2150 1672 2202
rect 1672 2150 1684 2202
rect 1684 2150 1698 2202
rect 1722 2150 1736 2202
rect 1736 2150 1748 2202
rect 1748 2150 1778 2202
rect 1802 2150 1812 2202
rect 1812 2150 1858 2202
rect 1562 2148 1618 2150
rect 1642 2148 1698 2150
rect 1722 2148 1778 2150
rect 1802 2148 1858 2150
rect 3112 2746 3168 2748
rect 3192 2746 3248 2748
rect 3272 2746 3328 2748
rect 3352 2746 3408 2748
rect 3112 2694 3158 2746
rect 3158 2694 3168 2746
rect 3192 2694 3222 2746
rect 3222 2694 3234 2746
rect 3234 2694 3248 2746
rect 3272 2694 3286 2746
rect 3286 2694 3298 2746
rect 3298 2694 3328 2746
rect 3352 2694 3362 2746
rect 3362 2694 3408 2746
rect 3112 2692 3168 2694
rect 3192 2692 3248 2694
rect 3272 2692 3328 2694
rect 3352 2692 3408 2694
rect 4662 10906 4718 10908
rect 4742 10906 4798 10908
rect 4822 10906 4878 10908
rect 4902 10906 4958 10908
rect 4662 10854 4708 10906
rect 4708 10854 4718 10906
rect 4742 10854 4772 10906
rect 4772 10854 4784 10906
rect 4784 10854 4798 10906
rect 4822 10854 4836 10906
rect 4836 10854 4848 10906
rect 4848 10854 4878 10906
rect 4902 10854 4912 10906
rect 4912 10854 4958 10906
rect 4662 10852 4718 10854
rect 4742 10852 4798 10854
rect 4822 10852 4878 10854
rect 4902 10852 4958 10854
rect 6212 12538 6268 12540
rect 6292 12538 6348 12540
rect 6372 12538 6428 12540
rect 6452 12538 6508 12540
rect 6212 12486 6258 12538
rect 6258 12486 6268 12538
rect 6292 12486 6322 12538
rect 6322 12486 6334 12538
rect 6334 12486 6348 12538
rect 6372 12486 6386 12538
rect 6386 12486 6398 12538
rect 6398 12486 6428 12538
rect 6452 12486 6462 12538
rect 6462 12486 6508 12538
rect 6212 12484 6268 12486
rect 6292 12484 6348 12486
rect 6372 12484 6428 12486
rect 6452 12484 6508 12486
rect 6212 11450 6268 11452
rect 6292 11450 6348 11452
rect 6372 11450 6428 11452
rect 6452 11450 6508 11452
rect 6212 11398 6258 11450
rect 6258 11398 6268 11450
rect 6292 11398 6322 11450
rect 6322 11398 6334 11450
rect 6334 11398 6348 11450
rect 6372 11398 6386 11450
rect 6386 11398 6398 11450
rect 6398 11398 6428 11450
rect 6452 11398 6462 11450
rect 6462 11398 6508 11450
rect 6212 11396 6268 11398
rect 6292 11396 6348 11398
rect 6372 11396 6428 11398
rect 6452 11396 6508 11398
rect 6212 10362 6268 10364
rect 6292 10362 6348 10364
rect 6372 10362 6428 10364
rect 6452 10362 6508 10364
rect 6212 10310 6258 10362
rect 6258 10310 6268 10362
rect 6292 10310 6322 10362
rect 6322 10310 6334 10362
rect 6334 10310 6348 10362
rect 6372 10310 6386 10362
rect 6386 10310 6398 10362
rect 6398 10310 6428 10362
rect 6452 10310 6462 10362
rect 6462 10310 6508 10362
rect 6212 10308 6268 10310
rect 6292 10308 6348 10310
rect 6372 10308 6428 10310
rect 6452 10308 6508 10310
rect 7762 15258 7818 15260
rect 7842 15258 7898 15260
rect 7922 15258 7978 15260
rect 8002 15258 8058 15260
rect 7762 15206 7808 15258
rect 7808 15206 7818 15258
rect 7842 15206 7872 15258
rect 7872 15206 7884 15258
rect 7884 15206 7898 15258
rect 7922 15206 7936 15258
rect 7936 15206 7948 15258
rect 7948 15206 7978 15258
rect 8002 15206 8012 15258
rect 8012 15206 8058 15258
rect 7762 15204 7818 15206
rect 7842 15204 7898 15206
rect 7922 15204 7978 15206
rect 8002 15204 8058 15206
rect 7762 14170 7818 14172
rect 7842 14170 7898 14172
rect 7922 14170 7978 14172
rect 8002 14170 8058 14172
rect 7762 14118 7808 14170
rect 7808 14118 7818 14170
rect 7842 14118 7872 14170
rect 7872 14118 7884 14170
rect 7884 14118 7898 14170
rect 7922 14118 7936 14170
rect 7936 14118 7948 14170
rect 7948 14118 7978 14170
rect 8002 14118 8012 14170
rect 8012 14118 8058 14170
rect 7762 14116 7818 14118
rect 7842 14116 7898 14118
rect 7922 14116 7978 14118
rect 8002 14116 8058 14118
rect 7762 13082 7818 13084
rect 7842 13082 7898 13084
rect 7922 13082 7978 13084
rect 8002 13082 8058 13084
rect 7762 13030 7808 13082
rect 7808 13030 7818 13082
rect 7842 13030 7872 13082
rect 7872 13030 7884 13082
rect 7884 13030 7898 13082
rect 7922 13030 7936 13082
rect 7936 13030 7948 13082
rect 7948 13030 7978 13082
rect 8002 13030 8012 13082
rect 8012 13030 8058 13082
rect 7762 13028 7818 13030
rect 7842 13028 7898 13030
rect 7922 13028 7978 13030
rect 8002 13028 8058 13030
rect 7762 11994 7818 11996
rect 7842 11994 7898 11996
rect 7922 11994 7978 11996
rect 8002 11994 8058 11996
rect 7762 11942 7808 11994
rect 7808 11942 7818 11994
rect 7842 11942 7872 11994
rect 7872 11942 7884 11994
rect 7884 11942 7898 11994
rect 7922 11942 7936 11994
rect 7936 11942 7948 11994
rect 7948 11942 7978 11994
rect 8002 11942 8012 11994
rect 8012 11942 8058 11994
rect 7762 11940 7818 11942
rect 7842 11940 7898 11942
rect 7922 11940 7978 11942
rect 8002 11940 8058 11942
rect 4662 9818 4718 9820
rect 4742 9818 4798 9820
rect 4822 9818 4878 9820
rect 4902 9818 4958 9820
rect 4662 9766 4708 9818
rect 4708 9766 4718 9818
rect 4742 9766 4772 9818
rect 4772 9766 4784 9818
rect 4784 9766 4798 9818
rect 4822 9766 4836 9818
rect 4836 9766 4848 9818
rect 4848 9766 4878 9818
rect 4902 9766 4912 9818
rect 4912 9766 4958 9818
rect 4662 9764 4718 9766
rect 4742 9764 4798 9766
rect 4822 9764 4878 9766
rect 4902 9764 4958 9766
rect 6212 9274 6268 9276
rect 6292 9274 6348 9276
rect 6372 9274 6428 9276
rect 6452 9274 6508 9276
rect 6212 9222 6258 9274
rect 6258 9222 6268 9274
rect 6292 9222 6322 9274
rect 6322 9222 6334 9274
rect 6334 9222 6348 9274
rect 6372 9222 6386 9274
rect 6386 9222 6398 9274
rect 6398 9222 6428 9274
rect 6452 9222 6462 9274
rect 6462 9222 6508 9274
rect 6212 9220 6268 9222
rect 6292 9220 6348 9222
rect 6372 9220 6428 9222
rect 6452 9220 6508 9222
rect 4662 8730 4718 8732
rect 4742 8730 4798 8732
rect 4822 8730 4878 8732
rect 4902 8730 4958 8732
rect 4662 8678 4708 8730
rect 4708 8678 4718 8730
rect 4742 8678 4772 8730
rect 4772 8678 4784 8730
rect 4784 8678 4798 8730
rect 4822 8678 4836 8730
rect 4836 8678 4848 8730
rect 4848 8678 4878 8730
rect 4902 8678 4912 8730
rect 4912 8678 4958 8730
rect 4662 8676 4718 8678
rect 4742 8676 4798 8678
rect 4822 8676 4878 8678
rect 4902 8676 4958 8678
rect 6212 8186 6268 8188
rect 6292 8186 6348 8188
rect 6372 8186 6428 8188
rect 6452 8186 6508 8188
rect 6212 8134 6258 8186
rect 6258 8134 6268 8186
rect 6292 8134 6322 8186
rect 6322 8134 6334 8186
rect 6334 8134 6348 8186
rect 6372 8134 6386 8186
rect 6386 8134 6398 8186
rect 6398 8134 6428 8186
rect 6452 8134 6462 8186
rect 6462 8134 6508 8186
rect 6212 8132 6268 8134
rect 6292 8132 6348 8134
rect 6372 8132 6428 8134
rect 6452 8132 6508 8134
rect 4662 7642 4718 7644
rect 4742 7642 4798 7644
rect 4822 7642 4878 7644
rect 4902 7642 4958 7644
rect 4662 7590 4708 7642
rect 4708 7590 4718 7642
rect 4742 7590 4772 7642
rect 4772 7590 4784 7642
rect 4784 7590 4798 7642
rect 4822 7590 4836 7642
rect 4836 7590 4848 7642
rect 4848 7590 4878 7642
rect 4902 7590 4912 7642
rect 4912 7590 4958 7642
rect 4662 7588 4718 7590
rect 4742 7588 4798 7590
rect 4822 7588 4878 7590
rect 4902 7588 4958 7590
rect 4662 6554 4718 6556
rect 4742 6554 4798 6556
rect 4822 6554 4878 6556
rect 4902 6554 4958 6556
rect 4662 6502 4708 6554
rect 4708 6502 4718 6554
rect 4742 6502 4772 6554
rect 4772 6502 4784 6554
rect 4784 6502 4798 6554
rect 4822 6502 4836 6554
rect 4836 6502 4848 6554
rect 4848 6502 4878 6554
rect 4902 6502 4912 6554
rect 4912 6502 4958 6554
rect 4662 6500 4718 6502
rect 4742 6500 4798 6502
rect 4822 6500 4878 6502
rect 4902 6500 4958 6502
rect 4662 5466 4718 5468
rect 4742 5466 4798 5468
rect 4822 5466 4878 5468
rect 4902 5466 4958 5468
rect 4662 5414 4708 5466
rect 4708 5414 4718 5466
rect 4742 5414 4772 5466
rect 4772 5414 4784 5466
rect 4784 5414 4798 5466
rect 4822 5414 4836 5466
rect 4836 5414 4848 5466
rect 4848 5414 4878 5466
rect 4902 5414 4912 5466
rect 4912 5414 4958 5466
rect 4662 5412 4718 5414
rect 4742 5412 4798 5414
rect 4822 5412 4878 5414
rect 4902 5412 4958 5414
rect 4662 4378 4718 4380
rect 4742 4378 4798 4380
rect 4822 4378 4878 4380
rect 4902 4378 4958 4380
rect 4662 4326 4708 4378
rect 4708 4326 4718 4378
rect 4742 4326 4772 4378
rect 4772 4326 4784 4378
rect 4784 4326 4798 4378
rect 4822 4326 4836 4378
rect 4836 4326 4848 4378
rect 4848 4326 4878 4378
rect 4902 4326 4912 4378
rect 4912 4326 4958 4378
rect 4662 4324 4718 4326
rect 4742 4324 4798 4326
rect 4822 4324 4878 4326
rect 4902 4324 4958 4326
rect 4662 3290 4718 3292
rect 4742 3290 4798 3292
rect 4822 3290 4878 3292
rect 4902 3290 4958 3292
rect 4662 3238 4708 3290
rect 4708 3238 4718 3290
rect 4742 3238 4772 3290
rect 4772 3238 4784 3290
rect 4784 3238 4798 3290
rect 4822 3238 4836 3290
rect 4836 3238 4848 3290
rect 4848 3238 4878 3290
rect 4902 3238 4912 3290
rect 4912 3238 4958 3290
rect 4662 3236 4718 3238
rect 4742 3236 4798 3238
rect 4822 3236 4878 3238
rect 4902 3236 4958 3238
rect 6212 7098 6268 7100
rect 6292 7098 6348 7100
rect 6372 7098 6428 7100
rect 6452 7098 6508 7100
rect 6212 7046 6258 7098
rect 6258 7046 6268 7098
rect 6292 7046 6322 7098
rect 6322 7046 6334 7098
rect 6334 7046 6348 7098
rect 6372 7046 6386 7098
rect 6386 7046 6398 7098
rect 6398 7046 6428 7098
rect 6452 7046 6462 7098
rect 6462 7046 6508 7098
rect 6212 7044 6268 7046
rect 6292 7044 6348 7046
rect 6372 7044 6428 7046
rect 6452 7044 6508 7046
rect 6212 6010 6268 6012
rect 6292 6010 6348 6012
rect 6372 6010 6428 6012
rect 6452 6010 6508 6012
rect 6212 5958 6258 6010
rect 6258 5958 6268 6010
rect 6292 5958 6322 6010
rect 6322 5958 6334 6010
rect 6334 5958 6348 6010
rect 6372 5958 6386 6010
rect 6386 5958 6398 6010
rect 6398 5958 6428 6010
rect 6452 5958 6462 6010
rect 6462 5958 6508 6010
rect 6212 5956 6268 5958
rect 6292 5956 6348 5958
rect 6372 5956 6428 5958
rect 6452 5956 6508 5958
rect 6212 4922 6268 4924
rect 6292 4922 6348 4924
rect 6372 4922 6428 4924
rect 6452 4922 6508 4924
rect 6212 4870 6258 4922
rect 6258 4870 6268 4922
rect 6292 4870 6322 4922
rect 6322 4870 6334 4922
rect 6334 4870 6348 4922
rect 6372 4870 6386 4922
rect 6386 4870 6398 4922
rect 6398 4870 6428 4922
rect 6452 4870 6462 4922
rect 6462 4870 6508 4922
rect 6212 4868 6268 4870
rect 6292 4868 6348 4870
rect 6372 4868 6428 4870
rect 6452 4868 6508 4870
rect 6212 3834 6268 3836
rect 6292 3834 6348 3836
rect 6372 3834 6428 3836
rect 6452 3834 6508 3836
rect 6212 3782 6258 3834
rect 6258 3782 6268 3834
rect 6292 3782 6322 3834
rect 6322 3782 6334 3834
rect 6334 3782 6348 3834
rect 6372 3782 6386 3834
rect 6386 3782 6398 3834
rect 6398 3782 6428 3834
rect 6452 3782 6462 3834
rect 6462 3782 6508 3834
rect 6212 3780 6268 3782
rect 6292 3780 6348 3782
rect 6372 3780 6428 3782
rect 6452 3780 6508 3782
rect 4662 2202 4718 2204
rect 4742 2202 4798 2204
rect 4822 2202 4878 2204
rect 4902 2202 4958 2204
rect 4662 2150 4708 2202
rect 4708 2150 4718 2202
rect 4742 2150 4772 2202
rect 4772 2150 4784 2202
rect 4784 2150 4798 2202
rect 4822 2150 4836 2202
rect 4836 2150 4848 2202
rect 4848 2150 4878 2202
rect 4902 2150 4912 2202
rect 4912 2150 4958 2202
rect 4662 2148 4718 2150
rect 4742 2148 4798 2150
rect 4822 2148 4878 2150
rect 4902 2148 4958 2150
rect 7762 10906 7818 10908
rect 7842 10906 7898 10908
rect 7922 10906 7978 10908
rect 8002 10906 8058 10908
rect 7762 10854 7808 10906
rect 7808 10854 7818 10906
rect 7842 10854 7872 10906
rect 7872 10854 7884 10906
rect 7884 10854 7898 10906
rect 7922 10854 7936 10906
rect 7936 10854 7948 10906
rect 7948 10854 7978 10906
rect 8002 10854 8012 10906
rect 8012 10854 8058 10906
rect 7762 10852 7818 10854
rect 7842 10852 7898 10854
rect 7922 10852 7978 10854
rect 8002 10852 8058 10854
rect 7762 9818 7818 9820
rect 7842 9818 7898 9820
rect 7922 9818 7978 9820
rect 8002 9818 8058 9820
rect 7762 9766 7808 9818
rect 7808 9766 7818 9818
rect 7842 9766 7872 9818
rect 7872 9766 7884 9818
rect 7884 9766 7898 9818
rect 7922 9766 7936 9818
rect 7936 9766 7948 9818
rect 7948 9766 7978 9818
rect 8002 9766 8012 9818
rect 8012 9766 8058 9818
rect 7762 9764 7818 9766
rect 7842 9764 7898 9766
rect 7922 9764 7978 9766
rect 8002 9764 8058 9766
rect 7762 8730 7818 8732
rect 7842 8730 7898 8732
rect 7922 8730 7978 8732
rect 8002 8730 8058 8732
rect 7762 8678 7808 8730
rect 7808 8678 7818 8730
rect 7842 8678 7872 8730
rect 7872 8678 7884 8730
rect 7884 8678 7898 8730
rect 7922 8678 7936 8730
rect 7936 8678 7948 8730
rect 7948 8678 7978 8730
rect 8002 8678 8012 8730
rect 8012 8678 8058 8730
rect 7762 8676 7818 8678
rect 7842 8676 7898 8678
rect 7922 8676 7978 8678
rect 8002 8676 8058 8678
rect 7762 7642 7818 7644
rect 7842 7642 7898 7644
rect 7922 7642 7978 7644
rect 8002 7642 8058 7644
rect 7762 7590 7808 7642
rect 7808 7590 7818 7642
rect 7842 7590 7872 7642
rect 7872 7590 7884 7642
rect 7884 7590 7898 7642
rect 7922 7590 7936 7642
rect 7936 7590 7948 7642
rect 7948 7590 7978 7642
rect 8002 7590 8012 7642
rect 8012 7590 8058 7642
rect 7762 7588 7818 7590
rect 7842 7588 7898 7590
rect 7922 7588 7978 7590
rect 8002 7588 8058 7590
rect 7762 6554 7818 6556
rect 7842 6554 7898 6556
rect 7922 6554 7978 6556
rect 8002 6554 8058 6556
rect 7762 6502 7808 6554
rect 7808 6502 7818 6554
rect 7842 6502 7872 6554
rect 7872 6502 7884 6554
rect 7884 6502 7898 6554
rect 7922 6502 7936 6554
rect 7936 6502 7948 6554
rect 7948 6502 7978 6554
rect 8002 6502 8012 6554
rect 8012 6502 8058 6554
rect 7762 6500 7818 6502
rect 7842 6500 7898 6502
rect 7922 6500 7978 6502
rect 8002 6500 8058 6502
rect 7762 5466 7818 5468
rect 7842 5466 7898 5468
rect 7922 5466 7978 5468
rect 8002 5466 8058 5468
rect 7762 5414 7808 5466
rect 7808 5414 7818 5466
rect 7842 5414 7872 5466
rect 7872 5414 7884 5466
rect 7884 5414 7898 5466
rect 7922 5414 7936 5466
rect 7936 5414 7948 5466
rect 7948 5414 7978 5466
rect 8002 5414 8012 5466
rect 8012 5414 8058 5466
rect 7762 5412 7818 5414
rect 7842 5412 7898 5414
rect 7922 5412 7978 5414
rect 8002 5412 8058 5414
rect 6212 2746 6268 2748
rect 6292 2746 6348 2748
rect 6372 2746 6428 2748
rect 6452 2746 6508 2748
rect 6212 2694 6258 2746
rect 6258 2694 6268 2746
rect 6292 2694 6322 2746
rect 6322 2694 6334 2746
rect 6334 2694 6348 2746
rect 6372 2694 6386 2746
rect 6386 2694 6398 2746
rect 6398 2694 6428 2746
rect 6452 2694 6462 2746
rect 6462 2694 6508 2746
rect 6212 2692 6268 2694
rect 6292 2692 6348 2694
rect 6372 2692 6428 2694
rect 6452 2692 6508 2694
rect 3112 1658 3168 1660
rect 3192 1658 3248 1660
rect 3272 1658 3328 1660
rect 3352 1658 3408 1660
rect 3112 1606 3158 1658
rect 3158 1606 3168 1658
rect 3192 1606 3222 1658
rect 3222 1606 3234 1658
rect 3234 1606 3248 1658
rect 3272 1606 3286 1658
rect 3286 1606 3298 1658
rect 3298 1606 3328 1658
rect 3352 1606 3362 1658
rect 3362 1606 3408 1658
rect 3112 1604 3168 1606
rect 3192 1604 3248 1606
rect 3272 1604 3328 1606
rect 3352 1604 3408 1606
rect 1562 1114 1618 1116
rect 1642 1114 1698 1116
rect 1722 1114 1778 1116
rect 1802 1114 1858 1116
rect 1562 1062 1608 1114
rect 1608 1062 1618 1114
rect 1642 1062 1672 1114
rect 1672 1062 1684 1114
rect 1684 1062 1698 1114
rect 1722 1062 1736 1114
rect 1736 1062 1748 1114
rect 1748 1062 1778 1114
rect 1802 1062 1812 1114
rect 1812 1062 1858 1114
rect 1562 1060 1618 1062
rect 1642 1060 1698 1062
rect 1722 1060 1778 1062
rect 1802 1060 1858 1062
rect 4662 1114 4718 1116
rect 4742 1114 4798 1116
rect 4822 1114 4878 1116
rect 4902 1114 4958 1116
rect 4662 1062 4708 1114
rect 4708 1062 4718 1114
rect 4742 1062 4772 1114
rect 4772 1062 4784 1114
rect 4784 1062 4798 1114
rect 4822 1062 4836 1114
rect 4836 1062 4848 1114
rect 4848 1062 4878 1114
rect 4902 1062 4912 1114
rect 4912 1062 4958 1114
rect 4662 1060 4718 1062
rect 4742 1060 4798 1062
rect 4822 1060 4878 1062
rect 4902 1060 4958 1062
rect 6212 1658 6268 1660
rect 6292 1658 6348 1660
rect 6372 1658 6428 1660
rect 6452 1658 6508 1660
rect 6212 1606 6258 1658
rect 6258 1606 6268 1658
rect 6292 1606 6322 1658
rect 6322 1606 6334 1658
rect 6334 1606 6348 1658
rect 6372 1606 6386 1658
rect 6386 1606 6398 1658
rect 6398 1606 6428 1658
rect 6452 1606 6462 1658
rect 6462 1606 6508 1658
rect 6212 1604 6268 1606
rect 6292 1604 6348 1606
rect 6372 1604 6428 1606
rect 6452 1604 6508 1606
rect 7762 4378 7818 4380
rect 7842 4378 7898 4380
rect 7922 4378 7978 4380
rect 8002 4378 8058 4380
rect 7762 4326 7808 4378
rect 7808 4326 7818 4378
rect 7842 4326 7872 4378
rect 7872 4326 7884 4378
rect 7884 4326 7898 4378
rect 7922 4326 7936 4378
rect 7936 4326 7948 4378
rect 7948 4326 7978 4378
rect 8002 4326 8012 4378
rect 8012 4326 8058 4378
rect 7762 4324 7818 4326
rect 7842 4324 7898 4326
rect 7922 4324 7978 4326
rect 8002 4324 8058 4326
rect 7762 3290 7818 3292
rect 7842 3290 7898 3292
rect 7922 3290 7978 3292
rect 8002 3290 8058 3292
rect 7762 3238 7808 3290
rect 7808 3238 7818 3290
rect 7842 3238 7872 3290
rect 7872 3238 7884 3290
rect 7884 3238 7898 3290
rect 7922 3238 7936 3290
rect 7936 3238 7948 3290
rect 7948 3238 7978 3290
rect 8002 3238 8012 3290
rect 8012 3238 8058 3290
rect 7762 3236 7818 3238
rect 7842 3236 7898 3238
rect 7922 3236 7978 3238
rect 8002 3236 8058 3238
rect 9312 15802 9368 15804
rect 9392 15802 9448 15804
rect 9472 15802 9528 15804
rect 9552 15802 9608 15804
rect 9312 15750 9358 15802
rect 9358 15750 9368 15802
rect 9392 15750 9422 15802
rect 9422 15750 9434 15802
rect 9434 15750 9448 15802
rect 9472 15750 9486 15802
rect 9486 15750 9498 15802
rect 9498 15750 9528 15802
rect 9552 15750 9562 15802
rect 9562 15750 9608 15802
rect 9312 15748 9368 15750
rect 9392 15748 9448 15750
rect 9472 15748 9528 15750
rect 9552 15748 9608 15750
rect 10862 17434 10918 17436
rect 10942 17434 10998 17436
rect 11022 17434 11078 17436
rect 11102 17434 11158 17436
rect 10862 17382 10908 17434
rect 10908 17382 10918 17434
rect 10942 17382 10972 17434
rect 10972 17382 10984 17434
rect 10984 17382 10998 17434
rect 11022 17382 11036 17434
rect 11036 17382 11048 17434
rect 11048 17382 11078 17434
rect 11102 17382 11112 17434
rect 11112 17382 11158 17434
rect 10862 17380 10918 17382
rect 10942 17380 10998 17382
rect 11022 17380 11078 17382
rect 11102 17380 11158 17382
rect 12412 17978 12468 17980
rect 12492 17978 12548 17980
rect 12572 17978 12628 17980
rect 12652 17978 12708 17980
rect 12412 17926 12458 17978
rect 12458 17926 12468 17978
rect 12492 17926 12522 17978
rect 12522 17926 12534 17978
rect 12534 17926 12548 17978
rect 12572 17926 12586 17978
rect 12586 17926 12598 17978
rect 12598 17926 12628 17978
rect 12652 17926 12662 17978
rect 12662 17926 12708 17978
rect 12412 17924 12468 17926
rect 12492 17924 12548 17926
rect 12572 17924 12628 17926
rect 12652 17924 12708 17926
rect 10862 16346 10918 16348
rect 10942 16346 10998 16348
rect 11022 16346 11078 16348
rect 11102 16346 11158 16348
rect 10862 16294 10908 16346
rect 10908 16294 10918 16346
rect 10942 16294 10972 16346
rect 10972 16294 10984 16346
rect 10984 16294 10998 16346
rect 11022 16294 11036 16346
rect 11036 16294 11048 16346
rect 11048 16294 11078 16346
rect 11102 16294 11112 16346
rect 11112 16294 11158 16346
rect 10862 16292 10918 16294
rect 10942 16292 10998 16294
rect 11022 16292 11078 16294
rect 11102 16292 11158 16294
rect 9312 14714 9368 14716
rect 9392 14714 9448 14716
rect 9472 14714 9528 14716
rect 9552 14714 9608 14716
rect 9312 14662 9358 14714
rect 9358 14662 9368 14714
rect 9392 14662 9422 14714
rect 9422 14662 9434 14714
rect 9434 14662 9448 14714
rect 9472 14662 9486 14714
rect 9486 14662 9498 14714
rect 9498 14662 9528 14714
rect 9552 14662 9562 14714
rect 9562 14662 9608 14714
rect 9312 14660 9368 14662
rect 9392 14660 9448 14662
rect 9472 14660 9528 14662
rect 9552 14660 9608 14662
rect 9312 13626 9368 13628
rect 9392 13626 9448 13628
rect 9472 13626 9528 13628
rect 9552 13626 9608 13628
rect 9312 13574 9358 13626
rect 9358 13574 9368 13626
rect 9392 13574 9422 13626
rect 9422 13574 9434 13626
rect 9434 13574 9448 13626
rect 9472 13574 9486 13626
rect 9486 13574 9498 13626
rect 9498 13574 9528 13626
rect 9552 13574 9562 13626
rect 9562 13574 9608 13626
rect 9312 13572 9368 13574
rect 9392 13572 9448 13574
rect 9472 13572 9528 13574
rect 9552 13572 9608 13574
rect 9312 12538 9368 12540
rect 9392 12538 9448 12540
rect 9472 12538 9528 12540
rect 9552 12538 9608 12540
rect 9312 12486 9358 12538
rect 9358 12486 9368 12538
rect 9392 12486 9422 12538
rect 9422 12486 9434 12538
rect 9434 12486 9448 12538
rect 9472 12486 9486 12538
rect 9486 12486 9498 12538
rect 9498 12486 9528 12538
rect 9552 12486 9562 12538
rect 9562 12486 9608 12538
rect 9312 12484 9368 12486
rect 9392 12484 9448 12486
rect 9472 12484 9528 12486
rect 9552 12484 9608 12486
rect 10862 15258 10918 15260
rect 10942 15258 10998 15260
rect 11022 15258 11078 15260
rect 11102 15258 11158 15260
rect 10862 15206 10908 15258
rect 10908 15206 10918 15258
rect 10942 15206 10972 15258
rect 10972 15206 10984 15258
rect 10984 15206 10998 15258
rect 11022 15206 11036 15258
rect 11036 15206 11048 15258
rect 11048 15206 11078 15258
rect 11102 15206 11112 15258
rect 11112 15206 11158 15258
rect 10862 15204 10918 15206
rect 10942 15204 10998 15206
rect 11022 15204 11078 15206
rect 11102 15204 11158 15206
rect 10862 14170 10918 14172
rect 10942 14170 10998 14172
rect 11022 14170 11078 14172
rect 11102 14170 11158 14172
rect 10862 14118 10908 14170
rect 10908 14118 10918 14170
rect 10942 14118 10972 14170
rect 10972 14118 10984 14170
rect 10984 14118 10998 14170
rect 11022 14118 11036 14170
rect 11036 14118 11048 14170
rect 11048 14118 11078 14170
rect 11102 14118 11112 14170
rect 11112 14118 11158 14170
rect 10862 14116 10918 14118
rect 10942 14116 10998 14118
rect 11022 14116 11078 14118
rect 11102 14116 11158 14118
rect 9312 11450 9368 11452
rect 9392 11450 9448 11452
rect 9472 11450 9528 11452
rect 9552 11450 9608 11452
rect 9312 11398 9358 11450
rect 9358 11398 9368 11450
rect 9392 11398 9422 11450
rect 9422 11398 9434 11450
rect 9434 11398 9448 11450
rect 9472 11398 9486 11450
rect 9486 11398 9498 11450
rect 9498 11398 9528 11450
rect 9552 11398 9562 11450
rect 9562 11398 9608 11450
rect 9312 11396 9368 11398
rect 9392 11396 9448 11398
rect 9472 11396 9528 11398
rect 9552 11396 9608 11398
rect 9312 10362 9368 10364
rect 9392 10362 9448 10364
rect 9472 10362 9528 10364
rect 9552 10362 9608 10364
rect 9312 10310 9358 10362
rect 9358 10310 9368 10362
rect 9392 10310 9422 10362
rect 9422 10310 9434 10362
rect 9434 10310 9448 10362
rect 9472 10310 9486 10362
rect 9486 10310 9498 10362
rect 9498 10310 9528 10362
rect 9552 10310 9562 10362
rect 9562 10310 9608 10362
rect 9312 10308 9368 10310
rect 9392 10308 9448 10310
rect 9472 10308 9528 10310
rect 9552 10308 9608 10310
rect 9312 9274 9368 9276
rect 9392 9274 9448 9276
rect 9472 9274 9528 9276
rect 9552 9274 9608 9276
rect 9312 9222 9358 9274
rect 9358 9222 9368 9274
rect 9392 9222 9422 9274
rect 9422 9222 9434 9274
rect 9434 9222 9448 9274
rect 9472 9222 9486 9274
rect 9486 9222 9498 9274
rect 9498 9222 9528 9274
rect 9552 9222 9562 9274
rect 9562 9222 9608 9274
rect 9312 9220 9368 9222
rect 9392 9220 9448 9222
rect 9472 9220 9528 9222
rect 9552 9220 9608 9222
rect 10862 13082 10918 13084
rect 10942 13082 10998 13084
rect 11022 13082 11078 13084
rect 11102 13082 11158 13084
rect 10862 13030 10908 13082
rect 10908 13030 10918 13082
rect 10942 13030 10972 13082
rect 10972 13030 10984 13082
rect 10984 13030 10998 13082
rect 11022 13030 11036 13082
rect 11036 13030 11048 13082
rect 11048 13030 11078 13082
rect 11102 13030 11112 13082
rect 11112 13030 11158 13082
rect 10862 13028 10918 13030
rect 10942 13028 10998 13030
rect 11022 13028 11078 13030
rect 11102 13028 11158 13030
rect 13962 18522 14018 18524
rect 14042 18522 14098 18524
rect 14122 18522 14178 18524
rect 14202 18522 14258 18524
rect 13962 18470 14008 18522
rect 14008 18470 14018 18522
rect 14042 18470 14072 18522
rect 14072 18470 14084 18522
rect 14084 18470 14098 18522
rect 14122 18470 14136 18522
rect 14136 18470 14148 18522
rect 14148 18470 14178 18522
rect 14202 18470 14212 18522
rect 14212 18470 14258 18522
rect 13962 18468 14018 18470
rect 14042 18468 14098 18470
rect 14122 18468 14178 18470
rect 14202 18468 14258 18470
rect 12412 16890 12468 16892
rect 12492 16890 12548 16892
rect 12572 16890 12628 16892
rect 12652 16890 12708 16892
rect 12412 16838 12458 16890
rect 12458 16838 12468 16890
rect 12492 16838 12522 16890
rect 12522 16838 12534 16890
rect 12534 16838 12548 16890
rect 12572 16838 12586 16890
rect 12586 16838 12598 16890
rect 12598 16838 12628 16890
rect 12652 16838 12662 16890
rect 12662 16838 12708 16890
rect 12412 16836 12468 16838
rect 12492 16836 12548 16838
rect 12572 16836 12628 16838
rect 12652 16836 12708 16838
rect 12412 15802 12468 15804
rect 12492 15802 12548 15804
rect 12572 15802 12628 15804
rect 12652 15802 12708 15804
rect 12412 15750 12458 15802
rect 12458 15750 12468 15802
rect 12492 15750 12522 15802
rect 12522 15750 12534 15802
rect 12534 15750 12548 15802
rect 12572 15750 12586 15802
rect 12586 15750 12598 15802
rect 12598 15750 12628 15802
rect 12652 15750 12662 15802
rect 12662 15750 12708 15802
rect 12412 15748 12468 15750
rect 12492 15748 12548 15750
rect 12572 15748 12628 15750
rect 12652 15748 12708 15750
rect 13358 16632 13414 16688
rect 13962 17434 14018 17436
rect 14042 17434 14098 17436
rect 14122 17434 14178 17436
rect 14202 17434 14258 17436
rect 13962 17382 14008 17434
rect 14008 17382 14018 17434
rect 14042 17382 14072 17434
rect 14072 17382 14084 17434
rect 14084 17382 14098 17434
rect 14122 17382 14136 17434
rect 14136 17382 14148 17434
rect 14148 17382 14178 17434
rect 14202 17382 14212 17434
rect 14212 17382 14258 17434
rect 13962 17380 14018 17382
rect 14042 17380 14098 17382
rect 14122 17380 14178 17382
rect 14202 17380 14258 17382
rect 12412 14714 12468 14716
rect 12492 14714 12548 14716
rect 12572 14714 12628 14716
rect 12652 14714 12708 14716
rect 12412 14662 12458 14714
rect 12458 14662 12468 14714
rect 12492 14662 12522 14714
rect 12522 14662 12534 14714
rect 12534 14662 12548 14714
rect 12572 14662 12586 14714
rect 12586 14662 12598 14714
rect 12598 14662 12628 14714
rect 12652 14662 12662 14714
rect 12662 14662 12708 14714
rect 12412 14660 12468 14662
rect 12492 14660 12548 14662
rect 12572 14660 12628 14662
rect 12652 14660 12708 14662
rect 12412 13626 12468 13628
rect 12492 13626 12548 13628
rect 12572 13626 12628 13628
rect 12652 13626 12708 13628
rect 12412 13574 12458 13626
rect 12458 13574 12468 13626
rect 12492 13574 12522 13626
rect 12522 13574 12534 13626
rect 12534 13574 12548 13626
rect 12572 13574 12586 13626
rect 12586 13574 12598 13626
rect 12598 13574 12628 13626
rect 12652 13574 12662 13626
rect 12662 13574 12708 13626
rect 12412 13572 12468 13574
rect 12492 13572 12548 13574
rect 12572 13572 12628 13574
rect 12652 13572 12708 13574
rect 10862 11994 10918 11996
rect 10942 11994 10998 11996
rect 11022 11994 11078 11996
rect 11102 11994 11158 11996
rect 10862 11942 10908 11994
rect 10908 11942 10918 11994
rect 10942 11942 10972 11994
rect 10972 11942 10984 11994
rect 10984 11942 10998 11994
rect 11022 11942 11036 11994
rect 11036 11942 11048 11994
rect 11048 11942 11078 11994
rect 11102 11942 11112 11994
rect 11112 11942 11158 11994
rect 10862 11940 10918 11942
rect 10942 11940 10998 11942
rect 11022 11940 11078 11942
rect 11102 11940 11158 11942
rect 12412 12538 12468 12540
rect 12492 12538 12548 12540
rect 12572 12538 12628 12540
rect 12652 12538 12708 12540
rect 12412 12486 12458 12538
rect 12458 12486 12468 12538
rect 12492 12486 12522 12538
rect 12522 12486 12534 12538
rect 12534 12486 12548 12538
rect 12572 12486 12586 12538
rect 12586 12486 12598 12538
rect 12598 12486 12628 12538
rect 12652 12486 12662 12538
rect 12662 12486 12708 12538
rect 12412 12484 12468 12486
rect 12492 12484 12548 12486
rect 12572 12484 12628 12486
rect 12652 12484 12708 12486
rect 9312 8186 9368 8188
rect 9392 8186 9448 8188
rect 9472 8186 9528 8188
rect 9552 8186 9608 8188
rect 9312 8134 9358 8186
rect 9358 8134 9368 8186
rect 9392 8134 9422 8186
rect 9422 8134 9434 8186
rect 9434 8134 9448 8186
rect 9472 8134 9486 8186
rect 9486 8134 9498 8186
rect 9498 8134 9528 8186
rect 9552 8134 9562 8186
rect 9562 8134 9608 8186
rect 9312 8132 9368 8134
rect 9392 8132 9448 8134
rect 9472 8132 9528 8134
rect 9552 8132 9608 8134
rect 10862 10906 10918 10908
rect 10942 10906 10998 10908
rect 11022 10906 11078 10908
rect 11102 10906 11158 10908
rect 10862 10854 10908 10906
rect 10908 10854 10918 10906
rect 10942 10854 10972 10906
rect 10972 10854 10984 10906
rect 10984 10854 10998 10906
rect 11022 10854 11036 10906
rect 11036 10854 11048 10906
rect 11048 10854 11078 10906
rect 11102 10854 11112 10906
rect 11112 10854 11158 10906
rect 10862 10852 10918 10854
rect 10942 10852 10998 10854
rect 11022 10852 11078 10854
rect 11102 10852 11158 10854
rect 10862 9818 10918 9820
rect 10942 9818 10998 9820
rect 11022 9818 11078 9820
rect 11102 9818 11158 9820
rect 10862 9766 10908 9818
rect 10908 9766 10918 9818
rect 10942 9766 10972 9818
rect 10972 9766 10984 9818
rect 10984 9766 10998 9818
rect 11022 9766 11036 9818
rect 11036 9766 11048 9818
rect 11048 9766 11078 9818
rect 11102 9766 11112 9818
rect 11112 9766 11158 9818
rect 10862 9764 10918 9766
rect 10942 9764 10998 9766
rect 11022 9764 11078 9766
rect 11102 9764 11158 9766
rect 9312 7098 9368 7100
rect 9392 7098 9448 7100
rect 9472 7098 9528 7100
rect 9552 7098 9608 7100
rect 9312 7046 9358 7098
rect 9358 7046 9368 7098
rect 9392 7046 9422 7098
rect 9422 7046 9434 7098
rect 9434 7046 9448 7098
rect 9472 7046 9486 7098
rect 9486 7046 9498 7098
rect 9498 7046 9528 7098
rect 9552 7046 9562 7098
rect 9562 7046 9608 7098
rect 9312 7044 9368 7046
rect 9392 7044 9448 7046
rect 9472 7044 9528 7046
rect 9552 7044 9608 7046
rect 9312 6010 9368 6012
rect 9392 6010 9448 6012
rect 9472 6010 9528 6012
rect 9552 6010 9608 6012
rect 9312 5958 9358 6010
rect 9358 5958 9368 6010
rect 9392 5958 9422 6010
rect 9422 5958 9434 6010
rect 9434 5958 9448 6010
rect 9472 5958 9486 6010
rect 9486 5958 9498 6010
rect 9498 5958 9528 6010
rect 9552 5958 9562 6010
rect 9562 5958 9608 6010
rect 9312 5956 9368 5958
rect 9392 5956 9448 5958
rect 9472 5956 9528 5958
rect 9552 5956 9608 5958
rect 9312 4922 9368 4924
rect 9392 4922 9448 4924
rect 9472 4922 9528 4924
rect 9552 4922 9608 4924
rect 9312 4870 9358 4922
rect 9358 4870 9368 4922
rect 9392 4870 9422 4922
rect 9422 4870 9434 4922
rect 9434 4870 9448 4922
rect 9472 4870 9486 4922
rect 9486 4870 9498 4922
rect 9498 4870 9528 4922
rect 9552 4870 9562 4922
rect 9562 4870 9608 4922
rect 9312 4868 9368 4870
rect 9392 4868 9448 4870
rect 9472 4868 9528 4870
rect 9552 4868 9608 4870
rect 9312 3834 9368 3836
rect 9392 3834 9448 3836
rect 9472 3834 9528 3836
rect 9552 3834 9608 3836
rect 9312 3782 9358 3834
rect 9358 3782 9368 3834
rect 9392 3782 9422 3834
rect 9422 3782 9434 3834
rect 9434 3782 9448 3834
rect 9472 3782 9486 3834
rect 9486 3782 9498 3834
rect 9498 3782 9528 3834
rect 9552 3782 9562 3834
rect 9562 3782 9608 3834
rect 9312 3780 9368 3782
rect 9392 3780 9448 3782
rect 9472 3780 9528 3782
rect 9552 3780 9608 3782
rect 9312 2746 9368 2748
rect 9392 2746 9448 2748
rect 9472 2746 9528 2748
rect 9552 2746 9608 2748
rect 9312 2694 9358 2746
rect 9358 2694 9368 2746
rect 9392 2694 9422 2746
rect 9422 2694 9434 2746
rect 9434 2694 9448 2746
rect 9472 2694 9486 2746
rect 9486 2694 9498 2746
rect 9498 2694 9528 2746
rect 9552 2694 9562 2746
rect 9562 2694 9608 2746
rect 9312 2692 9368 2694
rect 9392 2692 9448 2694
rect 9472 2692 9528 2694
rect 9552 2692 9608 2694
rect 7762 2202 7818 2204
rect 7842 2202 7898 2204
rect 7922 2202 7978 2204
rect 8002 2202 8058 2204
rect 7762 2150 7808 2202
rect 7808 2150 7818 2202
rect 7842 2150 7872 2202
rect 7872 2150 7884 2202
rect 7884 2150 7898 2202
rect 7922 2150 7936 2202
rect 7936 2150 7948 2202
rect 7948 2150 7978 2202
rect 8002 2150 8012 2202
rect 8012 2150 8058 2202
rect 7762 2148 7818 2150
rect 7842 2148 7898 2150
rect 7922 2148 7978 2150
rect 8002 2148 8058 2150
rect 10862 8730 10918 8732
rect 10942 8730 10998 8732
rect 11022 8730 11078 8732
rect 11102 8730 11158 8732
rect 10862 8678 10908 8730
rect 10908 8678 10918 8730
rect 10942 8678 10972 8730
rect 10972 8678 10984 8730
rect 10984 8678 10998 8730
rect 11022 8678 11036 8730
rect 11036 8678 11048 8730
rect 11048 8678 11078 8730
rect 11102 8678 11112 8730
rect 11112 8678 11158 8730
rect 10862 8676 10918 8678
rect 10942 8676 10998 8678
rect 11022 8676 11078 8678
rect 11102 8676 11158 8678
rect 12412 11450 12468 11452
rect 12492 11450 12548 11452
rect 12572 11450 12628 11452
rect 12652 11450 12708 11452
rect 12412 11398 12458 11450
rect 12458 11398 12468 11450
rect 12492 11398 12522 11450
rect 12522 11398 12534 11450
rect 12534 11398 12548 11450
rect 12572 11398 12586 11450
rect 12586 11398 12598 11450
rect 12598 11398 12628 11450
rect 12652 11398 12662 11450
rect 12662 11398 12708 11450
rect 12412 11396 12468 11398
rect 12492 11396 12548 11398
rect 12572 11396 12628 11398
rect 12652 11396 12708 11398
rect 12412 10362 12468 10364
rect 12492 10362 12548 10364
rect 12572 10362 12628 10364
rect 12652 10362 12708 10364
rect 12412 10310 12458 10362
rect 12458 10310 12468 10362
rect 12492 10310 12522 10362
rect 12522 10310 12534 10362
rect 12534 10310 12548 10362
rect 12572 10310 12586 10362
rect 12586 10310 12598 10362
rect 12598 10310 12628 10362
rect 12652 10310 12662 10362
rect 12662 10310 12708 10362
rect 12412 10308 12468 10310
rect 12492 10308 12548 10310
rect 12572 10308 12628 10310
rect 12652 10308 12708 10310
rect 12412 9274 12468 9276
rect 12492 9274 12548 9276
rect 12572 9274 12628 9276
rect 12652 9274 12708 9276
rect 12412 9222 12458 9274
rect 12458 9222 12468 9274
rect 12492 9222 12522 9274
rect 12522 9222 12534 9274
rect 12534 9222 12548 9274
rect 12572 9222 12586 9274
rect 12586 9222 12598 9274
rect 12598 9222 12628 9274
rect 12652 9222 12662 9274
rect 12662 9222 12708 9274
rect 12412 9220 12468 9222
rect 12492 9220 12548 9222
rect 12572 9220 12628 9222
rect 12652 9220 12708 9222
rect 10862 7642 10918 7644
rect 10942 7642 10998 7644
rect 11022 7642 11078 7644
rect 11102 7642 11158 7644
rect 10862 7590 10908 7642
rect 10908 7590 10918 7642
rect 10942 7590 10972 7642
rect 10972 7590 10984 7642
rect 10984 7590 10998 7642
rect 11022 7590 11036 7642
rect 11036 7590 11048 7642
rect 11048 7590 11078 7642
rect 11102 7590 11112 7642
rect 11112 7590 11158 7642
rect 10862 7588 10918 7590
rect 10942 7588 10998 7590
rect 11022 7588 11078 7590
rect 11102 7588 11158 7590
rect 12412 8186 12468 8188
rect 12492 8186 12548 8188
rect 12572 8186 12628 8188
rect 12652 8186 12708 8188
rect 12412 8134 12458 8186
rect 12458 8134 12468 8186
rect 12492 8134 12522 8186
rect 12522 8134 12534 8186
rect 12534 8134 12548 8186
rect 12572 8134 12586 8186
rect 12586 8134 12598 8186
rect 12598 8134 12628 8186
rect 12652 8134 12662 8186
rect 12662 8134 12708 8186
rect 12412 8132 12468 8134
rect 12492 8132 12548 8134
rect 12572 8132 12628 8134
rect 12652 8132 12708 8134
rect 10862 6554 10918 6556
rect 10942 6554 10998 6556
rect 11022 6554 11078 6556
rect 11102 6554 11158 6556
rect 10862 6502 10908 6554
rect 10908 6502 10918 6554
rect 10942 6502 10972 6554
rect 10972 6502 10984 6554
rect 10984 6502 10998 6554
rect 11022 6502 11036 6554
rect 11036 6502 11048 6554
rect 11048 6502 11078 6554
rect 11102 6502 11112 6554
rect 11112 6502 11158 6554
rect 10862 6500 10918 6502
rect 10942 6500 10998 6502
rect 11022 6500 11078 6502
rect 11102 6500 11158 6502
rect 10862 5466 10918 5468
rect 10942 5466 10998 5468
rect 11022 5466 11078 5468
rect 11102 5466 11158 5468
rect 10862 5414 10908 5466
rect 10908 5414 10918 5466
rect 10942 5414 10972 5466
rect 10972 5414 10984 5466
rect 10984 5414 10998 5466
rect 11022 5414 11036 5466
rect 11036 5414 11048 5466
rect 11048 5414 11078 5466
rect 11102 5414 11112 5466
rect 11112 5414 11158 5466
rect 10862 5412 10918 5414
rect 10942 5412 10998 5414
rect 11022 5412 11078 5414
rect 11102 5412 11158 5414
rect 14278 16632 14334 16688
rect 13962 16346 14018 16348
rect 14042 16346 14098 16348
rect 14122 16346 14178 16348
rect 14202 16346 14258 16348
rect 13962 16294 14008 16346
rect 14008 16294 14018 16346
rect 14042 16294 14072 16346
rect 14072 16294 14084 16346
rect 14084 16294 14098 16346
rect 14122 16294 14136 16346
rect 14136 16294 14148 16346
rect 14148 16294 14178 16346
rect 14202 16294 14212 16346
rect 14212 16294 14258 16346
rect 13962 16292 14018 16294
rect 14042 16292 14098 16294
rect 14122 16292 14178 16294
rect 14202 16292 14258 16294
rect 13962 15258 14018 15260
rect 14042 15258 14098 15260
rect 14122 15258 14178 15260
rect 14202 15258 14258 15260
rect 13962 15206 14008 15258
rect 14008 15206 14018 15258
rect 14042 15206 14072 15258
rect 14072 15206 14084 15258
rect 14084 15206 14098 15258
rect 14122 15206 14136 15258
rect 14136 15206 14148 15258
rect 14148 15206 14178 15258
rect 14202 15206 14212 15258
rect 14212 15206 14258 15258
rect 13962 15204 14018 15206
rect 14042 15204 14098 15206
rect 14122 15204 14178 15206
rect 14202 15204 14258 15206
rect 14738 16632 14794 16688
rect 13962 14170 14018 14172
rect 14042 14170 14098 14172
rect 14122 14170 14178 14172
rect 14202 14170 14258 14172
rect 13962 14118 14008 14170
rect 14008 14118 14018 14170
rect 14042 14118 14072 14170
rect 14072 14118 14084 14170
rect 14084 14118 14098 14170
rect 14122 14118 14136 14170
rect 14136 14118 14148 14170
rect 14148 14118 14178 14170
rect 14202 14118 14212 14170
rect 14212 14118 14258 14170
rect 13962 14116 14018 14118
rect 14042 14116 14098 14118
rect 14122 14116 14178 14118
rect 14202 14116 14258 14118
rect 12412 7098 12468 7100
rect 12492 7098 12548 7100
rect 12572 7098 12628 7100
rect 12652 7098 12708 7100
rect 12412 7046 12458 7098
rect 12458 7046 12468 7098
rect 12492 7046 12522 7098
rect 12522 7046 12534 7098
rect 12534 7046 12548 7098
rect 12572 7046 12586 7098
rect 12586 7046 12598 7098
rect 12598 7046 12628 7098
rect 12652 7046 12662 7098
rect 12662 7046 12708 7098
rect 12412 7044 12468 7046
rect 12492 7044 12548 7046
rect 12572 7044 12628 7046
rect 12652 7044 12708 7046
rect 12412 6010 12468 6012
rect 12492 6010 12548 6012
rect 12572 6010 12628 6012
rect 12652 6010 12708 6012
rect 12412 5958 12458 6010
rect 12458 5958 12468 6010
rect 12492 5958 12522 6010
rect 12522 5958 12534 6010
rect 12534 5958 12548 6010
rect 12572 5958 12586 6010
rect 12586 5958 12598 6010
rect 12598 5958 12628 6010
rect 12652 5958 12662 6010
rect 12662 5958 12708 6010
rect 12412 5956 12468 5958
rect 12492 5956 12548 5958
rect 12572 5956 12628 5958
rect 12652 5956 12708 5958
rect 12412 4922 12468 4924
rect 12492 4922 12548 4924
rect 12572 4922 12628 4924
rect 12652 4922 12708 4924
rect 12412 4870 12458 4922
rect 12458 4870 12468 4922
rect 12492 4870 12522 4922
rect 12522 4870 12534 4922
rect 12534 4870 12548 4922
rect 12572 4870 12586 4922
rect 12586 4870 12598 4922
rect 12598 4870 12628 4922
rect 12652 4870 12662 4922
rect 12662 4870 12708 4922
rect 12412 4868 12468 4870
rect 12492 4868 12548 4870
rect 12572 4868 12628 4870
rect 12652 4868 12708 4870
rect 13962 13082 14018 13084
rect 14042 13082 14098 13084
rect 14122 13082 14178 13084
rect 14202 13082 14258 13084
rect 13962 13030 14008 13082
rect 14008 13030 14018 13082
rect 14042 13030 14072 13082
rect 14072 13030 14084 13082
rect 14084 13030 14098 13082
rect 14122 13030 14136 13082
rect 14136 13030 14148 13082
rect 14148 13030 14178 13082
rect 14202 13030 14212 13082
rect 14212 13030 14258 13082
rect 13962 13028 14018 13030
rect 14042 13028 14098 13030
rect 14122 13028 14178 13030
rect 14202 13028 14258 13030
rect 13962 11994 14018 11996
rect 14042 11994 14098 11996
rect 14122 11994 14178 11996
rect 14202 11994 14258 11996
rect 13962 11942 14008 11994
rect 14008 11942 14018 11994
rect 14042 11942 14072 11994
rect 14072 11942 14084 11994
rect 14084 11942 14098 11994
rect 14122 11942 14136 11994
rect 14136 11942 14148 11994
rect 14148 11942 14178 11994
rect 14202 11942 14212 11994
rect 14212 11942 14258 11994
rect 13962 11940 14018 11942
rect 14042 11940 14098 11942
rect 14122 11940 14178 11942
rect 14202 11940 14258 11942
rect 13962 10906 14018 10908
rect 14042 10906 14098 10908
rect 14122 10906 14178 10908
rect 14202 10906 14258 10908
rect 13962 10854 14008 10906
rect 14008 10854 14018 10906
rect 14042 10854 14072 10906
rect 14072 10854 14084 10906
rect 14084 10854 14098 10906
rect 14122 10854 14136 10906
rect 14136 10854 14148 10906
rect 14148 10854 14178 10906
rect 14202 10854 14212 10906
rect 14212 10854 14258 10906
rect 13962 10852 14018 10854
rect 14042 10852 14098 10854
rect 14122 10852 14178 10854
rect 14202 10852 14258 10854
rect 13962 9818 14018 9820
rect 14042 9818 14098 9820
rect 14122 9818 14178 9820
rect 14202 9818 14258 9820
rect 13962 9766 14008 9818
rect 14008 9766 14018 9818
rect 14042 9766 14072 9818
rect 14072 9766 14084 9818
rect 14084 9766 14098 9818
rect 14122 9766 14136 9818
rect 14136 9766 14148 9818
rect 14148 9766 14178 9818
rect 14202 9766 14212 9818
rect 14212 9766 14258 9818
rect 13962 9764 14018 9766
rect 14042 9764 14098 9766
rect 14122 9764 14178 9766
rect 14202 9764 14258 9766
rect 13962 8730 14018 8732
rect 14042 8730 14098 8732
rect 14122 8730 14178 8732
rect 14202 8730 14258 8732
rect 13962 8678 14008 8730
rect 14008 8678 14018 8730
rect 14042 8678 14072 8730
rect 14072 8678 14084 8730
rect 14084 8678 14098 8730
rect 14122 8678 14136 8730
rect 14136 8678 14148 8730
rect 14148 8678 14178 8730
rect 14202 8678 14212 8730
rect 14212 8678 14258 8730
rect 13962 8676 14018 8678
rect 14042 8676 14098 8678
rect 14122 8676 14178 8678
rect 14202 8676 14258 8678
rect 13962 7642 14018 7644
rect 14042 7642 14098 7644
rect 14122 7642 14178 7644
rect 14202 7642 14258 7644
rect 13962 7590 14008 7642
rect 14008 7590 14018 7642
rect 14042 7590 14072 7642
rect 14072 7590 14084 7642
rect 14084 7590 14098 7642
rect 14122 7590 14136 7642
rect 14136 7590 14148 7642
rect 14148 7590 14178 7642
rect 14202 7590 14212 7642
rect 14212 7590 14258 7642
rect 13962 7588 14018 7590
rect 14042 7588 14098 7590
rect 14122 7588 14178 7590
rect 14202 7588 14258 7590
rect 13962 6554 14018 6556
rect 14042 6554 14098 6556
rect 14122 6554 14178 6556
rect 14202 6554 14258 6556
rect 13962 6502 14008 6554
rect 14008 6502 14018 6554
rect 14042 6502 14072 6554
rect 14072 6502 14084 6554
rect 14084 6502 14098 6554
rect 14122 6502 14136 6554
rect 14136 6502 14148 6554
rect 14148 6502 14178 6554
rect 14202 6502 14212 6554
rect 14212 6502 14258 6554
rect 13962 6500 14018 6502
rect 14042 6500 14098 6502
rect 14122 6500 14178 6502
rect 14202 6500 14258 6502
rect 13962 5466 14018 5468
rect 14042 5466 14098 5468
rect 14122 5466 14178 5468
rect 14202 5466 14258 5468
rect 13962 5414 14008 5466
rect 14008 5414 14018 5466
rect 14042 5414 14072 5466
rect 14072 5414 14084 5466
rect 14084 5414 14098 5466
rect 14122 5414 14136 5466
rect 14136 5414 14148 5466
rect 14148 5414 14178 5466
rect 14202 5414 14212 5466
rect 14212 5414 14258 5466
rect 13962 5412 14018 5414
rect 14042 5412 14098 5414
rect 14122 5412 14178 5414
rect 14202 5412 14258 5414
rect 18418 18536 18474 18592
rect 17062 18522 17118 18524
rect 17142 18522 17198 18524
rect 17222 18522 17278 18524
rect 17302 18522 17358 18524
rect 17062 18470 17108 18522
rect 17108 18470 17118 18522
rect 17142 18470 17172 18522
rect 17172 18470 17184 18522
rect 17184 18470 17198 18522
rect 17222 18470 17236 18522
rect 17236 18470 17248 18522
rect 17248 18470 17278 18522
rect 17302 18470 17312 18522
rect 17312 18470 17358 18522
rect 17062 18468 17118 18470
rect 17142 18468 17198 18470
rect 17222 18468 17278 18470
rect 17302 18468 17358 18470
rect 15512 17978 15568 17980
rect 15592 17978 15648 17980
rect 15672 17978 15728 17980
rect 15752 17978 15808 17980
rect 15512 17926 15558 17978
rect 15558 17926 15568 17978
rect 15592 17926 15622 17978
rect 15622 17926 15634 17978
rect 15634 17926 15648 17978
rect 15672 17926 15686 17978
rect 15686 17926 15698 17978
rect 15698 17926 15728 17978
rect 15752 17926 15762 17978
rect 15762 17926 15808 17978
rect 15512 17924 15568 17926
rect 15592 17924 15648 17926
rect 15672 17924 15728 17926
rect 15752 17924 15808 17926
rect 15512 16890 15568 16892
rect 15592 16890 15648 16892
rect 15672 16890 15728 16892
rect 15752 16890 15808 16892
rect 15512 16838 15558 16890
rect 15558 16838 15568 16890
rect 15592 16838 15622 16890
rect 15622 16838 15634 16890
rect 15634 16838 15648 16890
rect 15672 16838 15686 16890
rect 15686 16838 15698 16890
rect 15698 16838 15728 16890
rect 15752 16838 15762 16890
rect 15762 16838 15808 16890
rect 15512 16836 15568 16838
rect 15592 16836 15648 16838
rect 15672 16836 15728 16838
rect 15752 16836 15808 16838
rect 16302 16632 16358 16688
rect 15512 15802 15568 15804
rect 15592 15802 15648 15804
rect 15672 15802 15728 15804
rect 15752 15802 15808 15804
rect 15512 15750 15558 15802
rect 15558 15750 15568 15802
rect 15592 15750 15622 15802
rect 15622 15750 15634 15802
rect 15634 15750 15648 15802
rect 15672 15750 15686 15802
rect 15686 15750 15698 15802
rect 15698 15750 15728 15802
rect 15752 15750 15762 15802
rect 15762 15750 15808 15802
rect 15512 15748 15568 15750
rect 15592 15748 15648 15750
rect 15672 15748 15728 15750
rect 15752 15748 15808 15750
rect 15512 14714 15568 14716
rect 15592 14714 15648 14716
rect 15672 14714 15728 14716
rect 15752 14714 15808 14716
rect 15512 14662 15558 14714
rect 15558 14662 15568 14714
rect 15592 14662 15622 14714
rect 15622 14662 15634 14714
rect 15634 14662 15648 14714
rect 15672 14662 15686 14714
rect 15686 14662 15698 14714
rect 15698 14662 15728 14714
rect 15752 14662 15762 14714
rect 15762 14662 15808 14714
rect 15512 14660 15568 14662
rect 15592 14660 15648 14662
rect 15672 14660 15728 14662
rect 15752 14660 15808 14662
rect 15512 13626 15568 13628
rect 15592 13626 15648 13628
rect 15672 13626 15728 13628
rect 15752 13626 15808 13628
rect 15512 13574 15558 13626
rect 15558 13574 15568 13626
rect 15592 13574 15622 13626
rect 15622 13574 15634 13626
rect 15634 13574 15648 13626
rect 15672 13574 15686 13626
rect 15686 13574 15698 13626
rect 15698 13574 15728 13626
rect 15752 13574 15762 13626
rect 15762 13574 15808 13626
rect 15512 13572 15568 13574
rect 15592 13572 15648 13574
rect 15672 13572 15728 13574
rect 15752 13572 15808 13574
rect 15512 12538 15568 12540
rect 15592 12538 15648 12540
rect 15672 12538 15728 12540
rect 15752 12538 15808 12540
rect 15512 12486 15558 12538
rect 15558 12486 15568 12538
rect 15592 12486 15622 12538
rect 15622 12486 15634 12538
rect 15634 12486 15648 12538
rect 15672 12486 15686 12538
rect 15686 12486 15698 12538
rect 15698 12486 15728 12538
rect 15752 12486 15762 12538
rect 15762 12486 15808 12538
rect 15512 12484 15568 12486
rect 15592 12484 15648 12486
rect 15672 12484 15728 12486
rect 15752 12484 15808 12486
rect 15512 11450 15568 11452
rect 15592 11450 15648 11452
rect 15672 11450 15728 11452
rect 15752 11450 15808 11452
rect 15512 11398 15558 11450
rect 15558 11398 15568 11450
rect 15592 11398 15622 11450
rect 15622 11398 15634 11450
rect 15634 11398 15648 11450
rect 15672 11398 15686 11450
rect 15686 11398 15698 11450
rect 15698 11398 15728 11450
rect 15752 11398 15762 11450
rect 15762 11398 15808 11450
rect 15512 11396 15568 11398
rect 15592 11396 15648 11398
rect 15672 11396 15728 11398
rect 15752 11396 15808 11398
rect 15512 10362 15568 10364
rect 15592 10362 15648 10364
rect 15672 10362 15728 10364
rect 15752 10362 15808 10364
rect 15512 10310 15558 10362
rect 15558 10310 15568 10362
rect 15592 10310 15622 10362
rect 15622 10310 15634 10362
rect 15634 10310 15648 10362
rect 15672 10310 15686 10362
rect 15686 10310 15698 10362
rect 15698 10310 15728 10362
rect 15752 10310 15762 10362
rect 15762 10310 15808 10362
rect 15512 10308 15568 10310
rect 15592 10308 15648 10310
rect 15672 10308 15728 10310
rect 15752 10308 15808 10310
rect 15512 9274 15568 9276
rect 15592 9274 15648 9276
rect 15672 9274 15728 9276
rect 15752 9274 15808 9276
rect 15512 9222 15558 9274
rect 15558 9222 15568 9274
rect 15592 9222 15622 9274
rect 15622 9222 15634 9274
rect 15634 9222 15648 9274
rect 15672 9222 15686 9274
rect 15686 9222 15698 9274
rect 15698 9222 15728 9274
rect 15752 9222 15762 9274
rect 15762 9222 15808 9274
rect 15512 9220 15568 9222
rect 15592 9220 15648 9222
rect 15672 9220 15728 9222
rect 15752 9220 15808 9222
rect 15512 8186 15568 8188
rect 15592 8186 15648 8188
rect 15672 8186 15728 8188
rect 15752 8186 15808 8188
rect 15512 8134 15558 8186
rect 15558 8134 15568 8186
rect 15592 8134 15622 8186
rect 15622 8134 15634 8186
rect 15634 8134 15648 8186
rect 15672 8134 15686 8186
rect 15686 8134 15698 8186
rect 15698 8134 15728 8186
rect 15752 8134 15762 8186
rect 15762 8134 15808 8186
rect 15512 8132 15568 8134
rect 15592 8132 15648 8134
rect 15672 8132 15728 8134
rect 15752 8132 15808 8134
rect 17062 17434 17118 17436
rect 17142 17434 17198 17436
rect 17222 17434 17278 17436
rect 17302 17434 17358 17436
rect 17062 17382 17108 17434
rect 17108 17382 17118 17434
rect 17142 17382 17172 17434
rect 17172 17382 17184 17434
rect 17184 17382 17198 17434
rect 17222 17382 17236 17434
rect 17236 17382 17248 17434
rect 17248 17382 17278 17434
rect 17302 17382 17312 17434
rect 17312 17382 17358 17434
rect 17062 17380 17118 17382
rect 17142 17380 17198 17382
rect 17222 17380 17278 17382
rect 17302 17380 17358 17382
rect 17062 16346 17118 16348
rect 17142 16346 17198 16348
rect 17222 16346 17278 16348
rect 17302 16346 17358 16348
rect 17062 16294 17108 16346
rect 17108 16294 17118 16346
rect 17142 16294 17172 16346
rect 17172 16294 17184 16346
rect 17184 16294 17198 16346
rect 17222 16294 17236 16346
rect 17236 16294 17248 16346
rect 17248 16294 17278 16346
rect 17302 16294 17312 16346
rect 17312 16294 17358 16346
rect 17062 16292 17118 16294
rect 17142 16292 17198 16294
rect 17222 16292 17278 16294
rect 17302 16292 17358 16294
rect 17062 15258 17118 15260
rect 17142 15258 17198 15260
rect 17222 15258 17278 15260
rect 17302 15258 17358 15260
rect 17062 15206 17108 15258
rect 17108 15206 17118 15258
rect 17142 15206 17172 15258
rect 17172 15206 17184 15258
rect 17184 15206 17198 15258
rect 17222 15206 17236 15258
rect 17236 15206 17248 15258
rect 17248 15206 17278 15258
rect 17302 15206 17312 15258
rect 17312 15206 17358 15258
rect 17062 15204 17118 15206
rect 17142 15204 17198 15206
rect 17222 15204 17278 15206
rect 17302 15204 17358 15206
rect 18418 16124 18420 16144
rect 18420 16124 18472 16144
rect 18472 16124 18474 16144
rect 18418 16088 18474 16124
rect 10862 4378 10918 4380
rect 10942 4378 10998 4380
rect 11022 4378 11078 4380
rect 11102 4378 11158 4380
rect 10862 4326 10908 4378
rect 10908 4326 10918 4378
rect 10942 4326 10972 4378
rect 10972 4326 10984 4378
rect 10984 4326 10998 4378
rect 11022 4326 11036 4378
rect 11036 4326 11048 4378
rect 11048 4326 11078 4378
rect 11102 4326 11112 4378
rect 11112 4326 11158 4378
rect 10862 4324 10918 4326
rect 10942 4324 10998 4326
rect 11022 4324 11078 4326
rect 11102 4324 11158 4326
rect 12412 3834 12468 3836
rect 12492 3834 12548 3836
rect 12572 3834 12628 3836
rect 12652 3834 12708 3836
rect 12412 3782 12458 3834
rect 12458 3782 12468 3834
rect 12492 3782 12522 3834
rect 12522 3782 12534 3834
rect 12534 3782 12548 3834
rect 12572 3782 12586 3834
rect 12586 3782 12598 3834
rect 12598 3782 12628 3834
rect 12652 3782 12662 3834
rect 12662 3782 12708 3834
rect 12412 3780 12468 3782
rect 12492 3780 12548 3782
rect 12572 3780 12628 3782
rect 12652 3780 12708 3782
rect 10862 3290 10918 3292
rect 10942 3290 10998 3292
rect 11022 3290 11078 3292
rect 11102 3290 11158 3292
rect 10862 3238 10908 3290
rect 10908 3238 10918 3290
rect 10942 3238 10972 3290
rect 10972 3238 10984 3290
rect 10984 3238 10998 3290
rect 11022 3238 11036 3290
rect 11036 3238 11048 3290
rect 11048 3238 11078 3290
rect 11102 3238 11112 3290
rect 11112 3238 11158 3290
rect 10862 3236 10918 3238
rect 10942 3236 10998 3238
rect 11022 3236 11078 3238
rect 11102 3236 11158 3238
rect 10862 2202 10918 2204
rect 10942 2202 10998 2204
rect 11022 2202 11078 2204
rect 11102 2202 11158 2204
rect 10862 2150 10908 2202
rect 10908 2150 10918 2202
rect 10942 2150 10972 2202
rect 10972 2150 10984 2202
rect 10984 2150 10998 2202
rect 11022 2150 11036 2202
rect 11036 2150 11048 2202
rect 11048 2150 11078 2202
rect 11102 2150 11112 2202
rect 11112 2150 11158 2202
rect 10862 2148 10918 2150
rect 10942 2148 10998 2150
rect 11022 2148 11078 2150
rect 11102 2148 11158 2150
rect 12412 2746 12468 2748
rect 12492 2746 12548 2748
rect 12572 2746 12628 2748
rect 12652 2746 12708 2748
rect 12412 2694 12458 2746
rect 12458 2694 12468 2746
rect 12492 2694 12522 2746
rect 12522 2694 12534 2746
rect 12534 2694 12548 2746
rect 12572 2694 12586 2746
rect 12586 2694 12598 2746
rect 12598 2694 12628 2746
rect 12652 2694 12662 2746
rect 12662 2694 12708 2746
rect 12412 2692 12468 2694
rect 12492 2692 12548 2694
rect 12572 2692 12628 2694
rect 12652 2692 12708 2694
rect 9312 1658 9368 1660
rect 9392 1658 9448 1660
rect 9472 1658 9528 1660
rect 9552 1658 9608 1660
rect 9312 1606 9358 1658
rect 9358 1606 9368 1658
rect 9392 1606 9422 1658
rect 9422 1606 9434 1658
rect 9434 1606 9448 1658
rect 9472 1606 9486 1658
rect 9486 1606 9498 1658
rect 9498 1606 9528 1658
rect 9552 1606 9562 1658
rect 9562 1606 9608 1658
rect 9312 1604 9368 1606
rect 9392 1604 9448 1606
rect 9472 1604 9528 1606
rect 9552 1604 9608 1606
rect 7762 1114 7818 1116
rect 7842 1114 7898 1116
rect 7922 1114 7978 1116
rect 8002 1114 8058 1116
rect 7762 1062 7808 1114
rect 7808 1062 7818 1114
rect 7842 1062 7872 1114
rect 7872 1062 7884 1114
rect 7884 1062 7898 1114
rect 7922 1062 7936 1114
rect 7936 1062 7948 1114
rect 7948 1062 7978 1114
rect 8002 1062 8012 1114
rect 8012 1062 8058 1114
rect 7762 1060 7818 1062
rect 7842 1060 7898 1062
rect 7922 1060 7978 1062
rect 8002 1060 8058 1062
rect 10862 1114 10918 1116
rect 10942 1114 10998 1116
rect 11022 1114 11078 1116
rect 11102 1114 11158 1116
rect 10862 1062 10908 1114
rect 10908 1062 10918 1114
rect 10942 1062 10972 1114
rect 10972 1062 10984 1114
rect 10984 1062 10998 1114
rect 11022 1062 11036 1114
rect 11036 1062 11048 1114
rect 11048 1062 11078 1114
rect 11102 1062 11112 1114
rect 11112 1062 11158 1114
rect 10862 1060 10918 1062
rect 10942 1060 10998 1062
rect 11022 1060 11078 1062
rect 11102 1060 11158 1062
rect 12412 1658 12468 1660
rect 12492 1658 12548 1660
rect 12572 1658 12628 1660
rect 12652 1658 12708 1660
rect 12412 1606 12458 1658
rect 12458 1606 12468 1658
rect 12492 1606 12522 1658
rect 12522 1606 12534 1658
rect 12534 1606 12548 1658
rect 12572 1606 12586 1658
rect 12586 1606 12598 1658
rect 12598 1606 12628 1658
rect 12652 1606 12662 1658
rect 12662 1606 12708 1658
rect 12412 1604 12468 1606
rect 12492 1604 12548 1606
rect 12572 1604 12628 1606
rect 12652 1604 12708 1606
rect 13962 4378 14018 4380
rect 14042 4378 14098 4380
rect 14122 4378 14178 4380
rect 14202 4378 14258 4380
rect 13962 4326 14008 4378
rect 14008 4326 14018 4378
rect 14042 4326 14072 4378
rect 14072 4326 14084 4378
rect 14084 4326 14098 4378
rect 14122 4326 14136 4378
rect 14136 4326 14148 4378
rect 14148 4326 14178 4378
rect 14202 4326 14212 4378
rect 14212 4326 14258 4378
rect 13962 4324 14018 4326
rect 14042 4324 14098 4326
rect 14122 4324 14178 4326
rect 14202 4324 14258 4326
rect 13962 3290 14018 3292
rect 14042 3290 14098 3292
rect 14122 3290 14178 3292
rect 14202 3290 14258 3292
rect 13962 3238 14008 3290
rect 14008 3238 14018 3290
rect 14042 3238 14072 3290
rect 14072 3238 14084 3290
rect 14084 3238 14098 3290
rect 14122 3238 14136 3290
rect 14136 3238 14148 3290
rect 14148 3238 14178 3290
rect 14202 3238 14212 3290
rect 14212 3238 14258 3290
rect 13962 3236 14018 3238
rect 14042 3236 14098 3238
rect 14122 3236 14178 3238
rect 14202 3236 14258 3238
rect 13962 2202 14018 2204
rect 14042 2202 14098 2204
rect 14122 2202 14178 2204
rect 14202 2202 14258 2204
rect 13962 2150 14008 2202
rect 14008 2150 14018 2202
rect 14042 2150 14072 2202
rect 14072 2150 14084 2202
rect 14084 2150 14098 2202
rect 14122 2150 14136 2202
rect 14136 2150 14148 2202
rect 14148 2150 14178 2202
rect 14202 2150 14212 2202
rect 14212 2150 14258 2202
rect 13962 2148 14018 2150
rect 14042 2148 14098 2150
rect 14122 2148 14178 2150
rect 14202 2148 14258 2150
rect 15512 7098 15568 7100
rect 15592 7098 15648 7100
rect 15672 7098 15728 7100
rect 15752 7098 15808 7100
rect 15512 7046 15558 7098
rect 15558 7046 15568 7098
rect 15592 7046 15622 7098
rect 15622 7046 15634 7098
rect 15634 7046 15648 7098
rect 15672 7046 15686 7098
rect 15686 7046 15698 7098
rect 15698 7046 15728 7098
rect 15752 7046 15762 7098
rect 15762 7046 15808 7098
rect 15512 7044 15568 7046
rect 15592 7044 15648 7046
rect 15672 7044 15728 7046
rect 15752 7044 15808 7046
rect 17062 14170 17118 14172
rect 17142 14170 17198 14172
rect 17222 14170 17278 14172
rect 17302 14170 17358 14172
rect 17062 14118 17108 14170
rect 17108 14118 17118 14170
rect 17142 14118 17172 14170
rect 17172 14118 17184 14170
rect 17184 14118 17198 14170
rect 17222 14118 17236 14170
rect 17236 14118 17248 14170
rect 17248 14118 17278 14170
rect 17302 14118 17312 14170
rect 17312 14118 17358 14170
rect 17062 14116 17118 14118
rect 17142 14116 17198 14118
rect 17222 14116 17278 14118
rect 17302 14116 17358 14118
rect 17062 13082 17118 13084
rect 17142 13082 17198 13084
rect 17222 13082 17278 13084
rect 17302 13082 17358 13084
rect 17062 13030 17108 13082
rect 17108 13030 17118 13082
rect 17142 13030 17172 13082
rect 17172 13030 17184 13082
rect 17184 13030 17198 13082
rect 17222 13030 17236 13082
rect 17236 13030 17248 13082
rect 17248 13030 17278 13082
rect 17302 13030 17312 13082
rect 17312 13030 17358 13082
rect 17062 13028 17118 13030
rect 17142 13028 17198 13030
rect 17222 13028 17278 13030
rect 17302 13028 17358 13030
rect 17062 11994 17118 11996
rect 17142 11994 17198 11996
rect 17222 11994 17278 11996
rect 17302 11994 17358 11996
rect 17062 11942 17108 11994
rect 17108 11942 17118 11994
rect 17142 11942 17172 11994
rect 17172 11942 17184 11994
rect 17184 11942 17198 11994
rect 17222 11942 17236 11994
rect 17236 11942 17248 11994
rect 17248 11942 17278 11994
rect 17302 11942 17312 11994
rect 17312 11942 17358 11994
rect 17062 11940 17118 11942
rect 17142 11940 17198 11942
rect 17222 11940 17278 11942
rect 17302 11940 17358 11942
rect 17062 10906 17118 10908
rect 17142 10906 17198 10908
rect 17222 10906 17278 10908
rect 17302 10906 17358 10908
rect 17062 10854 17108 10906
rect 17108 10854 17118 10906
rect 17142 10854 17172 10906
rect 17172 10854 17184 10906
rect 17184 10854 17198 10906
rect 17222 10854 17236 10906
rect 17236 10854 17248 10906
rect 17248 10854 17278 10906
rect 17302 10854 17312 10906
rect 17312 10854 17358 10906
rect 17062 10852 17118 10854
rect 17142 10852 17198 10854
rect 17222 10852 17278 10854
rect 17302 10852 17358 10854
rect 17062 9818 17118 9820
rect 17142 9818 17198 9820
rect 17222 9818 17278 9820
rect 17302 9818 17358 9820
rect 17062 9766 17108 9818
rect 17108 9766 17118 9818
rect 17142 9766 17172 9818
rect 17172 9766 17184 9818
rect 17184 9766 17198 9818
rect 17222 9766 17236 9818
rect 17236 9766 17248 9818
rect 17248 9766 17278 9818
rect 17302 9766 17312 9818
rect 17312 9766 17358 9818
rect 17062 9764 17118 9766
rect 17142 9764 17198 9766
rect 17222 9764 17278 9766
rect 17302 9764 17358 9766
rect 15512 6010 15568 6012
rect 15592 6010 15648 6012
rect 15672 6010 15728 6012
rect 15752 6010 15808 6012
rect 15512 5958 15558 6010
rect 15558 5958 15568 6010
rect 15592 5958 15622 6010
rect 15622 5958 15634 6010
rect 15634 5958 15648 6010
rect 15672 5958 15686 6010
rect 15686 5958 15698 6010
rect 15698 5958 15728 6010
rect 15752 5958 15762 6010
rect 15762 5958 15808 6010
rect 15512 5956 15568 5958
rect 15592 5956 15648 5958
rect 15672 5956 15728 5958
rect 15752 5956 15808 5958
rect 15512 4922 15568 4924
rect 15592 4922 15648 4924
rect 15672 4922 15728 4924
rect 15752 4922 15808 4924
rect 15512 4870 15558 4922
rect 15558 4870 15568 4922
rect 15592 4870 15622 4922
rect 15622 4870 15634 4922
rect 15634 4870 15648 4922
rect 15672 4870 15686 4922
rect 15686 4870 15698 4922
rect 15698 4870 15728 4922
rect 15752 4870 15762 4922
rect 15762 4870 15808 4922
rect 15512 4868 15568 4870
rect 15592 4868 15648 4870
rect 15672 4868 15728 4870
rect 15752 4868 15808 4870
rect 15512 3834 15568 3836
rect 15592 3834 15648 3836
rect 15672 3834 15728 3836
rect 15752 3834 15808 3836
rect 15512 3782 15558 3834
rect 15558 3782 15568 3834
rect 15592 3782 15622 3834
rect 15622 3782 15634 3834
rect 15634 3782 15648 3834
rect 15672 3782 15686 3834
rect 15686 3782 15698 3834
rect 15698 3782 15728 3834
rect 15752 3782 15762 3834
rect 15762 3782 15808 3834
rect 15512 3780 15568 3782
rect 15592 3780 15648 3782
rect 15672 3780 15728 3782
rect 15752 3780 15808 3782
rect 15512 2746 15568 2748
rect 15592 2746 15648 2748
rect 15672 2746 15728 2748
rect 15752 2746 15808 2748
rect 15512 2694 15558 2746
rect 15558 2694 15568 2746
rect 15592 2694 15622 2746
rect 15622 2694 15634 2746
rect 15634 2694 15648 2746
rect 15672 2694 15686 2746
rect 15686 2694 15698 2746
rect 15698 2694 15728 2746
rect 15752 2694 15762 2746
rect 15762 2694 15808 2746
rect 15512 2692 15568 2694
rect 15592 2692 15648 2694
rect 15672 2692 15728 2694
rect 15752 2692 15808 2694
rect 17062 8730 17118 8732
rect 17142 8730 17198 8732
rect 17222 8730 17278 8732
rect 17302 8730 17358 8732
rect 17062 8678 17108 8730
rect 17108 8678 17118 8730
rect 17142 8678 17172 8730
rect 17172 8678 17184 8730
rect 17184 8678 17198 8730
rect 17222 8678 17236 8730
rect 17236 8678 17248 8730
rect 17248 8678 17278 8730
rect 17302 8678 17312 8730
rect 17312 8678 17358 8730
rect 17062 8676 17118 8678
rect 17142 8676 17198 8678
rect 17222 8676 17278 8678
rect 17302 8676 17358 8678
rect 17062 7642 17118 7644
rect 17142 7642 17198 7644
rect 17222 7642 17278 7644
rect 17302 7642 17358 7644
rect 17062 7590 17108 7642
rect 17108 7590 17118 7642
rect 17142 7590 17172 7642
rect 17172 7590 17184 7642
rect 17184 7590 17198 7642
rect 17222 7590 17236 7642
rect 17236 7590 17248 7642
rect 17248 7590 17278 7642
rect 17302 7590 17312 7642
rect 17312 7590 17358 7642
rect 17062 7588 17118 7590
rect 17142 7588 17198 7590
rect 17222 7588 17278 7590
rect 17302 7588 17358 7590
rect 17062 6554 17118 6556
rect 17142 6554 17198 6556
rect 17222 6554 17278 6556
rect 17302 6554 17358 6556
rect 17062 6502 17108 6554
rect 17108 6502 17118 6554
rect 17142 6502 17172 6554
rect 17172 6502 17184 6554
rect 17184 6502 17198 6554
rect 17222 6502 17236 6554
rect 17236 6502 17248 6554
rect 17248 6502 17278 6554
rect 17302 6502 17312 6554
rect 17312 6502 17358 6554
rect 17062 6500 17118 6502
rect 17142 6500 17198 6502
rect 17222 6500 17278 6502
rect 17302 6500 17358 6502
rect 17062 5466 17118 5468
rect 17142 5466 17198 5468
rect 17222 5466 17278 5468
rect 17302 5466 17358 5468
rect 17062 5414 17108 5466
rect 17108 5414 17118 5466
rect 17142 5414 17172 5466
rect 17172 5414 17184 5466
rect 17184 5414 17198 5466
rect 17222 5414 17236 5466
rect 17236 5414 17248 5466
rect 17248 5414 17278 5466
rect 17302 5414 17312 5466
rect 17312 5414 17358 5466
rect 17062 5412 17118 5414
rect 17142 5412 17198 5414
rect 17222 5412 17278 5414
rect 17302 5412 17358 5414
rect 17062 4378 17118 4380
rect 17142 4378 17198 4380
rect 17222 4378 17278 4380
rect 17302 4378 17358 4380
rect 17062 4326 17108 4378
rect 17108 4326 17118 4378
rect 17142 4326 17172 4378
rect 17172 4326 17184 4378
rect 17184 4326 17198 4378
rect 17222 4326 17236 4378
rect 17236 4326 17248 4378
rect 17248 4326 17278 4378
rect 17302 4326 17312 4378
rect 17312 4326 17358 4378
rect 17062 4324 17118 4326
rect 17142 4324 17198 4326
rect 17222 4324 17278 4326
rect 17302 4324 17358 4326
rect 15512 1658 15568 1660
rect 15592 1658 15648 1660
rect 15672 1658 15728 1660
rect 15752 1658 15808 1660
rect 15512 1606 15558 1658
rect 15558 1606 15568 1658
rect 15592 1606 15622 1658
rect 15622 1606 15634 1658
rect 15634 1606 15648 1658
rect 15672 1606 15686 1658
rect 15686 1606 15698 1658
rect 15698 1606 15728 1658
rect 15752 1606 15762 1658
rect 15762 1606 15808 1658
rect 15512 1604 15568 1606
rect 15592 1604 15648 1606
rect 15672 1604 15728 1606
rect 15752 1604 15808 1606
rect 17062 3290 17118 3292
rect 17142 3290 17198 3292
rect 17222 3290 17278 3292
rect 17302 3290 17358 3292
rect 17062 3238 17108 3290
rect 17108 3238 17118 3290
rect 17142 3238 17172 3290
rect 17172 3238 17184 3290
rect 17184 3238 17198 3290
rect 17222 3238 17236 3290
rect 17236 3238 17248 3290
rect 17248 3238 17278 3290
rect 17302 3238 17312 3290
rect 17312 3238 17358 3290
rect 17062 3236 17118 3238
rect 17142 3236 17198 3238
rect 17222 3236 17278 3238
rect 17302 3236 17358 3238
rect 18612 17978 18668 17980
rect 18692 17978 18748 17980
rect 18772 17978 18828 17980
rect 18852 17978 18908 17980
rect 18612 17926 18658 17978
rect 18658 17926 18668 17978
rect 18692 17926 18722 17978
rect 18722 17926 18734 17978
rect 18734 17926 18748 17978
rect 18772 17926 18786 17978
rect 18786 17926 18798 17978
rect 18798 17926 18828 17978
rect 18852 17926 18862 17978
rect 18862 17926 18908 17978
rect 18612 17924 18668 17926
rect 18692 17924 18748 17926
rect 18772 17924 18828 17926
rect 18852 17924 18908 17926
rect 18612 16890 18668 16892
rect 18692 16890 18748 16892
rect 18772 16890 18828 16892
rect 18852 16890 18908 16892
rect 18612 16838 18658 16890
rect 18658 16838 18668 16890
rect 18692 16838 18722 16890
rect 18722 16838 18734 16890
rect 18734 16838 18748 16890
rect 18772 16838 18786 16890
rect 18786 16838 18798 16890
rect 18798 16838 18828 16890
rect 18852 16838 18862 16890
rect 18862 16838 18908 16890
rect 18612 16836 18668 16838
rect 18692 16836 18748 16838
rect 18772 16836 18828 16838
rect 18852 16836 18908 16838
rect 18612 15802 18668 15804
rect 18692 15802 18748 15804
rect 18772 15802 18828 15804
rect 18852 15802 18908 15804
rect 18612 15750 18658 15802
rect 18658 15750 18668 15802
rect 18692 15750 18722 15802
rect 18722 15750 18734 15802
rect 18734 15750 18748 15802
rect 18772 15750 18786 15802
rect 18786 15750 18798 15802
rect 18798 15750 18828 15802
rect 18852 15750 18862 15802
rect 18862 15750 18908 15802
rect 18612 15748 18668 15750
rect 18692 15748 18748 15750
rect 18772 15748 18828 15750
rect 18852 15748 18908 15750
rect 18612 14714 18668 14716
rect 18692 14714 18748 14716
rect 18772 14714 18828 14716
rect 18852 14714 18908 14716
rect 18612 14662 18658 14714
rect 18658 14662 18668 14714
rect 18692 14662 18722 14714
rect 18722 14662 18734 14714
rect 18734 14662 18748 14714
rect 18772 14662 18786 14714
rect 18786 14662 18798 14714
rect 18798 14662 18828 14714
rect 18852 14662 18862 14714
rect 18862 14662 18908 14714
rect 18612 14660 18668 14662
rect 18692 14660 18748 14662
rect 18772 14660 18828 14662
rect 18852 14660 18908 14662
rect 19062 13640 19118 13696
rect 18612 13626 18668 13628
rect 18692 13626 18748 13628
rect 18772 13626 18828 13628
rect 18852 13626 18908 13628
rect 18612 13574 18658 13626
rect 18658 13574 18668 13626
rect 18692 13574 18722 13626
rect 18722 13574 18734 13626
rect 18734 13574 18748 13626
rect 18772 13574 18786 13626
rect 18786 13574 18798 13626
rect 18798 13574 18828 13626
rect 18852 13574 18862 13626
rect 18862 13574 18908 13626
rect 18612 13572 18668 13574
rect 18692 13572 18748 13574
rect 18772 13572 18828 13574
rect 18852 13572 18908 13574
rect 18612 12538 18668 12540
rect 18692 12538 18748 12540
rect 18772 12538 18828 12540
rect 18852 12538 18908 12540
rect 18612 12486 18658 12538
rect 18658 12486 18668 12538
rect 18692 12486 18722 12538
rect 18722 12486 18734 12538
rect 18734 12486 18748 12538
rect 18772 12486 18786 12538
rect 18786 12486 18798 12538
rect 18798 12486 18828 12538
rect 18852 12486 18862 12538
rect 18862 12486 18908 12538
rect 18612 12484 18668 12486
rect 18692 12484 18748 12486
rect 18772 12484 18828 12486
rect 18852 12484 18908 12486
rect 18612 11450 18668 11452
rect 18692 11450 18748 11452
rect 18772 11450 18828 11452
rect 18852 11450 18908 11452
rect 18612 11398 18658 11450
rect 18658 11398 18668 11450
rect 18692 11398 18722 11450
rect 18722 11398 18734 11450
rect 18734 11398 18748 11450
rect 18772 11398 18786 11450
rect 18786 11398 18798 11450
rect 18798 11398 18828 11450
rect 18852 11398 18862 11450
rect 18862 11398 18908 11450
rect 18612 11396 18668 11398
rect 18692 11396 18748 11398
rect 18772 11396 18828 11398
rect 18852 11396 18908 11398
rect 18418 11192 18474 11248
rect 18612 10362 18668 10364
rect 18692 10362 18748 10364
rect 18772 10362 18828 10364
rect 18852 10362 18908 10364
rect 18612 10310 18658 10362
rect 18658 10310 18668 10362
rect 18692 10310 18722 10362
rect 18722 10310 18734 10362
rect 18734 10310 18748 10362
rect 18772 10310 18786 10362
rect 18786 10310 18798 10362
rect 18798 10310 18828 10362
rect 18852 10310 18862 10362
rect 18862 10310 18908 10362
rect 18612 10308 18668 10310
rect 18692 10308 18748 10310
rect 18772 10308 18828 10310
rect 18852 10308 18908 10310
rect 18612 9274 18668 9276
rect 18692 9274 18748 9276
rect 18772 9274 18828 9276
rect 18852 9274 18908 9276
rect 18612 9222 18658 9274
rect 18658 9222 18668 9274
rect 18692 9222 18722 9274
rect 18722 9222 18734 9274
rect 18734 9222 18748 9274
rect 18772 9222 18786 9274
rect 18786 9222 18798 9274
rect 18798 9222 18828 9274
rect 18852 9222 18862 9274
rect 18862 9222 18908 9274
rect 18612 9220 18668 9222
rect 18692 9220 18748 9222
rect 18772 9220 18828 9222
rect 18852 9220 18908 9222
rect 18418 8744 18474 8800
rect 18612 8186 18668 8188
rect 18692 8186 18748 8188
rect 18772 8186 18828 8188
rect 18852 8186 18908 8188
rect 18612 8134 18658 8186
rect 18658 8134 18668 8186
rect 18692 8134 18722 8186
rect 18722 8134 18734 8186
rect 18734 8134 18748 8186
rect 18772 8134 18786 8186
rect 18786 8134 18798 8186
rect 18798 8134 18828 8186
rect 18852 8134 18862 8186
rect 18862 8134 18908 8186
rect 18612 8132 18668 8134
rect 18692 8132 18748 8134
rect 18772 8132 18828 8134
rect 18852 8132 18908 8134
rect 18612 7098 18668 7100
rect 18692 7098 18748 7100
rect 18772 7098 18828 7100
rect 18852 7098 18908 7100
rect 18612 7046 18658 7098
rect 18658 7046 18668 7098
rect 18692 7046 18722 7098
rect 18722 7046 18734 7098
rect 18734 7046 18748 7098
rect 18772 7046 18786 7098
rect 18786 7046 18798 7098
rect 18798 7046 18828 7098
rect 18852 7046 18862 7098
rect 18862 7046 18908 7098
rect 18612 7044 18668 7046
rect 18692 7044 18748 7046
rect 18772 7044 18828 7046
rect 18852 7044 18908 7046
rect 18418 6296 18474 6352
rect 18612 6010 18668 6012
rect 18692 6010 18748 6012
rect 18772 6010 18828 6012
rect 18852 6010 18908 6012
rect 18612 5958 18658 6010
rect 18658 5958 18668 6010
rect 18692 5958 18722 6010
rect 18722 5958 18734 6010
rect 18734 5958 18748 6010
rect 18772 5958 18786 6010
rect 18786 5958 18798 6010
rect 18798 5958 18828 6010
rect 18852 5958 18862 6010
rect 18862 5958 18908 6010
rect 18612 5956 18668 5958
rect 18692 5956 18748 5958
rect 18772 5956 18828 5958
rect 18852 5956 18908 5958
rect 18612 4922 18668 4924
rect 18692 4922 18748 4924
rect 18772 4922 18828 4924
rect 18852 4922 18908 4924
rect 18612 4870 18658 4922
rect 18658 4870 18668 4922
rect 18692 4870 18722 4922
rect 18722 4870 18734 4922
rect 18734 4870 18748 4922
rect 18772 4870 18786 4922
rect 18786 4870 18798 4922
rect 18798 4870 18828 4922
rect 18852 4870 18862 4922
rect 18862 4870 18908 4922
rect 18612 4868 18668 4870
rect 18692 4868 18748 4870
rect 18772 4868 18828 4870
rect 18852 4868 18908 4870
rect 19062 3848 19118 3904
rect 18612 3834 18668 3836
rect 18692 3834 18748 3836
rect 18772 3834 18828 3836
rect 18852 3834 18908 3836
rect 18612 3782 18658 3834
rect 18658 3782 18668 3834
rect 18692 3782 18722 3834
rect 18722 3782 18734 3834
rect 18734 3782 18748 3834
rect 18772 3782 18786 3834
rect 18786 3782 18798 3834
rect 18798 3782 18828 3834
rect 18852 3782 18862 3834
rect 18862 3782 18908 3834
rect 18612 3780 18668 3782
rect 18692 3780 18748 3782
rect 18772 3780 18828 3782
rect 18852 3780 18908 3782
rect 18612 2746 18668 2748
rect 18692 2746 18748 2748
rect 18772 2746 18828 2748
rect 18852 2746 18908 2748
rect 18612 2694 18658 2746
rect 18658 2694 18668 2746
rect 18692 2694 18722 2746
rect 18722 2694 18734 2746
rect 18734 2694 18748 2746
rect 18772 2694 18786 2746
rect 18786 2694 18798 2746
rect 18798 2694 18828 2746
rect 18852 2694 18862 2746
rect 18862 2694 18908 2746
rect 18612 2692 18668 2694
rect 18692 2692 18748 2694
rect 18772 2692 18828 2694
rect 18852 2692 18908 2694
rect 17062 2202 17118 2204
rect 17142 2202 17198 2204
rect 17222 2202 17278 2204
rect 17302 2202 17358 2204
rect 17062 2150 17108 2202
rect 17108 2150 17118 2202
rect 17142 2150 17172 2202
rect 17172 2150 17184 2202
rect 17184 2150 17198 2202
rect 17222 2150 17236 2202
rect 17236 2150 17248 2202
rect 17248 2150 17278 2202
rect 17302 2150 17312 2202
rect 17312 2150 17358 2202
rect 17062 2148 17118 2150
rect 17142 2148 17198 2150
rect 17222 2148 17278 2150
rect 17302 2148 17358 2150
rect 13962 1114 14018 1116
rect 14042 1114 14098 1116
rect 14122 1114 14178 1116
rect 14202 1114 14258 1116
rect 13962 1062 14008 1114
rect 14008 1062 14018 1114
rect 14042 1062 14072 1114
rect 14072 1062 14084 1114
rect 14084 1062 14098 1114
rect 14122 1062 14136 1114
rect 14136 1062 14148 1114
rect 14148 1062 14178 1114
rect 14202 1062 14212 1114
rect 14212 1062 14258 1114
rect 13962 1060 14018 1062
rect 14042 1060 14098 1062
rect 14122 1060 14178 1062
rect 14202 1060 14258 1062
rect 17062 1114 17118 1116
rect 17142 1114 17198 1116
rect 17222 1114 17278 1116
rect 17302 1114 17358 1116
rect 17062 1062 17108 1114
rect 17108 1062 17118 1114
rect 17142 1062 17172 1114
rect 17172 1062 17184 1114
rect 17184 1062 17198 1114
rect 17222 1062 17236 1114
rect 17236 1062 17248 1114
rect 17248 1062 17278 1114
rect 17302 1062 17312 1114
rect 17312 1062 17358 1114
rect 17062 1060 17118 1062
rect 17142 1060 17198 1062
rect 17222 1060 17278 1062
rect 17302 1060 17358 1062
rect 18612 1658 18668 1660
rect 18692 1658 18748 1660
rect 18772 1658 18828 1660
rect 18852 1658 18908 1660
rect 18612 1606 18658 1658
rect 18658 1606 18668 1658
rect 18692 1606 18722 1658
rect 18722 1606 18734 1658
rect 18734 1606 18748 1658
rect 18772 1606 18786 1658
rect 18786 1606 18798 1658
rect 18798 1606 18828 1658
rect 18852 1606 18862 1658
rect 18862 1606 18908 1658
rect 18612 1604 18668 1606
rect 18692 1604 18748 1606
rect 18772 1604 18828 1606
rect 18852 1604 18908 1606
rect 18418 1400 18474 1456
rect 3112 570 3168 572
rect 3192 570 3248 572
rect 3272 570 3328 572
rect 3352 570 3408 572
rect 3112 518 3158 570
rect 3158 518 3168 570
rect 3192 518 3222 570
rect 3222 518 3234 570
rect 3234 518 3248 570
rect 3272 518 3286 570
rect 3286 518 3298 570
rect 3298 518 3328 570
rect 3352 518 3362 570
rect 3362 518 3408 570
rect 3112 516 3168 518
rect 3192 516 3248 518
rect 3272 516 3328 518
rect 3352 516 3408 518
rect 6212 570 6268 572
rect 6292 570 6348 572
rect 6372 570 6428 572
rect 6452 570 6508 572
rect 6212 518 6258 570
rect 6258 518 6268 570
rect 6292 518 6322 570
rect 6322 518 6334 570
rect 6334 518 6348 570
rect 6372 518 6386 570
rect 6386 518 6398 570
rect 6398 518 6428 570
rect 6452 518 6462 570
rect 6462 518 6508 570
rect 6212 516 6268 518
rect 6292 516 6348 518
rect 6372 516 6428 518
rect 6452 516 6508 518
rect 9312 570 9368 572
rect 9392 570 9448 572
rect 9472 570 9528 572
rect 9552 570 9608 572
rect 9312 518 9358 570
rect 9358 518 9368 570
rect 9392 518 9422 570
rect 9422 518 9434 570
rect 9434 518 9448 570
rect 9472 518 9486 570
rect 9486 518 9498 570
rect 9498 518 9528 570
rect 9552 518 9562 570
rect 9562 518 9608 570
rect 9312 516 9368 518
rect 9392 516 9448 518
rect 9472 516 9528 518
rect 9552 516 9608 518
rect 12412 570 12468 572
rect 12492 570 12548 572
rect 12572 570 12628 572
rect 12652 570 12708 572
rect 12412 518 12458 570
rect 12458 518 12468 570
rect 12492 518 12522 570
rect 12522 518 12534 570
rect 12534 518 12548 570
rect 12572 518 12586 570
rect 12586 518 12598 570
rect 12598 518 12628 570
rect 12652 518 12662 570
rect 12662 518 12708 570
rect 12412 516 12468 518
rect 12492 516 12548 518
rect 12572 516 12628 518
rect 12652 516 12708 518
rect 15512 570 15568 572
rect 15592 570 15648 572
rect 15672 570 15728 572
rect 15752 570 15808 572
rect 15512 518 15558 570
rect 15558 518 15568 570
rect 15592 518 15622 570
rect 15622 518 15634 570
rect 15634 518 15648 570
rect 15672 518 15686 570
rect 15686 518 15698 570
rect 15698 518 15728 570
rect 15752 518 15762 570
rect 15762 518 15808 570
rect 15512 516 15568 518
rect 15592 516 15648 518
rect 15672 516 15728 518
rect 15752 516 15808 518
rect 18612 570 18668 572
rect 18692 570 18748 572
rect 18772 570 18828 572
rect 18852 570 18908 572
rect 18612 518 18658 570
rect 18658 518 18668 570
rect 18692 518 18722 570
rect 18722 518 18734 570
rect 18734 518 18748 570
rect 18772 518 18786 570
rect 18786 518 18798 570
rect 18798 518 18828 570
rect 18852 518 18862 570
rect 18862 518 18908 570
rect 18612 516 18668 518
rect 18692 516 18748 518
rect 18772 516 18828 518
rect 18852 516 18908 518
<< metal3 >>
rect 18413 18594 18479 18597
rect 19200 18594 20000 18624
rect 18413 18592 20000 18594
rect 18413 18536 18418 18592
rect 18474 18536 20000 18592
rect 18413 18534 20000 18536
rect 18413 18531 18479 18534
rect 1552 18528 1868 18529
rect 1552 18464 1558 18528
rect 1622 18464 1638 18528
rect 1702 18464 1718 18528
rect 1782 18464 1798 18528
rect 1862 18464 1868 18528
rect 1552 18463 1868 18464
rect 4652 18528 4968 18529
rect 4652 18464 4658 18528
rect 4722 18464 4738 18528
rect 4802 18464 4818 18528
rect 4882 18464 4898 18528
rect 4962 18464 4968 18528
rect 4652 18463 4968 18464
rect 7752 18528 8068 18529
rect 7752 18464 7758 18528
rect 7822 18464 7838 18528
rect 7902 18464 7918 18528
rect 7982 18464 7998 18528
rect 8062 18464 8068 18528
rect 7752 18463 8068 18464
rect 10852 18528 11168 18529
rect 10852 18464 10858 18528
rect 10922 18464 10938 18528
rect 11002 18464 11018 18528
rect 11082 18464 11098 18528
rect 11162 18464 11168 18528
rect 10852 18463 11168 18464
rect 13952 18528 14268 18529
rect 13952 18464 13958 18528
rect 14022 18464 14038 18528
rect 14102 18464 14118 18528
rect 14182 18464 14198 18528
rect 14262 18464 14268 18528
rect 13952 18463 14268 18464
rect 17052 18528 17368 18529
rect 17052 18464 17058 18528
rect 17122 18464 17138 18528
rect 17202 18464 17218 18528
rect 17282 18464 17298 18528
rect 17362 18464 17368 18528
rect 19200 18504 20000 18534
rect 17052 18463 17368 18464
rect 3102 17984 3418 17985
rect 3102 17920 3108 17984
rect 3172 17920 3188 17984
rect 3252 17920 3268 17984
rect 3332 17920 3348 17984
rect 3412 17920 3418 17984
rect 3102 17919 3418 17920
rect 6202 17984 6518 17985
rect 6202 17920 6208 17984
rect 6272 17920 6288 17984
rect 6352 17920 6368 17984
rect 6432 17920 6448 17984
rect 6512 17920 6518 17984
rect 6202 17919 6518 17920
rect 9302 17984 9618 17985
rect 9302 17920 9308 17984
rect 9372 17920 9388 17984
rect 9452 17920 9468 17984
rect 9532 17920 9548 17984
rect 9612 17920 9618 17984
rect 9302 17919 9618 17920
rect 12402 17984 12718 17985
rect 12402 17920 12408 17984
rect 12472 17920 12488 17984
rect 12552 17920 12568 17984
rect 12632 17920 12648 17984
rect 12712 17920 12718 17984
rect 12402 17919 12718 17920
rect 15502 17984 15818 17985
rect 15502 17920 15508 17984
rect 15572 17920 15588 17984
rect 15652 17920 15668 17984
rect 15732 17920 15748 17984
rect 15812 17920 15818 17984
rect 15502 17919 15818 17920
rect 18602 17984 18918 17985
rect 18602 17920 18608 17984
rect 18672 17920 18688 17984
rect 18752 17920 18768 17984
rect 18832 17920 18848 17984
rect 18912 17920 18918 17984
rect 18602 17919 18918 17920
rect 1552 17440 1868 17441
rect 1552 17376 1558 17440
rect 1622 17376 1638 17440
rect 1702 17376 1718 17440
rect 1782 17376 1798 17440
rect 1862 17376 1868 17440
rect 1552 17375 1868 17376
rect 4652 17440 4968 17441
rect 4652 17376 4658 17440
rect 4722 17376 4738 17440
rect 4802 17376 4818 17440
rect 4882 17376 4898 17440
rect 4962 17376 4968 17440
rect 4652 17375 4968 17376
rect 7752 17440 8068 17441
rect 7752 17376 7758 17440
rect 7822 17376 7838 17440
rect 7902 17376 7918 17440
rect 7982 17376 7998 17440
rect 8062 17376 8068 17440
rect 7752 17375 8068 17376
rect 10852 17440 11168 17441
rect 10852 17376 10858 17440
rect 10922 17376 10938 17440
rect 11002 17376 11018 17440
rect 11082 17376 11098 17440
rect 11162 17376 11168 17440
rect 10852 17375 11168 17376
rect 13952 17440 14268 17441
rect 13952 17376 13958 17440
rect 14022 17376 14038 17440
rect 14102 17376 14118 17440
rect 14182 17376 14198 17440
rect 14262 17376 14268 17440
rect 13952 17375 14268 17376
rect 17052 17440 17368 17441
rect 17052 17376 17058 17440
rect 17122 17376 17138 17440
rect 17202 17376 17218 17440
rect 17282 17376 17298 17440
rect 17362 17376 17368 17440
rect 17052 17375 17368 17376
rect 3102 16896 3418 16897
rect 3102 16832 3108 16896
rect 3172 16832 3188 16896
rect 3252 16832 3268 16896
rect 3332 16832 3348 16896
rect 3412 16832 3418 16896
rect 3102 16831 3418 16832
rect 6202 16896 6518 16897
rect 6202 16832 6208 16896
rect 6272 16832 6288 16896
rect 6352 16832 6368 16896
rect 6432 16832 6448 16896
rect 6512 16832 6518 16896
rect 6202 16831 6518 16832
rect 9302 16896 9618 16897
rect 9302 16832 9308 16896
rect 9372 16832 9388 16896
rect 9452 16832 9468 16896
rect 9532 16832 9548 16896
rect 9612 16832 9618 16896
rect 9302 16831 9618 16832
rect 12402 16896 12718 16897
rect 12402 16832 12408 16896
rect 12472 16832 12488 16896
rect 12552 16832 12568 16896
rect 12632 16832 12648 16896
rect 12712 16832 12718 16896
rect 12402 16831 12718 16832
rect 15502 16896 15818 16897
rect 15502 16832 15508 16896
rect 15572 16832 15588 16896
rect 15652 16832 15668 16896
rect 15732 16832 15748 16896
rect 15812 16832 15818 16896
rect 15502 16831 15818 16832
rect 18602 16896 18918 16897
rect 18602 16832 18608 16896
rect 18672 16832 18688 16896
rect 18752 16832 18768 16896
rect 18832 16832 18848 16896
rect 18912 16832 18918 16896
rect 18602 16831 18918 16832
rect 13353 16690 13419 16693
rect 14273 16690 14339 16693
rect 14733 16690 14799 16693
rect 16297 16690 16363 16693
rect 13353 16688 16363 16690
rect 13353 16632 13358 16688
rect 13414 16632 14278 16688
rect 14334 16632 14738 16688
rect 14794 16632 16302 16688
rect 16358 16632 16363 16688
rect 13353 16630 16363 16632
rect 13353 16627 13419 16630
rect 14273 16627 14339 16630
rect 14733 16627 14799 16630
rect 16297 16627 16363 16630
rect 1552 16352 1868 16353
rect 1552 16288 1558 16352
rect 1622 16288 1638 16352
rect 1702 16288 1718 16352
rect 1782 16288 1798 16352
rect 1862 16288 1868 16352
rect 1552 16287 1868 16288
rect 4652 16352 4968 16353
rect 4652 16288 4658 16352
rect 4722 16288 4738 16352
rect 4802 16288 4818 16352
rect 4882 16288 4898 16352
rect 4962 16288 4968 16352
rect 4652 16287 4968 16288
rect 7752 16352 8068 16353
rect 7752 16288 7758 16352
rect 7822 16288 7838 16352
rect 7902 16288 7918 16352
rect 7982 16288 7998 16352
rect 8062 16288 8068 16352
rect 7752 16287 8068 16288
rect 10852 16352 11168 16353
rect 10852 16288 10858 16352
rect 10922 16288 10938 16352
rect 11002 16288 11018 16352
rect 11082 16288 11098 16352
rect 11162 16288 11168 16352
rect 10852 16287 11168 16288
rect 13952 16352 14268 16353
rect 13952 16288 13958 16352
rect 14022 16288 14038 16352
rect 14102 16288 14118 16352
rect 14182 16288 14198 16352
rect 14262 16288 14268 16352
rect 13952 16287 14268 16288
rect 17052 16352 17368 16353
rect 17052 16288 17058 16352
rect 17122 16288 17138 16352
rect 17202 16288 17218 16352
rect 17282 16288 17298 16352
rect 17362 16288 17368 16352
rect 17052 16287 17368 16288
rect 18413 16146 18479 16149
rect 19200 16146 20000 16176
rect 18413 16144 20000 16146
rect 18413 16088 18418 16144
rect 18474 16088 20000 16144
rect 18413 16086 20000 16088
rect 18413 16083 18479 16086
rect 19200 16056 20000 16086
rect 3102 15808 3418 15809
rect 3102 15744 3108 15808
rect 3172 15744 3188 15808
rect 3252 15744 3268 15808
rect 3332 15744 3348 15808
rect 3412 15744 3418 15808
rect 3102 15743 3418 15744
rect 6202 15808 6518 15809
rect 6202 15744 6208 15808
rect 6272 15744 6288 15808
rect 6352 15744 6368 15808
rect 6432 15744 6448 15808
rect 6512 15744 6518 15808
rect 6202 15743 6518 15744
rect 9302 15808 9618 15809
rect 9302 15744 9308 15808
rect 9372 15744 9388 15808
rect 9452 15744 9468 15808
rect 9532 15744 9548 15808
rect 9612 15744 9618 15808
rect 9302 15743 9618 15744
rect 12402 15808 12718 15809
rect 12402 15744 12408 15808
rect 12472 15744 12488 15808
rect 12552 15744 12568 15808
rect 12632 15744 12648 15808
rect 12712 15744 12718 15808
rect 12402 15743 12718 15744
rect 15502 15808 15818 15809
rect 15502 15744 15508 15808
rect 15572 15744 15588 15808
rect 15652 15744 15668 15808
rect 15732 15744 15748 15808
rect 15812 15744 15818 15808
rect 15502 15743 15818 15744
rect 18602 15808 18918 15809
rect 18602 15744 18608 15808
rect 18672 15744 18688 15808
rect 18752 15744 18768 15808
rect 18832 15744 18848 15808
rect 18912 15744 18918 15808
rect 18602 15743 18918 15744
rect 1552 15264 1868 15265
rect 1552 15200 1558 15264
rect 1622 15200 1638 15264
rect 1702 15200 1718 15264
rect 1782 15200 1798 15264
rect 1862 15200 1868 15264
rect 1552 15199 1868 15200
rect 4652 15264 4968 15265
rect 4652 15200 4658 15264
rect 4722 15200 4738 15264
rect 4802 15200 4818 15264
rect 4882 15200 4898 15264
rect 4962 15200 4968 15264
rect 4652 15199 4968 15200
rect 7752 15264 8068 15265
rect 7752 15200 7758 15264
rect 7822 15200 7838 15264
rect 7902 15200 7918 15264
rect 7982 15200 7998 15264
rect 8062 15200 8068 15264
rect 7752 15199 8068 15200
rect 10852 15264 11168 15265
rect 10852 15200 10858 15264
rect 10922 15200 10938 15264
rect 11002 15200 11018 15264
rect 11082 15200 11098 15264
rect 11162 15200 11168 15264
rect 10852 15199 11168 15200
rect 13952 15264 14268 15265
rect 13952 15200 13958 15264
rect 14022 15200 14038 15264
rect 14102 15200 14118 15264
rect 14182 15200 14198 15264
rect 14262 15200 14268 15264
rect 13952 15199 14268 15200
rect 17052 15264 17368 15265
rect 17052 15200 17058 15264
rect 17122 15200 17138 15264
rect 17202 15200 17218 15264
rect 17282 15200 17298 15264
rect 17362 15200 17368 15264
rect 17052 15199 17368 15200
rect 3102 14720 3418 14721
rect 3102 14656 3108 14720
rect 3172 14656 3188 14720
rect 3252 14656 3268 14720
rect 3332 14656 3348 14720
rect 3412 14656 3418 14720
rect 3102 14655 3418 14656
rect 6202 14720 6518 14721
rect 6202 14656 6208 14720
rect 6272 14656 6288 14720
rect 6352 14656 6368 14720
rect 6432 14656 6448 14720
rect 6512 14656 6518 14720
rect 6202 14655 6518 14656
rect 9302 14720 9618 14721
rect 9302 14656 9308 14720
rect 9372 14656 9388 14720
rect 9452 14656 9468 14720
rect 9532 14656 9548 14720
rect 9612 14656 9618 14720
rect 9302 14655 9618 14656
rect 12402 14720 12718 14721
rect 12402 14656 12408 14720
rect 12472 14656 12488 14720
rect 12552 14656 12568 14720
rect 12632 14656 12648 14720
rect 12712 14656 12718 14720
rect 12402 14655 12718 14656
rect 15502 14720 15818 14721
rect 15502 14656 15508 14720
rect 15572 14656 15588 14720
rect 15652 14656 15668 14720
rect 15732 14656 15748 14720
rect 15812 14656 15818 14720
rect 15502 14655 15818 14656
rect 18602 14720 18918 14721
rect 18602 14656 18608 14720
rect 18672 14656 18688 14720
rect 18752 14656 18768 14720
rect 18832 14656 18848 14720
rect 18912 14656 18918 14720
rect 18602 14655 18918 14656
rect 1552 14176 1868 14177
rect 1552 14112 1558 14176
rect 1622 14112 1638 14176
rect 1702 14112 1718 14176
rect 1782 14112 1798 14176
rect 1862 14112 1868 14176
rect 1552 14111 1868 14112
rect 4652 14176 4968 14177
rect 4652 14112 4658 14176
rect 4722 14112 4738 14176
rect 4802 14112 4818 14176
rect 4882 14112 4898 14176
rect 4962 14112 4968 14176
rect 4652 14111 4968 14112
rect 7752 14176 8068 14177
rect 7752 14112 7758 14176
rect 7822 14112 7838 14176
rect 7902 14112 7918 14176
rect 7982 14112 7998 14176
rect 8062 14112 8068 14176
rect 7752 14111 8068 14112
rect 10852 14176 11168 14177
rect 10852 14112 10858 14176
rect 10922 14112 10938 14176
rect 11002 14112 11018 14176
rect 11082 14112 11098 14176
rect 11162 14112 11168 14176
rect 10852 14111 11168 14112
rect 13952 14176 14268 14177
rect 13952 14112 13958 14176
rect 14022 14112 14038 14176
rect 14102 14112 14118 14176
rect 14182 14112 14198 14176
rect 14262 14112 14268 14176
rect 13952 14111 14268 14112
rect 17052 14176 17368 14177
rect 17052 14112 17058 14176
rect 17122 14112 17138 14176
rect 17202 14112 17218 14176
rect 17282 14112 17298 14176
rect 17362 14112 17368 14176
rect 17052 14111 17368 14112
rect 19057 13698 19123 13701
rect 19200 13698 20000 13728
rect 19057 13696 20000 13698
rect 19057 13640 19062 13696
rect 19118 13640 20000 13696
rect 19057 13638 20000 13640
rect 19057 13635 19123 13638
rect 3102 13632 3418 13633
rect 3102 13568 3108 13632
rect 3172 13568 3188 13632
rect 3252 13568 3268 13632
rect 3332 13568 3348 13632
rect 3412 13568 3418 13632
rect 3102 13567 3418 13568
rect 6202 13632 6518 13633
rect 6202 13568 6208 13632
rect 6272 13568 6288 13632
rect 6352 13568 6368 13632
rect 6432 13568 6448 13632
rect 6512 13568 6518 13632
rect 6202 13567 6518 13568
rect 9302 13632 9618 13633
rect 9302 13568 9308 13632
rect 9372 13568 9388 13632
rect 9452 13568 9468 13632
rect 9532 13568 9548 13632
rect 9612 13568 9618 13632
rect 9302 13567 9618 13568
rect 12402 13632 12718 13633
rect 12402 13568 12408 13632
rect 12472 13568 12488 13632
rect 12552 13568 12568 13632
rect 12632 13568 12648 13632
rect 12712 13568 12718 13632
rect 12402 13567 12718 13568
rect 15502 13632 15818 13633
rect 15502 13568 15508 13632
rect 15572 13568 15588 13632
rect 15652 13568 15668 13632
rect 15732 13568 15748 13632
rect 15812 13568 15818 13632
rect 15502 13567 15818 13568
rect 18602 13632 18918 13633
rect 18602 13568 18608 13632
rect 18672 13568 18688 13632
rect 18752 13568 18768 13632
rect 18832 13568 18848 13632
rect 18912 13568 18918 13632
rect 19200 13608 20000 13638
rect 18602 13567 18918 13568
rect 1552 13088 1868 13089
rect 1552 13024 1558 13088
rect 1622 13024 1638 13088
rect 1702 13024 1718 13088
rect 1782 13024 1798 13088
rect 1862 13024 1868 13088
rect 1552 13023 1868 13024
rect 4652 13088 4968 13089
rect 4652 13024 4658 13088
rect 4722 13024 4738 13088
rect 4802 13024 4818 13088
rect 4882 13024 4898 13088
rect 4962 13024 4968 13088
rect 4652 13023 4968 13024
rect 7752 13088 8068 13089
rect 7752 13024 7758 13088
rect 7822 13024 7838 13088
rect 7902 13024 7918 13088
rect 7982 13024 7998 13088
rect 8062 13024 8068 13088
rect 7752 13023 8068 13024
rect 10852 13088 11168 13089
rect 10852 13024 10858 13088
rect 10922 13024 10938 13088
rect 11002 13024 11018 13088
rect 11082 13024 11098 13088
rect 11162 13024 11168 13088
rect 10852 13023 11168 13024
rect 13952 13088 14268 13089
rect 13952 13024 13958 13088
rect 14022 13024 14038 13088
rect 14102 13024 14118 13088
rect 14182 13024 14198 13088
rect 14262 13024 14268 13088
rect 13952 13023 14268 13024
rect 17052 13088 17368 13089
rect 17052 13024 17058 13088
rect 17122 13024 17138 13088
rect 17202 13024 17218 13088
rect 17282 13024 17298 13088
rect 17362 13024 17368 13088
rect 17052 13023 17368 13024
rect 3102 12544 3418 12545
rect 3102 12480 3108 12544
rect 3172 12480 3188 12544
rect 3252 12480 3268 12544
rect 3332 12480 3348 12544
rect 3412 12480 3418 12544
rect 3102 12479 3418 12480
rect 6202 12544 6518 12545
rect 6202 12480 6208 12544
rect 6272 12480 6288 12544
rect 6352 12480 6368 12544
rect 6432 12480 6448 12544
rect 6512 12480 6518 12544
rect 6202 12479 6518 12480
rect 9302 12544 9618 12545
rect 9302 12480 9308 12544
rect 9372 12480 9388 12544
rect 9452 12480 9468 12544
rect 9532 12480 9548 12544
rect 9612 12480 9618 12544
rect 9302 12479 9618 12480
rect 12402 12544 12718 12545
rect 12402 12480 12408 12544
rect 12472 12480 12488 12544
rect 12552 12480 12568 12544
rect 12632 12480 12648 12544
rect 12712 12480 12718 12544
rect 12402 12479 12718 12480
rect 15502 12544 15818 12545
rect 15502 12480 15508 12544
rect 15572 12480 15588 12544
rect 15652 12480 15668 12544
rect 15732 12480 15748 12544
rect 15812 12480 15818 12544
rect 15502 12479 15818 12480
rect 18602 12544 18918 12545
rect 18602 12480 18608 12544
rect 18672 12480 18688 12544
rect 18752 12480 18768 12544
rect 18832 12480 18848 12544
rect 18912 12480 18918 12544
rect 18602 12479 18918 12480
rect 1552 12000 1868 12001
rect 1552 11936 1558 12000
rect 1622 11936 1638 12000
rect 1702 11936 1718 12000
rect 1782 11936 1798 12000
rect 1862 11936 1868 12000
rect 1552 11935 1868 11936
rect 4652 12000 4968 12001
rect 4652 11936 4658 12000
rect 4722 11936 4738 12000
rect 4802 11936 4818 12000
rect 4882 11936 4898 12000
rect 4962 11936 4968 12000
rect 4652 11935 4968 11936
rect 7752 12000 8068 12001
rect 7752 11936 7758 12000
rect 7822 11936 7838 12000
rect 7902 11936 7918 12000
rect 7982 11936 7998 12000
rect 8062 11936 8068 12000
rect 7752 11935 8068 11936
rect 10852 12000 11168 12001
rect 10852 11936 10858 12000
rect 10922 11936 10938 12000
rect 11002 11936 11018 12000
rect 11082 11936 11098 12000
rect 11162 11936 11168 12000
rect 10852 11935 11168 11936
rect 13952 12000 14268 12001
rect 13952 11936 13958 12000
rect 14022 11936 14038 12000
rect 14102 11936 14118 12000
rect 14182 11936 14198 12000
rect 14262 11936 14268 12000
rect 13952 11935 14268 11936
rect 17052 12000 17368 12001
rect 17052 11936 17058 12000
rect 17122 11936 17138 12000
rect 17202 11936 17218 12000
rect 17282 11936 17298 12000
rect 17362 11936 17368 12000
rect 17052 11935 17368 11936
rect 3102 11456 3418 11457
rect 3102 11392 3108 11456
rect 3172 11392 3188 11456
rect 3252 11392 3268 11456
rect 3332 11392 3348 11456
rect 3412 11392 3418 11456
rect 3102 11391 3418 11392
rect 6202 11456 6518 11457
rect 6202 11392 6208 11456
rect 6272 11392 6288 11456
rect 6352 11392 6368 11456
rect 6432 11392 6448 11456
rect 6512 11392 6518 11456
rect 6202 11391 6518 11392
rect 9302 11456 9618 11457
rect 9302 11392 9308 11456
rect 9372 11392 9388 11456
rect 9452 11392 9468 11456
rect 9532 11392 9548 11456
rect 9612 11392 9618 11456
rect 9302 11391 9618 11392
rect 12402 11456 12718 11457
rect 12402 11392 12408 11456
rect 12472 11392 12488 11456
rect 12552 11392 12568 11456
rect 12632 11392 12648 11456
rect 12712 11392 12718 11456
rect 12402 11391 12718 11392
rect 15502 11456 15818 11457
rect 15502 11392 15508 11456
rect 15572 11392 15588 11456
rect 15652 11392 15668 11456
rect 15732 11392 15748 11456
rect 15812 11392 15818 11456
rect 15502 11391 15818 11392
rect 18602 11456 18918 11457
rect 18602 11392 18608 11456
rect 18672 11392 18688 11456
rect 18752 11392 18768 11456
rect 18832 11392 18848 11456
rect 18912 11392 18918 11456
rect 18602 11391 18918 11392
rect 18413 11250 18479 11253
rect 19200 11250 20000 11280
rect 18413 11248 20000 11250
rect 18413 11192 18418 11248
rect 18474 11192 20000 11248
rect 18413 11190 20000 11192
rect 18413 11187 18479 11190
rect 19200 11160 20000 11190
rect 1552 10912 1868 10913
rect 1552 10848 1558 10912
rect 1622 10848 1638 10912
rect 1702 10848 1718 10912
rect 1782 10848 1798 10912
rect 1862 10848 1868 10912
rect 1552 10847 1868 10848
rect 4652 10912 4968 10913
rect 4652 10848 4658 10912
rect 4722 10848 4738 10912
rect 4802 10848 4818 10912
rect 4882 10848 4898 10912
rect 4962 10848 4968 10912
rect 4652 10847 4968 10848
rect 7752 10912 8068 10913
rect 7752 10848 7758 10912
rect 7822 10848 7838 10912
rect 7902 10848 7918 10912
rect 7982 10848 7998 10912
rect 8062 10848 8068 10912
rect 7752 10847 8068 10848
rect 10852 10912 11168 10913
rect 10852 10848 10858 10912
rect 10922 10848 10938 10912
rect 11002 10848 11018 10912
rect 11082 10848 11098 10912
rect 11162 10848 11168 10912
rect 10852 10847 11168 10848
rect 13952 10912 14268 10913
rect 13952 10848 13958 10912
rect 14022 10848 14038 10912
rect 14102 10848 14118 10912
rect 14182 10848 14198 10912
rect 14262 10848 14268 10912
rect 13952 10847 14268 10848
rect 17052 10912 17368 10913
rect 17052 10848 17058 10912
rect 17122 10848 17138 10912
rect 17202 10848 17218 10912
rect 17282 10848 17298 10912
rect 17362 10848 17368 10912
rect 17052 10847 17368 10848
rect 3102 10368 3418 10369
rect 3102 10304 3108 10368
rect 3172 10304 3188 10368
rect 3252 10304 3268 10368
rect 3332 10304 3348 10368
rect 3412 10304 3418 10368
rect 3102 10303 3418 10304
rect 6202 10368 6518 10369
rect 6202 10304 6208 10368
rect 6272 10304 6288 10368
rect 6352 10304 6368 10368
rect 6432 10304 6448 10368
rect 6512 10304 6518 10368
rect 6202 10303 6518 10304
rect 9302 10368 9618 10369
rect 9302 10304 9308 10368
rect 9372 10304 9388 10368
rect 9452 10304 9468 10368
rect 9532 10304 9548 10368
rect 9612 10304 9618 10368
rect 9302 10303 9618 10304
rect 12402 10368 12718 10369
rect 12402 10304 12408 10368
rect 12472 10304 12488 10368
rect 12552 10304 12568 10368
rect 12632 10304 12648 10368
rect 12712 10304 12718 10368
rect 12402 10303 12718 10304
rect 15502 10368 15818 10369
rect 15502 10304 15508 10368
rect 15572 10304 15588 10368
rect 15652 10304 15668 10368
rect 15732 10304 15748 10368
rect 15812 10304 15818 10368
rect 15502 10303 15818 10304
rect 18602 10368 18918 10369
rect 18602 10304 18608 10368
rect 18672 10304 18688 10368
rect 18752 10304 18768 10368
rect 18832 10304 18848 10368
rect 18912 10304 18918 10368
rect 18602 10303 18918 10304
rect 0 10026 800 10056
rect 933 10026 999 10029
rect 0 10024 999 10026
rect 0 9968 938 10024
rect 994 9968 999 10024
rect 0 9966 999 9968
rect 0 9936 800 9966
rect 933 9963 999 9966
rect 1552 9824 1868 9825
rect 1552 9760 1558 9824
rect 1622 9760 1638 9824
rect 1702 9760 1718 9824
rect 1782 9760 1798 9824
rect 1862 9760 1868 9824
rect 1552 9759 1868 9760
rect 4652 9824 4968 9825
rect 4652 9760 4658 9824
rect 4722 9760 4738 9824
rect 4802 9760 4818 9824
rect 4882 9760 4898 9824
rect 4962 9760 4968 9824
rect 4652 9759 4968 9760
rect 7752 9824 8068 9825
rect 7752 9760 7758 9824
rect 7822 9760 7838 9824
rect 7902 9760 7918 9824
rect 7982 9760 7998 9824
rect 8062 9760 8068 9824
rect 7752 9759 8068 9760
rect 10852 9824 11168 9825
rect 10852 9760 10858 9824
rect 10922 9760 10938 9824
rect 11002 9760 11018 9824
rect 11082 9760 11098 9824
rect 11162 9760 11168 9824
rect 10852 9759 11168 9760
rect 13952 9824 14268 9825
rect 13952 9760 13958 9824
rect 14022 9760 14038 9824
rect 14102 9760 14118 9824
rect 14182 9760 14198 9824
rect 14262 9760 14268 9824
rect 13952 9759 14268 9760
rect 17052 9824 17368 9825
rect 17052 9760 17058 9824
rect 17122 9760 17138 9824
rect 17202 9760 17218 9824
rect 17282 9760 17298 9824
rect 17362 9760 17368 9824
rect 17052 9759 17368 9760
rect 3102 9280 3418 9281
rect 3102 9216 3108 9280
rect 3172 9216 3188 9280
rect 3252 9216 3268 9280
rect 3332 9216 3348 9280
rect 3412 9216 3418 9280
rect 3102 9215 3418 9216
rect 6202 9280 6518 9281
rect 6202 9216 6208 9280
rect 6272 9216 6288 9280
rect 6352 9216 6368 9280
rect 6432 9216 6448 9280
rect 6512 9216 6518 9280
rect 6202 9215 6518 9216
rect 9302 9280 9618 9281
rect 9302 9216 9308 9280
rect 9372 9216 9388 9280
rect 9452 9216 9468 9280
rect 9532 9216 9548 9280
rect 9612 9216 9618 9280
rect 9302 9215 9618 9216
rect 12402 9280 12718 9281
rect 12402 9216 12408 9280
rect 12472 9216 12488 9280
rect 12552 9216 12568 9280
rect 12632 9216 12648 9280
rect 12712 9216 12718 9280
rect 12402 9215 12718 9216
rect 15502 9280 15818 9281
rect 15502 9216 15508 9280
rect 15572 9216 15588 9280
rect 15652 9216 15668 9280
rect 15732 9216 15748 9280
rect 15812 9216 15818 9280
rect 15502 9215 15818 9216
rect 18602 9280 18918 9281
rect 18602 9216 18608 9280
rect 18672 9216 18688 9280
rect 18752 9216 18768 9280
rect 18832 9216 18848 9280
rect 18912 9216 18918 9280
rect 18602 9215 18918 9216
rect 18413 8802 18479 8805
rect 19200 8802 20000 8832
rect 18413 8800 20000 8802
rect 18413 8744 18418 8800
rect 18474 8744 20000 8800
rect 18413 8742 20000 8744
rect 18413 8739 18479 8742
rect 1552 8736 1868 8737
rect 1552 8672 1558 8736
rect 1622 8672 1638 8736
rect 1702 8672 1718 8736
rect 1782 8672 1798 8736
rect 1862 8672 1868 8736
rect 1552 8671 1868 8672
rect 4652 8736 4968 8737
rect 4652 8672 4658 8736
rect 4722 8672 4738 8736
rect 4802 8672 4818 8736
rect 4882 8672 4898 8736
rect 4962 8672 4968 8736
rect 4652 8671 4968 8672
rect 7752 8736 8068 8737
rect 7752 8672 7758 8736
rect 7822 8672 7838 8736
rect 7902 8672 7918 8736
rect 7982 8672 7998 8736
rect 8062 8672 8068 8736
rect 7752 8671 8068 8672
rect 10852 8736 11168 8737
rect 10852 8672 10858 8736
rect 10922 8672 10938 8736
rect 11002 8672 11018 8736
rect 11082 8672 11098 8736
rect 11162 8672 11168 8736
rect 10852 8671 11168 8672
rect 13952 8736 14268 8737
rect 13952 8672 13958 8736
rect 14022 8672 14038 8736
rect 14102 8672 14118 8736
rect 14182 8672 14198 8736
rect 14262 8672 14268 8736
rect 13952 8671 14268 8672
rect 17052 8736 17368 8737
rect 17052 8672 17058 8736
rect 17122 8672 17138 8736
rect 17202 8672 17218 8736
rect 17282 8672 17298 8736
rect 17362 8672 17368 8736
rect 19200 8712 20000 8742
rect 17052 8671 17368 8672
rect 3102 8192 3418 8193
rect 3102 8128 3108 8192
rect 3172 8128 3188 8192
rect 3252 8128 3268 8192
rect 3332 8128 3348 8192
rect 3412 8128 3418 8192
rect 3102 8127 3418 8128
rect 6202 8192 6518 8193
rect 6202 8128 6208 8192
rect 6272 8128 6288 8192
rect 6352 8128 6368 8192
rect 6432 8128 6448 8192
rect 6512 8128 6518 8192
rect 6202 8127 6518 8128
rect 9302 8192 9618 8193
rect 9302 8128 9308 8192
rect 9372 8128 9388 8192
rect 9452 8128 9468 8192
rect 9532 8128 9548 8192
rect 9612 8128 9618 8192
rect 9302 8127 9618 8128
rect 12402 8192 12718 8193
rect 12402 8128 12408 8192
rect 12472 8128 12488 8192
rect 12552 8128 12568 8192
rect 12632 8128 12648 8192
rect 12712 8128 12718 8192
rect 12402 8127 12718 8128
rect 15502 8192 15818 8193
rect 15502 8128 15508 8192
rect 15572 8128 15588 8192
rect 15652 8128 15668 8192
rect 15732 8128 15748 8192
rect 15812 8128 15818 8192
rect 15502 8127 15818 8128
rect 18602 8192 18918 8193
rect 18602 8128 18608 8192
rect 18672 8128 18688 8192
rect 18752 8128 18768 8192
rect 18832 8128 18848 8192
rect 18912 8128 18918 8192
rect 18602 8127 18918 8128
rect 1552 7648 1868 7649
rect 1552 7584 1558 7648
rect 1622 7584 1638 7648
rect 1702 7584 1718 7648
rect 1782 7584 1798 7648
rect 1862 7584 1868 7648
rect 1552 7583 1868 7584
rect 4652 7648 4968 7649
rect 4652 7584 4658 7648
rect 4722 7584 4738 7648
rect 4802 7584 4818 7648
rect 4882 7584 4898 7648
rect 4962 7584 4968 7648
rect 4652 7583 4968 7584
rect 7752 7648 8068 7649
rect 7752 7584 7758 7648
rect 7822 7584 7838 7648
rect 7902 7584 7918 7648
rect 7982 7584 7998 7648
rect 8062 7584 8068 7648
rect 7752 7583 8068 7584
rect 10852 7648 11168 7649
rect 10852 7584 10858 7648
rect 10922 7584 10938 7648
rect 11002 7584 11018 7648
rect 11082 7584 11098 7648
rect 11162 7584 11168 7648
rect 10852 7583 11168 7584
rect 13952 7648 14268 7649
rect 13952 7584 13958 7648
rect 14022 7584 14038 7648
rect 14102 7584 14118 7648
rect 14182 7584 14198 7648
rect 14262 7584 14268 7648
rect 13952 7583 14268 7584
rect 17052 7648 17368 7649
rect 17052 7584 17058 7648
rect 17122 7584 17138 7648
rect 17202 7584 17218 7648
rect 17282 7584 17298 7648
rect 17362 7584 17368 7648
rect 17052 7583 17368 7584
rect 3102 7104 3418 7105
rect 3102 7040 3108 7104
rect 3172 7040 3188 7104
rect 3252 7040 3268 7104
rect 3332 7040 3348 7104
rect 3412 7040 3418 7104
rect 3102 7039 3418 7040
rect 6202 7104 6518 7105
rect 6202 7040 6208 7104
rect 6272 7040 6288 7104
rect 6352 7040 6368 7104
rect 6432 7040 6448 7104
rect 6512 7040 6518 7104
rect 6202 7039 6518 7040
rect 9302 7104 9618 7105
rect 9302 7040 9308 7104
rect 9372 7040 9388 7104
rect 9452 7040 9468 7104
rect 9532 7040 9548 7104
rect 9612 7040 9618 7104
rect 9302 7039 9618 7040
rect 12402 7104 12718 7105
rect 12402 7040 12408 7104
rect 12472 7040 12488 7104
rect 12552 7040 12568 7104
rect 12632 7040 12648 7104
rect 12712 7040 12718 7104
rect 12402 7039 12718 7040
rect 15502 7104 15818 7105
rect 15502 7040 15508 7104
rect 15572 7040 15588 7104
rect 15652 7040 15668 7104
rect 15732 7040 15748 7104
rect 15812 7040 15818 7104
rect 15502 7039 15818 7040
rect 18602 7104 18918 7105
rect 18602 7040 18608 7104
rect 18672 7040 18688 7104
rect 18752 7040 18768 7104
rect 18832 7040 18848 7104
rect 18912 7040 18918 7104
rect 18602 7039 18918 7040
rect 1552 6560 1868 6561
rect 1552 6496 1558 6560
rect 1622 6496 1638 6560
rect 1702 6496 1718 6560
rect 1782 6496 1798 6560
rect 1862 6496 1868 6560
rect 1552 6495 1868 6496
rect 4652 6560 4968 6561
rect 4652 6496 4658 6560
rect 4722 6496 4738 6560
rect 4802 6496 4818 6560
rect 4882 6496 4898 6560
rect 4962 6496 4968 6560
rect 4652 6495 4968 6496
rect 7752 6560 8068 6561
rect 7752 6496 7758 6560
rect 7822 6496 7838 6560
rect 7902 6496 7918 6560
rect 7982 6496 7998 6560
rect 8062 6496 8068 6560
rect 7752 6495 8068 6496
rect 10852 6560 11168 6561
rect 10852 6496 10858 6560
rect 10922 6496 10938 6560
rect 11002 6496 11018 6560
rect 11082 6496 11098 6560
rect 11162 6496 11168 6560
rect 10852 6495 11168 6496
rect 13952 6560 14268 6561
rect 13952 6496 13958 6560
rect 14022 6496 14038 6560
rect 14102 6496 14118 6560
rect 14182 6496 14198 6560
rect 14262 6496 14268 6560
rect 13952 6495 14268 6496
rect 17052 6560 17368 6561
rect 17052 6496 17058 6560
rect 17122 6496 17138 6560
rect 17202 6496 17218 6560
rect 17282 6496 17298 6560
rect 17362 6496 17368 6560
rect 17052 6495 17368 6496
rect 18413 6354 18479 6357
rect 19200 6354 20000 6384
rect 18413 6352 20000 6354
rect 18413 6296 18418 6352
rect 18474 6296 20000 6352
rect 18413 6294 20000 6296
rect 18413 6291 18479 6294
rect 19200 6264 20000 6294
rect 3102 6016 3418 6017
rect 3102 5952 3108 6016
rect 3172 5952 3188 6016
rect 3252 5952 3268 6016
rect 3332 5952 3348 6016
rect 3412 5952 3418 6016
rect 3102 5951 3418 5952
rect 6202 6016 6518 6017
rect 6202 5952 6208 6016
rect 6272 5952 6288 6016
rect 6352 5952 6368 6016
rect 6432 5952 6448 6016
rect 6512 5952 6518 6016
rect 6202 5951 6518 5952
rect 9302 6016 9618 6017
rect 9302 5952 9308 6016
rect 9372 5952 9388 6016
rect 9452 5952 9468 6016
rect 9532 5952 9548 6016
rect 9612 5952 9618 6016
rect 9302 5951 9618 5952
rect 12402 6016 12718 6017
rect 12402 5952 12408 6016
rect 12472 5952 12488 6016
rect 12552 5952 12568 6016
rect 12632 5952 12648 6016
rect 12712 5952 12718 6016
rect 12402 5951 12718 5952
rect 15502 6016 15818 6017
rect 15502 5952 15508 6016
rect 15572 5952 15588 6016
rect 15652 5952 15668 6016
rect 15732 5952 15748 6016
rect 15812 5952 15818 6016
rect 15502 5951 15818 5952
rect 18602 6016 18918 6017
rect 18602 5952 18608 6016
rect 18672 5952 18688 6016
rect 18752 5952 18768 6016
rect 18832 5952 18848 6016
rect 18912 5952 18918 6016
rect 18602 5951 18918 5952
rect 1552 5472 1868 5473
rect 1552 5408 1558 5472
rect 1622 5408 1638 5472
rect 1702 5408 1718 5472
rect 1782 5408 1798 5472
rect 1862 5408 1868 5472
rect 1552 5407 1868 5408
rect 4652 5472 4968 5473
rect 4652 5408 4658 5472
rect 4722 5408 4738 5472
rect 4802 5408 4818 5472
rect 4882 5408 4898 5472
rect 4962 5408 4968 5472
rect 4652 5407 4968 5408
rect 7752 5472 8068 5473
rect 7752 5408 7758 5472
rect 7822 5408 7838 5472
rect 7902 5408 7918 5472
rect 7982 5408 7998 5472
rect 8062 5408 8068 5472
rect 7752 5407 8068 5408
rect 10852 5472 11168 5473
rect 10852 5408 10858 5472
rect 10922 5408 10938 5472
rect 11002 5408 11018 5472
rect 11082 5408 11098 5472
rect 11162 5408 11168 5472
rect 10852 5407 11168 5408
rect 13952 5472 14268 5473
rect 13952 5408 13958 5472
rect 14022 5408 14038 5472
rect 14102 5408 14118 5472
rect 14182 5408 14198 5472
rect 14262 5408 14268 5472
rect 13952 5407 14268 5408
rect 17052 5472 17368 5473
rect 17052 5408 17058 5472
rect 17122 5408 17138 5472
rect 17202 5408 17218 5472
rect 17282 5408 17298 5472
rect 17362 5408 17368 5472
rect 17052 5407 17368 5408
rect 3102 4928 3418 4929
rect 3102 4864 3108 4928
rect 3172 4864 3188 4928
rect 3252 4864 3268 4928
rect 3332 4864 3348 4928
rect 3412 4864 3418 4928
rect 3102 4863 3418 4864
rect 6202 4928 6518 4929
rect 6202 4864 6208 4928
rect 6272 4864 6288 4928
rect 6352 4864 6368 4928
rect 6432 4864 6448 4928
rect 6512 4864 6518 4928
rect 6202 4863 6518 4864
rect 9302 4928 9618 4929
rect 9302 4864 9308 4928
rect 9372 4864 9388 4928
rect 9452 4864 9468 4928
rect 9532 4864 9548 4928
rect 9612 4864 9618 4928
rect 9302 4863 9618 4864
rect 12402 4928 12718 4929
rect 12402 4864 12408 4928
rect 12472 4864 12488 4928
rect 12552 4864 12568 4928
rect 12632 4864 12648 4928
rect 12712 4864 12718 4928
rect 12402 4863 12718 4864
rect 15502 4928 15818 4929
rect 15502 4864 15508 4928
rect 15572 4864 15588 4928
rect 15652 4864 15668 4928
rect 15732 4864 15748 4928
rect 15812 4864 15818 4928
rect 15502 4863 15818 4864
rect 18602 4928 18918 4929
rect 18602 4864 18608 4928
rect 18672 4864 18688 4928
rect 18752 4864 18768 4928
rect 18832 4864 18848 4928
rect 18912 4864 18918 4928
rect 18602 4863 18918 4864
rect 1552 4384 1868 4385
rect 1552 4320 1558 4384
rect 1622 4320 1638 4384
rect 1702 4320 1718 4384
rect 1782 4320 1798 4384
rect 1862 4320 1868 4384
rect 1552 4319 1868 4320
rect 4652 4384 4968 4385
rect 4652 4320 4658 4384
rect 4722 4320 4738 4384
rect 4802 4320 4818 4384
rect 4882 4320 4898 4384
rect 4962 4320 4968 4384
rect 4652 4319 4968 4320
rect 7752 4384 8068 4385
rect 7752 4320 7758 4384
rect 7822 4320 7838 4384
rect 7902 4320 7918 4384
rect 7982 4320 7998 4384
rect 8062 4320 8068 4384
rect 7752 4319 8068 4320
rect 10852 4384 11168 4385
rect 10852 4320 10858 4384
rect 10922 4320 10938 4384
rect 11002 4320 11018 4384
rect 11082 4320 11098 4384
rect 11162 4320 11168 4384
rect 10852 4319 11168 4320
rect 13952 4384 14268 4385
rect 13952 4320 13958 4384
rect 14022 4320 14038 4384
rect 14102 4320 14118 4384
rect 14182 4320 14198 4384
rect 14262 4320 14268 4384
rect 13952 4319 14268 4320
rect 17052 4384 17368 4385
rect 17052 4320 17058 4384
rect 17122 4320 17138 4384
rect 17202 4320 17218 4384
rect 17282 4320 17298 4384
rect 17362 4320 17368 4384
rect 17052 4319 17368 4320
rect 19057 3906 19123 3909
rect 19200 3906 20000 3936
rect 19057 3904 20000 3906
rect 19057 3848 19062 3904
rect 19118 3848 20000 3904
rect 19057 3846 20000 3848
rect 19057 3843 19123 3846
rect 3102 3840 3418 3841
rect 3102 3776 3108 3840
rect 3172 3776 3188 3840
rect 3252 3776 3268 3840
rect 3332 3776 3348 3840
rect 3412 3776 3418 3840
rect 3102 3775 3418 3776
rect 6202 3840 6518 3841
rect 6202 3776 6208 3840
rect 6272 3776 6288 3840
rect 6352 3776 6368 3840
rect 6432 3776 6448 3840
rect 6512 3776 6518 3840
rect 6202 3775 6518 3776
rect 9302 3840 9618 3841
rect 9302 3776 9308 3840
rect 9372 3776 9388 3840
rect 9452 3776 9468 3840
rect 9532 3776 9548 3840
rect 9612 3776 9618 3840
rect 9302 3775 9618 3776
rect 12402 3840 12718 3841
rect 12402 3776 12408 3840
rect 12472 3776 12488 3840
rect 12552 3776 12568 3840
rect 12632 3776 12648 3840
rect 12712 3776 12718 3840
rect 12402 3775 12718 3776
rect 15502 3840 15818 3841
rect 15502 3776 15508 3840
rect 15572 3776 15588 3840
rect 15652 3776 15668 3840
rect 15732 3776 15748 3840
rect 15812 3776 15818 3840
rect 15502 3775 15818 3776
rect 18602 3840 18918 3841
rect 18602 3776 18608 3840
rect 18672 3776 18688 3840
rect 18752 3776 18768 3840
rect 18832 3776 18848 3840
rect 18912 3776 18918 3840
rect 19200 3816 20000 3846
rect 18602 3775 18918 3776
rect 1552 3296 1868 3297
rect 1552 3232 1558 3296
rect 1622 3232 1638 3296
rect 1702 3232 1718 3296
rect 1782 3232 1798 3296
rect 1862 3232 1868 3296
rect 1552 3231 1868 3232
rect 4652 3296 4968 3297
rect 4652 3232 4658 3296
rect 4722 3232 4738 3296
rect 4802 3232 4818 3296
rect 4882 3232 4898 3296
rect 4962 3232 4968 3296
rect 4652 3231 4968 3232
rect 7752 3296 8068 3297
rect 7752 3232 7758 3296
rect 7822 3232 7838 3296
rect 7902 3232 7918 3296
rect 7982 3232 7998 3296
rect 8062 3232 8068 3296
rect 7752 3231 8068 3232
rect 10852 3296 11168 3297
rect 10852 3232 10858 3296
rect 10922 3232 10938 3296
rect 11002 3232 11018 3296
rect 11082 3232 11098 3296
rect 11162 3232 11168 3296
rect 10852 3231 11168 3232
rect 13952 3296 14268 3297
rect 13952 3232 13958 3296
rect 14022 3232 14038 3296
rect 14102 3232 14118 3296
rect 14182 3232 14198 3296
rect 14262 3232 14268 3296
rect 13952 3231 14268 3232
rect 17052 3296 17368 3297
rect 17052 3232 17058 3296
rect 17122 3232 17138 3296
rect 17202 3232 17218 3296
rect 17282 3232 17298 3296
rect 17362 3232 17368 3296
rect 17052 3231 17368 3232
rect 3102 2752 3418 2753
rect 3102 2688 3108 2752
rect 3172 2688 3188 2752
rect 3252 2688 3268 2752
rect 3332 2688 3348 2752
rect 3412 2688 3418 2752
rect 3102 2687 3418 2688
rect 6202 2752 6518 2753
rect 6202 2688 6208 2752
rect 6272 2688 6288 2752
rect 6352 2688 6368 2752
rect 6432 2688 6448 2752
rect 6512 2688 6518 2752
rect 6202 2687 6518 2688
rect 9302 2752 9618 2753
rect 9302 2688 9308 2752
rect 9372 2688 9388 2752
rect 9452 2688 9468 2752
rect 9532 2688 9548 2752
rect 9612 2688 9618 2752
rect 9302 2687 9618 2688
rect 12402 2752 12718 2753
rect 12402 2688 12408 2752
rect 12472 2688 12488 2752
rect 12552 2688 12568 2752
rect 12632 2688 12648 2752
rect 12712 2688 12718 2752
rect 12402 2687 12718 2688
rect 15502 2752 15818 2753
rect 15502 2688 15508 2752
rect 15572 2688 15588 2752
rect 15652 2688 15668 2752
rect 15732 2688 15748 2752
rect 15812 2688 15818 2752
rect 15502 2687 15818 2688
rect 18602 2752 18918 2753
rect 18602 2688 18608 2752
rect 18672 2688 18688 2752
rect 18752 2688 18768 2752
rect 18832 2688 18848 2752
rect 18912 2688 18918 2752
rect 18602 2687 18918 2688
rect 1552 2208 1868 2209
rect 1552 2144 1558 2208
rect 1622 2144 1638 2208
rect 1702 2144 1718 2208
rect 1782 2144 1798 2208
rect 1862 2144 1868 2208
rect 1552 2143 1868 2144
rect 4652 2208 4968 2209
rect 4652 2144 4658 2208
rect 4722 2144 4738 2208
rect 4802 2144 4818 2208
rect 4882 2144 4898 2208
rect 4962 2144 4968 2208
rect 4652 2143 4968 2144
rect 7752 2208 8068 2209
rect 7752 2144 7758 2208
rect 7822 2144 7838 2208
rect 7902 2144 7918 2208
rect 7982 2144 7998 2208
rect 8062 2144 8068 2208
rect 7752 2143 8068 2144
rect 10852 2208 11168 2209
rect 10852 2144 10858 2208
rect 10922 2144 10938 2208
rect 11002 2144 11018 2208
rect 11082 2144 11098 2208
rect 11162 2144 11168 2208
rect 10852 2143 11168 2144
rect 13952 2208 14268 2209
rect 13952 2144 13958 2208
rect 14022 2144 14038 2208
rect 14102 2144 14118 2208
rect 14182 2144 14198 2208
rect 14262 2144 14268 2208
rect 13952 2143 14268 2144
rect 17052 2208 17368 2209
rect 17052 2144 17058 2208
rect 17122 2144 17138 2208
rect 17202 2144 17218 2208
rect 17282 2144 17298 2208
rect 17362 2144 17368 2208
rect 17052 2143 17368 2144
rect 3102 1664 3418 1665
rect 3102 1600 3108 1664
rect 3172 1600 3188 1664
rect 3252 1600 3268 1664
rect 3332 1600 3348 1664
rect 3412 1600 3418 1664
rect 3102 1599 3418 1600
rect 6202 1664 6518 1665
rect 6202 1600 6208 1664
rect 6272 1600 6288 1664
rect 6352 1600 6368 1664
rect 6432 1600 6448 1664
rect 6512 1600 6518 1664
rect 6202 1599 6518 1600
rect 9302 1664 9618 1665
rect 9302 1600 9308 1664
rect 9372 1600 9388 1664
rect 9452 1600 9468 1664
rect 9532 1600 9548 1664
rect 9612 1600 9618 1664
rect 9302 1599 9618 1600
rect 12402 1664 12718 1665
rect 12402 1600 12408 1664
rect 12472 1600 12488 1664
rect 12552 1600 12568 1664
rect 12632 1600 12648 1664
rect 12712 1600 12718 1664
rect 12402 1599 12718 1600
rect 15502 1664 15818 1665
rect 15502 1600 15508 1664
rect 15572 1600 15588 1664
rect 15652 1600 15668 1664
rect 15732 1600 15748 1664
rect 15812 1600 15818 1664
rect 15502 1599 15818 1600
rect 18602 1664 18918 1665
rect 18602 1600 18608 1664
rect 18672 1600 18688 1664
rect 18752 1600 18768 1664
rect 18832 1600 18848 1664
rect 18912 1600 18918 1664
rect 18602 1599 18918 1600
rect 18413 1458 18479 1461
rect 19200 1458 20000 1488
rect 18413 1456 20000 1458
rect 18413 1400 18418 1456
rect 18474 1400 20000 1456
rect 18413 1398 20000 1400
rect 18413 1395 18479 1398
rect 19200 1368 20000 1398
rect 1552 1120 1868 1121
rect 1552 1056 1558 1120
rect 1622 1056 1638 1120
rect 1702 1056 1718 1120
rect 1782 1056 1798 1120
rect 1862 1056 1868 1120
rect 1552 1055 1868 1056
rect 4652 1120 4968 1121
rect 4652 1056 4658 1120
rect 4722 1056 4738 1120
rect 4802 1056 4818 1120
rect 4882 1056 4898 1120
rect 4962 1056 4968 1120
rect 4652 1055 4968 1056
rect 7752 1120 8068 1121
rect 7752 1056 7758 1120
rect 7822 1056 7838 1120
rect 7902 1056 7918 1120
rect 7982 1056 7998 1120
rect 8062 1056 8068 1120
rect 7752 1055 8068 1056
rect 10852 1120 11168 1121
rect 10852 1056 10858 1120
rect 10922 1056 10938 1120
rect 11002 1056 11018 1120
rect 11082 1056 11098 1120
rect 11162 1056 11168 1120
rect 10852 1055 11168 1056
rect 13952 1120 14268 1121
rect 13952 1056 13958 1120
rect 14022 1056 14038 1120
rect 14102 1056 14118 1120
rect 14182 1056 14198 1120
rect 14262 1056 14268 1120
rect 13952 1055 14268 1056
rect 17052 1120 17368 1121
rect 17052 1056 17058 1120
rect 17122 1056 17138 1120
rect 17202 1056 17218 1120
rect 17282 1056 17298 1120
rect 17362 1056 17368 1120
rect 17052 1055 17368 1056
rect 3102 576 3418 577
rect 3102 512 3108 576
rect 3172 512 3188 576
rect 3252 512 3268 576
rect 3332 512 3348 576
rect 3412 512 3418 576
rect 3102 511 3418 512
rect 6202 576 6518 577
rect 6202 512 6208 576
rect 6272 512 6288 576
rect 6352 512 6368 576
rect 6432 512 6448 576
rect 6512 512 6518 576
rect 6202 511 6518 512
rect 9302 576 9618 577
rect 9302 512 9308 576
rect 9372 512 9388 576
rect 9452 512 9468 576
rect 9532 512 9548 576
rect 9612 512 9618 576
rect 9302 511 9618 512
rect 12402 576 12718 577
rect 12402 512 12408 576
rect 12472 512 12488 576
rect 12552 512 12568 576
rect 12632 512 12648 576
rect 12712 512 12718 576
rect 12402 511 12718 512
rect 15502 576 15818 577
rect 15502 512 15508 576
rect 15572 512 15588 576
rect 15652 512 15668 576
rect 15732 512 15748 576
rect 15812 512 15818 576
rect 15502 511 15818 512
rect 18602 576 18918 577
rect 18602 512 18608 576
rect 18672 512 18688 576
rect 18752 512 18768 576
rect 18832 512 18848 576
rect 18912 512 18918 576
rect 18602 511 18918 512
<< via3 >>
rect 1558 18524 1622 18528
rect 1558 18468 1562 18524
rect 1562 18468 1618 18524
rect 1618 18468 1622 18524
rect 1558 18464 1622 18468
rect 1638 18524 1702 18528
rect 1638 18468 1642 18524
rect 1642 18468 1698 18524
rect 1698 18468 1702 18524
rect 1638 18464 1702 18468
rect 1718 18524 1782 18528
rect 1718 18468 1722 18524
rect 1722 18468 1778 18524
rect 1778 18468 1782 18524
rect 1718 18464 1782 18468
rect 1798 18524 1862 18528
rect 1798 18468 1802 18524
rect 1802 18468 1858 18524
rect 1858 18468 1862 18524
rect 1798 18464 1862 18468
rect 4658 18524 4722 18528
rect 4658 18468 4662 18524
rect 4662 18468 4718 18524
rect 4718 18468 4722 18524
rect 4658 18464 4722 18468
rect 4738 18524 4802 18528
rect 4738 18468 4742 18524
rect 4742 18468 4798 18524
rect 4798 18468 4802 18524
rect 4738 18464 4802 18468
rect 4818 18524 4882 18528
rect 4818 18468 4822 18524
rect 4822 18468 4878 18524
rect 4878 18468 4882 18524
rect 4818 18464 4882 18468
rect 4898 18524 4962 18528
rect 4898 18468 4902 18524
rect 4902 18468 4958 18524
rect 4958 18468 4962 18524
rect 4898 18464 4962 18468
rect 7758 18524 7822 18528
rect 7758 18468 7762 18524
rect 7762 18468 7818 18524
rect 7818 18468 7822 18524
rect 7758 18464 7822 18468
rect 7838 18524 7902 18528
rect 7838 18468 7842 18524
rect 7842 18468 7898 18524
rect 7898 18468 7902 18524
rect 7838 18464 7902 18468
rect 7918 18524 7982 18528
rect 7918 18468 7922 18524
rect 7922 18468 7978 18524
rect 7978 18468 7982 18524
rect 7918 18464 7982 18468
rect 7998 18524 8062 18528
rect 7998 18468 8002 18524
rect 8002 18468 8058 18524
rect 8058 18468 8062 18524
rect 7998 18464 8062 18468
rect 10858 18524 10922 18528
rect 10858 18468 10862 18524
rect 10862 18468 10918 18524
rect 10918 18468 10922 18524
rect 10858 18464 10922 18468
rect 10938 18524 11002 18528
rect 10938 18468 10942 18524
rect 10942 18468 10998 18524
rect 10998 18468 11002 18524
rect 10938 18464 11002 18468
rect 11018 18524 11082 18528
rect 11018 18468 11022 18524
rect 11022 18468 11078 18524
rect 11078 18468 11082 18524
rect 11018 18464 11082 18468
rect 11098 18524 11162 18528
rect 11098 18468 11102 18524
rect 11102 18468 11158 18524
rect 11158 18468 11162 18524
rect 11098 18464 11162 18468
rect 13958 18524 14022 18528
rect 13958 18468 13962 18524
rect 13962 18468 14018 18524
rect 14018 18468 14022 18524
rect 13958 18464 14022 18468
rect 14038 18524 14102 18528
rect 14038 18468 14042 18524
rect 14042 18468 14098 18524
rect 14098 18468 14102 18524
rect 14038 18464 14102 18468
rect 14118 18524 14182 18528
rect 14118 18468 14122 18524
rect 14122 18468 14178 18524
rect 14178 18468 14182 18524
rect 14118 18464 14182 18468
rect 14198 18524 14262 18528
rect 14198 18468 14202 18524
rect 14202 18468 14258 18524
rect 14258 18468 14262 18524
rect 14198 18464 14262 18468
rect 17058 18524 17122 18528
rect 17058 18468 17062 18524
rect 17062 18468 17118 18524
rect 17118 18468 17122 18524
rect 17058 18464 17122 18468
rect 17138 18524 17202 18528
rect 17138 18468 17142 18524
rect 17142 18468 17198 18524
rect 17198 18468 17202 18524
rect 17138 18464 17202 18468
rect 17218 18524 17282 18528
rect 17218 18468 17222 18524
rect 17222 18468 17278 18524
rect 17278 18468 17282 18524
rect 17218 18464 17282 18468
rect 17298 18524 17362 18528
rect 17298 18468 17302 18524
rect 17302 18468 17358 18524
rect 17358 18468 17362 18524
rect 17298 18464 17362 18468
rect 3108 17980 3172 17984
rect 3108 17924 3112 17980
rect 3112 17924 3168 17980
rect 3168 17924 3172 17980
rect 3108 17920 3172 17924
rect 3188 17980 3252 17984
rect 3188 17924 3192 17980
rect 3192 17924 3248 17980
rect 3248 17924 3252 17980
rect 3188 17920 3252 17924
rect 3268 17980 3332 17984
rect 3268 17924 3272 17980
rect 3272 17924 3328 17980
rect 3328 17924 3332 17980
rect 3268 17920 3332 17924
rect 3348 17980 3412 17984
rect 3348 17924 3352 17980
rect 3352 17924 3408 17980
rect 3408 17924 3412 17980
rect 3348 17920 3412 17924
rect 6208 17980 6272 17984
rect 6208 17924 6212 17980
rect 6212 17924 6268 17980
rect 6268 17924 6272 17980
rect 6208 17920 6272 17924
rect 6288 17980 6352 17984
rect 6288 17924 6292 17980
rect 6292 17924 6348 17980
rect 6348 17924 6352 17980
rect 6288 17920 6352 17924
rect 6368 17980 6432 17984
rect 6368 17924 6372 17980
rect 6372 17924 6428 17980
rect 6428 17924 6432 17980
rect 6368 17920 6432 17924
rect 6448 17980 6512 17984
rect 6448 17924 6452 17980
rect 6452 17924 6508 17980
rect 6508 17924 6512 17980
rect 6448 17920 6512 17924
rect 9308 17980 9372 17984
rect 9308 17924 9312 17980
rect 9312 17924 9368 17980
rect 9368 17924 9372 17980
rect 9308 17920 9372 17924
rect 9388 17980 9452 17984
rect 9388 17924 9392 17980
rect 9392 17924 9448 17980
rect 9448 17924 9452 17980
rect 9388 17920 9452 17924
rect 9468 17980 9532 17984
rect 9468 17924 9472 17980
rect 9472 17924 9528 17980
rect 9528 17924 9532 17980
rect 9468 17920 9532 17924
rect 9548 17980 9612 17984
rect 9548 17924 9552 17980
rect 9552 17924 9608 17980
rect 9608 17924 9612 17980
rect 9548 17920 9612 17924
rect 12408 17980 12472 17984
rect 12408 17924 12412 17980
rect 12412 17924 12468 17980
rect 12468 17924 12472 17980
rect 12408 17920 12472 17924
rect 12488 17980 12552 17984
rect 12488 17924 12492 17980
rect 12492 17924 12548 17980
rect 12548 17924 12552 17980
rect 12488 17920 12552 17924
rect 12568 17980 12632 17984
rect 12568 17924 12572 17980
rect 12572 17924 12628 17980
rect 12628 17924 12632 17980
rect 12568 17920 12632 17924
rect 12648 17980 12712 17984
rect 12648 17924 12652 17980
rect 12652 17924 12708 17980
rect 12708 17924 12712 17980
rect 12648 17920 12712 17924
rect 15508 17980 15572 17984
rect 15508 17924 15512 17980
rect 15512 17924 15568 17980
rect 15568 17924 15572 17980
rect 15508 17920 15572 17924
rect 15588 17980 15652 17984
rect 15588 17924 15592 17980
rect 15592 17924 15648 17980
rect 15648 17924 15652 17980
rect 15588 17920 15652 17924
rect 15668 17980 15732 17984
rect 15668 17924 15672 17980
rect 15672 17924 15728 17980
rect 15728 17924 15732 17980
rect 15668 17920 15732 17924
rect 15748 17980 15812 17984
rect 15748 17924 15752 17980
rect 15752 17924 15808 17980
rect 15808 17924 15812 17980
rect 15748 17920 15812 17924
rect 18608 17980 18672 17984
rect 18608 17924 18612 17980
rect 18612 17924 18668 17980
rect 18668 17924 18672 17980
rect 18608 17920 18672 17924
rect 18688 17980 18752 17984
rect 18688 17924 18692 17980
rect 18692 17924 18748 17980
rect 18748 17924 18752 17980
rect 18688 17920 18752 17924
rect 18768 17980 18832 17984
rect 18768 17924 18772 17980
rect 18772 17924 18828 17980
rect 18828 17924 18832 17980
rect 18768 17920 18832 17924
rect 18848 17980 18912 17984
rect 18848 17924 18852 17980
rect 18852 17924 18908 17980
rect 18908 17924 18912 17980
rect 18848 17920 18912 17924
rect 1558 17436 1622 17440
rect 1558 17380 1562 17436
rect 1562 17380 1618 17436
rect 1618 17380 1622 17436
rect 1558 17376 1622 17380
rect 1638 17436 1702 17440
rect 1638 17380 1642 17436
rect 1642 17380 1698 17436
rect 1698 17380 1702 17436
rect 1638 17376 1702 17380
rect 1718 17436 1782 17440
rect 1718 17380 1722 17436
rect 1722 17380 1778 17436
rect 1778 17380 1782 17436
rect 1718 17376 1782 17380
rect 1798 17436 1862 17440
rect 1798 17380 1802 17436
rect 1802 17380 1858 17436
rect 1858 17380 1862 17436
rect 1798 17376 1862 17380
rect 4658 17436 4722 17440
rect 4658 17380 4662 17436
rect 4662 17380 4718 17436
rect 4718 17380 4722 17436
rect 4658 17376 4722 17380
rect 4738 17436 4802 17440
rect 4738 17380 4742 17436
rect 4742 17380 4798 17436
rect 4798 17380 4802 17436
rect 4738 17376 4802 17380
rect 4818 17436 4882 17440
rect 4818 17380 4822 17436
rect 4822 17380 4878 17436
rect 4878 17380 4882 17436
rect 4818 17376 4882 17380
rect 4898 17436 4962 17440
rect 4898 17380 4902 17436
rect 4902 17380 4958 17436
rect 4958 17380 4962 17436
rect 4898 17376 4962 17380
rect 7758 17436 7822 17440
rect 7758 17380 7762 17436
rect 7762 17380 7818 17436
rect 7818 17380 7822 17436
rect 7758 17376 7822 17380
rect 7838 17436 7902 17440
rect 7838 17380 7842 17436
rect 7842 17380 7898 17436
rect 7898 17380 7902 17436
rect 7838 17376 7902 17380
rect 7918 17436 7982 17440
rect 7918 17380 7922 17436
rect 7922 17380 7978 17436
rect 7978 17380 7982 17436
rect 7918 17376 7982 17380
rect 7998 17436 8062 17440
rect 7998 17380 8002 17436
rect 8002 17380 8058 17436
rect 8058 17380 8062 17436
rect 7998 17376 8062 17380
rect 10858 17436 10922 17440
rect 10858 17380 10862 17436
rect 10862 17380 10918 17436
rect 10918 17380 10922 17436
rect 10858 17376 10922 17380
rect 10938 17436 11002 17440
rect 10938 17380 10942 17436
rect 10942 17380 10998 17436
rect 10998 17380 11002 17436
rect 10938 17376 11002 17380
rect 11018 17436 11082 17440
rect 11018 17380 11022 17436
rect 11022 17380 11078 17436
rect 11078 17380 11082 17436
rect 11018 17376 11082 17380
rect 11098 17436 11162 17440
rect 11098 17380 11102 17436
rect 11102 17380 11158 17436
rect 11158 17380 11162 17436
rect 11098 17376 11162 17380
rect 13958 17436 14022 17440
rect 13958 17380 13962 17436
rect 13962 17380 14018 17436
rect 14018 17380 14022 17436
rect 13958 17376 14022 17380
rect 14038 17436 14102 17440
rect 14038 17380 14042 17436
rect 14042 17380 14098 17436
rect 14098 17380 14102 17436
rect 14038 17376 14102 17380
rect 14118 17436 14182 17440
rect 14118 17380 14122 17436
rect 14122 17380 14178 17436
rect 14178 17380 14182 17436
rect 14118 17376 14182 17380
rect 14198 17436 14262 17440
rect 14198 17380 14202 17436
rect 14202 17380 14258 17436
rect 14258 17380 14262 17436
rect 14198 17376 14262 17380
rect 17058 17436 17122 17440
rect 17058 17380 17062 17436
rect 17062 17380 17118 17436
rect 17118 17380 17122 17436
rect 17058 17376 17122 17380
rect 17138 17436 17202 17440
rect 17138 17380 17142 17436
rect 17142 17380 17198 17436
rect 17198 17380 17202 17436
rect 17138 17376 17202 17380
rect 17218 17436 17282 17440
rect 17218 17380 17222 17436
rect 17222 17380 17278 17436
rect 17278 17380 17282 17436
rect 17218 17376 17282 17380
rect 17298 17436 17362 17440
rect 17298 17380 17302 17436
rect 17302 17380 17358 17436
rect 17358 17380 17362 17436
rect 17298 17376 17362 17380
rect 3108 16892 3172 16896
rect 3108 16836 3112 16892
rect 3112 16836 3168 16892
rect 3168 16836 3172 16892
rect 3108 16832 3172 16836
rect 3188 16892 3252 16896
rect 3188 16836 3192 16892
rect 3192 16836 3248 16892
rect 3248 16836 3252 16892
rect 3188 16832 3252 16836
rect 3268 16892 3332 16896
rect 3268 16836 3272 16892
rect 3272 16836 3328 16892
rect 3328 16836 3332 16892
rect 3268 16832 3332 16836
rect 3348 16892 3412 16896
rect 3348 16836 3352 16892
rect 3352 16836 3408 16892
rect 3408 16836 3412 16892
rect 3348 16832 3412 16836
rect 6208 16892 6272 16896
rect 6208 16836 6212 16892
rect 6212 16836 6268 16892
rect 6268 16836 6272 16892
rect 6208 16832 6272 16836
rect 6288 16892 6352 16896
rect 6288 16836 6292 16892
rect 6292 16836 6348 16892
rect 6348 16836 6352 16892
rect 6288 16832 6352 16836
rect 6368 16892 6432 16896
rect 6368 16836 6372 16892
rect 6372 16836 6428 16892
rect 6428 16836 6432 16892
rect 6368 16832 6432 16836
rect 6448 16892 6512 16896
rect 6448 16836 6452 16892
rect 6452 16836 6508 16892
rect 6508 16836 6512 16892
rect 6448 16832 6512 16836
rect 9308 16892 9372 16896
rect 9308 16836 9312 16892
rect 9312 16836 9368 16892
rect 9368 16836 9372 16892
rect 9308 16832 9372 16836
rect 9388 16892 9452 16896
rect 9388 16836 9392 16892
rect 9392 16836 9448 16892
rect 9448 16836 9452 16892
rect 9388 16832 9452 16836
rect 9468 16892 9532 16896
rect 9468 16836 9472 16892
rect 9472 16836 9528 16892
rect 9528 16836 9532 16892
rect 9468 16832 9532 16836
rect 9548 16892 9612 16896
rect 9548 16836 9552 16892
rect 9552 16836 9608 16892
rect 9608 16836 9612 16892
rect 9548 16832 9612 16836
rect 12408 16892 12472 16896
rect 12408 16836 12412 16892
rect 12412 16836 12468 16892
rect 12468 16836 12472 16892
rect 12408 16832 12472 16836
rect 12488 16892 12552 16896
rect 12488 16836 12492 16892
rect 12492 16836 12548 16892
rect 12548 16836 12552 16892
rect 12488 16832 12552 16836
rect 12568 16892 12632 16896
rect 12568 16836 12572 16892
rect 12572 16836 12628 16892
rect 12628 16836 12632 16892
rect 12568 16832 12632 16836
rect 12648 16892 12712 16896
rect 12648 16836 12652 16892
rect 12652 16836 12708 16892
rect 12708 16836 12712 16892
rect 12648 16832 12712 16836
rect 15508 16892 15572 16896
rect 15508 16836 15512 16892
rect 15512 16836 15568 16892
rect 15568 16836 15572 16892
rect 15508 16832 15572 16836
rect 15588 16892 15652 16896
rect 15588 16836 15592 16892
rect 15592 16836 15648 16892
rect 15648 16836 15652 16892
rect 15588 16832 15652 16836
rect 15668 16892 15732 16896
rect 15668 16836 15672 16892
rect 15672 16836 15728 16892
rect 15728 16836 15732 16892
rect 15668 16832 15732 16836
rect 15748 16892 15812 16896
rect 15748 16836 15752 16892
rect 15752 16836 15808 16892
rect 15808 16836 15812 16892
rect 15748 16832 15812 16836
rect 18608 16892 18672 16896
rect 18608 16836 18612 16892
rect 18612 16836 18668 16892
rect 18668 16836 18672 16892
rect 18608 16832 18672 16836
rect 18688 16892 18752 16896
rect 18688 16836 18692 16892
rect 18692 16836 18748 16892
rect 18748 16836 18752 16892
rect 18688 16832 18752 16836
rect 18768 16892 18832 16896
rect 18768 16836 18772 16892
rect 18772 16836 18828 16892
rect 18828 16836 18832 16892
rect 18768 16832 18832 16836
rect 18848 16892 18912 16896
rect 18848 16836 18852 16892
rect 18852 16836 18908 16892
rect 18908 16836 18912 16892
rect 18848 16832 18912 16836
rect 1558 16348 1622 16352
rect 1558 16292 1562 16348
rect 1562 16292 1618 16348
rect 1618 16292 1622 16348
rect 1558 16288 1622 16292
rect 1638 16348 1702 16352
rect 1638 16292 1642 16348
rect 1642 16292 1698 16348
rect 1698 16292 1702 16348
rect 1638 16288 1702 16292
rect 1718 16348 1782 16352
rect 1718 16292 1722 16348
rect 1722 16292 1778 16348
rect 1778 16292 1782 16348
rect 1718 16288 1782 16292
rect 1798 16348 1862 16352
rect 1798 16292 1802 16348
rect 1802 16292 1858 16348
rect 1858 16292 1862 16348
rect 1798 16288 1862 16292
rect 4658 16348 4722 16352
rect 4658 16292 4662 16348
rect 4662 16292 4718 16348
rect 4718 16292 4722 16348
rect 4658 16288 4722 16292
rect 4738 16348 4802 16352
rect 4738 16292 4742 16348
rect 4742 16292 4798 16348
rect 4798 16292 4802 16348
rect 4738 16288 4802 16292
rect 4818 16348 4882 16352
rect 4818 16292 4822 16348
rect 4822 16292 4878 16348
rect 4878 16292 4882 16348
rect 4818 16288 4882 16292
rect 4898 16348 4962 16352
rect 4898 16292 4902 16348
rect 4902 16292 4958 16348
rect 4958 16292 4962 16348
rect 4898 16288 4962 16292
rect 7758 16348 7822 16352
rect 7758 16292 7762 16348
rect 7762 16292 7818 16348
rect 7818 16292 7822 16348
rect 7758 16288 7822 16292
rect 7838 16348 7902 16352
rect 7838 16292 7842 16348
rect 7842 16292 7898 16348
rect 7898 16292 7902 16348
rect 7838 16288 7902 16292
rect 7918 16348 7982 16352
rect 7918 16292 7922 16348
rect 7922 16292 7978 16348
rect 7978 16292 7982 16348
rect 7918 16288 7982 16292
rect 7998 16348 8062 16352
rect 7998 16292 8002 16348
rect 8002 16292 8058 16348
rect 8058 16292 8062 16348
rect 7998 16288 8062 16292
rect 10858 16348 10922 16352
rect 10858 16292 10862 16348
rect 10862 16292 10918 16348
rect 10918 16292 10922 16348
rect 10858 16288 10922 16292
rect 10938 16348 11002 16352
rect 10938 16292 10942 16348
rect 10942 16292 10998 16348
rect 10998 16292 11002 16348
rect 10938 16288 11002 16292
rect 11018 16348 11082 16352
rect 11018 16292 11022 16348
rect 11022 16292 11078 16348
rect 11078 16292 11082 16348
rect 11018 16288 11082 16292
rect 11098 16348 11162 16352
rect 11098 16292 11102 16348
rect 11102 16292 11158 16348
rect 11158 16292 11162 16348
rect 11098 16288 11162 16292
rect 13958 16348 14022 16352
rect 13958 16292 13962 16348
rect 13962 16292 14018 16348
rect 14018 16292 14022 16348
rect 13958 16288 14022 16292
rect 14038 16348 14102 16352
rect 14038 16292 14042 16348
rect 14042 16292 14098 16348
rect 14098 16292 14102 16348
rect 14038 16288 14102 16292
rect 14118 16348 14182 16352
rect 14118 16292 14122 16348
rect 14122 16292 14178 16348
rect 14178 16292 14182 16348
rect 14118 16288 14182 16292
rect 14198 16348 14262 16352
rect 14198 16292 14202 16348
rect 14202 16292 14258 16348
rect 14258 16292 14262 16348
rect 14198 16288 14262 16292
rect 17058 16348 17122 16352
rect 17058 16292 17062 16348
rect 17062 16292 17118 16348
rect 17118 16292 17122 16348
rect 17058 16288 17122 16292
rect 17138 16348 17202 16352
rect 17138 16292 17142 16348
rect 17142 16292 17198 16348
rect 17198 16292 17202 16348
rect 17138 16288 17202 16292
rect 17218 16348 17282 16352
rect 17218 16292 17222 16348
rect 17222 16292 17278 16348
rect 17278 16292 17282 16348
rect 17218 16288 17282 16292
rect 17298 16348 17362 16352
rect 17298 16292 17302 16348
rect 17302 16292 17358 16348
rect 17358 16292 17362 16348
rect 17298 16288 17362 16292
rect 3108 15804 3172 15808
rect 3108 15748 3112 15804
rect 3112 15748 3168 15804
rect 3168 15748 3172 15804
rect 3108 15744 3172 15748
rect 3188 15804 3252 15808
rect 3188 15748 3192 15804
rect 3192 15748 3248 15804
rect 3248 15748 3252 15804
rect 3188 15744 3252 15748
rect 3268 15804 3332 15808
rect 3268 15748 3272 15804
rect 3272 15748 3328 15804
rect 3328 15748 3332 15804
rect 3268 15744 3332 15748
rect 3348 15804 3412 15808
rect 3348 15748 3352 15804
rect 3352 15748 3408 15804
rect 3408 15748 3412 15804
rect 3348 15744 3412 15748
rect 6208 15804 6272 15808
rect 6208 15748 6212 15804
rect 6212 15748 6268 15804
rect 6268 15748 6272 15804
rect 6208 15744 6272 15748
rect 6288 15804 6352 15808
rect 6288 15748 6292 15804
rect 6292 15748 6348 15804
rect 6348 15748 6352 15804
rect 6288 15744 6352 15748
rect 6368 15804 6432 15808
rect 6368 15748 6372 15804
rect 6372 15748 6428 15804
rect 6428 15748 6432 15804
rect 6368 15744 6432 15748
rect 6448 15804 6512 15808
rect 6448 15748 6452 15804
rect 6452 15748 6508 15804
rect 6508 15748 6512 15804
rect 6448 15744 6512 15748
rect 9308 15804 9372 15808
rect 9308 15748 9312 15804
rect 9312 15748 9368 15804
rect 9368 15748 9372 15804
rect 9308 15744 9372 15748
rect 9388 15804 9452 15808
rect 9388 15748 9392 15804
rect 9392 15748 9448 15804
rect 9448 15748 9452 15804
rect 9388 15744 9452 15748
rect 9468 15804 9532 15808
rect 9468 15748 9472 15804
rect 9472 15748 9528 15804
rect 9528 15748 9532 15804
rect 9468 15744 9532 15748
rect 9548 15804 9612 15808
rect 9548 15748 9552 15804
rect 9552 15748 9608 15804
rect 9608 15748 9612 15804
rect 9548 15744 9612 15748
rect 12408 15804 12472 15808
rect 12408 15748 12412 15804
rect 12412 15748 12468 15804
rect 12468 15748 12472 15804
rect 12408 15744 12472 15748
rect 12488 15804 12552 15808
rect 12488 15748 12492 15804
rect 12492 15748 12548 15804
rect 12548 15748 12552 15804
rect 12488 15744 12552 15748
rect 12568 15804 12632 15808
rect 12568 15748 12572 15804
rect 12572 15748 12628 15804
rect 12628 15748 12632 15804
rect 12568 15744 12632 15748
rect 12648 15804 12712 15808
rect 12648 15748 12652 15804
rect 12652 15748 12708 15804
rect 12708 15748 12712 15804
rect 12648 15744 12712 15748
rect 15508 15804 15572 15808
rect 15508 15748 15512 15804
rect 15512 15748 15568 15804
rect 15568 15748 15572 15804
rect 15508 15744 15572 15748
rect 15588 15804 15652 15808
rect 15588 15748 15592 15804
rect 15592 15748 15648 15804
rect 15648 15748 15652 15804
rect 15588 15744 15652 15748
rect 15668 15804 15732 15808
rect 15668 15748 15672 15804
rect 15672 15748 15728 15804
rect 15728 15748 15732 15804
rect 15668 15744 15732 15748
rect 15748 15804 15812 15808
rect 15748 15748 15752 15804
rect 15752 15748 15808 15804
rect 15808 15748 15812 15804
rect 15748 15744 15812 15748
rect 18608 15804 18672 15808
rect 18608 15748 18612 15804
rect 18612 15748 18668 15804
rect 18668 15748 18672 15804
rect 18608 15744 18672 15748
rect 18688 15804 18752 15808
rect 18688 15748 18692 15804
rect 18692 15748 18748 15804
rect 18748 15748 18752 15804
rect 18688 15744 18752 15748
rect 18768 15804 18832 15808
rect 18768 15748 18772 15804
rect 18772 15748 18828 15804
rect 18828 15748 18832 15804
rect 18768 15744 18832 15748
rect 18848 15804 18912 15808
rect 18848 15748 18852 15804
rect 18852 15748 18908 15804
rect 18908 15748 18912 15804
rect 18848 15744 18912 15748
rect 1558 15260 1622 15264
rect 1558 15204 1562 15260
rect 1562 15204 1618 15260
rect 1618 15204 1622 15260
rect 1558 15200 1622 15204
rect 1638 15260 1702 15264
rect 1638 15204 1642 15260
rect 1642 15204 1698 15260
rect 1698 15204 1702 15260
rect 1638 15200 1702 15204
rect 1718 15260 1782 15264
rect 1718 15204 1722 15260
rect 1722 15204 1778 15260
rect 1778 15204 1782 15260
rect 1718 15200 1782 15204
rect 1798 15260 1862 15264
rect 1798 15204 1802 15260
rect 1802 15204 1858 15260
rect 1858 15204 1862 15260
rect 1798 15200 1862 15204
rect 4658 15260 4722 15264
rect 4658 15204 4662 15260
rect 4662 15204 4718 15260
rect 4718 15204 4722 15260
rect 4658 15200 4722 15204
rect 4738 15260 4802 15264
rect 4738 15204 4742 15260
rect 4742 15204 4798 15260
rect 4798 15204 4802 15260
rect 4738 15200 4802 15204
rect 4818 15260 4882 15264
rect 4818 15204 4822 15260
rect 4822 15204 4878 15260
rect 4878 15204 4882 15260
rect 4818 15200 4882 15204
rect 4898 15260 4962 15264
rect 4898 15204 4902 15260
rect 4902 15204 4958 15260
rect 4958 15204 4962 15260
rect 4898 15200 4962 15204
rect 7758 15260 7822 15264
rect 7758 15204 7762 15260
rect 7762 15204 7818 15260
rect 7818 15204 7822 15260
rect 7758 15200 7822 15204
rect 7838 15260 7902 15264
rect 7838 15204 7842 15260
rect 7842 15204 7898 15260
rect 7898 15204 7902 15260
rect 7838 15200 7902 15204
rect 7918 15260 7982 15264
rect 7918 15204 7922 15260
rect 7922 15204 7978 15260
rect 7978 15204 7982 15260
rect 7918 15200 7982 15204
rect 7998 15260 8062 15264
rect 7998 15204 8002 15260
rect 8002 15204 8058 15260
rect 8058 15204 8062 15260
rect 7998 15200 8062 15204
rect 10858 15260 10922 15264
rect 10858 15204 10862 15260
rect 10862 15204 10918 15260
rect 10918 15204 10922 15260
rect 10858 15200 10922 15204
rect 10938 15260 11002 15264
rect 10938 15204 10942 15260
rect 10942 15204 10998 15260
rect 10998 15204 11002 15260
rect 10938 15200 11002 15204
rect 11018 15260 11082 15264
rect 11018 15204 11022 15260
rect 11022 15204 11078 15260
rect 11078 15204 11082 15260
rect 11018 15200 11082 15204
rect 11098 15260 11162 15264
rect 11098 15204 11102 15260
rect 11102 15204 11158 15260
rect 11158 15204 11162 15260
rect 11098 15200 11162 15204
rect 13958 15260 14022 15264
rect 13958 15204 13962 15260
rect 13962 15204 14018 15260
rect 14018 15204 14022 15260
rect 13958 15200 14022 15204
rect 14038 15260 14102 15264
rect 14038 15204 14042 15260
rect 14042 15204 14098 15260
rect 14098 15204 14102 15260
rect 14038 15200 14102 15204
rect 14118 15260 14182 15264
rect 14118 15204 14122 15260
rect 14122 15204 14178 15260
rect 14178 15204 14182 15260
rect 14118 15200 14182 15204
rect 14198 15260 14262 15264
rect 14198 15204 14202 15260
rect 14202 15204 14258 15260
rect 14258 15204 14262 15260
rect 14198 15200 14262 15204
rect 17058 15260 17122 15264
rect 17058 15204 17062 15260
rect 17062 15204 17118 15260
rect 17118 15204 17122 15260
rect 17058 15200 17122 15204
rect 17138 15260 17202 15264
rect 17138 15204 17142 15260
rect 17142 15204 17198 15260
rect 17198 15204 17202 15260
rect 17138 15200 17202 15204
rect 17218 15260 17282 15264
rect 17218 15204 17222 15260
rect 17222 15204 17278 15260
rect 17278 15204 17282 15260
rect 17218 15200 17282 15204
rect 17298 15260 17362 15264
rect 17298 15204 17302 15260
rect 17302 15204 17358 15260
rect 17358 15204 17362 15260
rect 17298 15200 17362 15204
rect 3108 14716 3172 14720
rect 3108 14660 3112 14716
rect 3112 14660 3168 14716
rect 3168 14660 3172 14716
rect 3108 14656 3172 14660
rect 3188 14716 3252 14720
rect 3188 14660 3192 14716
rect 3192 14660 3248 14716
rect 3248 14660 3252 14716
rect 3188 14656 3252 14660
rect 3268 14716 3332 14720
rect 3268 14660 3272 14716
rect 3272 14660 3328 14716
rect 3328 14660 3332 14716
rect 3268 14656 3332 14660
rect 3348 14716 3412 14720
rect 3348 14660 3352 14716
rect 3352 14660 3408 14716
rect 3408 14660 3412 14716
rect 3348 14656 3412 14660
rect 6208 14716 6272 14720
rect 6208 14660 6212 14716
rect 6212 14660 6268 14716
rect 6268 14660 6272 14716
rect 6208 14656 6272 14660
rect 6288 14716 6352 14720
rect 6288 14660 6292 14716
rect 6292 14660 6348 14716
rect 6348 14660 6352 14716
rect 6288 14656 6352 14660
rect 6368 14716 6432 14720
rect 6368 14660 6372 14716
rect 6372 14660 6428 14716
rect 6428 14660 6432 14716
rect 6368 14656 6432 14660
rect 6448 14716 6512 14720
rect 6448 14660 6452 14716
rect 6452 14660 6508 14716
rect 6508 14660 6512 14716
rect 6448 14656 6512 14660
rect 9308 14716 9372 14720
rect 9308 14660 9312 14716
rect 9312 14660 9368 14716
rect 9368 14660 9372 14716
rect 9308 14656 9372 14660
rect 9388 14716 9452 14720
rect 9388 14660 9392 14716
rect 9392 14660 9448 14716
rect 9448 14660 9452 14716
rect 9388 14656 9452 14660
rect 9468 14716 9532 14720
rect 9468 14660 9472 14716
rect 9472 14660 9528 14716
rect 9528 14660 9532 14716
rect 9468 14656 9532 14660
rect 9548 14716 9612 14720
rect 9548 14660 9552 14716
rect 9552 14660 9608 14716
rect 9608 14660 9612 14716
rect 9548 14656 9612 14660
rect 12408 14716 12472 14720
rect 12408 14660 12412 14716
rect 12412 14660 12468 14716
rect 12468 14660 12472 14716
rect 12408 14656 12472 14660
rect 12488 14716 12552 14720
rect 12488 14660 12492 14716
rect 12492 14660 12548 14716
rect 12548 14660 12552 14716
rect 12488 14656 12552 14660
rect 12568 14716 12632 14720
rect 12568 14660 12572 14716
rect 12572 14660 12628 14716
rect 12628 14660 12632 14716
rect 12568 14656 12632 14660
rect 12648 14716 12712 14720
rect 12648 14660 12652 14716
rect 12652 14660 12708 14716
rect 12708 14660 12712 14716
rect 12648 14656 12712 14660
rect 15508 14716 15572 14720
rect 15508 14660 15512 14716
rect 15512 14660 15568 14716
rect 15568 14660 15572 14716
rect 15508 14656 15572 14660
rect 15588 14716 15652 14720
rect 15588 14660 15592 14716
rect 15592 14660 15648 14716
rect 15648 14660 15652 14716
rect 15588 14656 15652 14660
rect 15668 14716 15732 14720
rect 15668 14660 15672 14716
rect 15672 14660 15728 14716
rect 15728 14660 15732 14716
rect 15668 14656 15732 14660
rect 15748 14716 15812 14720
rect 15748 14660 15752 14716
rect 15752 14660 15808 14716
rect 15808 14660 15812 14716
rect 15748 14656 15812 14660
rect 18608 14716 18672 14720
rect 18608 14660 18612 14716
rect 18612 14660 18668 14716
rect 18668 14660 18672 14716
rect 18608 14656 18672 14660
rect 18688 14716 18752 14720
rect 18688 14660 18692 14716
rect 18692 14660 18748 14716
rect 18748 14660 18752 14716
rect 18688 14656 18752 14660
rect 18768 14716 18832 14720
rect 18768 14660 18772 14716
rect 18772 14660 18828 14716
rect 18828 14660 18832 14716
rect 18768 14656 18832 14660
rect 18848 14716 18912 14720
rect 18848 14660 18852 14716
rect 18852 14660 18908 14716
rect 18908 14660 18912 14716
rect 18848 14656 18912 14660
rect 1558 14172 1622 14176
rect 1558 14116 1562 14172
rect 1562 14116 1618 14172
rect 1618 14116 1622 14172
rect 1558 14112 1622 14116
rect 1638 14172 1702 14176
rect 1638 14116 1642 14172
rect 1642 14116 1698 14172
rect 1698 14116 1702 14172
rect 1638 14112 1702 14116
rect 1718 14172 1782 14176
rect 1718 14116 1722 14172
rect 1722 14116 1778 14172
rect 1778 14116 1782 14172
rect 1718 14112 1782 14116
rect 1798 14172 1862 14176
rect 1798 14116 1802 14172
rect 1802 14116 1858 14172
rect 1858 14116 1862 14172
rect 1798 14112 1862 14116
rect 4658 14172 4722 14176
rect 4658 14116 4662 14172
rect 4662 14116 4718 14172
rect 4718 14116 4722 14172
rect 4658 14112 4722 14116
rect 4738 14172 4802 14176
rect 4738 14116 4742 14172
rect 4742 14116 4798 14172
rect 4798 14116 4802 14172
rect 4738 14112 4802 14116
rect 4818 14172 4882 14176
rect 4818 14116 4822 14172
rect 4822 14116 4878 14172
rect 4878 14116 4882 14172
rect 4818 14112 4882 14116
rect 4898 14172 4962 14176
rect 4898 14116 4902 14172
rect 4902 14116 4958 14172
rect 4958 14116 4962 14172
rect 4898 14112 4962 14116
rect 7758 14172 7822 14176
rect 7758 14116 7762 14172
rect 7762 14116 7818 14172
rect 7818 14116 7822 14172
rect 7758 14112 7822 14116
rect 7838 14172 7902 14176
rect 7838 14116 7842 14172
rect 7842 14116 7898 14172
rect 7898 14116 7902 14172
rect 7838 14112 7902 14116
rect 7918 14172 7982 14176
rect 7918 14116 7922 14172
rect 7922 14116 7978 14172
rect 7978 14116 7982 14172
rect 7918 14112 7982 14116
rect 7998 14172 8062 14176
rect 7998 14116 8002 14172
rect 8002 14116 8058 14172
rect 8058 14116 8062 14172
rect 7998 14112 8062 14116
rect 10858 14172 10922 14176
rect 10858 14116 10862 14172
rect 10862 14116 10918 14172
rect 10918 14116 10922 14172
rect 10858 14112 10922 14116
rect 10938 14172 11002 14176
rect 10938 14116 10942 14172
rect 10942 14116 10998 14172
rect 10998 14116 11002 14172
rect 10938 14112 11002 14116
rect 11018 14172 11082 14176
rect 11018 14116 11022 14172
rect 11022 14116 11078 14172
rect 11078 14116 11082 14172
rect 11018 14112 11082 14116
rect 11098 14172 11162 14176
rect 11098 14116 11102 14172
rect 11102 14116 11158 14172
rect 11158 14116 11162 14172
rect 11098 14112 11162 14116
rect 13958 14172 14022 14176
rect 13958 14116 13962 14172
rect 13962 14116 14018 14172
rect 14018 14116 14022 14172
rect 13958 14112 14022 14116
rect 14038 14172 14102 14176
rect 14038 14116 14042 14172
rect 14042 14116 14098 14172
rect 14098 14116 14102 14172
rect 14038 14112 14102 14116
rect 14118 14172 14182 14176
rect 14118 14116 14122 14172
rect 14122 14116 14178 14172
rect 14178 14116 14182 14172
rect 14118 14112 14182 14116
rect 14198 14172 14262 14176
rect 14198 14116 14202 14172
rect 14202 14116 14258 14172
rect 14258 14116 14262 14172
rect 14198 14112 14262 14116
rect 17058 14172 17122 14176
rect 17058 14116 17062 14172
rect 17062 14116 17118 14172
rect 17118 14116 17122 14172
rect 17058 14112 17122 14116
rect 17138 14172 17202 14176
rect 17138 14116 17142 14172
rect 17142 14116 17198 14172
rect 17198 14116 17202 14172
rect 17138 14112 17202 14116
rect 17218 14172 17282 14176
rect 17218 14116 17222 14172
rect 17222 14116 17278 14172
rect 17278 14116 17282 14172
rect 17218 14112 17282 14116
rect 17298 14172 17362 14176
rect 17298 14116 17302 14172
rect 17302 14116 17358 14172
rect 17358 14116 17362 14172
rect 17298 14112 17362 14116
rect 3108 13628 3172 13632
rect 3108 13572 3112 13628
rect 3112 13572 3168 13628
rect 3168 13572 3172 13628
rect 3108 13568 3172 13572
rect 3188 13628 3252 13632
rect 3188 13572 3192 13628
rect 3192 13572 3248 13628
rect 3248 13572 3252 13628
rect 3188 13568 3252 13572
rect 3268 13628 3332 13632
rect 3268 13572 3272 13628
rect 3272 13572 3328 13628
rect 3328 13572 3332 13628
rect 3268 13568 3332 13572
rect 3348 13628 3412 13632
rect 3348 13572 3352 13628
rect 3352 13572 3408 13628
rect 3408 13572 3412 13628
rect 3348 13568 3412 13572
rect 6208 13628 6272 13632
rect 6208 13572 6212 13628
rect 6212 13572 6268 13628
rect 6268 13572 6272 13628
rect 6208 13568 6272 13572
rect 6288 13628 6352 13632
rect 6288 13572 6292 13628
rect 6292 13572 6348 13628
rect 6348 13572 6352 13628
rect 6288 13568 6352 13572
rect 6368 13628 6432 13632
rect 6368 13572 6372 13628
rect 6372 13572 6428 13628
rect 6428 13572 6432 13628
rect 6368 13568 6432 13572
rect 6448 13628 6512 13632
rect 6448 13572 6452 13628
rect 6452 13572 6508 13628
rect 6508 13572 6512 13628
rect 6448 13568 6512 13572
rect 9308 13628 9372 13632
rect 9308 13572 9312 13628
rect 9312 13572 9368 13628
rect 9368 13572 9372 13628
rect 9308 13568 9372 13572
rect 9388 13628 9452 13632
rect 9388 13572 9392 13628
rect 9392 13572 9448 13628
rect 9448 13572 9452 13628
rect 9388 13568 9452 13572
rect 9468 13628 9532 13632
rect 9468 13572 9472 13628
rect 9472 13572 9528 13628
rect 9528 13572 9532 13628
rect 9468 13568 9532 13572
rect 9548 13628 9612 13632
rect 9548 13572 9552 13628
rect 9552 13572 9608 13628
rect 9608 13572 9612 13628
rect 9548 13568 9612 13572
rect 12408 13628 12472 13632
rect 12408 13572 12412 13628
rect 12412 13572 12468 13628
rect 12468 13572 12472 13628
rect 12408 13568 12472 13572
rect 12488 13628 12552 13632
rect 12488 13572 12492 13628
rect 12492 13572 12548 13628
rect 12548 13572 12552 13628
rect 12488 13568 12552 13572
rect 12568 13628 12632 13632
rect 12568 13572 12572 13628
rect 12572 13572 12628 13628
rect 12628 13572 12632 13628
rect 12568 13568 12632 13572
rect 12648 13628 12712 13632
rect 12648 13572 12652 13628
rect 12652 13572 12708 13628
rect 12708 13572 12712 13628
rect 12648 13568 12712 13572
rect 15508 13628 15572 13632
rect 15508 13572 15512 13628
rect 15512 13572 15568 13628
rect 15568 13572 15572 13628
rect 15508 13568 15572 13572
rect 15588 13628 15652 13632
rect 15588 13572 15592 13628
rect 15592 13572 15648 13628
rect 15648 13572 15652 13628
rect 15588 13568 15652 13572
rect 15668 13628 15732 13632
rect 15668 13572 15672 13628
rect 15672 13572 15728 13628
rect 15728 13572 15732 13628
rect 15668 13568 15732 13572
rect 15748 13628 15812 13632
rect 15748 13572 15752 13628
rect 15752 13572 15808 13628
rect 15808 13572 15812 13628
rect 15748 13568 15812 13572
rect 18608 13628 18672 13632
rect 18608 13572 18612 13628
rect 18612 13572 18668 13628
rect 18668 13572 18672 13628
rect 18608 13568 18672 13572
rect 18688 13628 18752 13632
rect 18688 13572 18692 13628
rect 18692 13572 18748 13628
rect 18748 13572 18752 13628
rect 18688 13568 18752 13572
rect 18768 13628 18832 13632
rect 18768 13572 18772 13628
rect 18772 13572 18828 13628
rect 18828 13572 18832 13628
rect 18768 13568 18832 13572
rect 18848 13628 18912 13632
rect 18848 13572 18852 13628
rect 18852 13572 18908 13628
rect 18908 13572 18912 13628
rect 18848 13568 18912 13572
rect 1558 13084 1622 13088
rect 1558 13028 1562 13084
rect 1562 13028 1618 13084
rect 1618 13028 1622 13084
rect 1558 13024 1622 13028
rect 1638 13084 1702 13088
rect 1638 13028 1642 13084
rect 1642 13028 1698 13084
rect 1698 13028 1702 13084
rect 1638 13024 1702 13028
rect 1718 13084 1782 13088
rect 1718 13028 1722 13084
rect 1722 13028 1778 13084
rect 1778 13028 1782 13084
rect 1718 13024 1782 13028
rect 1798 13084 1862 13088
rect 1798 13028 1802 13084
rect 1802 13028 1858 13084
rect 1858 13028 1862 13084
rect 1798 13024 1862 13028
rect 4658 13084 4722 13088
rect 4658 13028 4662 13084
rect 4662 13028 4718 13084
rect 4718 13028 4722 13084
rect 4658 13024 4722 13028
rect 4738 13084 4802 13088
rect 4738 13028 4742 13084
rect 4742 13028 4798 13084
rect 4798 13028 4802 13084
rect 4738 13024 4802 13028
rect 4818 13084 4882 13088
rect 4818 13028 4822 13084
rect 4822 13028 4878 13084
rect 4878 13028 4882 13084
rect 4818 13024 4882 13028
rect 4898 13084 4962 13088
rect 4898 13028 4902 13084
rect 4902 13028 4958 13084
rect 4958 13028 4962 13084
rect 4898 13024 4962 13028
rect 7758 13084 7822 13088
rect 7758 13028 7762 13084
rect 7762 13028 7818 13084
rect 7818 13028 7822 13084
rect 7758 13024 7822 13028
rect 7838 13084 7902 13088
rect 7838 13028 7842 13084
rect 7842 13028 7898 13084
rect 7898 13028 7902 13084
rect 7838 13024 7902 13028
rect 7918 13084 7982 13088
rect 7918 13028 7922 13084
rect 7922 13028 7978 13084
rect 7978 13028 7982 13084
rect 7918 13024 7982 13028
rect 7998 13084 8062 13088
rect 7998 13028 8002 13084
rect 8002 13028 8058 13084
rect 8058 13028 8062 13084
rect 7998 13024 8062 13028
rect 10858 13084 10922 13088
rect 10858 13028 10862 13084
rect 10862 13028 10918 13084
rect 10918 13028 10922 13084
rect 10858 13024 10922 13028
rect 10938 13084 11002 13088
rect 10938 13028 10942 13084
rect 10942 13028 10998 13084
rect 10998 13028 11002 13084
rect 10938 13024 11002 13028
rect 11018 13084 11082 13088
rect 11018 13028 11022 13084
rect 11022 13028 11078 13084
rect 11078 13028 11082 13084
rect 11018 13024 11082 13028
rect 11098 13084 11162 13088
rect 11098 13028 11102 13084
rect 11102 13028 11158 13084
rect 11158 13028 11162 13084
rect 11098 13024 11162 13028
rect 13958 13084 14022 13088
rect 13958 13028 13962 13084
rect 13962 13028 14018 13084
rect 14018 13028 14022 13084
rect 13958 13024 14022 13028
rect 14038 13084 14102 13088
rect 14038 13028 14042 13084
rect 14042 13028 14098 13084
rect 14098 13028 14102 13084
rect 14038 13024 14102 13028
rect 14118 13084 14182 13088
rect 14118 13028 14122 13084
rect 14122 13028 14178 13084
rect 14178 13028 14182 13084
rect 14118 13024 14182 13028
rect 14198 13084 14262 13088
rect 14198 13028 14202 13084
rect 14202 13028 14258 13084
rect 14258 13028 14262 13084
rect 14198 13024 14262 13028
rect 17058 13084 17122 13088
rect 17058 13028 17062 13084
rect 17062 13028 17118 13084
rect 17118 13028 17122 13084
rect 17058 13024 17122 13028
rect 17138 13084 17202 13088
rect 17138 13028 17142 13084
rect 17142 13028 17198 13084
rect 17198 13028 17202 13084
rect 17138 13024 17202 13028
rect 17218 13084 17282 13088
rect 17218 13028 17222 13084
rect 17222 13028 17278 13084
rect 17278 13028 17282 13084
rect 17218 13024 17282 13028
rect 17298 13084 17362 13088
rect 17298 13028 17302 13084
rect 17302 13028 17358 13084
rect 17358 13028 17362 13084
rect 17298 13024 17362 13028
rect 3108 12540 3172 12544
rect 3108 12484 3112 12540
rect 3112 12484 3168 12540
rect 3168 12484 3172 12540
rect 3108 12480 3172 12484
rect 3188 12540 3252 12544
rect 3188 12484 3192 12540
rect 3192 12484 3248 12540
rect 3248 12484 3252 12540
rect 3188 12480 3252 12484
rect 3268 12540 3332 12544
rect 3268 12484 3272 12540
rect 3272 12484 3328 12540
rect 3328 12484 3332 12540
rect 3268 12480 3332 12484
rect 3348 12540 3412 12544
rect 3348 12484 3352 12540
rect 3352 12484 3408 12540
rect 3408 12484 3412 12540
rect 3348 12480 3412 12484
rect 6208 12540 6272 12544
rect 6208 12484 6212 12540
rect 6212 12484 6268 12540
rect 6268 12484 6272 12540
rect 6208 12480 6272 12484
rect 6288 12540 6352 12544
rect 6288 12484 6292 12540
rect 6292 12484 6348 12540
rect 6348 12484 6352 12540
rect 6288 12480 6352 12484
rect 6368 12540 6432 12544
rect 6368 12484 6372 12540
rect 6372 12484 6428 12540
rect 6428 12484 6432 12540
rect 6368 12480 6432 12484
rect 6448 12540 6512 12544
rect 6448 12484 6452 12540
rect 6452 12484 6508 12540
rect 6508 12484 6512 12540
rect 6448 12480 6512 12484
rect 9308 12540 9372 12544
rect 9308 12484 9312 12540
rect 9312 12484 9368 12540
rect 9368 12484 9372 12540
rect 9308 12480 9372 12484
rect 9388 12540 9452 12544
rect 9388 12484 9392 12540
rect 9392 12484 9448 12540
rect 9448 12484 9452 12540
rect 9388 12480 9452 12484
rect 9468 12540 9532 12544
rect 9468 12484 9472 12540
rect 9472 12484 9528 12540
rect 9528 12484 9532 12540
rect 9468 12480 9532 12484
rect 9548 12540 9612 12544
rect 9548 12484 9552 12540
rect 9552 12484 9608 12540
rect 9608 12484 9612 12540
rect 9548 12480 9612 12484
rect 12408 12540 12472 12544
rect 12408 12484 12412 12540
rect 12412 12484 12468 12540
rect 12468 12484 12472 12540
rect 12408 12480 12472 12484
rect 12488 12540 12552 12544
rect 12488 12484 12492 12540
rect 12492 12484 12548 12540
rect 12548 12484 12552 12540
rect 12488 12480 12552 12484
rect 12568 12540 12632 12544
rect 12568 12484 12572 12540
rect 12572 12484 12628 12540
rect 12628 12484 12632 12540
rect 12568 12480 12632 12484
rect 12648 12540 12712 12544
rect 12648 12484 12652 12540
rect 12652 12484 12708 12540
rect 12708 12484 12712 12540
rect 12648 12480 12712 12484
rect 15508 12540 15572 12544
rect 15508 12484 15512 12540
rect 15512 12484 15568 12540
rect 15568 12484 15572 12540
rect 15508 12480 15572 12484
rect 15588 12540 15652 12544
rect 15588 12484 15592 12540
rect 15592 12484 15648 12540
rect 15648 12484 15652 12540
rect 15588 12480 15652 12484
rect 15668 12540 15732 12544
rect 15668 12484 15672 12540
rect 15672 12484 15728 12540
rect 15728 12484 15732 12540
rect 15668 12480 15732 12484
rect 15748 12540 15812 12544
rect 15748 12484 15752 12540
rect 15752 12484 15808 12540
rect 15808 12484 15812 12540
rect 15748 12480 15812 12484
rect 18608 12540 18672 12544
rect 18608 12484 18612 12540
rect 18612 12484 18668 12540
rect 18668 12484 18672 12540
rect 18608 12480 18672 12484
rect 18688 12540 18752 12544
rect 18688 12484 18692 12540
rect 18692 12484 18748 12540
rect 18748 12484 18752 12540
rect 18688 12480 18752 12484
rect 18768 12540 18832 12544
rect 18768 12484 18772 12540
rect 18772 12484 18828 12540
rect 18828 12484 18832 12540
rect 18768 12480 18832 12484
rect 18848 12540 18912 12544
rect 18848 12484 18852 12540
rect 18852 12484 18908 12540
rect 18908 12484 18912 12540
rect 18848 12480 18912 12484
rect 1558 11996 1622 12000
rect 1558 11940 1562 11996
rect 1562 11940 1618 11996
rect 1618 11940 1622 11996
rect 1558 11936 1622 11940
rect 1638 11996 1702 12000
rect 1638 11940 1642 11996
rect 1642 11940 1698 11996
rect 1698 11940 1702 11996
rect 1638 11936 1702 11940
rect 1718 11996 1782 12000
rect 1718 11940 1722 11996
rect 1722 11940 1778 11996
rect 1778 11940 1782 11996
rect 1718 11936 1782 11940
rect 1798 11996 1862 12000
rect 1798 11940 1802 11996
rect 1802 11940 1858 11996
rect 1858 11940 1862 11996
rect 1798 11936 1862 11940
rect 4658 11996 4722 12000
rect 4658 11940 4662 11996
rect 4662 11940 4718 11996
rect 4718 11940 4722 11996
rect 4658 11936 4722 11940
rect 4738 11996 4802 12000
rect 4738 11940 4742 11996
rect 4742 11940 4798 11996
rect 4798 11940 4802 11996
rect 4738 11936 4802 11940
rect 4818 11996 4882 12000
rect 4818 11940 4822 11996
rect 4822 11940 4878 11996
rect 4878 11940 4882 11996
rect 4818 11936 4882 11940
rect 4898 11996 4962 12000
rect 4898 11940 4902 11996
rect 4902 11940 4958 11996
rect 4958 11940 4962 11996
rect 4898 11936 4962 11940
rect 7758 11996 7822 12000
rect 7758 11940 7762 11996
rect 7762 11940 7818 11996
rect 7818 11940 7822 11996
rect 7758 11936 7822 11940
rect 7838 11996 7902 12000
rect 7838 11940 7842 11996
rect 7842 11940 7898 11996
rect 7898 11940 7902 11996
rect 7838 11936 7902 11940
rect 7918 11996 7982 12000
rect 7918 11940 7922 11996
rect 7922 11940 7978 11996
rect 7978 11940 7982 11996
rect 7918 11936 7982 11940
rect 7998 11996 8062 12000
rect 7998 11940 8002 11996
rect 8002 11940 8058 11996
rect 8058 11940 8062 11996
rect 7998 11936 8062 11940
rect 10858 11996 10922 12000
rect 10858 11940 10862 11996
rect 10862 11940 10918 11996
rect 10918 11940 10922 11996
rect 10858 11936 10922 11940
rect 10938 11996 11002 12000
rect 10938 11940 10942 11996
rect 10942 11940 10998 11996
rect 10998 11940 11002 11996
rect 10938 11936 11002 11940
rect 11018 11996 11082 12000
rect 11018 11940 11022 11996
rect 11022 11940 11078 11996
rect 11078 11940 11082 11996
rect 11018 11936 11082 11940
rect 11098 11996 11162 12000
rect 11098 11940 11102 11996
rect 11102 11940 11158 11996
rect 11158 11940 11162 11996
rect 11098 11936 11162 11940
rect 13958 11996 14022 12000
rect 13958 11940 13962 11996
rect 13962 11940 14018 11996
rect 14018 11940 14022 11996
rect 13958 11936 14022 11940
rect 14038 11996 14102 12000
rect 14038 11940 14042 11996
rect 14042 11940 14098 11996
rect 14098 11940 14102 11996
rect 14038 11936 14102 11940
rect 14118 11996 14182 12000
rect 14118 11940 14122 11996
rect 14122 11940 14178 11996
rect 14178 11940 14182 11996
rect 14118 11936 14182 11940
rect 14198 11996 14262 12000
rect 14198 11940 14202 11996
rect 14202 11940 14258 11996
rect 14258 11940 14262 11996
rect 14198 11936 14262 11940
rect 17058 11996 17122 12000
rect 17058 11940 17062 11996
rect 17062 11940 17118 11996
rect 17118 11940 17122 11996
rect 17058 11936 17122 11940
rect 17138 11996 17202 12000
rect 17138 11940 17142 11996
rect 17142 11940 17198 11996
rect 17198 11940 17202 11996
rect 17138 11936 17202 11940
rect 17218 11996 17282 12000
rect 17218 11940 17222 11996
rect 17222 11940 17278 11996
rect 17278 11940 17282 11996
rect 17218 11936 17282 11940
rect 17298 11996 17362 12000
rect 17298 11940 17302 11996
rect 17302 11940 17358 11996
rect 17358 11940 17362 11996
rect 17298 11936 17362 11940
rect 3108 11452 3172 11456
rect 3108 11396 3112 11452
rect 3112 11396 3168 11452
rect 3168 11396 3172 11452
rect 3108 11392 3172 11396
rect 3188 11452 3252 11456
rect 3188 11396 3192 11452
rect 3192 11396 3248 11452
rect 3248 11396 3252 11452
rect 3188 11392 3252 11396
rect 3268 11452 3332 11456
rect 3268 11396 3272 11452
rect 3272 11396 3328 11452
rect 3328 11396 3332 11452
rect 3268 11392 3332 11396
rect 3348 11452 3412 11456
rect 3348 11396 3352 11452
rect 3352 11396 3408 11452
rect 3408 11396 3412 11452
rect 3348 11392 3412 11396
rect 6208 11452 6272 11456
rect 6208 11396 6212 11452
rect 6212 11396 6268 11452
rect 6268 11396 6272 11452
rect 6208 11392 6272 11396
rect 6288 11452 6352 11456
rect 6288 11396 6292 11452
rect 6292 11396 6348 11452
rect 6348 11396 6352 11452
rect 6288 11392 6352 11396
rect 6368 11452 6432 11456
rect 6368 11396 6372 11452
rect 6372 11396 6428 11452
rect 6428 11396 6432 11452
rect 6368 11392 6432 11396
rect 6448 11452 6512 11456
rect 6448 11396 6452 11452
rect 6452 11396 6508 11452
rect 6508 11396 6512 11452
rect 6448 11392 6512 11396
rect 9308 11452 9372 11456
rect 9308 11396 9312 11452
rect 9312 11396 9368 11452
rect 9368 11396 9372 11452
rect 9308 11392 9372 11396
rect 9388 11452 9452 11456
rect 9388 11396 9392 11452
rect 9392 11396 9448 11452
rect 9448 11396 9452 11452
rect 9388 11392 9452 11396
rect 9468 11452 9532 11456
rect 9468 11396 9472 11452
rect 9472 11396 9528 11452
rect 9528 11396 9532 11452
rect 9468 11392 9532 11396
rect 9548 11452 9612 11456
rect 9548 11396 9552 11452
rect 9552 11396 9608 11452
rect 9608 11396 9612 11452
rect 9548 11392 9612 11396
rect 12408 11452 12472 11456
rect 12408 11396 12412 11452
rect 12412 11396 12468 11452
rect 12468 11396 12472 11452
rect 12408 11392 12472 11396
rect 12488 11452 12552 11456
rect 12488 11396 12492 11452
rect 12492 11396 12548 11452
rect 12548 11396 12552 11452
rect 12488 11392 12552 11396
rect 12568 11452 12632 11456
rect 12568 11396 12572 11452
rect 12572 11396 12628 11452
rect 12628 11396 12632 11452
rect 12568 11392 12632 11396
rect 12648 11452 12712 11456
rect 12648 11396 12652 11452
rect 12652 11396 12708 11452
rect 12708 11396 12712 11452
rect 12648 11392 12712 11396
rect 15508 11452 15572 11456
rect 15508 11396 15512 11452
rect 15512 11396 15568 11452
rect 15568 11396 15572 11452
rect 15508 11392 15572 11396
rect 15588 11452 15652 11456
rect 15588 11396 15592 11452
rect 15592 11396 15648 11452
rect 15648 11396 15652 11452
rect 15588 11392 15652 11396
rect 15668 11452 15732 11456
rect 15668 11396 15672 11452
rect 15672 11396 15728 11452
rect 15728 11396 15732 11452
rect 15668 11392 15732 11396
rect 15748 11452 15812 11456
rect 15748 11396 15752 11452
rect 15752 11396 15808 11452
rect 15808 11396 15812 11452
rect 15748 11392 15812 11396
rect 18608 11452 18672 11456
rect 18608 11396 18612 11452
rect 18612 11396 18668 11452
rect 18668 11396 18672 11452
rect 18608 11392 18672 11396
rect 18688 11452 18752 11456
rect 18688 11396 18692 11452
rect 18692 11396 18748 11452
rect 18748 11396 18752 11452
rect 18688 11392 18752 11396
rect 18768 11452 18832 11456
rect 18768 11396 18772 11452
rect 18772 11396 18828 11452
rect 18828 11396 18832 11452
rect 18768 11392 18832 11396
rect 18848 11452 18912 11456
rect 18848 11396 18852 11452
rect 18852 11396 18908 11452
rect 18908 11396 18912 11452
rect 18848 11392 18912 11396
rect 1558 10908 1622 10912
rect 1558 10852 1562 10908
rect 1562 10852 1618 10908
rect 1618 10852 1622 10908
rect 1558 10848 1622 10852
rect 1638 10908 1702 10912
rect 1638 10852 1642 10908
rect 1642 10852 1698 10908
rect 1698 10852 1702 10908
rect 1638 10848 1702 10852
rect 1718 10908 1782 10912
rect 1718 10852 1722 10908
rect 1722 10852 1778 10908
rect 1778 10852 1782 10908
rect 1718 10848 1782 10852
rect 1798 10908 1862 10912
rect 1798 10852 1802 10908
rect 1802 10852 1858 10908
rect 1858 10852 1862 10908
rect 1798 10848 1862 10852
rect 4658 10908 4722 10912
rect 4658 10852 4662 10908
rect 4662 10852 4718 10908
rect 4718 10852 4722 10908
rect 4658 10848 4722 10852
rect 4738 10908 4802 10912
rect 4738 10852 4742 10908
rect 4742 10852 4798 10908
rect 4798 10852 4802 10908
rect 4738 10848 4802 10852
rect 4818 10908 4882 10912
rect 4818 10852 4822 10908
rect 4822 10852 4878 10908
rect 4878 10852 4882 10908
rect 4818 10848 4882 10852
rect 4898 10908 4962 10912
rect 4898 10852 4902 10908
rect 4902 10852 4958 10908
rect 4958 10852 4962 10908
rect 4898 10848 4962 10852
rect 7758 10908 7822 10912
rect 7758 10852 7762 10908
rect 7762 10852 7818 10908
rect 7818 10852 7822 10908
rect 7758 10848 7822 10852
rect 7838 10908 7902 10912
rect 7838 10852 7842 10908
rect 7842 10852 7898 10908
rect 7898 10852 7902 10908
rect 7838 10848 7902 10852
rect 7918 10908 7982 10912
rect 7918 10852 7922 10908
rect 7922 10852 7978 10908
rect 7978 10852 7982 10908
rect 7918 10848 7982 10852
rect 7998 10908 8062 10912
rect 7998 10852 8002 10908
rect 8002 10852 8058 10908
rect 8058 10852 8062 10908
rect 7998 10848 8062 10852
rect 10858 10908 10922 10912
rect 10858 10852 10862 10908
rect 10862 10852 10918 10908
rect 10918 10852 10922 10908
rect 10858 10848 10922 10852
rect 10938 10908 11002 10912
rect 10938 10852 10942 10908
rect 10942 10852 10998 10908
rect 10998 10852 11002 10908
rect 10938 10848 11002 10852
rect 11018 10908 11082 10912
rect 11018 10852 11022 10908
rect 11022 10852 11078 10908
rect 11078 10852 11082 10908
rect 11018 10848 11082 10852
rect 11098 10908 11162 10912
rect 11098 10852 11102 10908
rect 11102 10852 11158 10908
rect 11158 10852 11162 10908
rect 11098 10848 11162 10852
rect 13958 10908 14022 10912
rect 13958 10852 13962 10908
rect 13962 10852 14018 10908
rect 14018 10852 14022 10908
rect 13958 10848 14022 10852
rect 14038 10908 14102 10912
rect 14038 10852 14042 10908
rect 14042 10852 14098 10908
rect 14098 10852 14102 10908
rect 14038 10848 14102 10852
rect 14118 10908 14182 10912
rect 14118 10852 14122 10908
rect 14122 10852 14178 10908
rect 14178 10852 14182 10908
rect 14118 10848 14182 10852
rect 14198 10908 14262 10912
rect 14198 10852 14202 10908
rect 14202 10852 14258 10908
rect 14258 10852 14262 10908
rect 14198 10848 14262 10852
rect 17058 10908 17122 10912
rect 17058 10852 17062 10908
rect 17062 10852 17118 10908
rect 17118 10852 17122 10908
rect 17058 10848 17122 10852
rect 17138 10908 17202 10912
rect 17138 10852 17142 10908
rect 17142 10852 17198 10908
rect 17198 10852 17202 10908
rect 17138 10848 17202 10852
rect 17218 10908 17282 10912
rect 17218 10852 17222 10908
rect 17222 10852 17278 10908
rect 17278 10852 17282 10908
rect 17218 10848 17282 10852
rect 17298 10908 17362 10912
rect 17298 10852 17302 10908
rect 17302 10852 17358 10908
rect 17358 10852 17362 10908
rect 17298 10848 17362 10852
rect 3108 10364 3172 10368
rect 3108 10308 3112 10364
rect 3112 10308 3168 10364
rect 3168 10308 3172 10364
rect 3108 10304 3172 10308
rect 3188 10364 3252 10368
rect 3188 10308 3192 10364
rect 3192 10308 3248 10364
rect 3248 10308 3252 10364
rect 3188 10304 3252 10308
rect 3268 10364 3332 10368
rect 3268 10308 3272 10364
rect 3272 10308 3328 10364
rect 3328 10308 3332 10364
rect 3268 10304 3332 10308
rect 3348 10364 3412 10368
rect 3348 10308 3352 10364
rect 3352 10308 3408 10364
rect 3408 10308 3412 10364
rect 3348 10304 3412 10308
rect 6208 10364 6272 10368
rect 6208 10308 6212 10364
rect 6212 10308 6268 10364
rect 6268 10308 6272 10364
rect 6208 10304 6272 10308
rect 6288 10364 6352 10368
rect 6288 10308 6292 10364
rect 6292 10308 6348 10364
rect 6348 10308 6352 10364
rect 6288 10304 6352 10308
rect 6368 10364 6432 10368
rect 6368 10308 6372 10364
rect 6372 10308 6428 10364
rect 6428 10308 6432 10364
rect 6368 10304 6432 10308
rect 6448 10364 6512 10368
rect 6448 10308 6452 10364
rect 6452 10308 6508 10364
rect 6508 10308 6512 10364
rect 6448 10304 6512 10308
rect 9308 10364 9372 10368
rect 9308 10308 9312 10364
rect 9312 10308 9368 10364
rect 9368 10308 9372 10364
rect 9308 10304 9372 10308
rect 9388 10364 9452 10368
rect 9388 10308 9392 10364
rect 9392 10308 9448 10364
rect 9448 10308 9452 10364
rect 9388 10304 9452 10308
rect 9468 10364 9532 10368
rect 9468 10308 9472 10364
rect 9472 10308 9528 10364
rect 9528 10308 9532 10364
rect 9468 10304 9532 10308
rect 9548 10364 9612 10368
rect 9548 10308 9552 10364
rect 9552 10308 9608 10364
rect 9608 10308 9612 10364
rect 9548 10304 9612 10308
rect 12408 10364 12472 10368
rect 12408 10308 12412 10364
rect 12412 10308 12468 10364
rect 12468 10308 12472 10364
rect 12408 10304 12472 10308
rect 12488 10364 12552 10368
rect 12488 10308 12492 10364
rect 12492 10308 12548 10364
rect 12548 10308 12552 10364
rect 12488 10304 12552 10308
rect 12568 10364 12632 10368
rect 12568 10308 12572 10364
rect 12572 10308 12628 10364
rect 12628 10308 12632 10364
rect 12568 10304 12632 10308
rect 12648 10364 12712 10368
rect 12648 10308 12652 10364
rect 12652 10308 12708 10364
rect 12708 10308 12712 10364
rect 12648 10304 12712 10308
rect 15508 10364 15572 10368
rect 15508 10308 15512 10364
rect 15512 10308 15568 10364
rect 15568 10308 15572 10364
rect 15508 10304 15572 10308
rect 15588 10364 15652 10368
rect 15588 10308 15592 10364
rect 15592 10308 15648 10364
rect 15648 10308 15652 10364
rect 15588 10304 15652 10308
rect 15668 10364 15732 10368
rect 15668 10308 15672 10364
rect 15672 10308 15728 10364
rect 15728 10308 15732 10364
rect 15668 10304 15732 10308
rect 15748 10364 15812 10368
rect 15748 10308 15752 10364
rect 15752 10308 15808 10364
rect 15808 10308 15812 10364
rect 15748 10304 15812 10308
rect 18608 10364 18672 10368
rect 18608 10308 18612 10364
rect 18612 10308 18668 10364
rect 18668 10308 18672 10364
rect 18608 10304 18672 10308
rect 18688 10364 18752 10368
rect 18688 10308 18692 10364
rect 18692 10308 18748 10364
rect 18748 10308 18752 10364
rect 18688 10304 18752 10308
rect 18768 10364 18832 10368
rect 18768 10308 18772 10364
rect 18772 10308 18828 10364
rect 18828 10308 18832 10364
rect 18768 10304 18832 10308
rect 18848 10364 18912 10368
rect 18848 10308 18852 10364
rect 18852 10308 18908 10364
rect 18908 10308 18912 10364
rect 18848 10304 18912 10308
rect 1558 9820 1622 9824
rect 1558 9764 1562 9820
rect 1562 9764 1618 9820
rect 1618 9764 1622 9820
rect 1558 9760 1622 9764
rect 1638 9820 1702 9824
rect 1638 9764 1642 9820
rect 1642 9764 1698 9820
rect 1698 9764 1702 9820
rect 1638 9760 1702 9764
rect 1718 9820 1782 9824
rect 1718 9764 1722 9820
rect 1722 9764 1778 9820
rect 1778 9764 1782 9820
rect 1718 9760 1782 9764
rect 1798 9820 1862 9824
rect 1798 9764 1802 9820
rect 1802 9764 1858 9820
rect 1858 9764 1862 9820
rect 1798 9760 1862 9764
rect 4658 9820 4722 9824
rect 4658 9764 4662 9820
rect 4662 9764 4718 9820
rect 4718 9764 4722 9820
rect 4658 9760 4722 9764
rect 4738 9820 4802 9824
rect 4738 9764 4742 9820
rect 4742 9764 4798 9820
rect 4798 9764 4802 9820
rect 4738 9760 4802 9764
rect 4818 9820 4882 9824
rect 4818 9764 4822 9820
rect 4822 9764 4878 9820
rect 4878 9764 4882 9820
rect 4818 9760 4882 9764
rect 4898 9820 4962 9824
rect 4898 9764 4902 9820
rect 4902 9764 4958 9820
rect 4958 9764 4962 9820
rect 4898 9760 4962 9764
rect 7758 9820 7822 9824
rect 7758 9764 7762 9820
rect 7762 9764 7818 9820
rect 7818 9764 7822 9820
rect 7758 9760 7822 9764
rect 7838 9820 7902 9824
rect 7838 9764 7842 9820
rect 7842 9764 7898 9820
rect 7898 9764 7902 9820
rect 7838 9760 7902 9764
rect 7918 9820 7982 9824
rect 7918 9764 7922 9820
rect 7922 9764 7978 9820
rect 7978 9764 7982 9820
rect 7918 9760 7982 9764
rect 7998 9820 8062 9824
rect 7998 9764 8002 9820
rect 8002 9764 8058 9820
rect 8058 9764 8062 9820
rect 7998 9760 8062 9764
rect 10858 9820 10922 9824
rect 10858 9764 10862 9820
rect 10862 9764 10918 9820
rect 10918 9764 10922 9820
rect 10858 9760 10922 9764
rect 10938 9820 11002 9824
rect 10938 9764 10942 9820
rect 10942 9764 10998 9820
rect 10998 9764 11002 9820
rect 10938 9760 11002 9764
rect 11018 9820 11082 9824
rect 11018 9764 11022 9820
rect 11022 9764 11078 9820
rect 11078 9764 11082 9820
rect 11018 9760 11082 9764
rect 11098 9820 11162 9824
rect 11098 9764 11102 9820
rect 11102 9764 11158 9820
rect 11158 9764 11162 9820
rect 11098 9760 11162 9764
rect 13958 9820 14022 9824
rect 13958 9764 13962 9820
rect 13962 9764 14018 9820
rect 14018 9764 14022 9820
rect 13958 9760 14022 9764
rect 14038 9820 14102 9824
rect 14038 9764 14042 9820
rect 14042 9764 14098 9820
rect 14098 9764 14102 9820
rect 14038 9760 14102 9764
rect 14118 9820 14182 9824
rect 14118 9764 14122 9820
rect 14122 9764 14178 9820
rect 14178 9764 14182 9820
rect 14118 9760 14182 9764
rect 14198 9820 14262 9824
rect 14198 9764 14202 9820
rect 14202 9764 14258 9820
rect 14258 9764 14262 9820
rect 14198 9760 14262 9764
rect 17058 9820 17122 9824
rect 17058 9764 17062 9820
rect 17062 9764 17118 9820
rect 17118 9764 17122 9820
rect 17058 9760 17122 9764
rect 17138 9820 17202 9824
rect 17138 9764 17142 9820
rect 17142 9764 17198 9820
rect 17198 9764 17202 9820
rect 17138 9760 17202 9764
rect 17218 9820 17282 9824
rect 17218 9764 17222 9820
rect 17222 9764 17278 9820
rect 17278 9764 17282 9820
rect 17218 9760 17282 9764
rect 17298 9820 17362 9824
rect 17298 9764 17302 9820
rect 17302 9764 17358 9820
rect 17358 9764 17362 9820
rect 17298 9760 17362 9764
rect 3108 9276 3172 9280
rect 3108 9220 3112 9276
rect 3112 9220 3168 9276
rect 3168 9220 3172 9276
rect 3108 9216 3172 9220
rect 3188 9276 3252 9280
rect 3188 9220 3192 9276
rect 3192 9220 3248 9276
rect 3248 9220 3252 9276
rect 3188 9216 3252 9220
rect 3268 9276 3332 9280
rect 3268 9220 3272 9276
rect 3272 9220 3328 9276
rect 3328 9220 3332 9276
rect 3268 9216 3332 9220
rect 3348 9276 3412 9280
rect 3348 9220 3352 9276
rect 3352 9220 3408 9276
rect 3408 9220 3412 9276
rect 3348 9216 3412 9220
rect 6208 9276 6272 9280
rect 6208 9220 6212 9276
rect 6212 9220 6268 9276
rect 6268 9220 6272 9276
rect 6208 9216 6272 9220
rect 6288 9276 6352 9280
rect 6288 9220 6292 9276
rect 6292 9220 6348 9276
rect 6348 9220 6352 9276
rect 6288 9216 6352 9220
rect 6368 9276 6432 9280
rect 6368 9220 6372 9276
rect 6372 9220 6428 9276
rect 6428 9220 6432 9276
rect 6368 9216 6432 9220
rect 6448 9276 6512 9280
rect 6448 9220 6452 9276
rect 6452 9220 6508 9276
rect 6508 9220 6512 9276
rect 6448 9216 6512 9220
rect 9308 9276 9372 9280
rect 9308 9220 9312 9276
rect 9312 9220 9368 9276
rect 9368 9220 9372 9276
rect 9308 9216 9372 9220
rect 9388 9276 9452 9280
rect 9388 9220 9392 9276
rect 9392 9220 9448 9276
rect 9448 9220 9452 9276
rect 9388 9216 9452 9220
rect 9468 9276 9532 9280
rect 9468 9220 9472 9276
rect 9472 9220 9528 9276
rect 9528 9220 9532 9276
rect 9468 9216 9532 9220
rect 9548 9276 9612 9280
rect 9548 9220 9552 9276
rect 9552 9220 9608 9276
rect 9608 9220 9612 9276
rect 9548 9216 9612 9220
rect 12408 9276 12472 9280
rect 12408 9220 12412 9276
rect 12412 9220 12468 9276
rect 12468 9220 12472 9276
rect 12408 9216 12472 9220
rect 12488 9276 12552 9280
rect 12488 9220 12492 9276
rect 12492 9220 12548 9276
rect 12548 9220 12552 9276
rect 12488 9216 12552 9220
rect 12568 9276 12632 9280
rect 12568 9220 12572 9276
rect 12572 9220 12628 9276
rect 12628 9220 12632 9276
rect 12568 9216 12632 9220
rect 12648 9276 12712 9280
rect 12648 9220 12652 9276
rect 12652 9220 12708 9276
rect 12708 9220 12712 9276
rect 12648 9216 12712 9220
rect 15508 9276 15572 9280
rect 15508 9220 15512 9276
rect 15512 9220 15568 9276
rect 15568 9220 15572 9276
rect 15508 9216 15572 9220
rect 15588 9276 15652 9280
rect 15588 9220 15592 9276
rect 15592 9220 15648 9276
rect 15648 9220 15652 9276
rect 15588 9216 15652 9220
rect 15668 9276 15732 9280
rect 15668 9220 15672 9276
rect 15672 9220 15728 9276
rect 15728 9220 15732 9276
rect 15668 9216 15732 9220
rect 15748 9276 15812 9280
rect 15748 9220 15752 9276
rect 15752 9220 15808 9276
rect 15808 9220 15812 9276
rect 15748 9216 15812 9220
rect 18608 9276 18672 9280
rect 18608 9220 18612 9276
rect 18612 9220 18668 9276
rect 18668 9220 18672 9276
rect 18608 9216 18672 9220
rect 18688 9276 18752 9280
rect 18688 9220 18692 9276
rect 18692 9220 18748 9276
rect 18748 9220 18752 9276
rect 18688 9216 18752 9220
rect 18768 9276 18832 9280
rect 18768 9220 18772 9276
rect 18772 9220 18828 9276
rect 18828 9220 18832 9276
rect 18768 9216 18832 9220
rect 18848 9276 18912 9280
rect 18848 9220 18852 9276
rect 18852 9220 18908 9276
rect 18908 9220 18912 9276
rect 18848 9216 18912 9220
rect 1558 8732 1622 8736
rect 1558 8676 1562 8732
rect 1562 8676 1618 8732
rect 1618 8676 1622 8732
rect 1558 8672 1622 8676
rect 1638 8732 1702 8736
rect 1638 8676 1642 8732
rect 1642 8676 1698 8732
rect 1698 8676 1702 8732
rect 1638 8672 1702 8676
rect 1718 8732 1782 8736
rect 1718 8676 1722 8732
rect 1722 8676 1778 8732
rect 1778 8676 1782 8732
rect 1718 8672 1782 8676
rect 1798 8732 1862 8736
rect 1798 8676 1802 8732
rect 1802 8676 1858 8732
rect 1858 8676 1862 8732
rect 1798 8672 1862 8676
rect 4658 8732 4722 8736
rect 4658 8676 4662 8732
rect 4662 8676 4718 8732
rect 4718 8676 4722 8732
rect 4658 8672 4722 8676
rect 4738 8732 4802 8736
rect 4738 8676 4742 8732
rect 4742 8676 4798 8732
rect 4798 8676 4802 8732
rect 4738 8672 4802 8676
rect 4818 8732 4882 8736
rect 4818 8676 4822 8732
rect 4822 8676 4878 8732
rect 4878 8676 4882 8732
rect 4818 8672 4882 8676
rect 4898 8732 4962 8736
rect 4898 8676 4902 8732
rect 4902 8676 4958 8732
rect 4958 8676 4962 8732
rect 4898 8672 4962 8676
rect 7758 8732 7822 8736
rect 7758 8676 7762 8732
rect 7762 8676 7818 8732
rect 7818 8676 7822 8732
rect 7758 8672 7822 8676
rect 7838 8732 7902 8736
rect 7838 8676 7842 8732
rect 7842 8676 7898 8732
rect 7898 8676 7902 8732
rect 7838 8672 7902 8676
rect 7918 8732 7982 8736
rect 7918 8676 7922 8732
rect 7922 8676 7978 8732
rect 7978 8676 7982 8732
rect 7918 8672 7982 8676
rect 7998 8732 8062 8736
rect 7998 8676 8002 8732
rect 8002 8676 8058 8732
rect 8058 8676 8062 8732
rect 7998 8672 8062 8676
rect 10858 8732 10922 8736
rect 10858 8676 10862 8732
rect 10862 8676 10918 8732
rect 10918 8676 10922 8732
rect 10858 8672 10922 8676
rect 10938 8732 11002 8736
rect 10938 8676 10942 8732
rect 10942 8676 10998 8732
rect 10998 8676 11002 8732
rect 10938 8672 11002 8676
rect 11018 8732 11082 8736
rect 11018 8676 11022 8732
rect 11022 8676 11078 8732
rect 11078 8676 11082 8732
rect 11018 8672 11082 8676
rect 11098 8732 11162 8736
rect 11098 8676 11102 8732
rect 11102 8676 11158 8732
rect 11158 8676 11162 8732
rect 11098 8672 11162 8676
rect 13958 8732 14022 8736
rect 13958 8676 13962 8732
rect 13962 8676 14018 8732
rect 14018 8676 14022 8732
rect 13958 8672 14022 8676
rect 14038 8732 14102 8736
rect 14038 8676 14042 8732
rect 14042 8676 14098 8732
rect 14098 8676 14102 8732
rect 14038 8672 14102 8676
rect 14118 8732 14182 8736
rect 14118 8676 14122 8732
rect 14122 8676 14178 8732
rect 14178 8676 14182 8732
rect 14118 8672 14182 8676
rect 14198 8732 14262 8736
rect 14198 8676 14202 8732
rect 14202 8676 14258 8732
rect 14258 8676 14262 8732
rect 14198 8672 14262 8676
rect 17058 8732 17122 8736
rect 17058 8676 17062 8732
rect 17062 8676 17118 8732
rect 17118 8676 17122 8732
rect 17058 8672 17122 8676
rect 17138 8732 17202 8736
rect 17138 8676 17142 8732
rect 17142 8676 17198 8732
rect 17198 8676 17202 8732
rect 17138 8672 17202 8676
rect 17218 8732 17282 8736
rect 17218 8676 17222 8732
rect 17222 8676 17278 8732
rect 17278 8676 17282 8732
rect 17218 8672 17282 8676
rect 17298 8732 17362 8736
rect 17298 8676 17302 8732
rect 17302 8676 17358 8732
rect 17358 8676 17362 8732
rect 17298 8672 17362 8676
rect 3108 8188 3172 8192
rect 3108 8132 3112 8188
rect 3112 8132 3168 8188
rect 3168 8132 3172 8188
rect 3108 8128 3172 8132
rect 3188 8188 3252 8192
rect 3188 8132 3192 8188
rect 3192 8132 3248 8188
rect 3248 8132 3252 8188
rect 3188 8128 3252 8132
rect 3268 8188 3332 8192
rect 3268 8132 3272 8188
rect 3272 8132 3328 8188
rect 3328 8132 3332 8188
rect 3268 8128 3332 8132
rect 3348 8188 3412 8192
rect 3348 8132 3352 8188
rect 3352 8132 3408 8188
rect 3408 8132 3412 8188
rect 3348 8128 3412 8132
rect 6208 8188 6272 8192
rect 6208 8132 6212 8188
rect 6212 8132 6268 8188
rect 6268 8132 6272 8188
rect 6208 8128 6272 8132
rect 6288 8188 6352 8192
rect 6288 8132 6292 8188
rect 6292 8132 6348 8188
rect 6348 8132 6352 8188
rect 6288 8128 6352 8132
rect 6368 8188 6432 8192
rect 6368 8132 6372 8188
rect 6372 8132 6428 8188
rect 6428 8132 6432 8188
rect 6368 8128 6432 8132
rect 6448 8188 6512 8192
rect 6448 8132 6452 8188
rect 6452 8132 6508 8188
rect 6508 8132 6512 8188
rect 6448 8128 6512 8132
rect 9308 8188 9372 8192
rect 9308 8132 9312 8188
rect 9312 8132 9368 8188
rect 9368 8132 9372 8188
rect 9308 8128 9372 8132
rect 9388 8188 9452 8192
rect 9388 8132 9392 8188
rect 9392 8132 9448 8188
rect 9448 8132 9452 8188
rect 9388 8128 9452 8132
rect 9468 8188 9532 8192
rect 9468 8132 9472 8188
rect 9472 8132 9528 8188
rect 9528 8132 9532 8188
rect 9468 8128 9532 8132
rect 9548 8188 9612 8192
rect 9548 8132 9552 8188
rect 9552 8132 9608 8188
rect 9608 8132 9612 8188
rect 9548 8128 9612 8132
rect 12408 8188 12472 8192
rect 12408 8132 12412 8188
rect 12412 8132 12468 8188
rect 12468 8132 12472 8188
rect 12408 8128 12472 8132
rect 12488 8188 12552 8192
rect 12488 8132 12492 8188
rect 12492 8132 12548 8188
rect 12548 8132 12552 8188
rect 12488 8128 12552 8132
rect 12568 8188 12632 8192
rect 12568 8132 12572 8188
rect 12572 8132 12628 8188
rect 12628 8132 12632 8188
rect 12568 8128 12632 8132
rect 12648 8188 12712 8192
rect 12648 8132 12652 8188
rect 12652 8132 12708 8188
rect 12708 8132 12712 8188
rect 12648 8128 12712 8132
rect 15508 8188 15572 8192
rect 15508 8132 15512 8188
rect 15512 8132 15568 8188
rect 15568 8132 15572 8188
rect 15508 8128 15572 8132
rect 15588 8188 15652 8192
rect 15588 8132 15592 8188
rect 15592 8132 15648 8188
rect 15648 8132 15652 8188
rect 15588 8128 15652 8132
rect 15668 8188 15732 8192
rect 15668 8132 15672 8188
rect 15672 8132 15728 8188
rect 15728 8132 15732 8188
rect 15668 8128 15732 8132
rect 15748 8188 15812 8192
rect 15748 8132 15752 8188
rect 15752 8132 15808 8188
rect 15808 8132 15812 8188
rect 15748 8128 15812 8132
rect 18608 8188 18672 8192
rect 18608 8132 18612 8188
rect 18612 8132 18668 8188
rect 18668 8132 18672 8188
rect 18608 8128 18672 8132
rect 18688 8188 18752 8192
rect 18688 8132 18692 8188
rect 18692 8132 18748 8188
rect 18748 8132 18752 8188
rect 18688 8128 18752 8132
rect 18768 8188 18832 8192
rect 18768 8132 18772 8188
rect 18772 8132 18828 8188
rect 18828 8132 18832 8188
rect 18768 8128 18832 8132
rect 18848 8188 18912 8192
rect 18848 8132 18852 8188
rect 18852 8132 18908 8188
rect 18908 8132 18912 8188
rect 18848 8128 18912 8132
rect 1558 7644 1622 7648
rect 1558 7588 1562 7644
rect 1562 7588 1618 7644
rect 1618 7588 1622 7644
rect 1558 7584 1622 7588
rect 1638 7644 1702 7648
rect 1638 7588 1642 7644
rect 1642 7588 1698 7644
rect 1698 7588 1702 7644
rect 1638 7584 1702 7588
rect 1718 7644 1782 7648
rect 1718 7588 1722 7644
rect 1722 7588 1778 7644
rect 1778 7588 1782 7644
rect 1718 7584 1782 7588
rect 1798 7644 1862 7648
rect 1798 7588 1802 7644
rect 1802 7588 1858 7644
rect 1858 7588 1862 7644
rect 1798 7584 1862 7588
rect 4658 7644 4722 7648
rect 4658 7588 4662 7644
rect 4662 7588 4718 7644
rect 4718 7588 4722 7644
rect 4658 7584 4722 7588
rect 4738 7644 4802 7648
rect 4738 7588 4742 7644
rect 4742 7588 4798 7644
rect 4798 7588 4802 7644
rect 4738 7584 4802 7588
rect 4818 7644 4882 7648
rect 4818 7588 4822 7644
rect 4822 7588 4878 7644
rect 4878 7588 4882 7644
rect 4818 7584 4882 7588
rect 4898 7644 4962 7648
rect 4898 7588 4902 7644
rect 4902 7588 4958 7644
rect 4958 7588 4962 7644
rect 4898 7584 4962 7588
rect 7758 7644 7822 7648
rect 7758 7588 7762 7644
rect 7762 7588 7818 7644
rect 7818 7588 7822 7644
rect 7758 7584 7822 7588
rect 7838 7644 7902 7648
rect 7838 7588 7842 7644
rect 7842 7588 7898 7644
rect 7898 7588 7902 7644
rect 7838 7584 7902 7588
rect 7918 7644 7982 7648
rect 7918 7588 7922 7644
rect 7922 7588 7978 7644
rect 7978 7588 7982 7644
rect 7918 7584 7982 7588
rect 7998 7644 8062 7648
rect 7998 7588 8002 7644
rect 8002 7588 8058 7644
rect 8058 7588 8062 7644
rect 7998 7584 8062 7588
rect 10858 7644 10922 7648
rect 10858 7588 10862 7644
rect 10862 7588 10918 7644
rect 10918 7588 10922 7644
rect 10858 7584 10922 7588
rect 10938 7644 11002 7648
rect 10938 7588 10942 7644
rect 10942 7588 10998 7644
rect 10998 7588 11002 7644
rect 10938 7584 11002 7588
rect 11018 7644 11082 7648
rect 11018 7588 11022 7644
rect 11022 7588 11078 7644
rect 11078 7588 11082 7644
rect 11018 7584 11082 7588
rect 11098 7644 11162 7648
rect 11098 7588 11102 7644
rect 11102 7588 11158 7644
rect 11158 7588 11162 7644
rect 11098 7584 11162 7588
rect 13958 7644 14022 7648
rect 13958 7588 13962 7644
rect 13962 7588 14018 7644
rect 14018 7588 14022 7644
rect 13958 7584 14022 7588
rect 14038 7644 14102 7648
rect 14038 7588 14042 7644
rect 14042 7588 14098 7644
rect 14098 7588 14102 7644
rect 14038 7584 14102 7588
rect 14118 7644 14182 7648
rect 14118 7588 14122 7644
rect 14122 7588 14178 7644
rect 14178 7588 14182 7644
rect 14118 7584 14182 7588
rect 14198 7644 14262 7648
rect 14198 7588 14202 7644
rect 14202 7588 14258 7644
rect 14258 7588 14262 7644
rect 14198 7584 14262 7588
rect 17058 7644 17122 7648
rect 17058 7588 17062 7644
rect 17062 7588 17118 7644
rect 17118 7588 17122 7644
rect 17058 7584 17122 7588
rect 17138 7644 17202 7648
rect 17138 7588 17142 7644
rect 17142 7588 17198 7644
rect 17198 7588 17202 7644
rect 17138 7584 17202 7588
rect 17218 7644 17282 7648
rect 17218 7588 17222 7644
rect 17222 7588 17278 7644
rect 17278 7588 17282 7644
rect 17218 7584 17282 7588
rect 17298 7644 17362 7648
rect 17298 7588 17302 7644
rect 17302 7588 17358 7644
rect 17358 7588 17362 7644
rect 17298 7584 17362 7588
rect 3108 7100 3172 7104
rect 3108 7044 3112 7100
rect 3112 7044 3168 7100
rect 3168 7044 3172 7100
rect 3108 7040 3172 7044
rect 3188 7100 3252 7104
rect 3188 7044 3192 7100
rect 3192 7044 3248 7100
rect 3248 7044 3252 7100
rect 3188 7040 3252 7044
rect 3268 7100 3332 7104
rect 3268 7044 3272 7100
rect 3272 7044 3328 7100
rect 3328 7044 3332 7100
rect 3268 7040 3332 7044
rect 3348 7100 3412 7104
rect 3348 7044 3352 7100
rect 3352 7044 3408 7100
rect 3408 7044 3412 7100
rect 3348 7040 3412 7044
rect 6208 7100 6272 7104
rect 6208 7044 6212 7100
rect 6212 7044 6268 7100
rect 6268 7044 6272 7100
rect 6208 7040 6272 7044
rect 6288 7100 6352 7104
rect 6288 7044 6292 7100
rect 6292 7044 6348 7100
rect 6348 7044 6352 7100
rect 6288 7040 6352 7044
rect 6368 7100 6432 7104
rect 6368 7044 6372 7100
rect 6372 7044 6428 7100
rect 6428 7044 6432 7100
rect 6368 7040 6432 7044
rect 6448 7100 6512 7104
rect 6448 7044 6452 7100
rect 6452 7044 6508 7100
rect 6508 7044 6512 7100
rect 6448 7040 6512 7044
rect 9308 7100 9372 7104
rect 9308 7044 9312 7100
rect 9312 7044 9368 7100
rect 9368 7044 9372 7100
rect 9308 7040 9372 7044
rect 9388 7100 9452 7104
rect 9388 7044 9392 7100
rect 9392 7044 9448 7100
rect 9448 7044 9452 7100
rect 9388 7040 9452 7044
rect 9468 7100 9532 7104
rect 9468 7044 9472 7100
rect 9472 7044 9528 7100
rect 9528 7044 9532 7100
rect 9468 7040 9532 7044
rect 9548 7100 9612 7104
rect 9548 7044 9552 7100
rect 9552 7044 9608 7100
rect 9608 7044 9612 7100
rect 9548 7040 9612 7044
rect 12408 7100 12472 7104
rect 12408 7044 12412 7100
rect 12412 7044 12468 7100
rect 12468 7044 12472 7100
rect 12408 7040 12472 7044
rect 12488 7100 12552 7104
rect 12488 7044 12492 7100
rect 12492 7044 12548 7100
rect 12548 7044 12552 7100
rect 12488 7040 12552 7044
rect 12568 7100 12632 7104
rect 12568 7044 12572 7100
rect 12572 7044 12628 7100
rect 12628 7044 12632 7100
rect 12568 7040 12632 7044
rect 12648 7100 12712 7104
rect 12648 7044 12652 7100
rect 12652 7044 12708 7100
rect 12708 7044 12712 7100
rect 12648 7040 12712 7044
rect 15508 7100 15572 7104
rect 15508 7044 15512 7100
rect 15512 7044 15568 7100
rect 15568 7044 15572 7100
rect 15508 7040 15572 7044
rect 15588 7100 15652 7104
rect 15588 7044 15592 7100
rect 15592 7044 15648 7100
rect 15648 7044 15652 7100
rect 15588 7040 15652 7044
rect 15668 7100 15732 7104
rect 15668 7044 15672 7100
rect 15672 7044 15728 7100
rect 15728 7044 15732 7100
rect 15668 7040 15732 7044
rect 15748 7100 15812 7104
rect 15748 7044 15752 7100
rect 15752 7044 15808 7100
rect 15808 7044 15812 7100
rect 15748 7040 15812 7044
rect 18608 7100 18672 7104
rect 18608 7044 18612 7100
rect 18612 7044 18668 7100
rect 18668 7044 18672 7100
rect 18608 7040 18672 7044
rect 18688 7100 18752 7104
rect 18688 7044 18692 7100
rect 18692 7044 18748 7100
rect 18748 7044 18752 7100
rect 18688 7040 18752 7044
rect 18768 7100 18832 7104
rect 18768 7044 18772 7100
rect 18772 7044 18828 7100
rect 18828 7044 18832 7100
rect 18768 7040 18832 7044
rect 18848 7100 18912 7104
rect 18848 7044 18852 7100
rect 18852 7044 18908 7100
rect 18908 7044 18912 7100
rect 18848 7040 18912 7044
rect 1558 6556 1622 6560
rect 1558 6500 1562 6556
rect 1562 6500 1618 6556
rect 1618 6500 1622 6556
rect 1558 6496 1622 6500
rect 1638 6556 1702 6560
rect 1638 6500 1642 6556
rect 1642 6500 1698 6556
rect 1698 6500 1702 6556
rect 1638 6496 1702 6500
rect 1718 6556 1782 6560
rect 1718 6500 1722 6556
rect 1722 6500 1778 6556
rect 1778 6500 1782 6556
rect 1718 6496 1782 6500
rect 1798 6556 1862 6560
rect 1798 6500 1802 6556
rect 1802 6500 1858 6556
rect 1858 6500 1862 6556
rect 1798 6496 1862 6500
rect 4658 6556 4722 6560
rect 4658 6500 4662 6556
rect 4662 6500 4718 6556
rect 4718 6500 4722 6556
rect 4658 6496 4722 6500
rect 4738 6556 4802 6560
rect 4738 6500 4742 6556
rect 4742 6500 4798 6556
rect 4798 6500 4802 6556
rect 4738 6496 4802 6500
rect 4818 6556 4882 6560
rect 4818 6500 4822 6556
rect 4822 6500 4878 6556
rect 4878 6500 4882 6556
rect 4818 6496 4882 6500
rect 4898 6556 4962 6560
rect 4898 6500 4902 6556
rect 4902 6500 4958 6556
rect 4958 6500 4962 6556
rect 4898 6496 4962 6500
rect 7758 6556 7822 6560
rect 7758 6500 7762 6556
rect 7762 6500 7818 6556
rect 7818 6500 7822 6556
rect 7758 6496 7822 6500
rect 7838 6556 7902 6560
rect 7838 6500 7842 6556
rect 7842 6500 7898 6556
rect 7898 6500 7902 6556
rect 7838 6496 7902 6500
rect 7918 6556 7982 6560
rect 7918 6500 7922 6556
rect 7922 6500 7978 6556
rect 7978 6500 7982 6556
rect 7918 6496 7982 6500
rect 7998 6556 8062 6560
rect 7998 6500 8002 6556
rect 8002 6500 8058 6556
rect 8058 6500 8062 6556
rect 7998 6496 8062 6500
rect 10858 6556 10922 6560
rect 10858 6500 10862 6556
rect 10862 6500 10918 6556
rect 10918 6500 10922 6556
rect 10858 6496 10922 6500
rect 10938 6556 11002 6560
rect 10938 6500 10942 6556
rect 10942 6500 10998 6556
rect 10998 6500 11002 6556
rect 10938 6496 11002 6500
rect 11018 6556 11082 6560
rect 11018 6500 11022 6556
rect 11022 6500 11078 6556
rect 11078 6500 11082 6556
rect 11018 6496 11082 6500
rect 11098 6556 11162 6560
rect 11098 6500 11102 6556
rect 11102 6500 11158 6556
rect 11158 6500 11162 6556
rect 11098 6496 11162 6500
rect 13958 6556 14022 6560
rect 13958 6500 13962 6556
rect 13962 6500 14018 6556
rect 14018 6500 14022 6556
rect 13958 6496 14022 6500
rect 14038 6556 14102 6560
rect 14038 6500 14042 6556
rect 14042 6500 14098 6556
rect 14098 6500 14102 6556
rect 14038 6496 14102 6500
rect 14118 6556 14182 6560
rect 14118 6500 14122 6556
rect 14122 6500 14178 6556
rect 14178 6500 14182 6556
rect 14118 6496 14182 6500
rect 14198 6556 14262 6560
rect 14198 6500 14202 6556
rect 14202 6500 14258 6556
rect 14258 6500 14262 6556
rect 14198 6496 14262 6500
rect 17058 6556 17122 6560
rect 17058 6500 17062 6556
rect 17062 6500 17118 6556
rect 17118 6500 17122 6556
rect 17058 6496 17122 6500
rect 17138 6556 17202 6560
rect 17138 6500 17142 6556
rect 17142 6500 17198 6556
rect 17198 6500 17202 6556
rect 17138 6496 17202 6500
rect 17218 6556 17282 6560
rect 17218 6500 17222 6556
rect 17222 6500 17278 6556
rect 17278 6500 17282 6556
rect 17218 6496 17282 6500
rect 17298 6556 17362 6560
rect 17298 6500 17302 6556
rect 17302 6500 17358 6556
rect 17358 6500 17362 6556
rect 17298 6496 17362 6500
rect 3108 6012 3172 6016
rect 3108 5956 3112 6012
rect 3112 5956 3168 6012
rect 3168 5956 3172 6012
rect 3108 5952 3172 5956
rect 3188 6012 3252 6016
rect 3188 5956 3192 6012
rect 3192 5956 3248 6012
rect 3248 5956 3252 6012
rect 3188 5952 3252 5956
rect 3268 6012 3332 6016
rect 3268 5956 3272 6012
rect 3272 5956 3328 6012
rect 3328 5956 3332 6012
rect 3268 5952 3332 5956
rect 3348 6012 3412 6016
rect 3348 5956 3352 6012
rect 3352 5956 3408 6012
rect 3408 5956 3412 6012
rect 3348 5952 3412 5956
rect 6208 6012 6272 6016
rect 6208 5956 6212 6012
rect 6212 5956 6268 6012
rect 6268 5956 6272 6012
rect 6208 5952 6272 5956
rect 6288 6012 6352 6016
rect 6288 5956 6292 6012
rect 6292 5956 6348 6012
rect 6348 5956 6352 6012
rect 6288 5952 6352 5956
rect 6368 6012 6432 6016
rect 6368 5956 6372 6012
rect 6372 5956 6428 6012
rect 6428 5956 6432 6012
rect 6368 5952 6432 5956
rect 6448 6012 6512 6016
rect 6448 5956 6452 6012
rect 6452 5956 6508 6012
rect 6508 5956 6512 6012
rect 6448 5952 6512 5956
rect 9308 6012 9372 6016
rect 9308 5956 9312 6012
rect 9312 5956 9368 6012
rect 9368 5956 9372 6012
rect 9308 5952 9372 5956
rect 9388 6012 9452 6016
rect 9388 5956 9392 6012
rect 9392 5956 9448 6012
rect 9448 5956 9452 6012
rect 9388 5952 9452 5956
rect 9468 6012 9532 6016
rect 9468 5956 9472 6012
rect 9472 5956 9528 6012
rect 9528 5956 9532 6012
rect 9468 5952 9532 5956
rect 9548 6012 9612 6016
rect 9548 5956 9552 6012
rect 9552 5956 9608 6012
rect 9608 5956 9612 6012
rect 9548 5952 9612 5956
rect 12408 6012 12472 6016
rect 12408 5956 12412 6012
rect 12412 5956 12468 6012
rect 12468 5956 12472 6012
rect 12408 5952 12472 5956
rect 12488 6012 12552 6016
rect 12488 5956 12492 6012
rect 12492 5956 12548 6012
rect 12548 5956 12552 6012
rect 12488 5952 12552 5956
rect 12568 6012 12632 6016
rect 12568 5956 12572 6012
rect 12572 5956 12628 6012
rect 12628 5956 12632 6012
rect 12568 5952 12632 5956
rect 12648 6012 12712 6016
rect 12648 5956 12652 6012
rect 12652 5956 12708 6012
rect 12708 5956 12712 6012
rect 12648 5952 12712 5956
rect 15508 6012 15572 6016
rect 15508 5956 15512 6012
rect 15512 5956 15568 6012
rect 15568 5956 15572 6012
rect 15508 5952 15572 5956
rect 15588 6012 15652 6016
rect 15588 5956 15592 6012
rect 15592 5956 15648 6012
rect 15648 5956 15652 6012
rect 15588 5952 15652 5956
rect 15668 6012 15732 6016
rect 15668 5956 15672 6012
rect 15672 5956 15728 6012
rect 15728 5956 15732 6012
rect 15668 5952 15732 5956
rect 15748 6012 15812 6016
rect 15748 5956 15752 6012
rect 15752 5956 15808 6012
rect 15808 5956 15812 6012
rect 15748 5952 15812 5956
rect 18608 6012 18672 6016
rect 18608 5956 18612 6012
rect 18612 5956 18668 6012
rect 18668 5956 18672 6012
rect 18608 5952 18672 5956
rect 18688 6012 18752 6016
rect 18688 5956 18692 6012
rect 18692 5956 18748 6012
rect 18748 5956 18752 6012
rect 18688 5952 18752 5956
rect 18768 6012 18832 6016
rect 18768 5956 18772 6012
rect 18772 5956 18828 6012
rect 18828 5956 18832 6012
rect 18768 5952 18832 5956
rect 18848 6012 18912 6016
rect 18848 5956 18852 6012
rect 18852 5956 18908 6012
rect 18908 5956 18912 6012
rect 18848 5952 18912 5956
rect 1558 5468 1622 5472
rect 1558 5412 1562 5468
rect 1562 5412 1618 5468
rect 1618 5412 1622 5468
rect 1558 5408 1622 5412
rect 1638 5468 1702 5472
rect 1638 5412 1642 5468
rect 1642 5412 1698 5468
rect 1698 5412 1702 5468
rect 1638 5408 1702 5412
rect 1718 5468 1782 5472
rect 1718 5412 1722 5468
rect 1722 5412 1778 5468
rect 1778 5412 1782 5468
rect 1718 5408 1782 5412
rect 1798 5468 1862 5472
rect 1798 5412 1802 5468
rect 1802 5412 1858 5468
rect 1858 5412 1862 5468
rect 1798 5408 1862 5412
rect 4658 5468 4722 5472
rect 4658 5412 4662 5468
rect 4662 5412 4718 5468
rect 4718 5412 4722 5468
rect 4658 5408 4722 5412
rect 4738 5468 4802 5472
rect 4738 5412 4742 5468
rect 4742 5412 4798 5468
rect 4798 5412 4802 5468
rect 4738 5408 4802 5412
rect 4818 5468 4882 5472
rect 4818 5412 4822 5468
rect 4822 5412 4878 5468
rect 4878 5412 4882 5468
rect 4818 5408 4882 5412
rect 4898 5468 4962 5472
rect 4898 5412 4902 5468
rect 4902 5412 4958 5468
rect 4958 5412 4962 5468
rect 4898 5408 4962 5412
rect 7758 5468 7822 5472
rect 7758 5412 7762 5468
rect 7762 5412 7818 5468
rect 7818 5412 7822 5468
rect 7758 5408 7822 5412
rect 7838 5468 7902 5472
rect 7838 5412 7842 5468
rect 7842 5412 7898 5468
rect 7898 5412 7902 5468
rect 7838 5408 7902 5412
rect 7918 5468 7982 5472
rect 7918 5412 7922 5468
rect 7922 5412 7978 5468
rect 7978 5412 7982 5468
rect 7918 5408 7982 5412
rect 7998 5468 8062 5472
rect 7998 5412 8002 5468
rect 8002 5412 8058 5468
rect 8058 5412 8062 5468
rect 7998 5408 8062 5412
rect 10858 5468 10922 5472
rect 10858 5412 10862 5468
rect 10862 5412 10918 5468
rect 10918 5412 10922 5468
rect 10858 5408 10922 5412
rect 10938 5468 11002 5472
rect 10938 5412 10942 5468
rect 10942 5412 10998 5468
rect 10998 5412 11002 5468
rect 10938 5408 11002 5412
rect 11018 5468 11082 5472
rect 11018 5412 11022 5468
rect 11022 5412 11078 5468
rect 11078 5412 11082 5468
rect 11018 5408 11082 5412
rect 11098 5468 11162 5472
rect 11098 5412 11102 5468
rect 11102 5412 11158 5468
rect 11158 5412 11162 5468
rect 11098 5408 11162 5412
rect 13958 5468 14022 5472
rect 13958 5412 13962 5468
rect 13962 5412 14018 5468
rect 14018 5412 14022 5468
rect 13958 5408 14022 5412
rect 14038 5468 14102 5472
rect 14038 5412 14042 5468
rect 14042 5412 14098 5468
rect 14098 5412 14102 5468
rect 14038 5408 14102 5412
rect 14118 5468 14182 5472
rect 14118 5412 14122 5468
rect 14122 5412 14178 5468
rect 14178 5412 14182 5468
rect 14118 5408 14182 5412
rect 14198 5468 14262 5472
rect 14198 5412 14202 5468
rect 14202 5412 14258 5468
rect 14258 5412 14262 5468
rect 14198 5408 14262 5412
rect 17058 5468 17122 5472
rect 17058 5412 17062 5468
rect 17062 5412 17118 5468
rect 17118 5412 17122 5468
rect 17058 5408 17122 5412
rect 17138 5468 17202 5472
rect 17138 5412 17142 5468
rect 17142 5412 17198 5468
rect 17198 5412 17202 5468
rect 17138 5408 17202 5412
rect 17218 5468 17282 5472
rect 17218 5412 17222 5468
rect 17222 5412 17278 5468
rect 17278 5412 17282 5468
rect 17218 5408 17282 5412
rect 17298 5468 17362 5472
rect 17298 5412 17302 5468
rect 17302 5412 17358 5468
rect 17358 5412 17362 5468
rect 17298 5408 17362 5412
rect 3108 4924 3172 4928
rect 3108 4868 3112 4924
rect 3112 4868 3168 4924
rect 3168 4868 3172 4924
rect 3108 4864 3172 4868
rect 3188 4924 3252 4928
rect 3188 4868 3192 4924
rect 3192 4868 3248 4924
rect 3248 4868 3252 4924
rect 3188 4864 3252 4868
rect 3268 4924 3332 4928
rect 3268 4868 3272 4924
rect 3272 4868 3328 4924
rect 3328 4868 3332 4924
rect 3268 4864 3332 4868
rect 3348 4924 3412 4928
rect 3348 4868 3352 4924
rect 3352 4868 3408 4924
rect 3408 4868 3412 4924
rect 3348 4864 3412 4868
rect 6208 4924 6272 4928
rect 6208 4868 6212 4924
rect 6212 4868 6268 4924
rect 6268 4868 6272 4924
rect 6208 4864 6272 4868
rect 6288 4924 6352 4928
rect 6288 4868 6292 4924
rect 6292 4868 6348 4924
rect 6348 4868 6352 4924
rect 6288 4864 6352 4868
rect 6368 4924 6432 4928
rect 6368 4868 6372 4924
rect 6372 4868 6428 4924
rect 6428 4868 6432 4924
rect 6368 4864 6432 4868
rect 6448 4924 6512 4928
rect 6448 4868 6452 4924
rect 6452 4868 6508 4924
rect 6508 4868 6512 4924
rect 6448 4864 6512 4868
rect 9308 4924 9372 4928
rect 9308 4868 9312 4924
rect 9312 4868 9368 4924
rect 9368 4868 9372 4924
rect 9308 4864 9372 4868
rect 9388 4924 9452 4928
rect 9388 4868 9392 4924
rect 9392 4868 9448 4924
rect 9448 4868 9452 4924
rect 9388 4864 9452 4868
rect 9468 4924 9532 4928
rect 9468 4868 9472 4924
rect 9472 4868 9528 4924
rect 9528 4868 9532 4924
rect 9468 4864 9532 4868
rect 9548 4924 9612 4928
rect 9548 4868 9552 4924
rect 9552 4868 9608 4924
rect 9608 4868 9612 4924
rect 9548 4864 9612 4868
rect 12408 4924 12472 4928
rect 12408 4868 12412 4924
rect 12412 4868 12468 4924
rect 12468 4868 12472 4924
rect 12408 4864 12472 4868
rect 12488 4924 12552 4928
rect 12488 4868 12492 4924
rect 12492 4868 12548 4924
rect 12548 4868 12552 4924
rect 12488 4864 12552 4868
rect 12568 4924 12632 4928
rect 12568 4868 12572 4924
rect 12572 4868 12628 4924
rect 12628 4868 12632 4924
rect 12568 4864 12632 4868
rect 12648 4924 12712 4928
rect 12648 4868 12652 4924
rect 12652 4868 12708 4924
rect 12708 4868 12712 4924
rect 12648 4864 12712 4868
rect 15508 4924 15572 4928
rect 15508 4868 15512 4924
rect 15512 4868 15568 4924
rect 15568 4868 15572 4924
rect 15508 4864 15572 4868
rect 15588 4924 15652 4928
rect 15588 4868 15592 4924
rect 15592 4868 15648 4924
rect 15648 4868 15652 4924
rect 15588 4864 15652 4868
rect 15668 4924 15732 4928
rect 15668 4868 15672 4924
rect 15672 4868 15728 4924
rect 15728 4868 15732 4924
rect 15668 4864 15732 4868
rect 15748 4924 15812 4928
rect 15748 4868 15752 4924
rect 15752 4868 15808 4924
rect 15808 4868 15812 4924
rect 15748 4864 15812 4868
rect 18608 4924 18672 4928
rect 18608 4868 18612 4924
rect 18612 4868 18668 4924
rect 18668 4868 18672 4924
rect 18608 4864 18672 4868
rect 18688 4924 18752 4928
rect 18688 4868 18692 4924
rect 18692 4868 18748 4924
rect 18748 4868 18752 4924
rect 18688 4864 18752 4868
rect 18768 4924 18832 4928
rect 18768 4868 18772 4924
rect 18772 4868 18828 4924
rect 18828 4868 18832 4924
rect 18768 4864 18832 4868
rect 18848 4924 18912 4928
rect 18848 4868 18852 4924
rect 18852 4868 18908 4924
rect 18908 4868 18912 4924
rect 18848 4864 18912 4868
rect 1558 4380 1622 4384
rect 1558 4324 1562 4380
rect 1562 4324 1618 4380
rect 1618 4324 1622 4380
rect 1558 4320 1622 4324
rect 1638 4380 1702 4384
rect 1638 4324 1642 4380
rect 1642 4324 1698 4380
rect 1698 4324 1702 4380
rect 1638 4320 1702 4324
rect 1718 4380 1782 4384
rect 1718 4324 1722 4380
rect 1722 4324 1778 4380
rect 1778 4324 1782 4380
rect 1718 4320 1782 4324
rect 1798 4380 1862 4384
rect 1798 4324 1802 4380
rect 1802 4324 1858 4380
rect 1858 4324 1862 4380
rect 1798 4320 1862 4324
rect 4658 4380 4722 4384
rect 4658 4324 4662 4380
rect 4662 4324 4718 4380
rect 4718 4324 4722 4380
rect 4658 4320 4722 4324
rect 4738 4380 4802 4384
rect 4738 4324 4742 4380
rect 4742 4324 4798 4380
rect 4798 4324 4802 4380
rect 4738 4320 4802 4324
rect 4818 4380 4882 4384
rect 4818 4324 4822 4380
rect 4822 4324 4878 4380
rect 4878 4324 4882 4380
rect 4818 4320 4882 4324
rect 4898 4380 4962 4384
rect 4898 4324 4902 4380
rect 4902 4324 4958 4380
rect 4958 4324 4962 4380
rect 4898 4320 4962 4324
rect 7758 4380 7822 4384
rect 7758 4324 7762 4380
rect 7762 4324 7818 4380
rect 7818 4324 7822 4380
rect 7758 4320 7822 4324
rect 7838 4380 7902 4384
rect 7838 4324 7842 4380
rect 7842 4324 7898 4380
rect 7898 4324 7902 4380
rect 7838 4320 7902 4324
rect 7918 4380 7982 4384
rect 7918 4324 7922 4380
rect 7922 4324 7978 4380
rect 7978 4324 7982 4380
rect 7918 4320 7982 4324
rect 7998 4380 8062 4384
rect 7998 4324 8002 4380
rect 8002 4324 8058 4380
rect 8058 4324 8062 4380
rect 7998 4320 8062 4324
rect 10858 4380 10922 4384
rect 10858 4324 10862 4380
rect 10862 4324 10918 4380
rect 10918 4324 10922 4380
rect 10858 4320 10922 4324
rect 10938 4380 11002 4384
rect 10938 4324 10942 4380
rect 10942 4324 10998 4380
rect 10998 4324 11002 4380
rect 10938 4320 11002 4324
rect 11018 4380 11082 4384
rect 11018 4324 11022 4380
rect 11022 4324 11078 4380
rect 11078 4324 11082 4380
rect 11018 4320 11082 4324
rect 11098 4380 11162 4384
rect 11098 4324 11102 4380
rect 11102 4324 11158 4380
rect 11158 4324 11162 4380
rect 11098 4320 11162 4324
rect 13958 4380 14022 4384
rect 13958 4324 13962 4380
rect 13962 4324 14018 4380
rect 14018 4324 14022 4380
rect 13958 4320 14022 4324
rect 14038 4380 14102 4384
rect 14038 4324 14042 4380
rect 14042 4324 14098 4380
rect 14098 4324 14102 4380
rect 14038 4320 14102 4324
rect 14118 4380 14182 4384
rect 14118 4324 14122 4380
rect 14122 4324 14178 4380
rect 14178 4324 14182 4380
rect 14118 4320 14182 4324
rect 14198 4380 14262 4384
rect 14198 4324 14202 4380
rect 14202 4324 14258 4380
rect 14258 4324 14262 4380
rect 14198 4320 14262 4324
rect 17058 4380 17122 4384
rect 17058 4324 17062 4380
rect 17062 4324 17118 4380
rect 17118 4324 17122 4380
rect 17058 4320 17122 4324
rect 17138 4380 17202 4384
rect 17138 4324 17142 4380
rect 17142 4324 17198 4380
rect 17198 4324 17202 4380
rect 17138 4320 17202 4324
rect 17218 4380 17282 4384
rect 17218 4324 17222 4380
rect 17222 4324 17278 4380
rect 17278 4324 17282 4380
rect 17218 4320 17282 4324
rect 17298 4380 17362 4384
rect 17298 4324 17302 4380
rect 17302 4324 17358 4380
rect 17358 4324 17362 4380
rect 17298 4320 17362 4324
rect 3108 3836 3172 3840
rect 3108 3780 3112 3836
rect 3112 3780 3168 3836
rect 3168 3780 3172 3836
rect 3108 3776 3172 3780
rect 3188 3836 3252 3840
rect 3188 3780 3192 3836
rect 3192 3780 3248 3836
rect 3248 3780 3252 3836
rect 3188 3776 3252 3780
rect 3268 3836 3332 3840
rect 3268 3780 3272 3836
rect 3272 3780 3328 3836
rect 3328 3780 3332 3836
rect 3268 3776 3332 3780
rect 3348 3836 3412 3840
rect 3348 3780 3352 3836
rect 3352 3780 3408 3836
rect 3408 3780 3412 3836
rect 3348 3776 3412 3780
rect 6208 3836 6272 3840
rect 6208 3780 6212 3836
rect 6212 3780 6268 3836
rect 6268 3780 6272 3836
rect 6208 3776 6272 3780
rect 6288 3836 6352 3840
rect 6288 3780 6292 3836
rect 6292 3780 6348 3836
rect 6348 3780 6352 3836
rect 6288 3776 6352 3780
rect 6368 3836 6432 3840
rect 6368 3780 6372 3836
rect 6372 3780 6428 3836
rect 6428 3780 6432 3836
rect 6368 3776 6432 3780
rect 6448 3836 6512 3840
rect 6448 3780 6452 3836
rect 6452 3780 6508 3836
rect 6508 3780 6512 3836
rect 6448 3776 6512 3780
rect 9308 3836 9372 3840
rect 9308 3780 9312 3836
rect 9312 3780 9368 3836
rect 9368 3780 9372 3836
rect 9308 3776 9372 3780
rect 9388 3836 9452 3840
rect 9388 3780 9392 3836
rect 9392 3780 9448 3836
rect 9448 3780 9452 3836
rect 9388 3776 9452 3780
rect 9468 3836 9532 3840
rect 9468 3780 9472 3836
rect 9472 3780 9528 3836
rect 9528 3780 9532 3836
rect 9468 3776 9532 3780
rect 9548 3836 9612 3840
rect 9548 3780 9552 3836
rect 9552 3780 9608 3836
rect 9608 3780 9612 3836
rect 9548 3776 9612 3780
rect 12408 3836 12472 3840
rect 12408 3780 12412 3836
rect 12412 3780 12468 3836
rect 12468 3780 12472 3836
rect 12408 3776 12472 3780
rect 12488 3836 12552 3840
rect 12488 3780 12492 3836
rect 12492 3780 12548 3836
rect 12548 3780 12552 3836
rect 12488 3776 12552 3780
rect 12568 3836 12632 3840
rect 12568 3780 12572 3836
rect 12572 3780 12628 3836
rect 12628 3780 12632 3836
rect 12568 3776 12632 3780
rect 12648 3836 12712 3840
rect 12648 3780 12652 3836
rect 12652 3780 12708 3836
rect 12708 3780 12712 3836
rect 12648 3776 12712 3780
rect 15508 3836 15572 3840
rect 15508 3780 15512 3836
rect 15512 3780 15568 3836
rect 15568 3780 15572 3836
rect 15508 3776 15572 3780
rect 15588 3836 15652 3840
rect 15588 3780 15592 3836
rect 15592 3780 15648 3836
rect 15648 3780 15652 3836
rect 15588 3776 15652 3780
rect 15668 3836 15732 3840
rect 15668 3780 15672 3836
rect 15672 3780 15728 3836
rect 15728 3780 15732 3836
rect 15668 3776 15732 3780
rect 15748 3836 15812 3840
rect 15748 3780 15752 3836
rect 15752 3780 15808 3836
rect 15808 3780 15812 3836
rect 15748 3776 15812 3780
rect 18608 3836 18672 3840
rect 18608 3780 18612 3836
rect 18612 3780 18668 3836
rect 18668 3780 18672 3836
rect 18608 3776 18672 3780
rect 18688 3836 18752 3840
rect 18688 3780 18692 3836
rect 18692 3780 18748 3836
rect 18748 3780 18752 3836
rect 18688 3776 18752 3780
rect 18768 3836 18832 3840
rect 18768 3780 18772 3836
rect 18772 3780 18828 3836
rect 18828 3780 18832 3836
rect 18768 3776 18832 3780
rect 18848 3836 18912 3840
rect 18848 3780 18852 3836
rect 18852 3780 18908 3836
rect 18908 3780 18912 3836
rect 18848 3776 18912 3780
rect 1558 3292 1622 3296
rect 1558 3236 1562 3292
rect 1562 3236 1618 3292
rect 1618 3236 1622 3292
rect 1558 3232 1622 3236
rect 1638 3292 1702 3296
rect 1638 3236 1642 3292
rect 1642 3236 1698 3292
rect 1698 3236 1702 3292
rect 1638 3232 1702 3236
rect 1718 3292 1782 3296
rect 1718 3236 1722 3292
rect 1722 3236 1778 3292
rect 1778 3236 1782 3292
rect 1718 3232 1782 3236
rect 1798 3292 1862 3296
rect 1798 3236 1802 3292
rect 1802 3236 1858 3292
rect 1858 3236 1862 3292
rect 1798 3232 1862 3236
rect 4658 3292 4722 3296
rect 4658 3236 4662 3292
rect 4662 3236 4718 3292
rect 4718 3236 4722 3292
rect 4658 3232 4722 3236
rect 4738 3292 4802 3296
rect 4738 3236 4742 3292
rect 4742 3236 4798 3292
rect 4798 3236 4802 3292
rect 4738 3232 4802 3236
rect 4818 3292 4882 3296
rect 4818 3236 4822 3292
rect 4822 3236 4878 3292
rect 4878 3236 4882 3292
rect 4818 3232 4882 3236
rect 4898 3292 4962 3296
rect 4898 3236 4902 3292
rect 4902 3236 4958 3292
rect 4958 3236 4962 3292
rect 4898 3232 4962 3236
rect 7758 3292 7822 3296
rect 7758 3236 7762 3292
rect 7762 3236 7818 3292
rect 7818 3236 7822 3292
rect 7758 3232 7822 3236
rect 7838 3292 7902 3296
rect 7838 3236 7842 3292
rect 7842 3236 7898 3292
rect 7898 3236 7902 3292
rect 7838 3232 7902 3236
rect 7918 3292 7982 3296
rect 7918 3236 7922 3292
rect 7922 3236 7978 3292
rect 7978 3236 7982 3292
rect 7918 3232 7982 3236
rect 7998 3292 8062 3296
rect 7998 3236 8002 3292
rect 8002 3236 8058 3292
rect 8058 3236 8062 3292
rect 7998 3232 8062 3236
rect 10858 3292 10922 3296
rect 10858 3236 10862 3292
rect 10862 3236 10918 3292
rect 10918 3236 10922 3292
rect 10858 3232 10922 3236
rect 10938 3292 11002 3296
rect 10938 3236 10942 3292
rect 10942 3236 10998 3292
rect 10998 3236 11002 3292
rect 10938 3232 11002 3236
rect 11018 3292 11082 3296
rect 11018 3236 11022 3292
rect 11022 3236 11078 3292
rect 11078 3236 11082 3292
rect 11018 3232 11082 3236
rect 11098 3292 11162 3296
rect 11098 3236 11102 3292
rect 11102 3236 11158 3292
rect 11158 3236 11162 3292
rect 11098 3232 11162 3236
rect 13958 3292 14022 3296
rect 13958 3236 13962 3292
rect 13962 3236 14018 3292
rect 14018 3236 14022 3292
rect 13958 3232 14022 3236
rect 14038 3292 14102 3296
rect 14038 3236 14042 3292
rect 14042 3236 14098 3292
rect 14098 3236 14102 3292
rect 14038 3232 14102 3236
rect 14118 3292 14182 3296
rect 14118 3236 14122 3292
rect 14122 3236 14178 3292
rect 14178 3236 14182 3292
rect 14118 3232 14182 3236
rect 14198 3292 14262 3296
rect 14198 3236 14202 3292
rect 14202 3236 14258 3292
rect 14258 3236 14262 3292
rect 14198 3232 14262 3236
rect 17058 3292 17122 3296
rect 17058 3236 17062 3292
rect 17062 3236 17118 3292
rect 17118 3236 17122 3292
rect 17058 3232 17122 3236
rect 17138 3292 17202 3296
rect 17138 3236 17142 3292
rect 17142 3236 17198 3292
rect 17198 3236 17202 3292
rect 17138 3232 17202 3236
rect 17218 3292 17282 3296
rect 17218 3236 17222 3292
rect 17222 3236 17278 3292
rect 17278 3236 17282 3292
rect 17218 3232 17282 3236
rect 17298 3292 17362 3296
rect 17298 3236 17302 3292
rect 17302 3236 17358 3292
rect 17358 3236 17362 3292
rect 17298 3232 17362 3236
rect 3108 2748 3172 2752
rect 3108 2692 3112 2748
rect 3112 2692 3168 2748
rect 3168 2692 3172 2748
rect 3108 2688 3172 2692
rect 3188 2748 3252 2752
rect 3188 2692 3192 2748
rect 3192 2692 3248 2748
rect 3248 2692 3252 2748
rect 3188 2688 3252 2692
rect 3268 2748 3332 2752
rect 3268 2692 3272 2748
rect 3272 2692 3328 2748
rect 3328 2692 3332 2748
rect 3268 2688 3332 2692
rect 3348 2748 3412 2752
rect 3348 2692 3352 2748
rect 3352 2692 3408 2748
rect 3408 2692 3412 2748
rect 3348 2688 3412 2692
rect 6208 2748 6272 2752
rect 6208 2692 6212 2748
rect 6212 2692 6268 2748
rect 6268 2692 6272 2748
rect 6208 2688 6272 2692
rect 6288 2748 6352 2752
rect 6288 2692 6292 2748
rect 6292 2692 6348 2748
rect 6348 2692 6352 2748
rect 6288 2688 6352 2692
rect 6368 2748 6432 2752
rect 6368 2692 6372 2748
rect 6372 2692 6428 2748
rect 6428 2692 6432 2748
rect 6368 2688 6432 2692
rect 6448 2748 6512 2752
rect 6448 2692 6452 2748
rect 6452 2692 6508 2748
rect 6508 2692 6512 2748
rect 6448 2688 6512 2692
rect 9308 2748 9372 2752
rect 9308 2692 9312 2748
rect 9312 2692 9368 2748
rect 9368 2692 9372 2748
rect 9308 2688 9372 2692
rect 9388 2748 9452 2752
rect 9388 2692 9392 2748
rect 9392 2692 9448 2748
rect 9448 2692 9452 2748
rect 9388 2688 9452 2692
rect 9468 2748 9532 2752
rect 9468 2692 9472 2748
rect 9472 2692 9528 2748
rect 9528 2692 9532 2748
rect 9468 2688 9532 2692
rect 9548 2748 9612 2752
rect 9548 2692 9552 2748
rect 9552 2692 9608 2748
rect 9608 2692 9612 2748
rect 9548 2688 9612 2692
rect 12408 2748 12472 2752
rect 12408 2692 12412 2748
rect 12412 2692 12468 2748
rect 12468 2692 12472 2748
rect 12408 2688 12472 2692
rect 12488 2748 12552 2752
rect 12488 2692 12492 2748
rect 12492 2692 12548 2748
rect 12548 2692 12552 2748
rect 12488 2688 12552 2692
rect 12568 2748 12632 2752
rect 12568 2692 12572 2748
rect 12572 2692 12628 2748
rect 12628 2692 12632 2748
rect 12568 2688 12632 2692
rect 12648 2748 12712 2752
rect 12648 2692 12652 2748
rect 12652 2692 12708 2748
rect 12708 2692 12712 2748
rect 12648 2688 12712 2692
rect 15508 2748 15572 2752
rect 15508 2692 15512 2748
rect 15512 2692 15568 2748
rect 15568 2692 15572 2748
rect 15508 2688 15572 2692
rect 15588 2748 15652 2752
rect 15588 2692 15592 2748
rect 15592 2692 15648 2748
rect 15648 2692 15652 2748
rect 15588 2688 15652 2692
rect 15668 2748 15732 2752
rect 15668 2692 15672 2748
rect 15672 2692 15728 2748
rect 15728 2692 15732 2748
rect 15668 2688 15732 2692
rect 15748 2748 15812 2752
rect 15748 2692 15752 2748
rect 15752 2692 15808 2748
rect 15808 2692 15812 2748
rect 15748 2688 15812 2692
rect 18608 2748 18672 2752
rect 18608 2692 18612 2748
rect 18612 2692 18668 2748
rect 18668 2692 18672 2748
rect 18608 2688 18672 2692
rect 18688 2748 18752 2752
rect 18688 2692 18692 2748
rect 18692 2692 18748 2748
rect 18748 2692 18752 2748
rect 18688 2688 18752 2692
rect 18768 2748 18832 2752
rect 18768 2692 18772 2748
rect 18772 2692 18828 2748
rect 18828 2692 18832 2748
rect 18768 2688 18832 2692
rect 18848 2748 18912 2752
rect 18848 2692 18852 2748
rect 18852 2692 18908 2748
rect 18908 2692 18912 2748
rect 18848 2688 18912 2692
rect 1558 2204 1622 2208
rect 1558 2148 1562 2204
rect 1562 2148 1618 2204
rect 1618 2148 1622 2204
rect 1558 2144 1622 2148
rect 1638 2204 1702 2208
rect 1638 2148 1642 2204
rect 1642 2148 1698 2204
rect 1698 2148 1702 2204
rect 1638 2144 1702 2148
rect 1718 2204 1782 2208
rect 1718 2148 1722 2204
rect 1722 2148 1778 2204
rect 1778 2148 1782 2204
rect 1718 2144 1782 2148
rect 1798 2204 1862 2208
rect 1798 2148 1802 2204
rect 1802 2148 1858 2204
rect 1858 2148 1862 2204
rect 1798 2144 1862 2148
rect 4658 2204 4722 2208
rect 4658 2148 4662 2204
rect 4662 2148 4718 2204
rect 4718 2148 4722 2204
rect 4658 2144 4722 2148
rect 4738 2204 4802 2208
rect 4738 2148 4742 2204
rect 4742 2148 4798 2204
rect 4798 2148 4802 2204
rect 4738 2144 4802 2148
rect 4818 2204 4882 2208
rect 4818 2148 4822 2204
rect 4822 2148 4878 2204
rect 4878 2148 4882 2204
rect 4818 2144 4882 2148
rect 4898 2204 4962 2208
rect 4898 2148 4902 2204
rect 4902 2148 4958 2204
rect 4958 2148 4962 2204
rect 4898 2144 4962 2148
rect 7758 2204 7822 2208
rect 7758 2148 7762 2204
rect 7762 2148 7818 2204
rect 7818 2148 7822 2204
rect 7758 2144 7822 2148
rect 7838 2204 7902 2208
rect 7838 2148 7842 2204
rect 7842 2148 7898 2204
rect 7898 2148 7902 2204
rect 7838 2144 7902 2148
rect 7918 2204 7982 2208
rect 7918 2148 7922 2204
rect 7922 2148 7978 2204
rect 7978 2148 7982 2204
rect 7918 2144 7982 2148
rect 7998 2204 8062 2208
rect 7998 2148 8002 2204
rect 8002 2148 8058 2204
rect 8058 2148 8062 2204
rect 7998 2144 8062 2148
rect 10858 2204 10922 2208
rect 10858 2148 10862 2204
rect 10862 2148 10918 2204
rect 10918 2148 10922 2204
rect 10858 2144 10922 2148
rect 10938 2204 11002 2208
rect 10938 2148 10942 2204
rect 10942 2148 10998 2204
rect 10998 2148 11002 2204
rect 10938 2144 11002 2148
rect 11018 2204 11082 2208
rect 11018 2148 11022 2204
rect 11022 2148 11078 2204
rect 11078 2148 11082 2204
rect 11018 2144 11082 2148
rect 11098 2204 11162 2208
rect 11098 2148 11102 2204
rect 11102 2148 11158 2204
rect 11158 2148 11162 2204
rect 11098 2144 11162 2148
rect 13958 2204 14022 2208
rect 13958 2148 13962 2204
rect 13962 2148 14018 2204
rect 14018 2148 14022 2204
rect 13958 2144 14022 2148
rect 14038 2204 14102 2208
rect 14038 2148 14042 2204
rect 14042 2148 14098 2204
rect 14098 2148 14102 2204
rect 14038 2144 14102 2148
rect 14118 2204 14182 2208
rect 14118 2148 14122 2204
rect 14122 2148 14178 2204
rect 14178 2148 14182 2204
rect 14118 2144 14182 2148
rect 14198 2204 14262 2208
rect 14198 2148 14202 2204
rect 14202 2148 14258 2204
rect 14258 2148 14262 2204
rect 14198 2144 14262 2148
rect 17058 2204 17122 2208
rect 17058 2148 17062 2204
rect 17062 2148 17118 2204
rect 17118 2148 17122 2204
rect 17058 2144 17122 2148
rect 17138 2204 17202 2208
rect 17138 2148 17142 2204
rect 17142 2148 17198 2204
rect 17198 2148 17202 2204
rect 17138 2144 17202 2148
rect 17218 2204 17282 2208
rect 17218 2148 17222 2204
rect 17222 2148 17278 2204
rect 17278 2148 17282 2204
rect 17218 2144 17282 2148
rect 17298 2204 17362 2208
rect 17298 2148 17302 2204
rect 17302 2148 17358 2204
rect 17358 2148 17362 2204
rect 17298 2144 17362 2148
rect 3108 1660 3172 1664
rect 3108 1604 3112 1660
rect 3112 1604 3168 1660
rect 3168 1604 3172 1660
rect 3108 1600 3172 1604
rect 3188 1660 3252 1664
rect 3188 1604 3192 1660
rect 3192 1604 3248 1660
rect 3248 1604 3252 1660
rect 3188 1600 3252 1604
rect 3268 1660 3332 1664
rect 3268 1604 3272 1660
rect 3272 1604 3328 1660
rect 3328 1604 3332 1660
rect 3268 1600 3332 1604
rect 3348 1660 3412 1664
rect 3348 1604 3352 1660
rect 3352 1604 3408 1660
rect 3408 1604 3412 1660
rect 3348 1600 3412 1604
rect 6208 1660 6272 1664
rect 6208 1604 6212 1660
rect 6212 1604 6268 1660
rect 6268 1604 6272 1660
rect 6208 1600 6272 1604
rect 6288 1660 6352 1664
rect 6288 1604 6292 1660
rect 6292 1604 6348 1660
rect 6348 1604 6352 1660
rect 6288 1600 6352 1604
rect 6368 1660 6432 1664
rect 6368 1604 6372 1660
rect 6372 1604 6428 1660
rect 6428 1604 6432 1660
rect 6368 1600 6432 1604
rect 6448 1660 6512 1664
rect 6448 1604 6452 1660
rect 6452 1604 6508 1660
rect 6508 1604 6512 1660
rect 6448 1600 6512 1604
rect 9308 1660 9372 1664
rect 9308 1604 9312 1660
rect 9312 1604 9368 1660
rect 9368 1604 9372 1660
rect 9308 1600 9372 1604
rect 9388 1660 9452 1664
rect 9388 1604 9392 1660
rect 9392 1604 9448 1660
rect 9448 1604 9452 1660
rect 9388 1600 9452 1604
rect 9468 1660 9532 1664
rect 9468 1604 9472 1660
rect 9472 1604 9528 1660
rect 9528 1604 9532 1660
rect 9468 1600 9532 1604
rect 9548 1660 9612 1664
rect 9548 1604 9552 1660
rect 9552 1604 9608 1660
rect 9608 1604 9612 1660
rect 9548 1600 9612 1604
rect 12408 1660 12472 1664
rect 12408 1604 12412 1660
rect 12412 1604 12468 1660
rect 12468 1604 12472 1660
rect 12408 1600 12472 1604
rect 12488 1660 12552 1664
rect 12488 1604 12492 1660
rect 12492 1604 12548 1660
rect 12548 1604 12552 1660
rect 12488 1600 12552 1604
rect 12568 1660 12632 1664
rect 12568 1604 12572 1660
rect 12572 1604 12628 1660
rect 12628 1604 12632 1660
rect 12568 1600 12632 1604
rect 12648 1660 12712 1664
rect 12648 1604 12652 1660
rect 12652 1604 12708 1660
rect 12708 1604 12712 1660
rect 12648 1600 12712 1604
rect 15508 1660 15572 1664
rect 15508 1604 15512 1660
rect 15512 1604 15568 1660
rect 15568 1604 15572 1660
rect 15508 1600 15572 1604
rect 15588 1660 15652 1664
rect 15588 1604 15592 1660
rect 15592 1604 15648 1660
rect 15648 1604 15652 1660
rect 15588 1600 15652 1604
rect 15668 1660 15732 1664
rect 15668 1604 15672 1660
rect 15672 1604 15728 1660
rect 15728 1604 15732 1660
rect 15668 1600 15732 1604
rect 15748 1660 15812 1664
rect 15748 1604 15752 1660
rect 15752 1604 15808 1660
rect 15808 1604 15812 1660
rect 15748 1600 15812 1604
rect 18608 1660 18672 1664
rect 18608 1604 18612 1660
rect 18612 1604 18668 1660
rect 18668 1604 18672 1660
rect 18608 1600 18672 1604
rect 18688 1660 18752 1664
rect 18688 1604 18692 1660
rect 18692 1604 18748 1660
rect 18748 1604 18752 1660
rect 18688 1600 18752 1604
rect 18768 1660 18832 1664
rect 18768 1604 18772 1660
rect 18772 1604 18828 1660
rect 18828 1604 18832 1660
rect 18768 1600 18832 1604
rect 18848 1660 18912 1664
rect 18848 1604 18852 1660
rect 18852 1604 18908 1660
rect 18908 1604 18912 1660
rect 18848 1600 18912 1604
rect 1558 1116 1622 1120
rect 1558 1060 1562 1116
rect 1562 1060 1618 1116
rect 1618 1060 1622 1116
rect 1558 1056 1622 1060
rect 1638 1116 1702 1120
rect 1638 1060 1642 1116
rect 1642 1060 1698 1116
rect 1698 1060 1702 1116
rect 1638 1056 1702 1060
rect 1718 1116 1782 1120
rect 1718 1060 1722 1116
rect 1722 1060 1778 1116
rect 1778 1060 1782 1116
rect 1718 1056 1782 1060
rect 1798 1116 1862 1120
rect 1798 1060 1802 1116
rect 1802 1060 1858 1116
rect 1858 1060 1862 1116
rect 1798 1056 1862 1060
rect 4658 1116 4722 1120
rect 4658 1060 4662 1116
rect 4662 1060 4718 1116
rect 4718 1060 4722 1116
rect 4658 1056 4722 1060
rect 4738 1116 4802 1120
rect 4738 1060 4742 1116
rect 4742 1060 4798 1116
rect 4798 1060 4802 1116
rect 4738 1056 4802 1060
rect 4818 1116 4882 1120
rect 4818 1060 4822 1116
rect 4822 1060 4878 1116
rect 4878 1060 4882 1116
rect 4818 1056 4882 1060
rect 4898 1116 4962 1120
rect 4898 1060 4902 1116
rect 4902 1060 4958 1116
rect 4958 1060 4962 1116
rect 4898 1056 4962 1060
rect 7758 1116 7822 1120
rect 7758 1060 7762 1116
rect 7762 1060 7818 1116
rect 7818 1060 7822 1116
rect 7758 1056 7822 1060
rect 7838 1116 7902 1120
rect 7838 1060 7842 1116
rect 7842 1060 7898 1116
rect 7898 1060 7902 1116
rect 7838 1056 7902 1060
rect 7918 1116 7982 1120
rect 7918 1060 7922 1116
rect 7922 1060 7978 1116
rect 7978 1060 7982 1116
rect 7918 1056 7982 1060
rect 7998 1116 8062 1120
rect 7998 1060 8002 1116
rect 8002 1060 8058 1116
rect 8058 1060 8062 1116
rect 7998 1056 8062 1060
rect 10858 1116 10922 1120
rect 10858 1060 10862 1116
rect 10862 1060 10918 1116
rect 10918 1060 10922 1116
rect 10858 1056 10922 1060
rect 10938 1116 11002 1120
rect 10938 1060 10942 1116
rect 10942 1060 10998 1116
rect 10998 1060 11002 1116
rect 10938 1056 11002 1060
rect 11018 1116 11082 1120
rect 11018 1060 11022 1116
rect 11022 1060 11078 1116
rect 11078 1060 11082 1116
rect 11018 1056 11082 1060
rect 11098 1116 11162 1120
rect 11098 1060 11102 1116
rect 11102 1060 11158 1116
rect 11158 1060 11162 1116
rect 11098 1056 11162 1060
rect 13958 1116 14022 1120
rect 13958 1060 13962 1116
rect 13962 1060 14018 1116
rect 14018 1060 14022 1116
rect 13958 1056 14022 1060
rect 14038 1116 14102 1120
rect 14038 1060 14042 1116
rect 14042 1060 14098 1116
rect 14098 1060 14102 1116
rect 14038 1056 14102 1060
rect 14118 1116 14182 1120
rect 14118 1060 14122 1116
rect 14122 1060 14178 1116
rect 14178 1060 14182 1116
rect 14118 1056 14182 1060
rect 14198 1116 14262 1120
rect 14198 1060 14202 1116
rect 14202 1060 14258 1116
rect 14258 1060 14262 1116
rect 14198 1056 14262 1060
rect 17058 1116 17122 1120
rect 17058 1060 17062 1116
rect 17062 1060 17118 1116
rect 17118 1060 17122 1116
rect 17058 1056 17122 1060
rect 17138 1116 17202 1120
rect 17138 1060 17142 1116
rect 17142 1060 17198 1116
rect 17198 1060 17202 1116
rect 17138 1056 17202 1060
rect 17218 1116 17282 1120
rect 17218 1060 17222 1116
rect 17222 1060 17278 1116
rect 17278 1060 17282 1116
rect 17218 1056 17282 1060
rect 17298 1116 17362 1120
rect 17298 1060 17302 1116
rect 17302 1060 17358 1116
rect 17358 1060 17362 1116
rect 17298 1056 17362 1060
rect 3108 572 3172 576
rect 3108 516 3112 572
rect 3112 516 3168 572
rect 3168 516 3172 572
rect 3108 512 3172 516
rect 3188 572 3252 576
rect 3188 516 3192 572
rect 3192 516 3248 572
rect 3248 516 3252 572
rect 3188 512 3252 516
rect 3268 572 3332 576
rect 3268 516 3272 572
rect 3272 516 3328 572
rect 3328 516 3332 572
rect 3268 512 3332 516
rect 3348 572 3412 576
rect 3348 516 3352 572
rect 3352 516 3408 572
rect 3408 516 3412 572
rect 3348 512 3412 516
rect 6208 572 6272 576
rect 6208 516 6212 572
rect 6212 516 6268 572
rect 6268 516 6272 572
rect 6208 512 6272 516
rect 6288 572 6352 576
rect 6288 516 6292 572
rect 6292 516 6348 572
rect 6348 516 6352 572
rect 6288 512 6352 516
rect 6368 572 6432 576
rect 6368 516 6372 572
rect 6372 516 6428 572
rect 6428 516 6432 572
rect 6368 512 6432 516
rect 6448 572 6512 576
rect 6448 516 6452 572
rect 6452 516 6508 572
rect 6508 516 6512 572
rect 6448 512 6512 516
rect 9308 572 9372 576
rect 9308 516 9312 572
rect 9312 516 9368 572
rect 9368 516 9372 572
rect 9308 512 9372 516
rect 9388 572 9452 576
rect 9388 516 9392 572
rect 9392 516 9448 572
rect 9448 516 9452 572
rect 9388 512 9452 516
rect 9468 572 9532 576
rect 9468 516 9472 572
rect 9472 516 9528 572
rect 9528 516 9532 572
rect 9468 512 9532 516
rect 9548 572 9612 576
rect 9548 516 9552 572
rect 9552 516 9608 572
rect 9608 516 9612 572
rect 9548 512 9612 516
rect 12408 572 12472 576
rect 12408 516 12412 572
rect 12412 516 12468 572
rect 12468 516 12472 572
rect 12408 512 12472 516
rect 12488 572 12552 576
rect 12488 516 12492 572
rect 12492 516 12548 572
rect 12548 516 12552 572
rect 12488 512 12552 516
rect 12568 572 12632 576
rect 12568 516 12572 572
rect 12572 516 12628 572
rect 12628 516 12632 572
rect 12568 512 12632 516
rect 12648 572 12712 576
rect 12648 516 12652 572
rect 12652 516 12708 572
rect 12708 516 12712 572
rect 12648 512 12712 516
rect 15508 572 15572 576
rect 15508 516 15512 572
rect 15512 516 15568 572
rect 15568 516 15572 572
rect 15508 512 15572 516
rect 15588 572 15652 576
rect 15588 516 15592 572
rect 15592 516 15648 572
rect 15648 516 15652 572
rect 15588 512 15652 516
rect 15668 572 15732 576
rect 15668 516 15672 572
rect 15672 516 15728 572
rect 15728 516 15732 572
rect 15668 512 15732 516
rect 15748 572 15812 576
rect 15748 516 15752 572
rect 15752 516 15808 572
rect 15808 516 15812 572
rect 15748 512 15812 516
rect 18608 572 18672 576
rect 18608 516 18612 572
rect 18612 516 18668 572
rect 18668 516 18672 572
rect 18608 512 18672 516
rect 18688 572 18752 576
rect 18688 516 18692 572
rect 18692 516 18748 572
rect 18748 516 18752 572
rect 18688 512 18752 516
rect 18768 572 18832 576
rect 18768 516 18772 572
rect 18772 516 18828 572
rect 18828 516 18832 572
rect 18768 512 18832 516
rect 18848 572 18912 576
rect 18848 516 18852 572
rect 18852 516 18908 572
rect 18908 516 18912 572
rect 18848 512 18912 516
<< metal4 >>
rect 1550 18528 1870 18544
rect 1550 18464 1558 18528
rect 1622 18464 1638 18528
rect 1702 18464 1718 18528
rect 1782 18464 1798 18528
rect 1862 18464 1870 18528
rect 1550 17440 1870 18464
rect 1550 17376 1558 17440
rect 1622 17376 1638 17440
rect 1702 17376 1718 17440
rect 1782 17376 1798 17440
rect 1862 17376 1870 17440
rect 1550 16352 1870 17376
rect 1550 16288 1558 16352
rect 1622 16288 1638 16352
rect 1702 16288 1718 16352
rect 1782 16288 1798 16352
rect 1862 16288 1870 16352
rect 1550 15264 1870 16288
rect 1550 15200 1558 15264
rect 1622 15200 1638 15264
rect 1702 15200 1718 15264
rect 1782 15200 1798 15264
rect 1862 15200 1870 15264
rect 1550 14176 1870 15200
rect 1550 14112 1558 14176
rect 1622 14112 1638 14176
rect 1702 14112 1718 14176
rect 1782 14112 1798 14176
rect 1862 14112 1870 14176
rect 1550 13088 1870 14112
rect 1550 13024 1558 13088
rect 1622 13024 1638 13088
rect 1702 13024 1718 13088
rect 1782 13024 1798 13088
rect 1862 13024 1870 13088
rect 1550 12000 1870 13024
rect 1550 11936 1558 12000
rect 1622 11936 1638 12000
rect 1702 11936 1718 12000
rect 1782 11936 1798 12000
rect 1862 11936 1870 12000
rect 1550 10912 1870 11936
rect 1550 10848 1558 10912
rect 1622 10848 1638 10912
rect 1702 10848 1718 10912
rect 1782 10848 1798 10912
rect 1862 10848 1870 10912
rect 1550 9824 1870 10848
rect 1550 9760 1558 9824
rect 1622 9760 1638 9824
rect 1702 9760 1718 9824
rect 1782 9760 1798 9824
rect 1862 9760 1870 9824
rect 1550 8736 1870 9760
rect 1550 8672 1558 8736
rect 1622 8672 1638 8736
rect 1702 8672 1718 8736
rect 1782 8672 1798 8736
rect 1862 8672 1870 8736
rect 1550 7648 1870 8672
rect 1550 7584 1558 7648
rect 1622 7584 1638 7648
rect 1702 7584 1718 7648
rect 1782 7584 1798 7648
rect 1862 7584 1870 7648
rect 1550 6560 1870 7584
rect 1550 6496 1558 6560
rect 1622 6496 1638 6560
rect 1702 6496 1718 6560
rect 1782 6496 1798 6560
rect 1862 6496 1870 6560
rect 1550 5472 1870 6496
rect 1550 5408 1558 5472
rect 1622 5408 1638 5472
rect 1702 5408 1718 5472
rect 1782 5408 1798 5472
rect 1862 5408 1870 5472
rect 1550 4384 1870 5408
rect 1550 4320 1558 4384
rect 1622 4320 1638 4384
rect 1702 4320 1718 4384
rect 1782 4320 1798 4384
rect 1862 4320 1870 4384
rect 1550 3296 1870 4320
rect 1550 3232 1558 3296
rect 1622 3232 1638 3296
rect 1702 3232 1718 3296
rect 1782 3232 1798 3296
rect 1862 3232 1870 3296
rect 1550 2208 1870 3232
rect 1550 2144 1558 2208
rect 1622 2144 1638 2208
rect 1702 2144 1718 2208
rect 1782 2144 1798 2208
rect 1862 2144 1870 2208
rect 1550 1120 1870 2144
rect 1550 1056 1558 1120
rect 1622 1056 1638 1120
rect 1702 1056 1718 1120
rect 1782 1056 1798 1120
rect 1862 1056 1870 1120
rect 1550 496 1870 1056
rect 3100 17984 3420 18544
rect 3100 17920 3108 17984
rect 3172 17920 3188 17984
rect 3252 17920 3268 17984
rect 3332 17920 3348 17984
rect 3412 17920 3420 17984
rect 3100 16896 3420 17920
rect 3100 16832 3108 16896
rect 3172 16832 3188 16896
rect 3252 16832 3268 16896
rect 3332 16832 3348 16896
rect 3412 16832 3420 16896
rect 3100 15808 3420 16832
rect 3100 15744 3108 15808
rect 3172 15744 3188 15808
rect 3252 15744 3268 15808
rect 3332 15744 3348 15808
rect 3412 15744 3420 15808
rect 3100 14720 3420 15744
rect 3100 14656 3108 14720
rect 3172 14656 3188 14720
rect 3252 14656 3268 14720
rect 3332 14656 3348 14720
rect 3412 14656 3420 14720
rect 3100 13632 3420 14656
rect 3100 13568 3108 13632
rect 3172 13568 3188 13632
rect 3252 13568 3268 13632
rect 3332 13568 3348 13632
rect 3412 13568 3420 13632
rect 3100 12544 3420 13568
rect 3100 12480 3108 12544
rect 3172 12480 3188 12544
rect 3252 12480 3268 12544
rect 3332 12480 3348 12544
rect 3412 12480 3420 12544
rect 3100 11456 3420 12480
rect 3100 11392 3108 11456
rect 3172 11392 3188 11456
rect 3252 11392 3268 11456
rect 3332 11392 3348 11456
rect 3412 11392 3420 11456
rect 3100 10368 3420 11392
rect 3100 10304 3108 10368
rect 3172 10304 3188 10368
rect 3252 10304 3268 10368
rect 3332 10304 3348 10368
rect 3412 10304 3420 10368
rect 3100 9280 3420 10304
rect 3100 9216 3108 9280
rect 3172 9216 3188 9280
rect 3252 9216 3268 9280
rect 3332 9216 3348 9280
rect 3412 9216 3420 9280
rect 3100 8192 3420 9216
rect 3100 8128 3108 8192
rect 3172 8128 3188 8192
rect 3252 8128 3268 8192
rect 3332 8128 3348 8192
rect 3412 8128 3420 8192
rect 3100 7104 3420 8128
rect 3100 7040 3108 7104
rect 3172 7040 3188 7104
rect 3252 7040 3268 7104
rect 3332 7040 3348 7104
rect 3412 7040 3420 7104
rect 3100 6016 3420 7040
rect 3100 5952 3108 6016
rect 3172 5952 3188 6016
rect 3252 5952 3268 6016
rect 3332 5952 3348 6016
rect 3412 5952 3420 6016
rect 3100 4928 3420 5952
rect 3100 4864 3108 4928
rect 3172 4864 3188 4928
rect 3252 4864 3268 4928
rect 3332 4864 3348 4928
rect 3412 4864 3420 4928
rect 3100 3840 3420 4864
rect 3100 3776 3108 3840
rect 3172 3776 3188 3840
rect 3252 3776 3268 3840
rect 3332 3776 3348 3840
rect 3412 3776 3420 3840
rect 3100 2752 3420 3776
rect 3100 2688 3108 2752
rect 3172 2688 3188 2752
rect 3252 2688 3268 2752
rect 3332 2688 3348 2752
rect 3412 2688 3420 2752
rect 3100 1664 3420 2688
rect 3100 1600 3108 1664
rect 3172 1600 3188 1664
rect 3252 1600 3268 1664
rect 3332 1600 3348 1664
rect 3412 1600 3420 1664
rect 3100 576 3420 1600
rect 3100 512 3108 576
rect 3172 512 3188 576
rect 3252 512 3268 576
rect 3332 512 3348 576
rect 3412 512 3420 576
rect 3100 496 3420 512
rect 4650 18528 4970 18544
rect 4650 18464 4658 18528
rect 4722 18464 4738 18528
rect 4802 18464 4818 18528
rect 4882 18464 4898 18528
rect 4962 18464 4970 18528
rect 4650 17440 4970 18464
rect 4650 17376 4658 17440
rect 4722 17376 4738 17440
rect 4802 17376 4818 17440
rect 4882 17376 4898 17440
rect 4962 17376 4970 17440
rect 4650 16352 4970 17376
rect 4650 16288 4658 16352
rect 4722 16288 4738 16352
rect 4802 16288 4818 16352
rect 4882 16288 4898 16352
rect 4962 16288 4970 16352
rect 4650 15264 4970 16288
rect 4650 15200 4658 15264
rect 4722 15200 4738 15264
rect 4802 15200 4818 15264
rect 4882 15200 4898 15264
rect 4962 15200 4970 15264
rect 4650 14176 4970 15200
rect 4650 14112 4658 14176
rect 4722 14112 4738 14176
rect 4802 14112 4818 14176
rect 4882 14112 4898 14176
rect 4962 14112 4970 14176
rect 4650 13088 4970 14112
rect 4650 13024 4658 13088
rect 4722 13024 4738 13088
rect 4802 13024 4818 13088
rect 4882 13024 4898 13088
rect 4962 13024 4970 13088
rect 4650 12000 4970 13024
rect 4650 11936 4658 12000
rect 4722 11936 4738 12000
rect 4802 11936 4818 12000
rect 4882 11936 4898 12000
rect 4962 11936 4970 12000
rect 4650 10912 4970 11936
rect 4650 10848 4658 10912
rect 4722 10848 4738 10912
rect 4802 10848 4818 10912
rect 4882 10848 4898 10912
rect 4962 10848 4970 10912
rect 4650 9824 4970 10848
rect 4650 9760 4658 9824
rect 4722 9760 4738 9824
rect 4802 9760 4818 9824
rect 4882 9760 4898 9824
rect 4962 9760 4970 9824
rect 4650 8736 4970 9760
rect 4650 8672 4658 8736
rect 4722 8672 4738 8736
rect 4802 8672 4818 8736
rect 4882 8672 4898 8736
rect 4962 8672 4970 8736
rect 4650 7648 4970 8672
rect 4650 7584 4658 7648
rect 4722 7584 4738 7648
rect 4802 7584 4818 7648
rect 4882 7584 4898 7648
rect 4962 7584 4970 7648
rect 4650 6560 4970 7584
rect 4650 6496 4658 6560
rect 4722 6496 4738 6560
rect 4802 6496 4818 6560
rect 4882 6496 4898 6560
rect 4962 6496 4970 6560
rect 4650 5472 4970 6496
rect 4650 5408 4658 5472
rect 4722 5408 4738 5472
rect 4802 5408 4818 5472
rect 4882 5408 4898 5472
rect 4962 5408 4970 5472
rect 4650 4384 4970 5408
rect 4650 4320 4658 4384
rect 4722 4320 4738 4384
rect 4802 4320 4818 4384
rect 4882 4320 4898 4384
rect 4962 4320 4970 4384
rect 4650 3296 4970 4320
rect 4650 3232 4658 3296
rect 4722 3232 4738 3296
rect 4802 3232 4818 3296
rect 4882 3232 4898 3296
rect 4962 3232 4970 3296
rect 4650 2208 4970 3232
rect 4650 2144 4658 2208
rect 4722 2144 4738 2208
rect 4802 2144 4818 2208
rect 4882 2144 4898 2208
rect 4962 2144 4970 2208
rect 4650 1120 4970 2144
rect 4650 1056 4658 1120
rect 4722 1056 4738 1120
rect 4802 1056 4818 1120
rect 4882 1056 4898 1120
rect 4962 1056 4970 1120
rect 4650 496 4970 1056
rect 6200 17984 6520 18544
rect 6200 17920 6208 17984
rect 6272 17920 6288 17984
rect 6352 17920 6368 17984
rect 6432 17920 6448 17984
rect 6512 17920 6520 17984
rect 6200 16896 6520 17920
rect 6200 16832 6208 16896
rect 6272 16832 6288 16896
rect 6352 16832 6368 16896
rect 6432 16832 6448 16896
rect 6512 16832 6520 16896
rect 6200 15808 6520 16832
rect 6200 15744 6208 15808
rect 6272 15744 6288 15808
rect 6352 15744 6368 15808
rect 6432 15744 6448 15808
rect 6512 15744 6520 15808
rect 6200 14720 6520 15744
rect 6200 14656 6208 14720
rect 6272 14656 6288 14720
rect 6352 14656 6368 14720
rect 6432 14656 6448 14720
rect 6512 14656 6520 14720
rect 6200 13632 6520 14656
rect 6200 13568 6208 13632
rect 6272 13568 6288 13632
rect 6352 13568 6368 13632
rect 6432 13568 6448 13632
rect 6512 13568 6520 13632
rect 6200 12544 6520 13568
rect 6200 12480 6208 12544
rect 6272 12480 6288 12544
rect 6352 12480 6368 12544
rect 6432 12480 6448 12544
rect 6512 12480 6520 12544
rect 6200 11456 6520 12480
rect 6200 11392 6208 11456
rect 6272 11392 6288 11456
rect 6352 11392 6368 11456
rect 6432 11392 6448 11456
rect 6512 11392 6520 11456
rect 6200 10368 6520 11392
rect 6200 10304 6208 10368
rect 6272 10304 6288 10368
rect 6352 10304 6368 10368
rect 6432 10304 6448 10368
rect 6512 10304 6520 10368
rect 6200 9280 6520 10304
rect 6200 9216 6208 9280
rect 6272 9216 6288 9280
rect 6352 9216 6368 9280
rect 6432 9216 6448 9280
rect 6512 9216 6520 9280
rect 6200 8192 6520 9216
rect 6200 8128 6208 8192
rect 6272 8128 6288 8192
rect 6352 8128 6368 8192
rect 6432 8128 6448 8192
rect 6512 8128 6520 8192
rect 6200 7104 6520 8128
rect 6200 7040 6208 7104
rect 6272 7040 6288 7104
rect 6352 7040 6368 7104
rect 6432 7040 6448 7104
rect 6512 7040 6520 7104
rect 6200 6016 6520 7040
rect 6200 5952 6208 6016
rect 6272 5952 6288 6016
rect 6352 5952 6368 6016
rect 6432 5952 6448 6016
rect 6512 5952 6520 6016
rect 6200 4928 6520 5952
rect 6200 4864 6208 4928
rect 6272 4864 6288 4928
rect 6352 4864 6368 4928
rect 6432 4864 6448 4928
rect 6512 4864 6520 4928
rect 6200 3840 6520 4864
rect 6200 3776 6208 3840
rect 6272 3776 6288 3840
rect 6352 3776 6368 3840
rect 6432 3776 6448 3840
rect 6512 3776 6520 3840
rect 6200 2752 6520 3776
rect 6200 2688 6208 2752
rect 6272 2688 6288 2752
rect 6352 2688 6368 2752
rect 6432 2688 6448 2752
rect 6512 2688 6520 2752
rect 6200 1664 6520 2688
rect 6200 1600 6208 1664
rect 6272 1600 6288 1664
rect 6352 1600 6368 1664
rect 6432 1600 6448 1664
rect 6512 1600 6520 1664
rect 6200 576 6520 1600
rect 6200 512 6208 576
rect 6272 512 6288 576
rect 6352 512 6368 576
rect 6432 512 6448 576
rect 6512 512 6520 576
rect 6200 496 6520 512
rect 7750 18528 8070 18544
rect 7750 18464 7758 18528
rect 7822 18464 7838 18528
rect 7902 18464 7918 18528
rect 7982 18464 7998 18528
rect 8062 18464 8070 18528
rect 7750 17440 8070 18464
rect 7750 17376 7758 17440
rect 7822 17376 7838 17440
rect 7902 17376 7918 17440
rect 7982 17376 7998 17440
rect 8062 17376 8070 17440
rect 7750 16352 8070 17376
rect 7750 16288 7758 16352
rect 7822 16288 7838 16352
rect 7902 16288 7918 16352
rect 7982 16288 7998 16352
rect 8062 16288 8070 16352
rect 7750 15264 8070 16288
rect 7750 15200 7758 15264
rect 7822 15200 7838 15264
rect 7902 15200 7918 15264
rect 7982 15200 7998 15264
rect 8062 15200 8070 15264
rect 7750 14176 8070 15200
rect 7750 14112 7758 14176
rect 7822 14112 7838 14176
rect 7902 14112 7918 14176
rect 7982 14112 7998 14176
rect 8062 14112 8070 14176
rect 7750 13088 8070 14112
rect 7750 13024 7758 13088
rect 7822 13024 7838 13088
rect 7902 13024 7918 13088
rect 7982 13024 7998 13088
rect 8062 13024 8070 13088
rect 7750 12000 8070 13024
rect 7750 11936 7758 12000
rect 7822 11936 7838 12000
rect 7902 11936 7918 12000
rect 7982 11936 7998 12000
rect 8062 11936 8070 12000
rect 7750 10912 8070 11936
rect 7750 10848 7758 10912
rect 7822 10848 7838 10912
rect 7902 10848 7918 10912
rect 7982 10848 7998 10912
rect 8062 10848 8070 10912
rect 7750 9824 8070 10848
rect 7750 9760 7758 9824
rect 7822 9760 7838 9824
rect 7902 9760 7918 9824
rect 7982 9760 7998 9824
rect 8062 9760 8070 9824
rect 7750 8736 8070 9760
rect 7750 8672 7758 8736
rect 7822 8672 7838 8736
rect 7902 8672 7918 8736
rect 7982 8672 7998 8736
rect 8062 8672 8070 8736
rect 7750 7648 8070 8672
rect 7750 7584 7758 7648
rect 7822 7584 7838 7648
rect 7902 7584 7918 7648
rect 7982 7584 7998 7648
rect 8062 7584 8070 7648
rect 7750 6560 8070 7584
rect 7750 6496 7758 6560
rect 7822 6496 7838 6560
rect 7902 6496 7918 6560
rect 7982 6496 7998 6560
rect 8062 6496 8070 6560
rect 7750 5472 8070 6496
rect 7750 5408 7758 5472
rect 7822 5408 7838 5472
rect 7902 5408 7918 5472
rect 7982 5408 7998 5472
rect 8062 5408 8070 5472
rect 7750 4384 8070 5408
rect 7750 4320 7758 4384
rect 7822 4320 7838 4384
rect 7902 4320 7918 4384
rect 7982 4320 7998 4384
rect 8062 4320 8070 4384
rect 7750 3296 8070 4320
rect 7750 3232 7758 3296
rect 7822 3232 7838 3296
rect 7902 3232 7918 3296
rect 7982 3232 7998 3296
rect 8062 3232 8070 3296
rect 7750 2208 8070 3232
rect 7750 2144 7758 2208
rect 7822 2144 7838 2208
rect 7902 2144 7918 2208
rect 7982 2144 7998 2208
rect 8062 2144 8070 2208
rect 7750 1120 8070 2144
rect 7750 1056 7758 1120
rect 7822 1056 7838 1120
rect 7902 1056 7918 1120
rect 7982 1056 7998 1120
rect 8062 1056 8070 1120
rect 7750 496 8070 1056
rect 9300 17984 9620 18544
rect 9300 17920 9308 17984
rect 9372 17920 9388 17984
rect 9452 17920 9468 17984
rect 9532 17920 9548 17984
rect 9612 17920 9620 17984
rect 9300 16896 9620 17920
rect 9300 16832 9308 16896
rect 9372 16832 9388 16896
rect 9452 16832 9468 16896
rect 9532 16832 9548 16896
rect 9612 16832 9620 16896
rect 9300 15808 9620 16832
rect 9300 15744 9308 15808
rect 9372 15744 9388 15808
rect 9452 15744 9468 15808
rect 9532 15744 9548 15808
rect 9612 15744 9620 15808
rect 9300 14720 9620 15744
rect 9300 14656 9308 14720
rect 9372 14656 9388 14720
rect 9452 14656 9468 14720
rect 9532 14656 9548 14720
rect 9612 14656 9620 14720
rect 9300 13632 9620 14656
rect 9300 13568 9308 13632
rect 9372 13568 9388 13632
rect 9452 13568 9468 13632
rect 9532 13568 9548 13632
rect 9612 13568 9620 13632
rect 9300 12544 9620 13568
rect 9300 12480 9308 12544
rect 9372 12480 9388 12544
rect 9452 12480 9468 12544
rect 9532 12480 9548 12544
rect 9612 12480 9620 12544
rect 9300 11456 9620 12480
rect 9300 11392 9308 11456
rect 9372 11392 9388 11456
rect 9452 11392 9468 11456
rect 9532 11392 9548 11456
rect 9612 11392 9620 11456
rect 9300 10368 9620 11392
rect 9300 10304 9308 10368
rect 9372 10304 9388 10368
rect 9452 10304 9468 10368
rect 9532 10304 9548 10368
rect 9612 10304 9620 10368
rect 9300 9280 9620 10304
rect 9300 9216 9308 9280
rect 9372 9216 9388 9280
rect 9452 9216 9468 9280
rect 9532 9216 9548 9280
rect 9612 9216 9620 9280
rect 9300 8192 9620 9216
rect 9300 8128 9308 8192
rect 9372 8128 9388 8192
rect 9452 8128 9468 8192
rect 9532 8128 9548 8192
rect 9612 8128 9620 8192
rect 9300 7104 9620 8128
rect 9300 7040 9308 7104
rect 9372 7040 9388 7104
rect 9452 7040 9468 7104
rect 9532 7040 9548 7104
rect 9612 7040 9620 7104
rect 9300 6016 9620 7040
rect 9300 5952 9308 6016
rect 9372 5952 9388 6016
rect 9452 5952 9468 6016
rect 9532 5952 9548 6016
rect 9612 5952 9620 6016
rect 9300 4928 9620 5952
rect 9300 4864 9308 4928
rect 9372 4864 9388 4928
rect 9452 4864 9468 4928
rect 9532 4864 9548 4928
rect 9612 4864 9620 4928
rect 9300 3840 9620 4864
rect 9300 3776 9308 3840
rect 9372 3776 9388 3840
rect 9452 3776 9468 3840
rect 9532 3776 9548 3840
rect 9612 3776 9620 3840
rect 9300 2752 9620 3776
rect 9300 2688 9308 2752
rect 9372 2688 9388 2752
rect 9452 2688 9468 2752
rect 9532 2688 9548 2752
rect 9612 2688 9620 2752
rect 9300 1664 9620 2688
rect 9300 1600 9308 1664
rect 9372 1600 9388 1664
rect 9452 1600 9468 1664
rect 9532 1600 9548 1664
rect 9612 1600 9620 1664
rect 9300 576 9620 1600
rect 9300 512 9308 576
rect 9372 512 9388 576
rect 9452 512 9468 576
rect 9532 512 9548 576
rect 9612 512 9620 576
rect 9300 496 9620 512
rect 10850 18528 11170 18544
rect 10850 18464 10858 18528
rect 10922 18464 10938 18528
rect 11002 18464 11018 18528
rect 11082 18464 11098 18528
rect 11162 18464 11170 18528
rect 10850 17440 11170 18464
rect 10850 17376 10858 17440
rect 10922 17376 10938 17440
rect 11002 17376 11018 17440
rect 11082 17376 11098 17440
rect 11162 17376 11170 17440
rect 10850 16352 11170 17376
rect 10850 16288 10858 16352
rect 10922 16288 10938 16352
rect 11002 16288 11018 16352
rect 11082 16288 11098 16352
rect 11162 16288 11170 16352
rect 10850 15264 11170 16288
rect 10850 15200 10858 15264
rect 10922 15200 10938 15264
rect 11002 15200 11018 15264
rect 11082 15200 11098 15264
rect 11162 15200 11170 15264
rect 10850 14176 11170 15200
rect 10850 14112 10858 14176
rect 10922 14112 10938 14176
rect 11002 14112 11018 14176
rect 11082 14112 11098 14176
rect 11162 14112 11170 14176
rect 10850 13088 11170 14112
rect 10850 13024 10858 13088
rect 10922 13024 10938 13088
rect 11002 13024 11018 13088
rect 11082 13024 11098 13088
rect 11162 13024 11170 13088
rect 10850 12000 11170 13024
rect 10850 11936 10858 12000
rect 10922 11936 10938 12000
rect 11002 11936 11018 12000
rect 11082 11936 11098 12000
rect 11162 11936 11170 12000
rect 10850 10912 11170 11936
rect 10850 10848 10858 10912
rect 10922 10848 10938 10912
rect 11002 10848 11018 10912
rect 11082 10848 11098 10912
rect 11162 10848 11170 10912
rect 10850 9824 11170 10848
rect 10850 9760 10858 9824
rect 10922 9760 10938 9824
rect 11002 9760 11018 9824
rect 11082 9760 11098 9824
rect 11162 9760 11170 9824
rect 10850 8736 11170 9760
rect 10850 8672 10858 8736
rect 10922 8672 10938 8736
rect 11002 8672 11018 8736
rect 11082 8672 11098 8736
rect 11162 8672 11170 8736
rect 10850 7648 11170 8672
rect 10850 7584 10858 7648
rect 10922 7584 10938 7648
rect 11002 7584 11018 7648
rect 11082 7584 11098 7648
rect 11162 7584 11170 7648
rect 10850 6560 11170 7584
rect 10850 6496 10858 6560
rect 10922 6496 10938 6560
rect 11002 6496 11018 6560
rect 11082 6496 11098 6560
rect 11162 6496 11170 6560
rect 10850 5472 11170 6496
rect 10850 5408 10858 5472
rect 10922 5408 10938 5472
rect 11002 5408 11018 5472
rect 11082 5408 11098 5472
rect 11162 5408 11170 5472
rect 10850 4384 11170 5408
rect 10850 4320 10858 4384
rect 10922 4320 10938 4384
rect 11002 4320 11018 4384
rect 11082 4320 11098 4384
rect 11162 4320 11170 4384
rect 10850 3296 11170 4320
rect 10850 3232 10858 3296
rect 10922 3232 10938 3296
rect 11002 3232 11018 3296
rect 11082 3232 11098 3296
rect 11162 3232 11170 3296
rect 10850 2208 11170 3232
rect 10850 2144 10858 2208
rect 10922 2144 10938 2208
rect 11002 2144 11018 2208
rect 11082 2144 11098 2208
rect 11162 2144 11170 2208
rect 10850 1120 11170 2144
rect 10850 1056 10858 1120
rect 10922 1056 10938 1120
rect 11002 1056 11018 1120
rect 11082 1056 11098 1120
rect 11162 1056 11170 1120
rect 10850 496 11170 1056
rect 12400 17984 12720 18544
rect 12400 17920 12408 17984
rect 12472 17920 12488 17984
rect 12552 17920 12568 17984
rect 12632 17920 12648 17984
rect 12712 17920 12720 17984
rect 12400 16896 12720 17920
rect 12400 16832 12408 16896
rect 12472 16832 12488 16896
rect 12552 16832 12568 16896
rect 12632 16832 12648 16896
rect 12712 16832 12720 16896
rect 12400 15808 12720 16832
rect 12400 15744 12408 15808
rect 12472 15744 12488 15808
rect 12552 15744 12568 15808
rect 12632 15744 12648 15808
rect 12712 15744 12720 15808
rect 12400 14720 12720 15744
rect 12400 14656 12408 14720
rect 12472 14656 12488 14720
rect 12552 14656 12568 14720
rect 12632 14656 12648 14720
rect 12712 14656 12720 14720
rect 12400 13632 12720 14656
rect 12400 13568 12408 13632
rect 12472 13568 12488 13632
rect 12552 13568 12568 13632
rect 12632 13568 12648 13632
rect 12712 13568 12720 13632
rect 12400 12544 12720 13568
rect 12400 12480 12408 12544
rect 12472 12480 12488 12544
rect 12552 12480 12568 12544
rect 12632 12480 12648 12544
rect 12712 12480 12720 12544
rect 12400 11456 12720 12480
rect 12400 11392 12408 11456
rect 12472 11392 12488 11456
rect 12552 11392 12568 11456
rect 12632 11392 12648 11456
rect 12712 11392 12720 11456
rect 12400 10368 12720 11392
rect 12400 10304 12408 10368
rect 12472 10304 12488 10368
rect 12552 10304 12568 10368
rect 12632 10304 12648 10368
rect 12712 10304 12720 10368
rect 12400 9280 12720 10304
rect 12400 9216 12408 9280
rect 12472 9216 12488 9280
rect 12552 9216 12568 9280
rect 12632 9216 12648 9280
rect 12712 9216 12720 9280
rect 12400 8192 12720 9216
rect 12400 8128 12408 8192
rect 12472 8128 12488 8192
rect 12552 8128 12568 8192
rect 12632 8128 12648 8192
rect 12712 8128 12720 8192
rect 12400 7104 12720 8128
rect 12400 7040 12408 7104
rect 12472 7040 12488 7104
rect 12552 7040 12568 7104
rect 12632 7040 12648 7104
rect 12712 7040 12720 7104
rect 12400 6016 12720 7040
rect 12400 5952 12408 6016
rect 12472 5952 12488 6016
rect 12552 5952 12568 6016
rect 12632 5952 12648 6016
rect 12712 5952 12720 6016
rect 12400 4928 12720 5952
rect 12400 4864 12408 4928
rect 12472 4864 12488 4928
rect 12552 4864 12568 4928
rect 12632 4864 12648 4928
rect 12712 4864 12720 4928
rect 12400 3840 12720 4864
rect 12400 3776 12408 3840
rect 12472 3776 12488 3840
rect 12552 3776 12568 3840
rect 12632 3776 12648 3840
rect 12712 3776 12720 3840
rect 12400 2752 12720 3776
rect 12400 2688 12408 2752
rect 12472 2688 12488 2752
rect 12552 2688 12568 2752
rect 12632 2688 12648 2752
rect 12712 2688 12720 2752
rect 12400 1664 12720 2688
rect 12400 1600 12408 1664
rect 12472 1600 12488 1664
rect 12552 1600 12568 1664
rect 12632 1600 12648 1664
rect 12712 1600 12720 1664
rect 12400 576 12720 1600
rect 12400 512 12408 576
rect 12472 512 12488 576
rect 12552 512 12568 576
rect 12632 512 12648 576
rect 12712 512 12720 576
rect 12400 496 12720 512
rect 13950 18528 14270 18544
rect 13950 18464 13958 18528
rect 14022 18464 14038 18528
rect 14102 18464 14118 18528
rect 14182 18464 14198 18528
rect 14262 18464 14270 18528
rect 13950 17440 14270 18464
rect 13950 17376 13958 17440
rect 14022 17376 14038 17440
rect 14102 17376 14118 17440
rect 14182 17376 14198 17440
rect 14262 17376 14270 17440
rect 13950 16352 14270 17376
rect 13950 16288 13958 16352
rect 14022 16288 14038 16352
rect 14102 16288 14118 16352
rect 14182 16288 14198 16352
rect 14262 16288 14270 16352
rect 13950 15264 14270 16288
rect 13950 15200 13958 15264
rect 14022 15200 14038 15264
rect 14102 15200 14118 15264
rect 14182 15200 14198 15264
rect 14262 15200 14270 15264
rect 13950 14176 14270 15200
rect 13950 14112 13958 14176
rect 14022 14112 14038 14176
rect 14102 14112 14118 14176
rect 14182 14112 14198 14176
rect 14262 14112 14270 14176
rect 13950 13088 14270 14112
rect 13950 13024 13958 13088
rect 14022 13024 14038 13088
rect 14102 13024 14118 13088
rect 14182 13024 14198 13088
rect 14262 13024 14270 13088
rect 13950 12000 14270 13024
rect 13950 11936 13958 12000
rect 14022 11936 14038 12000
rect 14102 11936 14118 12000
rect 14182 11936 14198 12000
rect 14262 11936 14270 12000
rect 13950 10912 14270 11936
rect 13950 10848 13958 10912
rect 14022 10848 14038 10912
rect 14102 10848 14118 10912
rect 14182 10848 14198 10912
rect 14262 10848 14270 10912
rect 13950 9824 14270 10848
rect 13950 9760 13958 9824
rect 14022 9760 14038 9824
rect 14102 9760 14118 9824
rect 14182 9760 14198 9824
rect 14262 9760 14270 9824
rect 13950 8736 14270 9760
rect 13950 8672 13958 8736
rect 14022 8672 14038 8736
rect 14102 8672 14118 8736
rect 14182 8672 14198 8736
rect 14262 8672 14270 8736
rect 13950 7648 14270 8672
rect 13950 7584 13958 7648
rect 14022 7584 14038 7648
rect 14102 7584 14118 7648
rect 14182 7584 14198 7648
rect 14262 7584 14270 7648
rect 13950 6560 14270 7584
rect 13950 6496 13958 6560
rect 14022 6496 14038 6560
rect 14102 6496 14118 6560
rect 14182 6496 14198 6560
rect 14262 6496 14270 6560
rect 13950 5472 14270 6496
rect 13950 5408 13958 5472
rect 14022 5408 14038 5472
rect 14102 5408 14118 5472
rect 14182 5408 14198 5472
rect 14262 5408 14270 5472
rect 13950 4384 14270 5408
rect 13950 4320 13958 4384
rect 14022 4320 14038 4384
rect 14102 4320 14118 4384
rect 14182 4320 14198 4384
rect 14262 4320 14270 4384
rect 13950 3296 14270 4320
rect 13950 3232 13958 3296
rect 14022 3232 14038 3296
rect 14102 3232 14118 3296
rect 14182 3232 14198 3296
rect 14262 3232 14270 3296
rect 13950 2208 14270 3232
rect 13950 2144 13958 2208
rect 14022 2144 14038 2208
rect 14102 2144 14118 2208
rect 14182 2144 14198 2208
rect 14262 2144 14270 2208
rect 13950 1120 14270 2144
rect 13950 1056 13958 1120
rect 14022 1056 14038 1120
rect 14102 1056 14118 1120
rect 14182 1056 14198 1120
rect 14262 1056 14270 1120
rect 13950 496 14270 1056
rect 15500 17984 15820 18544
rect 15500 17920 15508 17984
rect 15572 17920 15588 17984
rect 15652 17920 15668 17984
rect 15732 17920 15748 17984
rect 15812 17920 15820 17984
rect 15500 16896 15820 17920
rect 15500 16832 15508 16896
rect 15572 16832 15588 16896
rect 15652 16832 15668 16896
rect 15732 16832 15748 16896
rect 15812 16832 15820 16896
rect 15500 15808 15820 16832
rect 15500 15744 15508 15808
rect 15572 15744 15588 15808
rect 15652 15744 15668 15808
rect 15732 15744 15748 15808
rect 15812 15744 15820 15808
rect 15500 14720 15820 15744
rect 15500 14656 15508 14720
rect 15572 14656 15588 14720
rect 15652 14656 15668 14720
rect 15732 14656 15748 14720
rect 15812 14656 15820 14720
rect 15500 13632 15820 14656
rect 15500 13568 15508 13632
rect 15572 13568 15588 13632
rect 15652 13568 15668 13632
rect 15732 13568 15748 13632
rect 15812 13568 15820 13632
rect 15500 12544 15820 13568
rect 15500 12480 15508 12544
rect 15572 12480 15588 12544
rect 15652 12480 15668 12544
rect 15732 12480 15748 12544
rect 15812 12480 15820 12544
rect 15500 11456 15820 12480
rect 15500 11392 15508 11456
rect 15572 11392 15588 11456
rect 15652 11392 15668 11456
rect 15732 11392 15748 11456
rect 15812 11392 15820 11456
rect 15500 10368 15820 11392
rect 15500 10304 15508 10368
rect 15572 10304 15588 10368
rect 15652 10304 15668 10368
rect 15732 10304 15748 10368
rect 15812 10304 15820 10368
rect 15500 9280 15820 10304
rect 15500 9216 15508 9280
rect 15572 9216 15588 9280
rect 15652 9216 15668 9280
rect 15732 9216 15748 9280
rect 15812 9216 15820 9280
rect 15500 8192 15820 9216
rect 15500 8128 15508 8192
rect 15572 8128 15588 8192
rect 15652 8128 15668 8192
rect 15732 8128 15748 8192
rect 15812 8128 15820 8192
rect 15500 7104 15820 8128
rect 15500 7040 15508 7104
rect 15572 7040 15588 7104
rect 15652 7040 15668 7104
rect 15732 7040 15748 7104
rect 15812 7040 15820 7104
rect 15500 6016 15820 7040
rect 15500 5952 15508 6016
rect 15572 5952 15588 6016
rect 15652 5952 15668 6016
rect 15732 5952 15748 6016
rect 15812 5952 15820 6016
rect 15500 4928 15820 5952
rect 15500 4864 15508 4928
rect 15572 4864 15588 4928
rect 15652 4864 15668 4928
rect 15732 4864 15748 4928
rect 15812 4864 15820 4928
rect 15500 3840 15820 4864
rect 15500 3776 15508 3840
rect 15572 3776 15588 3840
rect 15652 3776 15668 3840
rect 15732 3776 15748 3840
rect 15812 3776 15820 3840
rect 15500 2752 15820 3776
rect 15500 2688 15508 2752
rect 15572 2688 15588 2752
rect 15652 2688 15668 2752
rect 15732 2688 15748 2752
rect 15812 2688 15820 2752
rect 15500 1664 15820 2688
rect 15500 1600 15508 1664
rect 15572 1600 15588 1664
rect 15652 1600 15668 1664
rect 15732 1600 15748 1664
rect 15812 1600 15820 1664
rect 15500 576 15820 1600
rect 15500 512 15508 576
rect 15572 512 15588 576
rect 15652 512 15668 576
rect 15732 512 15748 576
rect 15812 512 15820 576
rect 15500 496 15820 512
rect 17050 18528 17370 18544
rect 17050 18464 17058 18528
rect 17122 18464 17138 18528
rect 17202 18464 17218 18528
rect 17282 18464 17298 18528
rect 17362 18464 17370 18528
rect 17050 17440 17370 18464
rect 17050 17376 17058 17440
rect 17122 17376 17138 17440
rect 17202 17376 17218 17440
rect 17282 17376 17298 17440
rect 17362 17376 17370 17440
rect 17050 16352 17370 17376
rect 17050 16288 17058 16352
rect 17122 16288 17138 16352
rect 17202 16288 17218 16352
rect 17282 16288 17298 16352
rect 17362 16288 17370 16352
rect 17050 15264 17370 16288
rect 17050 15200 17058 15264
rect 17122 15200 17138 15264
rect 17202 15200 17218 15264
rect 17282 15200 17298 15264
rect 17362 15200 17370 15264
rect 17050 14176 17370 15200
rect 17050 14112 17058 14176
rect 17122 14112 17138 14176
rect 17202 14112 17218 14176
rect 17282 14112 17298 14176
rect 17362 14112 17370 14176
rect 17050 13088 17370 14112
rect 17050 13024 17058 13088
rect 17122 13024 17138 13088
rect 17202 13024 17218 13088
rect 17282 13024 17298 13088
rect 17362 13024 17370 13088
rect 17050 12000 17370 13024
rect 17050 11936 17058 12000
rect 17122 11936 17138 12000
rect 17202 11936 17218 12000
rect 17282 11936 17298 12000
rect 17362 11936 17370 12000
rect 17050 10912 17370 11936
rect 17050 10848 17058 10912
rect 17122 10848 17138 10912
rect 17202 10848 17218 10912
rect 17282 10848 17298 10912
rect 17362 10848 17370 10912
rect 17050 9824 17370 10848
rect 17050 9760 17058 9824
rect 17122 9760 17138 9824
rect 17202 9760 17218 9824
rect 17282 9760 17298 9824
rect 17362 9760 17370 9824
rect 17050 8736 17370 9760
rect 17050 8672 17058 8736
rect 17122 8672 17138 8736
rect 17202 8672 17218 8736
rect 17282 8672 17298 8736
rect 17362 8672 17370 8736
rect 17050 7648 17370 8672
rect 17050 7584 17058 7648
rect 17122 7584 17138 7648
rect 17202 7584 17218 7648
rect 17282 7584 17298 7648
rect 17362 7584 17370 7648
rect 17050 6560 17370 7584
rect 17050 6496 17058 6560
rect 17122 6496 17138 6560
rect 17202 6496 17218 6560
rect 17282 6496 17298 6560
rect 17362 6496 17370 6560
rect 17050 5472 17370 6496
rect 17050 5408 17058 5472
rect 17122 5408 17138 5472
rect 17202 5408 17218 5472
rect 17282 5408 17298 5472
rect 17362 5408 17370 5472
rect 17050 4384 17370 5408
rect 17050 4320 17058 4384
rect 17122 4320 17138 4384
rect 17202 4320 17218 4384
rect 17282 4320 17298 4384
rect 17362 4320 17370 4384
rect 17050 3296 17370 4320
rect 17050 3232 17058 3296
rect 17122 3232 17138 3296
rect 17202 3232 17218 3296
rect 17282 3232 17298 3296
rect 17362 3232 17370 3296
rect 17050 2208 17370 3232
rect 17050 2144 17058 2208
rect 17122 2144 17138 2208
rect 17202 2144 17218 2208
rect 17282 2144 17298 2208
rect 17362 2144 17370 2208
rect 17050 1120 17370 2144
rect 17050 1056 17058 1120
rect 17122 1056 17138 1120
rect 17202 1056 17218 1120
rect 17282 1056 17298 1120
rect 17362 1056 17370 1120
rect 17050 496 17370 1056
rect 18600 17984 18920 18544
rect 18600 17920 18608 17984
rect 18672 17920 18688 17984
rect 18752 17920 18768 17984
rect 18832 17920 18848 17984
rect 18912 17920 18920 17984
rect 18600 16896 18920 17920
rect 18600 16832 18608 16896
rect 18672 16832 18688 16896
rect 18752 16832 18768 16896
rect 18832 16832 18848 16896
rect 18912 16832 18920 16896
rect 18600 15808 18920 16832
rect 18600 15744 18608 15808
rect 18672 15744 18688 15808
rect 18752 15744 18768 15808
rect 18832 15744 18848 15808
rect 18912 15744 18920 15808
rect 18600 14720 18920 15744
rect 18600 14656 18608 14720
rect 18672 14656 18688 14720
rect 18752 14656 18768 14720
rect 18832 14656 18848 14720
rect 18912 14656 18920 14720
rect 18600 13632 18920 14656
rect 18600 13568 18608 13632
rect 18672 13568 18688 13632
rect 18752 13568 18768 13632
rect 18832 13568 18848 13632
rect 18912 13568 18920 13632
rect 18600 12544 18920 13568
rect 18600 12480 18608 12544
rect 18672 12480 18688 12544
rect 18752 12480 18768 12544
rect 18832 12480 18848 12544
rect 18912 12480 18920 12544
rect 18600 11456 18920 12480
rect 18600 11392 18608 11456
rect 18672 11392 18688 11456
rect 18752 11392 18768 11456
rect 18832 11392 18848 11456
rect 18912 11392 18920 11456
rect 18600 10368 18920 11392
rect 18600 10304 18608 10368
rect 18672 10304 18688 10368
rect 18752 10304 18768 10368
rect 18832 10304 18848 10368
rect 18912 10304 18920 10368
rect 18600 9280 18920 10304
rect 18600 9216 18608 9280
rect 18672 9216 18688 9280
rect 18752 9216 18768 9280
rect 18832 9216 18848 9280
rect 18912 9216 18920 9280
rect 18600 8192 18920 9216
rect 18600 8128 18608 8192
rect 18672 8128 18688 8192
rect 18752 8128 18768 8192
rect 18832 8128 18848 8192
rect 18912 8128 18920 8192
rect 18600 7104 18920 8128
rect 18600 7040 18608 7104
rect 18672 7040 18688 7104
rect 18752 7040 18768 7104
rect 18832 7040 18848 7104
rect 18912 7040 18920 7104
rect 18600 6016 18920 7040
rect 18600 5952 18608 6016
rect 18672 5952 18688 6016
rect 18752 5952 18768 6016
rect 18832 5952 18848 6016
rect 18912 5952 18920 6016
rect 18600 4928 18920 5952
rect 18600 4864 18608 4928
rect 18672 4864 18688 4928
rect 18752 4864 18768 4928
rect 18832 4864 18848 4928
rect 18912 4864 18920 4928
rect 18600 3840 18920 4864
rect 18600 3776 18608 3840
rect 18672 3776 18688 3840
rect 18752 3776 18768 3840
rect 18832 3776 18848 3840
rect 18912 3776 18920 3840
rect 18600 2752 18920 3776
rect 18600 2688 18608 2752
rect 18672 2688 18688 2752
rect 18752 2688 18768 2752
rect 18832 2688 18848 2752
rect 18912 2688 18920 2752
rect 18600 1664 18920 2688
rect 18600 1600 18608 1664
rect 18672 1600 18688 1664
rect 18752 1600 18768 1664
rect 18832 1600 18848 1664
rect 18912 1600 18920 1664
rect 18600 576 18920 1600
rect 18600 512 18608 576
rect 18672 512 18688 576
rect 18752 512 18768 576
rect 18832 512 18848 576
rect 18912 512 18920 576
rect 18600 496 18920 512
use sky130_fd_sc_hd__diode_2  ANTENNA__234__A1 swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 16652 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__235__A1
timestamp 1673029049
transform -1 0 15640 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__236__A1
timestamp 1673029049
transform 1 0 12512 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__239__A1
timestamp 1673029049
transform 1 0 14720 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__240__A1
timestamp 1673029049
transform 1 0 13984 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__241__A1
timestamp 1673029049
transform -1 0 12512 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__242__A1
timestamp 1673029049
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__243__A1
timestamp 1673029049
transform -1 0 17296 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__244__A1
timestamp 1673029049
transform -1 0 18492 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__268__A1
timestamp 1673029049
transform 1 0 15088 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__268__A2
timestamp 1673029049
transform 1 0 14720 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__270__A2
timestamp 1673029049
transform -1 0 18032 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__328__A
timestamp 1673029049
transform 1 0 13524 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__330__A
timestamp 1673029049
transform 1 0 14168 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__330__B
timestamp 1673029049
transform 1 0 13984 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__331__B1
timestamp 1673029049
transform 1 0 12880 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__345__A1
timestamp 1673029049
transform 1 0 14260 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__345__A2
timestamp 1673029049
transform 1 0 14076 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__381__A_N
timestamp 1673029049
transform 1 0 16928 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__382__B
timestamp 1673029049
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__384__A
timestamp 1673029049
transform 1 0 16376 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__385__A
timestamp 1673029049
transform 1 0 14536 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__417__D
timestamp 1673029049
transform 1 0 7084 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__417__RESET_B
timestamp 1673029049
transform 1 0 5060 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__425__RESET_B
timestamp 1673029049
transform 1 0 7636 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__426__RESET_B
timestamp 1673029049
transform 1 0 2760 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__427__SET_B
timestamp 1673029049
transform 1 0 3496 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__428__RESET_B
timestamp 1673029049
transform 1 0 4048 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__429__SET_B
timestamp 1673029049
transform 1 0 4968 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__430__RESET_B
timestamp 1673029049
transform 1 0 2576 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__432__RESET_B
timestamp 1673029049
transform 1 0 2760 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__433__RESET_B
timestamp 1673029049
transform 1 0 8556 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__434__SET_B
timestamp 1673029049
transform 1 0 6164 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__435__RESET_B
timestamp 1673029049
transform 1 0 8924 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__439__D
timestamp 1673029049
transform -1 0 10120 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__440__SET_B
timestamp 1673029049
transform 1 0 7084 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__441__RESET_B
timestamp 1673029049
transform 1 0 7360 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__442__RESET_B
timestamp 1673029049
transform 1 0 7728 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__444__RESET_B
timestamp 1673029049
transform 1 0 8280 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__447__D
timestamp 1673029049
transform 1 0 17112 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__448__D
timestamp 1673029049
transform 1 0 14168 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__461__SET_B
timestamp 1673029049
transform 1 0 7084 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_ext_clk_A
timestamp 1673029049
transform -1 0 2944 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_pll_clk90_A
timestamp 1673029049
transform 1 0 15548 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_pll_clk_A
timestamp 1673029049
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout26_A
timestamp 1673029049
transform 1 0 2852 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout27_A
timestamp 1673029049
transform -1 0 1288 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout28_A
timestamp 1673029049
transform 1 0 10672 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout29_A
timestamp 1673029049
transform -1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1673029049
transform 1 0 18308 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1673029049
transform 1 0 18308 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1673029049
transform -1 0 1196 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1673029049
transform -1 0 920 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1673029049
transform -1 0 18492 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1673029049
transform -1 0 18032 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1673029049
transform -1 0 18492 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1673029049
transform -1 0 18032 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1673029049
transform -1 0 18032 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1673029049
transform -1 0 18032 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3 swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 460 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11 swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 1196 0 1 544
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14 swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 1472 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27
timestamp 1673029049
transform 1 0 2668 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40
timestamp 1673029049
transform 1 0 3864 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53
timestamp 1673029049
transform 1 0 5060 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59 swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 5612 0 1 544
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66
timestamp 1673029049
transform 1 0 6256 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79
timestamp 1673029049
transform 1 0 7452 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92
timestamp 1673029049
transform 1 0 8648 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105
timestamp 1673029049
transform 1 0 9844 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_118 swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 11040 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_125 swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 11684 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_129 swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 12052 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_131
timestamp 1673029049
transform 1 0 12236 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_144
timestamp 1673029049
transform 1 0 13432 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_157
timestamp 1673029049
transform 1 0 14628 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_170
timestamp 1673029049
transform 1 0 15824 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_183
timestamp 1673029049
transform 1 0 17020 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_186
timestamp 1673029049
transform 1 0 17296 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_190
timestamp 1673029049
transform 1 0 17664 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_194
timestamp 1673029049
transform 1 0 18032 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_196
timestamp 1673029049
transform 1 0 18216 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_199
timestamp 1673029049
transform 1 0 18492 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1673029049
transform 1 0 460 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_15
timestamp 1673029049
transform 1 0 1564 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_23
timestamp 1673029049
transform 1 0 2300 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_27
timestamp 1673029049
transform 1 0 2668 0 -1 1632
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_36
timestamp 1673029049
transform 1 0 3496 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_48
timestamp 1673029049
transform 1 0 4600 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_53
timestamp 1673029049
transform 1 0 5060 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_57
timestamp 1673029049
transform 1 0 5428 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_63
timestamp 1673029049
transform 1 0 5980 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_69
timestamp 1673029049
transform 1 0 6532 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_77
timestamp 1673029049
transform 1 0 7268 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_79
timestamp 1673029049
transform 1 0 7452 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_87
timestamp 1673029049
transform 1 0 8188 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_95
timestamp 1673029049
transform 1 0 8924 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_103
timestamp 1673029049
transform 1 0 9660 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_105
timestamp 1673029049
transform 1 0 9844 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_110
timestamp 1673029049
transform 1 0 10304 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_114
timestamp 1673029049
transform 1 0 10672 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_119
timestamp 1673029049
transform 1 0 11132 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_126
timestamp 1673029049
transform 1 0 11776 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_131
timestamp 1673029049
transform 1 0 12236 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_134
timestamp 1673029049
transform 1 0 12512 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_140
timestamp 1673029049
transform 1 0 13064 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_148
timestamp 1673029049
transform 1 0 13800 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_157
timestamp 1673029049
transform 1 0 14628 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_165
timestamp 1673029049
transform 1 0 15364 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_178
timestamp 1673029049
transform 1 0 16560 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_183
timestamp 1673029049
transform 1 0 17020 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_193
timestamp 1673029049
transform 1 0 17940 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_198
timestamp 1673029049
transform 1 0 18400 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_3
timestamp 1673029049
transform 1 0 460 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_11
timestamp 1673029049
transform 1 0 1196 0 1 1632
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_14
timestamp 1673029049
transform 1 0 1472 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_26
timestamp 1673029049
transform 1 0 2576 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_38
timestamp 1673029049
transform 1 0 3680 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_40
timestamp 1673029049
transform 1 0 3864 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_51
timestamp 1673029049
transform 1 0 4876 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_58
timestamp 1673029049
transform 1 0 5520 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_64
timestamp 1673029049
transform 1 0 6072 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_66
timestamp 1673029049
transform 1 0 6256 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_76
timestamp 1673029049
transform 1 0 7176 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_80
timestamp 1673029049
transform 1 0 7544 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_90
timestamp 1673029049
transform 1 0 8464 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_92
timestamp 1673029049
transform 1 0 8648 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_101
timestamp 1673029049
transform 1 0 9476 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_108
timestamp 1673029049
transform 1 0 10120 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_114
timestamp 1673029049
transform 1 0 10672 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_118
timestamp 1673029049
transform 1 0 11040 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_122
timestamp 1673029049
transform 1 0 11408 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_132
timestamp 1673029049
transform 1 0 12328 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_142
timestamp 1673029049
transform 1 0 13248 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_144
timestamp 1673029049
transform 1 0 13432 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_156
timestamp 1673029049
transform 1 0 14536 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_160
timestamp 1673029049
transform 1 0 14904 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_168
timestamp 1673029049
transform 1 0 15640 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_170
timestamp 1673029049
transform 1 0 15824 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_180
timestamp 1673029049
transform 1 0 16744 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_191
timestamp 1673029049
transform 1 0 17756 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_196
timestamp 1673029049
transform 1 0 18216 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_199
timestamp 1673029049
transform 1 0 18492 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3
timestamp 1673029049
transform 1 0 460 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_18
timestamp 1673029049
transform 1 0 1840 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_24
timestamp 1673029049
transform 1 0 2392 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_27
timestamp 1673029049
transform 1 0 2668 0 -1 2720
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_38
timestamp 1673029049
transform 1 0 3680 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_50
timestamp 1673029049
transform 1 0 4784 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_53
timestamp 1673029049
transform 1 0 5060 0 -1 2720
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_65
timestamp 1673029049
transform 1 0 6164 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_77
timestamp 1673029049
transform 1 0 7268 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_79
timestamp 1673029049
transform 1 0 7452 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_96
timestamp 1673029049
transform 1 0 9016 0 -1 2720
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_105
timestamp 1673029049
transform 1 0 9844 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_117
timestamp 1673029049
transform 1 0 10948 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_129
timestamp 1673029049
transform 1 0 12052 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_131
timestamp 1673029049
transform 1 0 12236 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_134
timestamp 1673029049
transform 1 0 12512 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_146
timestamp 1673029049
transform 1 0 13616 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_150
timestamp 1673029049
transform 1 0 13984 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_153
timestamp 1673029049
transform 1 0 14260 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_157
timestamp 1673029049
transform 1 0 14628 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_167
timestamp 1673029049
transform 1 0 15548 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_179
timestamp 1673029049
transform 1 0 16652 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_183
timestamp 1673029049
transform 1 0 17020 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_188
timestamp 1673029049
transform 1 0 17480 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_199
timestamp 1673029049
transform 1 0 18492 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_3
timestamp 1673029049
transform 1 0 460 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_11
timestamp 1673029049
transform 1 0 1196 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_14
timestamp 1673029049
transform 1 0 1472 0 1 2720
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_26
timestamp 1673029049
transform 1 0 2576 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_38
timestamp 1673029049
transform 1 0 3680 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_40
timestamp 1673029049
transform 1 0 3864 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_52
timestamp 1673029049
transform 1 0 4968 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_56
timestamp 1673029049
transform 1 0 5336 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_64
timestamp 1673029049
transform 1 0 6072 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_66
timestamp 1673029049
transform 1 0 6256 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_83
timestamp 1673029049
transform 1 0 7820 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_92
timestamp 1673029049
transform 1 0 8648 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_100
timestamp 1673029049
transform 1 0 9384 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_110
timestamp 1673029049
transform 1 0 10304 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_116
timestamp 1673029049
transform 1 0 10856 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_118
timestamp 1673029049
transform 1 0 11040 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_129
timestamp 1673029049
transform 1 0 12052 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_142
timestamp 1673029049
transform 1 0 13248 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_144
timestamp 1673029049
transform 1 0 13432 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_148
timestamp 1673029049
transform 1 0 13800 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_152
timestamp 1673029049
transform 1 0 14168 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_167
timestamp 1673029049
transform 1 0 15548 0 1 2720
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_170
timestamp 1673029049
transform 1 0 15824 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_182
timestamp 1673029049
transform 1 0 16928 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_194
timestamp 1673029049
transform 1 0 18032 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_196
timestamp 1673029049
transform 1 0 18216 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_5_3
timestamp 1673029049
transform 1 0 460 0 -1 3808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_9
timestamp 1673029049
transform 1 0 1012 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_21
timestamp 1673029049
transform 1 0 2116 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_25
timestamp 1673029049
transform 1 0 2484 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1673029049
transform 1 0 2668 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_39
timestamp 1673029049
transform 1 0 3772 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_48
timestamp 1673029049
transform 1 0 4600 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_53
timestamp 1673029049
transform 1 0 5060 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_63
timestamp 1673029049
transform 1 0 5980 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_75
timestamp 1673029049
transform 1 0 7084 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_79
timestamp 1673029049
transform 1 0 7452 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_89
timestamp 1673029049
transform 1 0 8372 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_101
timestamp 1673029049
transform 1 0 9476 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_105
timestamp 1673029049
transform 1 0 9844 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_115
timestamp 1673029049
transform 1 0 10764 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_123
timestamp 1673029049
transform 1 0 11500 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_129
timestamp 1673029049
transform 1 0 12052 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_131
timestamp 1673029049
transform 1 0 12236 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_143
timestamp 1673029049
transform 1 0 13340 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_151
timestamp 1673029049
transform 1 0 14076 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_155
timestamp 1673029049
transform 1 0 14444 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_157
timestamp 1673029049
transform 1 0 14628 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_167
timestamp 1673029049
transform 1 0 15548 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_171
timestamp 1673029049
transform 1 0 15916 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_181
timestamp 1673029049
transform 1 0 16836 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_183
timestamp 1673029049
transform 1 0 17020 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_190
timestamp 1673029049
transform 1 0 17664 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_194
timestamp 1673029049
transform 1 0 18032 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_199
timestamp 1673029049
transform 1 0 18492 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_3
timestamp 1673029049
transform 1 0 460 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_10
timestamp 1673029049
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_14
timestamp 1673029049
transform 1 0 1472 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_21
timestamp 1673029049
transform 1 0 2116 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_33
timestamp 1673029049
transform 1 0 3220 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_37
timestamp 1673029049
transform 1 0 3588 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_40
timestamp 1673029049
transform 1 0 3864 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_58
timestamp 1673029049
transform 1 0 5520 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_64
timestamp 1673029049
transform 1 0 6072 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_66
timestamp 1673029049
transform 1 0 6256 0 1 3808
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_76
timestamp 1673029049
transform 1 0 7176 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_88
timestamp 1673029049
transform 1 0 8280 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_92
timestamp 1673029049
transform 1 0 8648 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1673029049
transform 1 0 9108 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_109
timestamp 1673029049
transform 1 0 10212 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_118
timestamp 1673029049
transform 1 0 11040 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_126
timestamp 1673029049
transform 1 0 11776 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_140
timestamp 1673029049
transform 1 0 13064 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_144
timestamp 1673029049
transform 1 0 13432 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_150
timestamp 1673029049
transform 1 0 13984 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_155
timestamp 1673029049
transform 1 0 14444 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_159
timestamp 1673029049
transform 1 0 14812 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_167
timestamp 1673029049
transform 1 0 15548 0 1 3808
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_170
timestamp 1673029049
transform 1 0 15824 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_187
timestamp 1673029049
transform 1 0 17388 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_194
timestamp 1673029049
transform 1 0 18032 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_196
timestamp 1673029049
transform 1 0 18216 0 1 3808
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1673029049
transform 1 0 460 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_15
timestamp 1673029049
transform 1 0 1564 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_21
timestamp 1673029049
transform 1 0 2116 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_25
timestamp 1673029049
transform 1 0 2484 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_27
timestamp 1673029049
transform 1 0 2668 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_35
timestamp 1673029049
transform 1 0 3404 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_42
timestamp 1673029049
transform 1 0 4048 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_46
timestamp 1673029049
transform 1 0 4416 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_51
timestamp 1673029049
transform 1 0 4876 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_53
timestamp 1673029049
transform 1 0 5060 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_65
timestamp 1673029049
transform 1 0 6164 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_77
timestamp 1673029049
transform 1 0 7268 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_79
timestamp 1673029049
transform 1 0 7452 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_85
timestamp 1673029049
transform 1 0 8004 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_91
timestamp 1673029049
transform 1 0 8556 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_101
timestamp 1673029049
transform 1 0 9476 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_105
timestamp 1673029049
transform 1 0 9844 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_129
timestamp 1673029049
transform 1 0 12052 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_131
timestamp 1673029049
transform 1 0 12236 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_139
timestamp 1673029049
transform 1 0 12972 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_151
timestamp 1673029049
transform 1 0 14076 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_155
timestamp 1673029049
transform 1 0 14444 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_157
timestamp 1673029049
transform 1 0 14628 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_160
timestamp 1673029049
transform 1 0 14904 0 -1 4896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_164
timestamp 1673029049
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_176
timestamp 1673029049
transform 1 0 16376 0 -1 4896
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_183
timestamp 1673029049
transform 1 0 17020 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_195
timestamp 1673029049
transform 1 0 18124 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_199
timestamp 1673029049
transform 1 0 18492 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_3
timestamp 1673029049
transform 1 0 460 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_11
timestamp 1673029049
transform 1 0 1196 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_14
timestamp 1673029049
transform 1 0 1472 0 1 4896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_25
timestamp 1673029049
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_37
timestamp 1673029049
transform 1 0 3588 0 1 4896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_40
timestamp 1673029049
transform 1 0 3864 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_52
timestamp 1673029049
transform 1 0 4968 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_64
timestamp 1673029049
transform 1 0 6072 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_66
timestamp 1673029049
transform 1 0 6256 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_77
timestamp 1673029049
transform 1 0 7268 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_83
timestamp 1673029049
transform 1 0 7820 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_88
timestamp 1673029049
transform 1 0 8280 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_92
timestamp 1673029049
transform 1 0 8648 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_113
timestamp 1673029049
transform 1 0 10580 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_118
timestamp 1673029049
transform 1 0 11040 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_141
timestamp 1673029049
transform 1 0 13156 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_144
timestamp 1673029049
transform 1 0 13432 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_168
timestamp 1673029049
transform 1 0 15640 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_170
timestamp 1673029049
transform 1 0 15824 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_192
timestamp 1673029049
transform 1 0 17848 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_196
timestamp 1673029049
transform 1 0 18216 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3
timestamp 1673029049
transform 1 0 460 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_24
timestamp 1673029049
transform 1 0 2392 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_27
timestamp 1673029049
transform 1 0 2668 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_30
timestamp 1673029049
transform 1 0 2944 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_38
timestamp 1673029049
transform 1 0 3680 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_44
timestamp 1673029049
transform 1 0 4232 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_51
timestamp 1673029049
transform 1 0 4876 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_53
timestamp 1673029049
transform 1 0 5060 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_61
timestamp 1673029049
transform 1 0 5796 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_67
timestamp 1673029049
transform 1 0 6348 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_75
timestamp 1673029049
transform 1 0 7084 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_79
timestamp 1673029049
transform 1 0 7452 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_85
timestamp 1673029049
transform 1 0 8004 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_89
timestamp 1673029049
transform 1 0 8372 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_93
timestamp 1673029049
transform 1 0 8740 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_97
timestamp 1673029049
transform 1 0 9108 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_103
timestamp 1673029049
transform 1 0 9660 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_105
timestamp 1673029049
transform 1 0 9844 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_117
timestamp 1673029049
transform 1 0 10948 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_129
timestamp 1673029049
transform 1 0 12052 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_131
timestamp 1673029049
transform 1 0 12236 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_143
timestamp 1673029049
transform 1 0 13340 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_155
timestamp 1673029049
transform 1 0 14444 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_157
timestamp 1673029049
transform 1 0 14628 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_181
timestamp 1673029049
transform 1 0 16836 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_183
timestamp 1673029049
transform 1 0 17020 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_191
timestamp 1673029049
transform 1 0 17756 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_199
timestamp 1673029049
transform 1 0 18492 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_3
timestamp 1673029049
transform 1 0 460 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_11
timestamp 1673029049
transform 1 0 1196 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_14
timestamp 1673029049
transform 1 0 1472 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_36
timestamp 1673029049
transform 1 0 3496 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_40
timestamp 1673029049
transform 1 0 3864 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_64
timestamp 1673029049
transform 1 0 6072 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_66
timestamp 1673029049
transform 1 0 6256 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_88
timestamp 1673029049
transform 1 0 8280 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_92
timestamp 1673029049
transform 1 0 8648 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_116
timestamp 1673029049
transform 1 0 10856 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_118
timestamp 1673029049
transform 1 0 11040 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_130
timestamp 1673029049
transform 1 0 12144 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_141
timestamp 1673029049
transform 1 0 13156 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_144
timestamp 1673029049
transform 1 0 13432 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_147
timestamp 1673029049
transform 1 0 13708 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_155
timestamp 1673029049
transform 1 0 14444 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_158
timestamp 1673029049
transform 1 0 14720 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_166
timestamp 1673029049
transform 1 0 15456 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_170
timestamp 1673029049
transform 1 0 15824 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_192
timestamp 1673029049
transform 1 0 17848 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_196
timestamp 1673029049
transform 1 0 18216 0 1 5984
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1673029049
transform 1 0 460 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_15
timestamp 1673029049
transform 1 0 1564 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_21
timestamp 1673029049
transform 1 0 2116 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_25
timestamp 1673029049
transform 1 0 2484 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1673029049
transform 1 0 2668 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1673029049
transform 1 0 3772 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_51
timestamp 1673029049
transform 1 0 4876 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_53
timestamp 1673029049
transform 1 0 5060 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_61
timestamp 1673029049
transform 1 0 5796 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_73
timestamp 1673029049
transform 1 0 6900 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_77
timestamp 1673029049
transform 1 0 7268 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_79
timestamp 1673029049
transform 1 0 7452 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_91
timestamp 1673029049
transform 1 0 8556 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_103
timestamp 1673029049
transform 1 0 9660 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_105
timestamp 1673029049
transform 1 0 9844 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_128
timestamp 1673029049
transform 1 0 11960 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_131
timestamp 1673029049
transform 1 0 12236 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_150
timestamp 1673029049
transform 1 0 13984 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_154
timestamp 1673029049
transform 1 0 14352 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_157
timestamp 1673029049
transform 1 0 14628 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_163
timestamp 1673029049
transform 1 0 15180 0 -1 7072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1673029049
transform 1 0 15732 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_181
timestamp 1673029049
transform 1 0 16836 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_183
timestamp 1673029049
transform 1 0 17020 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_191
timestamp 1673029049
transform 1 0 17756 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_194
timestamp 1673029049
transform 1 0 18032 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_199
timestamp 1673029049
transform 1 0 18492 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_3
timestamp 1673029049
transform 1 0 460 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_11
timestamp 1673029049
transform 1 0 1196 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_14
timestamp 1673029049
transform 1 0 1472 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_24
timestamp 1673029049
transform 1 0 2392 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_28
timestamp 1673029049
transform 1 0 2760 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_38
timestamp 1673029049
transform 1 0 3680 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_40
timestamp 1673029049
transform 1 0 3864 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_50
timestamp 1673029049
transform 1 0 4784 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_54
timestamp 1673029049
transform 1 0 5152 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_62
timestamp 1673029049
transform 1 0 5888 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_66
timestamp 1673029049
transform 1 0 6256 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_74
timestamp 1673029049
transform 1 0 6992 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_86
timestamp 1673029049
transform 1 0 8096 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_90
timestamp 1673029049
transform 1 0 8464 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_92
timestamp 1673029049
transform 1 0 8648 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_100
timestamp 1673029049
transform 1 0 9384 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_108
timestamp 1673029049
transform 1 0 10120 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_112
timestamp 1673029049
transform 1 0 10488 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_116
timestamp 1673029049
transform 1 0 10856 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_118
timestamp 1673029049
transform 1 0 11040 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_128
timestamp 1673029049
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_139
timestamp 1673029049
transform 1 0 12972 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_144
timestamp 1673029049
transform 1 0 13432 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_168
timestamp 1673029049
transform 1 0 15640 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_170
timestamp 1673029049
transform 1 0 15824 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_174
timestamp 1673029049
transform 1 0 16192 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_178
timestamp 1673029049
transform 1 0 16560 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_184
timestamp 1673029049
transform 1 0 17112 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_191
timestamp 1673029049
transform 1 0 17756 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_196
timestamp 1673029049
transform 1 0 18216 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1673029049
transform 1 0 460 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_25
timestamp 1673029049
transform 1 0 2484 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_27
timestamp 1673029049
transform 1 0 2668 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_48
timestamp 1673029049
transform 1 0 4600 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_53
timestamp 1673029049
transform 1 0 5060 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_75
timestamp 1673029049
transform 1 0 7084 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_79
timestamp 1673029049
transform 1 0 7452 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_89
timestamp 1673029049
transform 1 0 8372 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_97
timestamp 1673029049
transform 1 0 9108 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_103
timestamp 1673029049
transform 1 0 9660 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_105
timestamp 1673029049
transform 1 0 9844 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_112
timestamp 1673029049
transform 1 0 10488 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_122
timestamp 1673029049
transform 1 0 11408 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_131
timestamp 1673029049
transform 1 0 12236 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_155
timestamp 1673029049
transform 1 0 14444 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_157
timestamp 1673029049
transform 1 0 14628 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_165
timestamp 1673029049
transform 1 0 15364 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_173
timestamp 1673029049
transform 1 0 16100 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_177
timestamp 1673029049
transform 1 0 16468 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_181
timestamp 1673029049
transform 1 0 16836 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_183
timestamp 1673029049
transform 1 0 17020 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_192
timestamp 1673029049
transform 1 0 17848 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_3
timestamp 1673029049
transform 1 0 460 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_11
timestamp 1673029049
transform 1 0 1196 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_14
timestamp 1673029049
transform 1 0 1472 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_22
timestamp 1673029049
transform 1 0 2208 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_31
timestamp 1673029049
transform 1 0 3036 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_36
timestamp 1673029049
transform 1 0 3496 0 1 8160
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_40
timestamp 1673029049
transform 1 0 3864 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_52
timestamp 1673029049
transform 1 0 4968 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_60
timestamp 1673029049
transform 1 0 5704 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_64
timestamp 1673029049
transform 1 0 6072 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_66
timestamp 1673029049
transform 1 0 6256 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_75
timestamp 1673029049
transform 1 0 7084 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1673029049
transform 1 0 7820 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_88
timestamp 1673029049
transform 1 0 8280 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_92
timestamp 1673029049
transform 1 0 8648 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_99
timestamp 1673029049
transform 1 0 9292 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_111
timestamp 1673029049
transform 1 0 10396 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_116
timestamp 1673029049
transform 1 0 10856 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_118
timestamp 1673029049
transform 1 0 11040 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_128
timestamp 1673029049
transform 1 0 11960 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_140
timestamp 1673029049
transform 1 0 13064 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_144
timestamp 1673029049
transform 1 0 13432 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_148
timestamp 1673029049
transform 1 0 13800 0 1 8160
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_152
timestamp 1673029049
transform 1 0 14168 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_164
timestamp 1673029049
transform 1 0 15272 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_168
timestamp 1673029049
transform 1 0 15640 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_170
timestamp 1673029049
transform 1 0 15824 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_194
timestamp 1673029049
transform 1 0 18032 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_196
timestamp 1673029049
transform 1 0 18216 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_3
timestamp 1673029049
transform 1 0 460 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_24
timestamp 1673029049
transform 1 0 2392 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_27
timestamp 1673029049
transform 1 0 2668 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_30
timestamp 1673029049
transform 1 0 2944 0 -1 9248
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_38
timestamp 1673029049
transform 1 0 3680 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_50
timestamp 1673029049
transform 1 0 4784 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_53
timestamp 1673029049
transform 1 0 5060 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_70
timestamp 1673029049
transform 1 0 6624 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_74
timestamp 1673029049
transform 1 0 6992 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_77
timestamp 1673029049
transform 1 0 7268 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_79
timestamp 1673029049
transform 1 0 7452 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_101
timestamp 1673029049
transform 1 0 9476 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_105
timestamp 1673029049
transform 1 0 9844 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_127
timestamp 1673029049
transform 1 0 11868 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_131
timestamp 1673029049
transform 1 0 12236 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_144
timestamp 1673029049
transform 1 0 13432 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_150
timestamp 1673029049
transform 1 0 13984 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_154
timestamp 1673029049
transform 1 0 14352 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_157
timestamp 1673029049
transform 1 0 14628 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_179
timestamp 1673029049
transform 1 0 16652 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_183
timestamp 1673029049
transform 1 0 17020 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_191
timestamp 1673029049
transform 1 0 17756 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_194
timestamp 1673029049
transform 1 0 18032 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_199
timestamp 1673029049
transform 1 0 18492 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_3
timestamp 1673029049
transform 1 0 460 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_11
timestamp 1673029049
transform 1 0 1196 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_14
timestamp 1673029049
transform 1 0 1472 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_24
timestamp 1673029049
transform 1 0 2392 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_28
timestamp 1673029049
transform 1 0 2760 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_34
timestamp 1673029049
transform 1 0 3312 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_38
timestamp 1673029049
transform 1 0 3680 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_40
timestamp 1673029049
transform 1 0 3864 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_50
timestamp 1673029049
transform 1 0 4784 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_62
timestamp 1673029049
transform 1 0 5888 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_66
timestamp 1673029049
transform 1 0 6256 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_77
timestamp 1673029049
transform 1 0 7268 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_83
timestamp 1673029049
transform 1 0 7820 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_92
timestamp 1673029049
transform 1 0 8648 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_97
timestamp 1673029049
transform 1 0 9108 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_105
timestamp 1673029049
transform 1 0 9844 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_112
timestamp 1673029049
transform 1 0 10488 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_116
timestamp 1673029049
transform 1 0 10856 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_118
timestamp 1673029049
transform 1 0 11040 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_133
timestamp 1673029049
transform 1 0 12420 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_137
timestamp 1673029049
transform 1 0 12788 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_140
timestamp 1673029049
transform 1 0 13064 0 1 9248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_144
timestamp 1673029049
transform 1 0 13432 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_156
timestamp 1673029049
transform 1 0 14536 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_160
timestamp 1673029049
transform 1 0 14904 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_165
timestamp 1673029049
transform 1 0 15364 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_170
timestamp 1673029049
transform 1 0 15824 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_175
timestamp 1673029049
transform 1 0 16284 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_194
timestamp 1673029049
transform 1 0 18032 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_196
timestamp 1673029049
transform 1 0 18216 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_3
timestamp 1673029049
transform 1 0 460 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_7
timestamp 1673029049
transform 1 0 828 0 -1 10336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_11
timestamp 1673029049
transform 1 0 1196 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_23
timestamp 1673029049
transform 1 0 2300 0 -1 10336
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1673029049
transform 1 0 2668 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_43
timestamp 1673029049
transform 1 0 4140 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_51
timestamp 1673029049
transform 1 0 4876 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_53
timestamp 1673029049
transform 1 0 5060 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_57
timestamp 1673029049
transform 1 0 5428 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_64
timestamp 1673029049
transform 1 0 6072 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_70
timestamp 1673029049
transform 1 0 6624 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_77
timestamp 1673029049
transform 1 0 7268 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_79
timestamp 1673029049
transform 1 0 7452 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_103
timestamp 1673029049
transform 1 0 9660 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_105
timestamp 1673029049
transform 1 0 9844 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_113
timestamp 1673029049
transform 1 0 10580 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_122
timestamp 1673029049
transform 1 0 11408 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_129
timestamp 1673029049
transform 1 0 12052 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_131
timestamp 1673029049
transform 1 0 12236 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_138
timestamp 1673029049
transform 1 0 12880 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_146
timestamp 1673029049
transform 1 0 13616 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_154
timestamp 1673029049
transform 1 0 14352 0 -1 10336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_157
timestamp 1673029049
transform 1 0 14628 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1673029049
transform 1 0 15732 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_181
timestamp 1673029049
transform 1 0 16836 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_183
timestamp 1673029049
transform 1 0 17020 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_191
timestamp 1673029049
transform 1 0 17756 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_199
timestamp 1673029049
transform 1 0 18492 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_3
timestamp 1673029049
transform 1 0 460 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_11
timestamp 1673029049
transform 1 0 1196 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_14
timestamp 1673029049
transform 1 0 1472 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_25
timestamp 1673029049
transform 1 0 2484 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_36
timestamp 1673029049
transform 1 0 3496 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_40
timestamp 1673029049
transform 1 0 3864 0 1 10336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_48
timestamp 1673029049
transform 1 0 4600 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_60
timestamp 1673029049
transform 1 0 5704 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_64
timestamp 1673029049
transform 1 0 6072 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_66
timestamp 1673029049
transform 1 0 6256 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_74
timestamp 1673029049
transform 1 0 6992 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_87
timestamp 1673029049
transform 1 0 8188 0 1 10336
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_92
timestamp 1673029049
transform 1 0 8648 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_104
timestamp 1673029049
transform 1 0 9752 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_116
timestamp 1673029049
transform 1 0 10856 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_118
timestamp 1673029049
transform 1 0 11040 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_128
timestamp 1673029049
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_139
timestamp 1673029049
transform 1 0 12972 0 1 10336
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_144
timestamp 1673029049
transform 1 0 13432 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_156
timestamp 1673029049
transform 1 0 14536 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_164
timestamp 1673029049
transform 1 0 15272 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_168
timestamp 1673029049
transform 1 0 15640 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_170
timestamp 1673029049
transform 1 0 15824 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_184
timestamp 1673029049
transform 1 0 17112 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_188
timestamp 1673029049
transform 1 0 17480 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_191
timestamp 1673029049
transform 1 0 17756 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_196
timestamp 1673029049
transform 1 0 18216 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_3
timestamp 1673029049
transform 1 0 460 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_11
timestamp 1673029049
transform 1 0 1196 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_21
timestamp 1673029049
transform 1 0 2116 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_25
timestamp 1673029049
transform 1 0 2484 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1673029049
transform 1 0 2668 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_42
timestamp 1673029049
transform 1 0 4048 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_50
timestamp 1673029049
transform 1 0 4784 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_53
timestamp 1673029049
transform 1 0 5060 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_59
timestamp 1673029049
transform 1 0 5612 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_71
timestamp 1673029049
transform 1 0 6716 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_77
timestamp 1673029049
transform 1 0 7268 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_79
timestamp 1673029049
transform 1 0 7452 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_103
timestamp 1673029049
transform 1 0 9660 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_105
timestamp 1673029049
transform 1 0 9844 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_126
timestamp 1673029049
transform 1 0 11776 0 -1 11424
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_131
timestamp 1673029049
transform 1 0 12236 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_143
timestamp 1673029049
transform 1 0 13340 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_149
timestamp 1673029049
transform 1 0 13892 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_153
timestamp 1673029049
transform 1 0 14260 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_157
timestamp 1673029049
transform 1 0 14628 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_179
timestamp 1673029049
transform 1 0 16652 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_183
timestamp 1673029049
transform 1 0 17020 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_189
timestamp 1673029049
transform 1 0 17572 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_196
timestamp 1673029049
transform 1 0 18216 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_3
timestamp 1673029049
transform 1 0 460 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_11
timestamp 1673029049
transform 1 0 1196 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_14
timestamp 1673029049
transform 1 0 1472 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_36
timestamp 1673029049
transform 1 0 3496 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_40
timestamp 1673029049
transform 1 0 3864 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_64
timestamp 1673029049
transform 1 0 6072 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_66
timestamp 1673029049
transform 1 0 6256 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_69
timestamp 1673029049
transform 1 0 6532 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_83
timestamp 1673029049
transform 1 0 7820 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_88
timestamp 1673029049
transform 1 0 8280 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_92
timestamp 1673029049
transform 1 0 8648 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_114
timestamp 1673029049
transform 1 0 10672 0 1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_118
timestamp 1673029049
transform 1 0 11040 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_130
timestamp 1673029049
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1673029049
transform 1 0 13156 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_144
timestamp 1673029049
transform 1 0 13432 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_168
timestamp 1673029049
transform 1 0 15640 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_170
timestamp 1673029049
transform 1 0 15824 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_176
timestamp 1673029049
transform 1 0 16376 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_194
timestamp 1673029049
transform 1 0 18032 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_196
timestamp 1673029049
transform 1 0 18216 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_199
timestamp 1673029049
transform 1 0 18492 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1673029049
transform 1 0 460 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_15
timestamp 1673029049
transform 1 0 1564 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_21
timestamp 1673029049
transform 1 0 2116 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_25
timestamp 1673029049
transform 1 0 2484 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_27
timestamp 1673029049
transform 1 0 2668 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_33
timestamp 1673029049
transform 1 0 3220 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_50
timestamp 1673029049
transform 1 0 4784 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_53
timestamp 1673029049
transform 1 0 5060 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_60
timestamp 1673029049
transform 1 0 5704 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_66
timestamp 1673029049
transform 1 0 6256 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_74
timestamp 1673029049
transform 1 0 6992 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_77
timestamp 1673029049
transform 1 0 7268 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_79
timestamp 1673029049
transform 1 0 7452 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_103
timestamp 1673029049
transform 1 0 9660 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_105
timestamp 1673029049
transform 1 0 9844 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_117
timestamp 1673029049
transform 1 0 10948 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_123
timestamp 1673029049
transform 1 0 11500 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_129
timestamp 1673029049
transform 1 0 12052 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_131
timestamp 1673029049
transform 1 0 12236 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_137
timestamp 1673029049
transform 1 0 12788 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_145
timestamp 1673029049
transform 1 0 13524 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_154
timestamp 1673029049
transform 1 0 14352 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_157
timestamp 1673029049
transform 1 0 14628 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_165
timestamp 1673029049
transform 1 0 15364 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1673029049
transform 1 0 15732 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_176
timestamp 1673029049
transform 1 0 16376 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_181
timestamp 1673029049
transform 1 0 16836 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_183
timestamp 1673029049
transform 1 0 17020 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_186
timestamp 1673029049
transform 1 0 17296 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_191
timestamp 1673029049
transform 1 0 17756 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_195
timestamp 1673029049
transform 1 0 18124 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_199
timestamp 1673029049
transform 1 0 18492 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_3
timestamp 1673029049
transform 1 0 460 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_11
timestamp 1673029049
transform 1 0 1196 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_14
timestamp 1673029049
transform 1 0 1472 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_24
timestamp 1673029049
transform 1 0 2392 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_37
timestamp 1673029049
transform 1 0 3588 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_40
timestamp 1673029049
transform 1 0 3864 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_22_62
timestamp 1673029049
transform 1 0 5888 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_66
timestamp 1673029049
transform 1 0 6256 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_74
timestamp 1673029049
transform 1 0 6992 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_77
timestamp 1673029049
transform 1 0 7268 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_88
timestamp 1673029049
transform 1 0 8280 0 1 12512
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_92
timestamp 1673029049
transform 1 0 8648 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_104
timestamp 1673029049
transform 1 0 9752 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_116
timestamp 1673029049
transform 1 0 10856 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_118
timestamp 1673029049
transform 1 0 11040 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_123
timestamp 1673029049
transform 1 0 11500 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_131
timestamp 1673029049
transform 1 0 12236 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_138
timestamp 1673029049
transform 1 0 12880 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_142
timestamp 1673029049
transform 1 0 13248 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_144
timestamp 1673029049
transform 1 0 13432 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_148
timestamp 1673029049
transform 1 0 13800 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_166
timestamp 1673029049
transform 1 0 15456 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_170
timestamp 1673029049
transform 1 0 15824 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_181
timestamp 1673029049
transform 1 0 16836 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_190
timestamp 1673029049
transform 1 0 17664 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_194
timestamp 1673029049
transform 1 0 18032 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_196
timestamp 1673029049
transform 1 0 18216 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_3
timestamp 1673029049
transform 1 0 460 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_25
timestamp 1673029049
transform 1 0 2484 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_27
timestamp 1673029049
transform 1 0 2668 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_48
timestamp 1673029049
transform 1 0 4600 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_53
timestamp 1673029049
transform 1 0 5060 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_75
timestamp 1673029049
transform 1 0 7084 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_79
timestamp 1673029049
transform 1 0 7452 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_100
timestamp 1673029049
transform 1 0 9384 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_105
timestamp 1673029049
transform 1 0 9844 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_129
timestamp 1673029049
transform 1 0 12052 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_131
timestamp 1673029049
transform 1 0 12236 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_155
timestamp 1673029049
transform 1 0 14444 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_157
timestamp 1673029049
transform 1 0 14628 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_181
timestamp 1673029049
transform 1 0 16836 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_183
timestamp 1673029049
transform 1 0 17020 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_195
timestamp 1673029049
transform 1 0 18124 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_199
timestamp 1673029049
transform 1 0 18492 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_3
timestamp 1673029049
transform 1 0 460 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_11
timestamp 1673029049
transform 1 0 1196 0 1 13600
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_14
timestamp 1673029049
transform 1 0 1472 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_26
timestamp 1673029049
transform 1 0 2576 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_24_33
timestamp 1673029049
transform 1 0 3220 0 1 13600
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_40
timestamp 1673029049
transform 1 0 3864 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_52
timestamp 1673029049
transform 1 0 4968 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_55
timestamp 1673029049
transform 1 0 5244 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_63
timestamp 1673029049
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_66
timestamp 1673029049
transform 1 0 6256 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_75
timestamp 1673029049
transform 1 0 7084 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_80
timestamp 1673029049
transform 1 0 7544 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_84
timestamp 1673029049
transform 1 0 7912 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_90
timestamp 1673029049
transform 1 0 8464 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_92
timestamp 1673029049
transform 1 0 8648 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_114
timestamp 1673029049
transform 1 0 10672 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_118
timestamp 1673029049
transform 1 0 11040 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_122
timestamp 1673029049
transform 1 0 11408 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_134
timestamp 1673029049
transform 1 0 12512 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_142
timestamp 1673029049
transform 1 0 13248 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_144
timestamp 1673029049
transform 1 0 13432 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_154
timestamp 1673029049
transform 1 0 14352 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_160
timestamp 1673029049
transform 1 0 14904 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_168
timestamp 1673029049
transform 1 0 15640 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_170
timestamp 1673029049
transform 1 0 15824 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_194
timestamp 1673029049
transform 1 0 18032 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_196
timestamp 1673029049
transform 1 0 18216 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_3
timestamp 1673029049
transform 1 0 460 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_24
timestamp 1673029049
transform 1 0 2392 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_27
timestamp 1673029049
transform 1 0 2668 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_37
timestamp 1673029049
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_43
timestamp 1673029049
transform 1 0 4140 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_47
timestamp 1673029049
transform 1 0 4508 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_51
timestamp 1673029049
transform 1 0 4876 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_53
timestamp 1673029049
transform 1 0 5060 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_75
timestamp 1673029049
transform 1 0 7084 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_79
timestamp 1673029049
transform 1 0 7452 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_101
timestamp 1673029049
transform 1 0 9476 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_105
timestamp 1673029049
transform 1 0 9844 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_108
timestamp 1673029049
transform 1 0 10120 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_116
timestamp 1673029049
transform 1 0 10856 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_122
timestamp 1673029049
transform 1 0 11408 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_129
timestamp 1673029049
transform 1 0 12052 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_131
timestamp 1673029049
transform 1 0 12236 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_136
timestamp 1673029049
transform 1 0 12696 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_143
timestamp 1673029049
transform 1 0 13340 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_154
timestamp 1673029049
transform 1 0 14352 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_157
timestamp 1673029049
transform 1 0 14628 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_164
timestamp 1673029049
transform 1 0 15272 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_171
timestamp 1673029049
transform 1 0 15916 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_177
timestamp 1673029049
transform 1 0 16468 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_181
timestamp 1673029049
transform 1 0 16836 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_183
timestamp 1673029049
transform 1 0 17020 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_192
timestamp 1673029049
transform 1 0 17848 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_198
timestamp 1673029049
transform 1 0 18400 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_3
timestamp 1673029049
transform 1 0 460 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_11
timestamp 1673029049
transform 1 0 1196 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_14
timestamp 1673029049
transform 1 0 1472 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_24
timestamp 1673029049
transform 1 0 2392 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_33
timestamp 1673029049
transform 1 0 3220 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_38
timestamp 1673029049
transform 1 0 3680 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_40
timestamp 1673029049
transform 1 0 3864 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_50
timestamp 1673029049
transform 1 0 4784 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_56
timestamp 1673029049
transform 1 0 5336 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_64
timestamp 1673029049
transform 1 0 6072 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_66
timestamp 1673029049
transform 1 0 6256 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_87
timestamp 1673029049
transform 1 0 8188 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_92
timestamp 1673029049
transform 1 0 8648 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_113
timestamp 1673029049
transform 1 0 10580 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_118
timestamp 1673029049
transform 1 0 11040 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_124
timestamp 1673029049
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_129
timestamp 1673029049
transform 1 0 12052 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_137
timestamp 1673029049
transform 1 0 12788 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_142
timestamp 1673029049
transform 1 0 13248 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_144
timestamp 1673029049
transform 1 0 13432 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_155
timestamp 1673029049
transform 1 0 14444 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_167
timestamp 1673029049
transform 1 0 15548 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_170
timestamp 1673029049
transform 1 0 15824 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_194
timestamp 1673029049
transform 1 0 18032 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_196
timestamp 1673029049
transform 1 0 18216 0 1 14688
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1673029049
transform 1 0 460 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_15
timestamp 1673029049
transform 1 0 1564 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_23
timestamp 1673029049
transform 1 0 2300 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_27
timestamp 1673029049
transform 1 0 2668 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_48
timestamp 1673029049
transform 1 0 4600 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_53
timestamp 1673029049
transform 1 0 5060 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_75
timestamp 1673029049
transform 1 0 7084 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_79
timestamp 1673029049
transform 1 0 7452 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_102
timestamp 1673029049
transform 1 0 9568 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_105
timestamp 1673029049
transform 1 0 9844 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_129
timestamp 1673029049
transform 1 0 12052 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_131
timestamp 1673029049
transform 1 0 12236 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_141
timestamp 1673029049
transform 1 0 13156 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_145
timestamp 1673029049
transform 1 0 13524 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_155
timestamp 1673029049
transform 1 0 14444 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_157
timestamp 1673029049
transform 1 0 14628 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_178
timestamp 1673029049
transform 1 0 16560 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_183
timestamp 1673029049
transform 1 0 17020 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_191
timestamp 1673029049
transform 1 0 17756 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_194
timestamp 1673029049
transform 1 0 18032 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_199
timestamp 1673029049
transform 1 0 18492 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_3
timestamp 1673029049
transform 1 0 460 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_11
timestamp 1673029049
transform 1 0 1196 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_14
timestamp 1673029049
transform 1 0 1472 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_22
timestamp 1673029049
transform 1 0 2208 0 1 15776
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_27
timestamp 1673029049
transform 1 0 2668 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_40
timestamp 1673029049
transform 1 0 3864 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_63
timestamp 1673029049
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_66
timestamp 1673029049
transform 1 0 6256 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_90
timestamp 1673029049
transform 1 0 8464 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_92
timestamp 1673029049
transform 1 0 8648 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_113
timestamp 1673029049
transform 1 0 10580 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_118
timestamp 1673029049
transform 1 0 11040 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_139
timestamp 1673029049
transform 1 0 12972 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_144
timestamp 1673029049
transform 1 0 13432 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_165
timestamp 1673029049
transform 1 0 15364 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_28_170
timestamp 1673029049
transform 1 0 15824 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_194
timestamp 1673029049
transform 1 0 18032 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_196
timestamp 1673029049
transform 1 0 18216 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_199
timestamp 1673029049
transform 1 0 18492 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_3
timestamp 1673029049
transform 1 0 460 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_11
timestamp 1673029049
transform 1 0 1196 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_18
timestamp 1673029049
transform 1 0 1840 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_25
timestamp 1673029049
transform 1 0 2484 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_27
timestamp 1673029049
transform 1 0 2668 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_31
timestamp 1673029049
transform 1 0 3036 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_39
timestamp 1673029049
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_51
timestamp 1673029049
transform 1 0 4876 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_53
timestamp 1673029049
transform 1 0 5060 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_75
timestamp 1673029049
transform 1 0 7084 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_79
timestamp 1673029049
transform 1 0 7452 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_29_103
timestamp 1673029049
transform 1 0 9660 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_105
timestamp 1673029049
transform 1 0 9844 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_126
timestamp 1673029049
transform 1 0 11776 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_131
timestamp 1673029049
transform 1 0 12236 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_139
timestamp 1673029049
transform 1 0 12972 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_146
timestamp 1673029049
transform 1 0 13616 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_155
timestamp 1673029049
transform 1 0 14444 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_157
timestamp 1673029049
transform 1 0 14628 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_29_181
timestamp 1673029049
transform 1 0 16836 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_183
timestamp 1673029049
transform 1 0 17020 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_192
timestamp 1673029049
transform 1 0 17848 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_199
timestamp 1673029049
transform 1 0 18492 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_3
timestamp 1673029049
transform 1 0 460 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_12
timestamp 1673029049
transform 1 0 1288 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_14
timestamp 1673029049
transform 1 0 1472 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_20
timestamp 1673029049
transform 1 0 2024 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_28
timestamp 1673029049
transform 1 0 2760 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_38
timestamp 1673029049
transform 1 0 3680 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_40
timestamp 1673029049
transform 1 0 3864 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_64
timestamp 1673029049
transform 1 0 6072 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_66
timestamp 1673029049
transform 1 0 6256 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_89
timestamp 1673029049
transform 1 0 8372 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_92
timestamp 1673029049
transform 1 0 8648 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_114
timestamp 1673029049
transform 1 0 10672 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_118
timestamp 1673029049
transform 1 0 11040 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_130
timestamp 1673029049
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_142
timestamp 1673029049
transform 1 0 13248 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_144
timestamp 1673029049
transform 1 0 13432 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_168
timestamp 1673029049
transform 1 0 15640 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_170
timestamp 1673029049
transform 1 0 15824 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_30_194
timestamp 1673029049
transform 1 0 18032 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_196
timestamp 1673029049
transform 1 0 18216 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_3
timestamp 1673029049
transform 1 0 460 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_24
timestamp 1673029049
transform 1 0 2392 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_27
timestamp 1673029049
transform 1 0 2668 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_33
timestamp 1673029049
transform 1 0 3220 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_51
timestamp 1673029049
transform 1 0 4876 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_53
timestamp 1673029049
transform 1 0 5060 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_74
timestamp 1673029049
transform 1 0 6992 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_79
timestamp 1673029049
transform 1 0 7452 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_103
timestamp 1673029049
transform 1 0 9660 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_105
timestamp 1673029049
transform 1 0 9844 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_126
timestamp 1673029049
transform 1 0 11776 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_131
timestamp 1673029049
transform 1 0 12236 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_136
timestamp 1673029049
transform 1 0 12696 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_154
timestamp 1673029049
transform 1 0 14352 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_157
timestamp 1673029049
transform 1 0 14628 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_179
timestamp 1673029049
transform 1 0 16652 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_183
timestamp 1673029049
transform 1 0 17020 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_188
timestamp 1673029049
transform 1 0 17480 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_3
timestamp 1673029049
transform 1 0 460 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_8
timestamp 1673029049
transform 1 0 920 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_12
timestamp 1673029049
transform 1 0 1288 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_14
timestamp 1673029049
transform 1 0 1472 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_18
timestamp 1673029049
transform 1 0 1840 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_25
timestamp 1673029049
transform 1 0 2484 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1673029049
transform 1 0 2668 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_30
timestamp 1673029049
transform 1 0 2944 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_38
timestamp 1673029049
transform 1 0 3680 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_40
timestamp 1673029049
transform 1 0 3864 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_49
timestamp 1673029049
transform 1 0 4692 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_53
timestamp 1673029049
transform 1 0 5060 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_64
timestamp 1673029049
transform 1 0 6072 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_66
timestamp 1673029049
transform 1 0 6256 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_69
timestamp 1673029049
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_77
timestamp 1673029049
transform 1 0 7268 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_79
timestamp 1673029049
transform 1 0 7452 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_89
timestamp 1673029049
transform 1 0 8372 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_92
timestamp 1673029049
transform 1 0 8648 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_101
timestamp 1673029049
transform 1 0 9476 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_32_105
timestamp 1673029049
transform 1 0 9844 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_115
timestamp 1673029049
transform 1 0 10764 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_118
timestamp 1673029049
transform 1 0 11040 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_127
timestamp 1673029049
transform 1 0 11868 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_32_131
timestamp 1673029049
transform 1 0 12236 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_139
timestamp 1673029049
transform 1 0 12972 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_144
timestamp 1673029049
transform 1 0 13432 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_32_153
timestamp 1673029049
transform 1 0 14260 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_157
timestamp 1673029049
transform 1 0 14628 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_164
timestamp 1673029049
transform 1 0 15272 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_168
timestamp 1673029049
transform 1 0 15640 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_170
timestamp 1673029049
transform 1 0 15824 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_179
timestamp 1673029049
transform 1 0 16652 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_183
timestamp 1673029049
transform 1 0 17020 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_194
timestamp 1673029049
transform 1 0 18032 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_196
timestamp 1673029049
transform 1 0 18216 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_199
timestamp 1673029049
transform 1 0 18492 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1673029049
transform 1 0 184 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1673029049
transform -1 0 18860 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1673029049
transform 1 0 184 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1673029049
transform -1 0 18860 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1673029049
transform 1 0 184 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1673029049
transform -1 0 18860 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1673029049
transform 1 0 184 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1673029049
transform -1 0 18860 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1673029049
transform 1 0 184 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1673029049
transform -1 0 18860 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1673029049
transform 1 0 184 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1673029049
transform -1 0 18860 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1673029049
transform 1 0 184 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1673029049
transform -1 0 18860 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1673029049
transform 1 0 184 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1673029049
transform -1 0 18860 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1673029049
transform 1 0 184 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1673029049
transform -1 0 18860 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1673029049
transform 1 0 184 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1673029049
transform -1 0 18860 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1673029049
transform 1 0 184 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1673029049
transform -1 0 18860 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1673029049
transform 1 0 184 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1673029049
transform -1 0 18860 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1673029049
transform 1 0 184 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1673029049
transform -1 0 18860 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1673029049
transform 1 0 184 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1673029049
transform -1 0 18860 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1673029049
transform 1 0 184 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1673029049
transform -1 0 18860 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1673029049
transform 1 0 184 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1673029049
transform -1 0 18860 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1673029049
transform 1 0 184 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1673029049
transform -1 0 18860 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1673029049
transform 1 0 184 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1673029049
transform -1 0 18860 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1673029049
transform 1 0 184 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1673029049
transform -1 0 18860 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1673029049
transform 1 0 184 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1673029049
transform -1 0 18860 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1673029049
transform 1 0 184 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1673029049
transform -1 0 18860 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1673029049
transform 1 0 184 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1673029049
transform -1 0 18860 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1673029049
transform 1 0 184 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1673029049
transform -1 0 18860 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1673029049
transform 1 0 184 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1673029049
transform -1 0 18860 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1673029049
transform 1 0 184 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1673029049
transform -1 0 18860 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1673029049
transform 1 0 184 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1673029049
transform -1 0 18860 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1673029049
transform 1 0 184 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1673029049
transform -1 0 18860 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1673029049
transform 1 0 184 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1673029049
transform -1 0 18860 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1673029049
transform 1 0 184 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1673029049
transform -1 0 18860 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1673029049
transform 1 0 184 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1673029049
transform -1 0 18860 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1673029049
transform 1 0 184 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1673029049
transform -1 0 18860 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1673029049
transform 1 0 184 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1673029049
transform -1 0 18860 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1673029049
transform 1 0 184 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1673029049
transform -1 0 18860 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66 swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 1380 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1673029049
transform 1 0 2576 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1673029049
transform 1 0 3772 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1673029049
transform 1 0 4968 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1673029049
transform 1 0 6164 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1673029049
transform 1 0 7360 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1673029049
transform 1 0 8556 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1673029049
transform 1 0 9752 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1673029049
transform 1 0 10948 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1673029049
transform 1 0 12144 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1673029049
transform 1 0 13340 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1673029049
transform 1 0 14536 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1673029049
transform 1 0 15732 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1673029049
transform 1 0 16928 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1673029049
transform 1 0 18124 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1673029049
transform 1 0 2576 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1673029049
transform 1 0 4968 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1673029049
transform 1 0 7360 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1673029049
transform 1 0 9752 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1673029049
transform 1 0 12144 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1673029049
transform 1 0 14536 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1673029049
transform 1 0 16928 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1673029049
transform 1 0 1380 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1673029049
transform 1 0 3772 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1673029049
transform 1 0 6164 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1673029049
transform 1 0 8556 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1673029049
transform 1 0 10948 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1673029049
transform 1 0 13340 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1673029049
transform 1 0 15732 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1673029049
transform 1 0 18124 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1673029049
transform 1 0 2576 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1673029049
transform 1 0 4968 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1673029049
transform 1 0 7360 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1673029049
transform 1 0 9752 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1673029049
transform 1 0 12144 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1673029049
transform 1 0 14536 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1673029049
transform 1 0 16928 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1673029049
transform 1 0 1380 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1673029049
transform 1 0 3772 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1673029049
transform 1 0 6164 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1673029049
transform 1 0 8556 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1673029049
transform 1 0 10948 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1673029049
transform 1 0 13340 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1673029049
transform 1 0 15732 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1673029049
transform 1 0 18124 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1673029049
transform 1 0 2576 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1673029049
transform 1 0 4968 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1673029049
transform 1 0 7360 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1673029049
transform 1 0 9752 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1673029049
transform 1 0 12144 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1673029049
transform 1 0 14536 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1673029049
transform 1 0 16928 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1673029049
transform 1 0 1380 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1673029049
transform 1 0 3772 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1673029049
transform 1 0 6164 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1673029049
transform 1 0 8556 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1673029049
transform 1 0 10948 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1673029049
transform 1 0 13340 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1673029049
transform 1 0 15732 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1673029049
transform 1 0 18124 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1673029049
transform 1 0 2576 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1673029049
transform 1 0 4968 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1673029049
transform 1 0 7360 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1673029049
transform 1 0 9752 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1673029049
transform 1 0 12144 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1673029049
transform 1 0 14536 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1673029049
transform 1 0 16928 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1673029049
transform 1 0 1380 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1673029049
transform 1 0 3772 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1673029049
transform 1 0 6164 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1673029049
transform 1 0 8556 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1673029049
transform 1 0 10948 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1673029049
transform 1 0 13340 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1673029049
transform 1 0 15732 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1673029049
transform 1 0 18124 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1673029049
transform 1 0 2576 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1673029049
transform 1 0 4968 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1673029049
transform 1 0 7360 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1673029049
transform 1 0 9752 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1673029049
transform 1 0 12144 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1673029049
transform 1 0 14536 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1673029049
transform 1 0 16928 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1673029049
transform 1 0 1380 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1673029049
transform 1 0 3772 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1673029049
transform 1 0 6164 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1673029049
transform 1 0 8556 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1673029049
transform 1 0 10948 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1673029049
transform 1 0 13340 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1673029049
transform 1 0 15732 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1673029049
transform 1 0 18124 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1673029049
transform 1 0 2576 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1673029049
transform 1 0 4968 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1673029049
transform 1 0 7360 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1673029049
transform 1 0 9752 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1673029049
transform 1 0 12144 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1673029049
transform 1 0 14536 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1673029049
transform 1 0 16928 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1673029049
transform 1 0 1380 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1673029049
transform 1 0 3772 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1673029049
transform 1 0 6164 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1673029049
transform 1 0 8556 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1673029049
transform 1 0 10948 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1673029049
transform 1 0 13340 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1673029049
transform 1 0 15732 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1673029049
transform 1 0 18124 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1673029049
transform 1 0 2576 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1673029049
transform 1 0 4968 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1673029049
transform 1 0 7360 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1673029049
transform 1 0 9752 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1673029049
transform 1 0 12144 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1673029049
transform 1 0 14536 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1673029049
transform 1 0 16928 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1673029049
transform 1 0 1380 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1673029049
transform 1 0 3772 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1673029049
transform 1 0 6164 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1673029049
transform 1 0 8556 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1673029049
transform 1 0 10948 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1673029049
transform 1 0 13340 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1673029049
transform 1 0 15732 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1673029049
transform 1 0 18124 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1673029049
transform 1 0 2576 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1673029049
transform 1 0 4968 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1673029049
transform 1 0 7360 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1673029049
transform 1 0 9752 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1673029049
transform 1 0 12144 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1673029049
transform 1 0 14536 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1673029049
transform 1 0 16928 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1673029049
transform 1 0 1380 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1673029049
transform 1 0 3772 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1673029049
transform 1 0 6164 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1673029049
transform 1 0 8556 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1673029049
transform 1 0 10948 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1673029049
transform 1 0 13340 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1673029049
transform 1 0 15732 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1673029049
transform 1 0 18124 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1673029049
transform 1 0 2576 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1673029049
transform 1 0 4968 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1673029049
transform 1 0 7360 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1673029049
transform 1 0 9752 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1673029049
transform 1 0 12144 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1673029049
transform 1 0 14536 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1673029049
transform 1 0 16928 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1673029049
transform 1 0 1380 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1673029049
transform 1 0 3772 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1673029049
transform 1 0 6164 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1673029049
transform 1 0 8556 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1673029049
transform 1 0 10948 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1673029049
transform 1 0 13340 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1673029049
transform 1 0 15732 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1673029049
transform 1 0 18124 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1673029049
transform 1 0 2576 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1673029049
transform 1 0 4968 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1673029049
transform 1 0 7360 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1673029049
transform 1 0 9752 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1673029049
transform 1 0 12144 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1673029049
transform 1 0 14536 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1673029049
transform 1 0 16928 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1673029049
transform 1 0 1380 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1673029049
transform 1 0 3772 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1673029049
transform 1 0 6164 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1673029049
transform 1 0 8556 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1673029049
transform 1 0 10948 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1673029049
transform 1 0 13340 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1673029049
transform 1 0 15732 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1673029049
transform 1 0 18124 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1673029049
transform 1 0 2576 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1673029049
transform 1 0 4968 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1673029049
transform 1 0 7360 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1673029049
transform 1 0 9752 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1673029049
transform 1 0 12144 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1673029049
transform 1 0 14536 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1673029049
transform 1 0 16928 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1673029049
transform 1 0 1380 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1673029049
transform 1 0 3772 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1673029049
transform 1 0 6164 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1673029049
transform 1 0 8556 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1673029049
transform 1 0 10948 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1673029049
transform 1 0 13340 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1673029049
transform 1 0 15732 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1673029049
transform 1 0 18124 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1673029049
transform 1 0 2576 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1673029049
transform 1 0 4968 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1673029049
transform 1 0 7360 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1673029049
transform 1 0 9752 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1673029049
transform 1 0 12144 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1673029049
transform 1 0 14536 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1673029049
transform 1 0 16928 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1673029049
transform 1 0 1380 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1673029049
transform 1 0 3772 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1673029049
transform 1 0 6164 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1673029049
transform 1 0 8556 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1673029049
transform 1 0 10948 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1673029049
transform 1 0 13340 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1673029049
transform 1 0 15732 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1673029049
transform 1 0 18124 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1673029049
transform 1 0 2576 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1673029049
transform 1 0 4968 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1673029049
transform 1 0 7360 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1673029049
transform 1 0 9752 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1673029049
transform 1 0 12144 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1673029049
transform 1 0 14536 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1673029049
transform 1 0 16928 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1673029049
transform 1 0 1380 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1673029049
transform 1 0 3772 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1673029049
transform 1 0 6164 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1673029049
transform 1 0 8556 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1673029049
transform 1 0 10948 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1673029049
transform 1 0 13340 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1673029049
transform 1 0 15732 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1673029049
transform 1 0 18124 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1673029049
transform 1 0 2576 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1673029049
transform 1 0 4968 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1673029049
transform 1 0 7360 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1673029049
transform 1 0 9752 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1673029049
transform 1 0 12144 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1673029049
transform 1 0 14536 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1673029049
transform 1 0 16928 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1673029049
transform 1 0 1380 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1673029049
transform 1 0 3772 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1673029049
transform 1 0 6164 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1673029049
transform 1 0 8556 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1673029049
transform 1 0 10948 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1673029049
transform 1 0 13340 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1673029049
transform 1 0 15732 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1673029049
transform 1 0 18124 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1673029049
transform 1 0 2576 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1673029049
transform 1 0 4968 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1673029049
transform 1 0 7360 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1673029049
transform 1 0 9752 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1673029049
transform 1 0 12144 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1673029049
transform 1 0 14536 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1673029049
transform 1 0 16928 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1673029049
transform 1 0 1380 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1673029049
transform 1 0 3772 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1673029049
transform 1 0 6164 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1673029049
transform 1 0 8556 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1673029049
transform 1 0 10948 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1673029049
transform 1 0 13340 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1673029049
transform 1 0 15732 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1673029049
transform 1 0 18124 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1673029049
transform 1 0 2576 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1673029049
transform 1 0 4968 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1673029049
transform 1 0 7360 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1673029049
transform 1 0 9752 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1673029049
transform 1 0 12144 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1673029049
transform 1 0 14536 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1673029049
transform 1 0 16928 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1673029049
transform 1 0 1380 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1673029049
transform 1 0 2576 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1673029049
transform 1 0 3772 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1673029049
transform 1 0 4968 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1673029049
transform 1 0 6164 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1673029049
transform 1 0 7360 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1673029049
transform 1 0 8556 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1673029049
transform 1 0 9752 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1673029049
transform 1 0 10948 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1673029049
transform 1 0 12144 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1673029049
transform 1 0 13340 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1673029049
transform 1 0 14536 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1673029049
transform 1 0 15732 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1673029049
transform 1 0 16928 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1673029049
transform 1 0 18124 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _204_ swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 1656 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _205_
timestamp 1673029049
transform 1 0 12328 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _206_
timestamp 1673029049
transform -1 0 8280 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _207_
timestamp 1673029049
transform -1 0 6072 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _208_
timestamp 1673029049
transform 1 0 7544 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _209_
timestamp 1673029049
transform 1 0 17296 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _210_
timestamp 1673029049
transform 1 0 9936 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _211_
timestamp 1673029049
transform 1 0 3956 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _212_
timestamp 1673029049
transform 1 0 2668 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _213_
timestamp 1673029049
transform 1 0 3956 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _214_
timestamp 1673029049
transform 1 0 1748 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _215_
timestamp 1673029049
transform 1 0 1012 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _216_
timestamp 1673029049
transform -1 0 3680 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _217_
timestamp 1673029049
transform 1 0 2852 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _218_
timestamp 1673029049
transform 1 0 6348 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _219_
timestamp 1673029049
transform 1 0 5336 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _220_
timestamp 1673029049
transform 1 0 8188 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _221_
timestamp 1673029049
transform 1 0 7544 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _222_
timestamp 1673029049
transform 1 0 7636 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _223_
timestamp 1673029049
transform 1 0 6992 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _224_
timestamp 1673029049
transform -1 0 10304 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _225_
timestamp 1673029049
transform 1 0 9936 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _226_
timestamp 1673029049
transform 1 0 2760 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _227_
timestamp 1673029049
transform 1 0 2760 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _228_
timestamp 1673029049
transform 1 0 12144 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _229_
timestamp 1673029049
transform 1 0 12604 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _230_
timestamp 1673029049
transform 1 0 12144 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _231_
timestamp 1673029049
transform -1 0 14352 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _232_
timestamp 1673029049
transform 1 0 13524 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _233_
timestamp 1673029049
transform -1 0 14444 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _234_
timestamp 1673029049
transform 1 0 14720 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _235_
timestamp 1673029049
transform -1 0 12144 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _236_
timestamp 1673029049
transform 1 0 12328 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _237_
timestamp 1673029049
transform -1 0 15548 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _238_
timestamp 1673029049
transform 1 0 14720 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _239_
timestamp 1673029049
transform 1 0 13708 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _240_
timestamp 1673029049
transform 1 0 12420 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _241_
timestamp 1673029049
transform 1 0 11500 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _242_
timestamp 1673029049
transform 1 0 11224 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _243_
timestamp 1673029049
transform 1 0 17112 0 -1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _244_
timestamp 1673029049
transform 1 0 16928 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _245_ swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 15640 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_4  _246_ swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 6992 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_2  _247_ swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 2852 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _248_
timestamp 1673029049
transform 1 0 3220 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _249_
timestamp 1673029049
transform -1 0 2392 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_4  _250_
timestamp 1673029049
transform -1 0 8924 0 -1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _251_
timestamp 1673029049
transform 1 0 18124 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _252_
timestamp 1673029049
transform -1 0 10856 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _253_
timestamp 1673029049
transform -1 0 14904 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_4  _254_
timestamp 1673029049
transform -1 0 15364 0 -1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  _255_
timestamp 1673029049
transform 1 0 17848 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  _256_
timestamp 1673029049
transform 1 0 12328 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__inv_4  _257__7 swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 13616 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _258_
timestamp 1673029049
transform -1 0 1012 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_4  _259__4
timestamp 1673029049
transform -1 0 2116 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _260_
timestamp 1673029049
transform -1 0 5336 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _261_
timestamp 1673029049
transform -1 0 11408 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_4  _262__1
timestamp 1673029049
transform -1 0 15272 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _263_
timestamp 1673029049
transform -1 0 12052 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _264_
timestamp 1673029049
transform 1 0 11132 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__nor3b_2  _265_ swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 12328 0 1 16864
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_2  _266_ swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 12052 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _267_ swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 17756 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_2  _268_ swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 14904 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _269_ swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 16468 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__o211ai_4  _270_ swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 15456 0 1 12512
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _271_
timestamp 1673029049
transform 1 0 12512 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _272_ swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 14720 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__a41oi_1  _273_ swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 14352 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _274_ swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 13984 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _275_ swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 11132 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__nand2b_1  _276_ swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 12880 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _277_
timestamp 1673029049
transform 1 0 12972 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2ai_1  _278_ swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 14444 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _279_
timestamp 1673029049
transform -1 0 2116 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _280_
timestamp 1673029049
transform -1 0 4876 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nor3b_2  _281_
timestamp 1673029049
transform -1 0 4876 0 1 1632
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_2  _282_
timestamp 1673029049
transform 1 0 2852 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _283_
timestamp 1673029049
transform 1 0 8004 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _284_ swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 6532 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_2  _285_ swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 7728 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_4  _286_
timestamp 1673029049
transform -1 0 5520 0 1 3808
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _287_
timestamp 1673029049
transform 1 0 1840 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__o2111a_1  _288_ swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 5980 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _289_
timestamp 1673029049
transform 1 0 5704 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__nand2b_1  _290_
timestamp 1673029049
transform -1 0 4048 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _291_
timestamp 1673029049
transform 1 0 5152 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2ai_1  _292_
timestamp 1673029049
transform 1 0 5152 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _293_
timestamp 1673029049
transform -1 0 3588 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2ai_1  _294_
timestamp 1673029049
transform 1 0 2760 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _295_
timestamp 1673029049
transform 1 0 2392 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _296_
timestamp 1673029049
transform -1 0 3680 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _297_
timestamp 1673029049
transform 1 0 7544 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _298_
timestamp 1673029049
transform -1 0 8372 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_2  _299_ swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 9476 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_1  _300_ swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 17480 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__nand2b_1  _301_
timestamp 1673029049
transform 1 0 15456 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _302_
timestamp 1673029049
transform -1 0 13800 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_2  _303_
timestamp 1673029049
transform 1 0 12512 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__nand2b_2  _304_ swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 7544 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _305_ swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 6808 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _306_
timestamp 1673029049
transform -1 0 7268 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__o31ai_2  _307_ swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 6900 0 1 11424
box -38 -48 958 592
use sky130_fd_sc_hd__nand2b_2  _308_
timestamp 1673029049
transform -1 0 17664 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _309_
timestamp 1673029049
transform 1 0 15916 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _310_
timestamp 1673029049
transform 1 0 16560 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__o31ai_2  _311_
timestamp 1673029049
transform 1 0 15916 0 1 12512
box -38 -48 958 592
use sky130_fd_sc_hd__xnor2_1  _312_ swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 3036 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _313_
timestamp 1673029049
transform 1 0 1840 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _314_
timestamp 1673029049
transform 1 0 3772 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _315_
timestamp 1673029049
transform 1 0 4048 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _316_
timestamp 1673029049
transform -1 0 4048 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _317_
timestamp 1673029049
transform -1 0 3036 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _318_ swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 3680 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _319_
timestamp 1673029049
transform 1 0 2852 0 -1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _320_
timestamp 1673029049
transform -1 0 5520 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _321_
timestamp 1673029049
transform 1 0 5244 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__nand2b_1  _322_
timestamp 1673029049
transform 1 0 5520 0 -1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _323_
timestamp 1673029049
transform 1 0 6624 0 -1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _324_
timestamp 1673029049
transform 1 0 9936 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _325_
timestamp 1673029049
transform 1 0 10304 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__nand2b_1  _326_
timestamp 1673029049
transform -1 0 10120 0 1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _327_
timestamp 1673029049
transform 1 0 2576 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _328_
timestamp 1673029049
transform -1 0 13156 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _329_
timestamp 1673029049
transform 1 0 11776 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _330_
timestamp 1673029049
transform 1 0 13616 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _331_
timestamp 1673029049
transform 1 0 13064 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _332_
timestamp 1673029049
transform 1 0 13524 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _333_
timestamp 1673029049
transform -1 0 11408 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _334_
timestamp 1673029049
transform -1 0 12880 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _335_
timestamp 1673029049
transform -1 0 14444 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _336_
timestamp 1673029049
transform 1 0 17112 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _337_
timestamp 1673029049
transform -1 0 12696 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__nand2b_1  _338_
timestamp 1673029049
transform -1 0 12052 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _339_
timestamp 1673029049
transform 1 0 13156 0 -1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _340_
timestamp 1673029049
transform 1 0 11316 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _341_
timestamp 1673029049
transform 1 0 10764 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__nand2b_1  _342_
timestamp 1673029049
transform 1 0 11316 0 -1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _343_
timestamp 1673029049
transform 1 0 15916 0 -1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _344_ swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 2116 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__o2111ai_2  _345_ swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 14444 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__a21oi_1  _346_
timestamp 1673029049
transform 1 0 15916 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _347_
timestamp 1673029049
transform -1 0 15364 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__nand4bb_1  _348_ swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 3956 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _349_
timestamp 1673029049
transform 1 0 3772 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _350_
timestamp 1673029049
transform 1 0 4600 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _351_
timestamp 1673029049
transform 1 0 5152 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _352_
timestamp 1673029049
transform 1 0 5244 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _353_ swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 5888 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _354_
timestamp 1673029049
transform -1 0 5428 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _355_
timestamp 1673029049
transform 1 0 5612 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _356_
timestamp 1673029049
transform 1 0 6256 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _357_ swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 6992 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_1  _358_ swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 2116 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _359_
timestamp 1673029049
transform 1 0 736 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__nand3b_1  _360_
timestamp 1673029049
transform 1 0 4048 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _361_
timestamp 1673029049
transform -1 0 4876 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _362_
timestamp 1673029049
transform 1 0 1564 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _363_
timestamp 1673029049
transform 1 0 1564 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _364_
timestamp 1673029049
transform 1 0 6808 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _365_
timestamp 1673029049
transform -1 0 9108 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _366_
timestamp 1673029049
transform -1 0 8280 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _367_ swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 6532 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _368_
timestamp 1673029049
transform -1 0 8556 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _369_
timestamp 1673029049
transform 1 0 8740 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _370_
timestamp 1673029049
transform 1 0 1564 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _371_
timestamp 1673029049
transform 1 0 1564 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__nor4_1  _372_ swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 2024 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__o31ai_1  _373_ swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 1840 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _374_
timestamp 1673029049
transform -1 0 1288 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_2  _375_ swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 4876 0 -1 16864
box -38 -48 958 592
use sky130_fd_sc_hd__o21ba_2  _376_ swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 4692 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_1  _377_
timestamp 1673029049
transform -1 0 17756 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__nand3b_1  _378_
timestamp 1673029049
transform -1 0 17756 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _379_ swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 17848 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _380_
timestamp 1673029049
transform -1 0 16836 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _381_
timestamp 1673029049
transform 1 0 17112 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _382_
timestamp 1673029049
transform 1 0 17756 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _383_
timestamp 1673029049
transform -1 0 17756 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _384_
timestamp 1673029049
transform 1 0 15916 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _385_
timestamp 1673029049
transform 1 0 14720 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _386_
timestamp 1673029049
transform -1 0 15732 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _387_
timestamp 1673029049
transform 1 0 14720 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_1  _388_
timestamp 1673029049
transform -1 0 12880 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _389_
timestamp 1673029049
transform 1 0 11132 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__nand3b_1  _390_
timestamp 1673029049
transform -1 0 12788 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _391_
timestamp 1673029049
transform -1 0 11408 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _392_
timestamp 1673029049
transform 1 0 11132 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _393_
timestamp 1673029049
transform 1 0 11132 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _394_
timestamp 1673029049
transform 1 0 14076 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _395_
timestamp 1673029049
transform 1 0 13708 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__o21bai_1  _396_ swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 12512 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _397_ swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 12328 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__o21bai_1  _398_
timestamp 1673029049
transform 1 0 10948 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _399_
timestamp 1673029049
transform 1 0 11132 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__o2111ai_1  _400_ swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 8740 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _401_
timestamp 1673029049
transform 1 0 8740 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _402_
timestamp 1673029049
transform 1 0 7912 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _403_
timestamp 1673029049
transform 1 0 16008 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _404_
timestamp 1673029049
transform 1 0 15916 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__nor4_1  _405_
timestamp 1673029049
transform -1 0 17388 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__o31ai_1  _406_
timestamp 1673029049
transform 1 0 17112 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _407_
timestamp 1673029049
transform 1 0 17572 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  _408__8
timestamp 1673029049
transform -1 0 11592 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  _409__9
timestamp 1673029049
transform 1 0 5612 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  _410__5
timestamp 1673029049
transform -1 0 5704 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  _411__6
timestamp 1673029049
transform -1 0 2116 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  _412__2
timestamp 1673029049
transform -1 0 16376 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  _413__3
timestamp 1673029049
transform -1 0 10488 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__dfstp_1  _414_ swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 10672 0 1 16864
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _415_
timestamp 1673029049
transform -1 0 9660 0 -1 16864
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _416__31 swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 2208 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  _416_
timestamp 1673029049
transform 1 0 6440 0 1 16864
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _417_ swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 7084 0 -1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _418_
timestamp 1673029049
transform 1 0 6348 0 1 14688
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _419_
timestamp 1673029049
transform 1 0 14720 0 -1 9248
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _420_
timestamp 1673029049
transform 1 0 4140 0 1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _421_ swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 4416 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _422_
timestamp 1673029049
transform 1 0 3312 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _423_
timestamp 1673029049
transform -1 0 6624 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfstp_1  _424_
timestamp 1673029049
transform 1 0 5152 0 -1 14688
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _425_
timestamp 1673029049
transform 1 0 7820 0 -1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtn_1  _426_ swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 552 0 -1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_2  _427_ swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 1564 0 1 5984
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtn_1  _428_
timestamp 1673029049
transform 1 0 4232 0 1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _429_
timestamp 1673029049
transform 1 0 5152 0 -1 8160
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtn_1  _430_
timestamp 1673029049
transform 1 0 644 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _431_
timestamp 1673029049
transform 1 0 1564 0 1 11424
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtn_1  _432_
timestamp 1673029049
transform 1 0 552 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _433_ swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 8740 0 1 5984
box -38 -48 2154 592
use sky130_fd_sc_hd__dfstp_2  _434_
timestamp 1673029049
transform 1 0 6348 0 1 5984
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _435_
timestamp 1673029049
transform 1 0 8740 0 1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_2  _436_
timestamp 1673029049
transform 1 0 552 0 -1 13600
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _437_
timestamp 1673029049
transform 1 0 552 0 -1 14688
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _438_
timestamp 1673029049
transform 1 0 552 0 -1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _439_
timestamp 1673029049
transform -1 0 9476 0 -1 14688
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _440_
timestamp 1673029049
transform -1 0 9660 0 -1 12512
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _441_
timestamp 1673029049
transform -1 0 9384 0 -1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _442_
timestamp 1673029049
transform 1 0 7728 0 -1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _443_
timestamp 1673029049
transform 1 0 8740 0 1 11424
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _444_ swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 8740 0 1 13600
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_1  _445_
timestamp 1673029049
transform -1 0 4876 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _446_
timestamp 1673029049
transform 1 0 16560 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _447_
timestamp 1673029049
transform 1 0 16560 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _448_
timestamp 1673029049
transform 1 0 12512 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfstp_1  _449_
timestamp 1673029049
transform 1 0 16100 0 1 8160
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _450_
timestamp 1673029049
transform 1 0 13800 0 1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtn_1  _451_
timestamp 1673029049
transform 1 0 10212 0 -1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _452_
timestamp 1673029049
transform 1 0 14720 0 -1 17952
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtn_1  _453_
timestamp 1673029049
transform 1 0 10212 0 -1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _454_
timestamp 1673029049
transform 1 0 14720 0 -1 11424
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtn_1  _455_
timestamp 1673029049
transform 1 0 10120 0 -1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _456_
timestamp 1673029049
transform 1 0 9936 0 -1 9248
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtn_1  _457_
timestamp 1673029049
transform 1 0 9936 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _458_
timestamp 1673029049
transform 1 0 13524 0 1 4896
box -38 -48 2154 592
use sky130_fd_sc_hd__dfstp_1  _459_
timestamp 1673029049
transform -1 0 13156 0 1 4896
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _460_
timestamp 1673029049
transform 1 0 10212 0 -1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _461_
timestamp 1673029049
transform 1 0 7544 0 -1 9248
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_2  _462_
timestamp 1673029049
transform 1 0 15916 0 1 5984
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _463_
timestamp 1673029049
transform 1 0 15916 0 1 4896
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _464_
timestamp 1673029049
transform 1 0 14996 0 -1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _465_
timestamp 1673029049
transform 1 0 16192 0 1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _466_
timestamp 1673029049
transform 1 0 16100 0 1 16864
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _467_
timestamp 1673029049
transform 1 0 13800 0 1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _468_
timestamp 1673029049
transform 1 0 16192 0 1 14688
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _469_
timestamp 1673029049
transform 1 0 16100 0 1 15776
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _470_
timestamp 1673029049
transform 1 0 14904 0 -1 16864
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__037_ swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 9936 0 -1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_divider.out
timestamp 1673029049
transform 1 0 8740 0 1 14688
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_divider2.out
timestamp 1673029049
transform -1 0 16560 0 -1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_ext_clk
timestamp 1673029049
transform 1 0 5152 0 -1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_net11
timestamp 1673029049
transform 1 0 7820 0 -1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_pll_clk90
timestamp 1673029049
transform -1 0 15640 0 1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_pll_clk
timestamp 1673029049
transform -1 0 6072 0 1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__037_
timestamp 1673029049
transform -1 0 7084 0 -1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_divider.out
timestamp 1673029049
transform -1 0 9660 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_divider2.out
timestamp 1673029049
transform -1 0 15364 0 1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_ext_clk
timestamp 1673029049
transform -1 0 4600 0 -1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_net11
timestamp 1673029049
transform -1 0 7084 0 -1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_pll_clk90
timestamp 1673029049
transform -1 0 14444 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_pll_clk
timestamp 1673029049
transform -1 0 4600 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__037_
timestamp 1673029049
transform 1 0 11132 0 1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_divider.out
timestamp 1673029049
transform 1 0 8740 0 1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_divider2.out
timestamp 1673029049
transform 1 0 14996 0 -1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_ext_clk
timestamp 1673029049
transform 1 0 4232 0 1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_net11
timestamp 1673029049
transform 1 0 6624 0 1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_pll_clk90
timestamp 1673029049
transform -1 0 14444 0 -1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_pll_clk
timestamp 1673029049
transform -1 0 4600 0 -1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_4  fanout14 swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 12972 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout15 swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 14260 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout16
timestamp 1673029049
transform -1 0 15272 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout17 swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 18400 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout18
timestamp 1673029049
transform -1 0 10120 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout19
timestamp 1673029049
transform -1 0 10488 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout20
timestamp 1673029049
transform -1 0 9108 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout21
timestamp 1673029049
transform -1 0 5336 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout22
timestamp 1673029049
transform 1 0 15548 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout23
timestamp 1673029049
transform -1 0 15640 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout24 swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 7452 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout25
timestamp 1673029049
transform -1 0 9292 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout26
timestamp 1673029049
transform 1 0 3220 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout27
timestamp 1673029049
transform -1 0 3680 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout28
timestamp 1673029049
transform 1 0 10856 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout29
timestamp 1673029049
transform 1 0 6716 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout30
timestamp 1673029049
transform 1 0 2852 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 11868 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1673029049
transform 1 0 2944 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1673029049
transform -1 0 16652 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1673029049
transform -1 0 17848 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1673029049
transform -1 0 17848 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1673029049
transform 1 0 6348 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1673029049
transform 1 0 8740 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1 swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 18032 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1673029049
transform 1 0 17756 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1673029049
transform -1 0 828 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1673029049
transform -1 0 1840 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1673029049
transform 1 0 18216 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1673029049
transform 1 0 18216 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1673029049
transform 1 0 18216 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1673029049
transform 1 0 18216 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1673029049
transform 1 0 18216 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1673029049
transform 1 0 18216 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  output12 swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 12880 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  user_clk_out_buffer
timestamp 1673029049
transform 1 0 9936 0 -1 16864
box -38 -48 1878 592
<< labels >>
flabel metal4 s 3100 496 3420 18544 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 6200 496 6520 18544 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 9300 496 9620 18544 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 12400 496 12720 18544 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 15500 496 15820 18544 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 18600 496 18920 18544 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 1550 496 1870 18544 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 4650 496 4970 18544 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 7750 496 8070 18544 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 10850 496 11170 18544 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 13950 496 14270 18544 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 17050 496 17370 18544 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 7102 19200 7158 20000 0 FreeSans 224 90 0 0 core_clk
port 2 nsew signal tristate
flabel metal2 s 4250 19200 4306 20000 0 FreeSans 224 90 0 0 ext_clk
port 3 nsew signal input
flabel metal3 s 19200 1368 20000 1488 0 FreeSans 480 0 0 0 ext_clk_sel
port 4 nsew signal input
flabel metal3 s 19200 18504 20000 18624 0 FreeSans 480 0 0 0 ext_reset
port 5 nsew signal input
flabel metal2 s 15658 19200 15714 20000 0 FreeSans 224 90 0 0 pll_clk
port 6 nsew signal input
flabel metal2 s 18510 19200 18566 20000 0 FreeSans 224 90 0 0 pll_clk90
port 7 nsew signal input
flabel metal3 s 0 9936 800 10056 0 FreeSans 480 0 0 0 porb
port 8 nsew signal input
flabel metal2 s 1398 19200 1454 20000 0 FreeSans 224 90 0 0 resetb
port 9 nsew signal input
flabel metal2 s 12806 19200 12862 20000 0 FreeSans 224 90 0 0 resetb_sync
port 10 nsew signal tristate
flabel metal3 s 19200 11160 20000 11280 0 FreeSans 480 0 0 0 sel2[0]
port 11 nsew signal input
flabel metal3 s 19200 13608 20000 13728 0 FreeSans 480 0 0 0 sel2[1]
port 12 nsew signal input
flabel metal3 s 19200 16056 20000 16176 0 FreeSans 480 0 0 0 sel2[2]
port 13 nsew signal input
flabel metal3 s 19200 3816 20000 3936 0 FreeSans 480 0 0 0 sel[0]
port 14 nsew signal input
flabel metal3 s 19200 6264 20000 6384 0 FreeSans 480 0 0 0 sel[1]
port 15 nsew signal input
flabel metal3 s 19200 8712 20000 8832 0 FreeSans 480 0 0 0 sel[2]
port 16 nsew signal input
flabel metal2 s 9954 19200 10010 20000 0 FreeSans 224 90 0 0 user_clk
port 17 nsew signal tristate
rlabel metal1 9552 17952 9552 17952 0 VGND
rlabel metal1 9522 18496 9522 18496 0 VPWR
rlabel metal1 15502 14246 15502 14246 0 _000_
rlabel metal1 7084 5134 7084 5134 0 _001_
rlabel metal2 11822 11084 11822 11084 0 _002_
rlabel metal1 1932 5338 1932 5338 0 _003_
rlabel metal1 2806 12648 2806 12648 0 _004_
rlabel metal2 2714 14722 2714 14722 0 _005_
rlabel metal1 1012 2618 1012 2618 0 _006_
rlabel metal1 2852 2618 2852 2618 0 _007_
rlabel metal1 5336 2618 5336 2618 0 _008_
rlabel metal2 7590 3910 7590 3910 0 _009_
rlabel metal1 7084 3162 7084 3162 0 _010_
rlabel metal2 9982 4182 9982 4182 0 _011_
rlabel metal1 4002 7208 4002 7208 0 _012_
rlabel metal2 2714 10948 2714 10948 0 _013_
rlabel metal1 4002 9384 4002 9384 0 _014_
rlabel metal1 17020 1530 17020 1530 0 _015_
rlabel metal1 16974 1768 16974 1768 0 _016_
rlabel metal2 13570 14042 13570 14042 0 _017_
rlabel metal1 14582 14926 14582 14926 0 _018_
rlabel metal1 12190 14926 12190 14926 0 _019_
rlabel metal2 14766 3910 14766 3910 0 _020_
rlabel metal1 12650 3162 12650 3162 0 _021_
rlabel metal1 11316 3162 11316 3162 0 _022_
rlabel metal1 11914 7174 11914 7174 0 _023_
rlabel metal2 12650 8670 12650 8670 0 _024_
rlabel metal1 11914 10438 11914 10438 0 _025_
rlabel metal1 7544 12818 7544 12818 0 _026_
rlabel metal1 17756 13294 17756 13294 0 _027_
rlabel metal1 3496 14382 3496 14382 0 _028_
rlabel metal2 1978 4998 1978 4998 0 _029_
rlabel metal1 4784 1734 4784 1734 0 _030_
rlabel metal1 9292 2414 9292 2414 0 _031_
rlabel metal1 17480 1938 17480 1938 0 _032_
rlabel metal2 12926 11900 12926 11900 0 _033_
rlabel metal2 13846 14569 13846 14569 0 _034_
rlabel metal2 14398 2176 14398 2176 0 _035_
rlabel metal1 8188 12614 8188 12614 0 _036_
rlabel metal1 9936 17782 9936 17782 0 _037_
rlabel metal1 17342 12818 17342 12818 0 _038_
rlabel metal1 3864 8330 3864 8330 0 _039_
rlabel metal1 4462 7412 4462 7412 0 _040_
rlabel metal1 2438 10472 2438 10472 0 _041_
rlabel metal2 3174 10812 3174 10812 0 _042_
rlabel metal1 4002 9146 4002 9146 0 _043_
rlabel metal2 4094 9996 4094 9996 0 _044_
rlabel metal2 2162 2720 2162 2720 0 _045_
rlabel metal1 1610 2618 1610 2618 0 _046_
rlabel metal1 3496 1530 3496 1530 0 _047_
rlabel metal2 3634 2278 3634 2278 0 _048_
rlabel metal1 6348 1530 6348 1530 0 _049_
rlabel metal2 6394 2278 6394 2278 0 _050_
rlabel metal1 8832 2618 8832 2618 0 _051_
rlabel metal1 8096 3570 8096 3570 0 _052_
rlabel metal1 7636 1530 7636 1530 0 _053_
rlabel metal1 7544 2074 7544 2074 0 _054_
rlabel metal2 9890 2448 9890 2448 0 _055_
rlabel metal2 10258 3366 10258 3366 0 _056_
rlabel metal1 3128 12818 3128 12818 0 _057_
rlabel metal1 3128 14586 3128 14586 0 _058_
rlabel metal1 12742 7310 12742 7310 0 _059_
rlabel metal1 12742 6426 12742 6426 0 _060_
rlabel metal1 12926 9146 12926 9146 0 _061_
rlabel metal1 13340 8602 13340 8602 0 _062_
rlabel metal2 12834 10370 12834 10370 0 _063_
rlabel metal1 13156 9894 13156 9894 0 _064_
rlabel metal1 14260 13770 14260 13770 0 _065_
rlabel metal2 14306 14246 14306 14246 0 _066_
rlabel metal1 14168 15674 14168 15674 0 _067_
rlabel metal1 14996 14926 14996 14926 0 _068_
rlabel metal1 11684 14586 11684 14586 0 _069_
rlabel metal1 12788 15674 12788 15674 0 _070_
rlabel metal1 14444 2618 14444 2618 0 _071_
rlabel metal1 15456 2618 15456 2618 0 _072_
rlabel metal1 13938 1258 13938 1258 0 _073_
rlabel metal1 13294 2074 13294 2074 0 _074_
rlabel metal1 11822 1530 11822 1530 0 _075_
rlabel metal1 11592 2074 11592 2074 0 _076_
rlabel metal2 17526 2006 17526 2006 0 _077_
rlabel metal2 17342 1496 17342 1496 0 _078_
rlabel metal2 15134 9180 15134 9180 0 _088_
rlabel metal1 5152 14382 5152 14382 0 _089_
rlabel metal2 8142 10302 8142 10302 0 _090_
rlabel metal1 1012 3978 1012 3978 0 _091_
rlabel metal1 3036 4794 3036 4794 0 _092_
rlabel metal2 4554 5474 4554 5474 0 _093_
rlabel metal1 5658 6698 5658 6698 0 _094_
rlabel metal1 1288 7514 1288 7514 0 _095_
rlabel metal2 2070 11492 2070 11492 0 _096_
rlabel metal2 874 9214 874 9214 0 _097_
rlabel metal1 8878 3910 8878 3910 0 _098_
rlabel metal1 6670 5338 6670 5338 0 _099_
rlabel metal2 8786 4760 8786 4760 0 _100_
rlabel metal1 1288 12954 1288 12954 0 _101_
rlabel metal2 874 14654 874 14654 0 _102_
rlabel metal2 874 17442 874 17442 0 _103_
rlabel metal1 4512 17782 4512 17782 0 _104_
rlabel metal2 16606 8228 16606 8228 0 _105_
rlabel metal1 14444 7378 14444 7378 0 _106_
rlabel metal1 10994 12682 10994 12682 0 _107_
rlabel metal1 14582 15130 14582 15130 0 _108_
rlabel metal1 11316 14586 11316 14586 0 _109_
rlabel metal1 14628 11118 14628 11118 0 _110_
rlabel metal1 10803 6630 10803 6630 0 _111_
rlabel metal1 10764 8602 10764 8602 0 _112_
rlabel metal1 10718 10778 10718 10778 0 _113_
rlabel metal1 13938 4794 13938 4794 0 _114_
rlabel metal2 12834 4964 12834 4964 0 _115_
rlabel metal1 11224 4114 11224 4114 0 _116_
rlabel metal2 8142 8772 8142 8772 0 _117_
rlabel metal1 16192 3706 16192 3706 0 _118_
rlabel metal1 16100 2074 16100 2074 0 _119_
rlabel metal1 17388 4250 17388 4250 0 _120_
rlabel metal2 15226 11492 15226 11492 0 _121_
rlabel metal1 5796 6834 5796 6834 0 _122_
rlabel metal1 828 3706 828 3706 0 _123_
rlabel metal2 5198 3910 5198 3910 0 _124_
rlabel metal2 11224 12750 11224 12750 0 _125_
rlabel metal2 11362 14620 11362 14620 0 _126_
rlabel metal1 14122 12750 14122 12750 0 _127_
rlabel metal1 15318 7786 15318 7786 0 _128_
rlabel metal1 16192 14246 16192 14246 0 _129_
rlabel metal2 12558 12682 12558 12682 0 _130_
rlabel metal1 14352 11186 14352 11186 0 _131_
rlabel metal1 14030 11220 14030 11220 0 _132_
rlabel metal1 11316 12954 11316 12954 0 _133_
rlabel metal1 13800 14586 13800 14586 0 _134_
rlabel metal1 13846 14960 13846 14960 0 _135_
rlabel metal1 5566 5644 5566 5644 0 _136_
rlabel metal1 3082 9010 3082 9010 0 _137_
rlabel metal1 6486 4182 6486 4182 0 _138_
rlabel metal1 7728 7786 7728 7786 0 _139_
rlabel metal1 1794 4080 1794 4080 0 _140_
rlabel metal1 5796 3706 5796 3706 0 _141_
rlabel metal1 1817 4250 1817 4250 0 _142_
rlabel metal1 3910 4794 3910 4794 0 _143_
rlabel metal1 5244 5882 5244 5882 0 _144_
rlabel metal1 3404 4250 3404 4250 0 _145_
rlabel metal2 3634 15402 3634 15402 0 _146_
rlabel metal2 8326 6460 8326 6460 0 _147_
rlabel metal1 14490 2992 14490 2992 0 _148_
rlabel metal1 7728 10778 7728 10778 0 _149_
rlabel metal1 7314 10234 7314 10234 0 _150_
rlabel metal2 7130 10608 7130 10608 0 _151_
rlabel metal1 17066 12682 17066 12682 0 _152_
rlabel metal1 16376 12750 16376 12750 0 _153_
rlabel metal1 16054 12716 16054 12716 0 _154_
rlabel metal2 3818 10710 3818 10710 0 _155_
rlabel metal1 3220 8602 3220 8602 0 _156_
rlabel metal2 5566 1564 5566 1564 0 _157_
rlabel metal1 5566 986 5566 986 0 _158_
rlabel metal2 10074 1700 10074 1700 0 _159_
rlabel viali 9981 1870 9981 1870 0 _160_
rlabel metal1 13708 8398 13708 8398 0 _161_
rlabel metal1 12650 10132 12650 10132 0 _162_
rlabel metal2 13754 14688 13754 14688 0 _163_
rlabel metal2 11914 15980 11914 15980 0 _164_
rlabel metal2 11362 1190 11362 1190 0 _165_
rlabel viali 11454 1394 11454 1394 0 _166_
rlabel metal2 15272 9486 15272 9486 0 _167_
rlabel metal1 15042 9588 15042 9588 0 _168_
rlabel metal2 4830 14620 4830 14620 0 _169_
rlabel metal1 4646 14484 4646 14484 0 _170_
rlabel metal2 5566 11764 5566 11764 0 _171_
rlabel metal1 5888 12274 5888 12274 0 _172_
rlabel metal2 6762 11322 6762 11322 0 _173_
rlabel metal1 6302 10132 6302 10132 0 _174_
rlabel metal1 6210 9894 6210 9894 0 _175_
rlabel metal2 6578 10404 6578 10404 0 _176_
rlabel metal1 1334 4114 1334 4114 0 _177_
rlabel metal2 4554 4148 4554 4148 0 _178_
rlabel metal1 8786 4046 8786 4046 0 _179_
rlabel metal1 6854 5168 6854 5168 0 _180_
rlabel metal1 9062 4692 9062 4692 0 _181_
rlabel metal1 1702 16762 1702 16762 0 _182_
rlabel metal1 1288 16694 1288 16694 0 _183_
rlabel metal1 4600 16558 4600 16558 0 _184_
rlabel metal2 17434 6596 17434 6596 0 _185_
rlabel metal1 16928 7514 16928 7514 0 _186_
rlabel metal1 16974 7922 16974 7922 0 _187_
rlabel metal2 17434 10540 17434 10540 0 _188_
rlabel metal2 17526 10608 17526 10608 0 _189_
rlabel metal1 14950 7888 14950 7888 0 _190_
rlabel metal1 15870 6834 15870 6834 0 _191_
rlabel metal1 15364 6698 15364 6698 0 _192_
rlabel metal1 15318 6970 15318 6970 0 _193_
rlabel metal1 11914 12818 11914 12818 0 _194_
rlabel metal1 11684 14382 11684 14382 0 _195_
rlabel metal2 14306 4420 14306 4420 0 _196_
rlabel metal2 12742 4284 12742 4284 0 _197_
rlabel metal1 11408 3706 11408 3706 0 _198_
rlabel metal1 8510 8534 8510 8534 0 _199_
rlabel metal2 8234 9044 8234 9044 0 _200_
rlabel metal1 17618 3978 17618 3978 0 _201_
rlabel metal1 17664 3706 17664 3706 0 _202_
rlabel metal2 11178 15810 11178 15810 0 clknet_0__037_
rlabel metal1 9568 14790 9568 14790 0 clknet_0_divider.out
rlabel metal1 15134 15334 15134 15334 0 clknet_0_divider2.out
rlabel metal1 4370 17102 4370 17102 0 clknet_0_ext_clk
rlabel metal2 7038 17102 7038 17102 0 clknet_0_net11
rlabel metal2 4554 9758 4554 9758 0 clknet_0_pll_clk
rlabel metal1 14352 11526 14352 11526 0 clknet_0_pll_clk90
rlabel metal1 7406 18190 7406 18190 0 clknet_1_0__leaf__037_
rlabel via1 9338 13277 9338 13277 0 clknet_1_0__leaf_divider.out
rlabel metal2 13846 17646 13846 17646 0 clknet_1_0__leaf_divider2.out
rlabel metal2 4094 16150 4094 16150 0 clknet_1_0__leaf_ext_clk
rlabel metal1 1334 6902 1334 6902 0 clknet_1_0__leaf_pll_clk
rlabel metal1 16238 8466 16238 8466 0 clknet_1_0__leaf_pll_clk90
rlabel metal2 10350 17136 10350 17136 0 clknet_1_1__leaf__037_
rlabel metal1 7774 15572 7774 15572 0 clknet_1_1__leaf_divider.out
rlabel metal2 16238 13668 16238 13668 0 clknet_1_1__leaf_divider2.out
rlabel metal2 5658 17680 5658 17680 0 clknet_1_1__leaf_ext_clk
rlabel metal1 13294 16592 13294 16592 0 clknet_1_1__leaf_net11
rlabel metal2 598 13906 598 13906 0 clknet_1_1__leaf_pll_clk
rlabel metal1 14030 13498 14030 13498 0 clknet_1_1__leaf_pll_clk90
rlabel metal1 6440 16490 6440 16490 0 core_clk
rlabel metal2 9522 15198 9522 15198 0 divider.even_0.N\[0\]
rlabel via1 3629 12274 3629 12274 0 divider.even_0.N\[1\]
rlabel metal1 8924 14042 8924 14042 0 divider.even_0.N\[2\]
rlabel metal1 1886 16422 1886 16422 0 divider.even_0.counter\[0\]
rlabel metal1 2001 16490 2001 16490 0 divider.even_0.counter\[1\]
rlabel metal2 2070 17068 2070 17068 0 divider.even_0.counter\[2\]
rlabel via1 7015 14246 7015 14246 0 divider.even_0.out_counter
rlabel metal2 2714 17510 2714 17510 0 divider.even_0.resetb
rlabel metal1 1886 4012 1886 4012 0 divider.odd_0.counter2\[0\]
rlabel metal1 4738 1836 4738 1836 0 divider.odd_0.counter2\[1\]
rlabel metal2 4830 5916 4830 5916 0 divider.odd_0.counter2\[2\]
rlabel metal1 10626 2074 10626 2074 0 divider.odd_0.counter\[0\]
rlabel metal1 9292 1870 9292 1870 0 divider.odd_0.counter\[1\]
rlabel metal1 9154 1904 9154 1904 0 divider.odd_0.counter\[2\]
rlabel metal2 2622 9622 2622 9622 0 divider.odd_0.initial_begin\[0\]
rlabel metal2 1702 11424 1702 11424 0 divider.odd_0.initial_begin\[1\]
rlabel metal1 2116 9486 2116 9486 0 divider.odd_0.initial_begin\[2\]
rlabel metal1 5888 12342 5888 12342 0 divider.odd_0.old_N\[0\]
rlabel metal1 5014 12274 5014 12274 0 divider.odd_0.old_N\[1\]
rlabel metal2 5382 9622 5382 9622 0 divider.odd_0.old_N\[2\]
rlabel metal2 7222 9792 7222 9792 0 divider.odd_0.out_counter
rlabel metal1 6923 7718 6923 7718 0 divider.odd_0.out_counter2
rlabel metal2 9154 9146 9154 9146 0 divider.odd_0.rst_pulse
rlabel metal1 7774 14790 7774 14790 0 divider.out
rlabel metal2 7682 15028 7682 15028 0 divider.syncNp\[0\]
rlabel metal1 9016 11662 9016 11662 0 divider.syncNp\[1\]
rlabel metal1 8004 13498 8004 13498 0 divider.syncNp\[2\]
rlabel metal1 16698 14518 16698 14518 0 divider2.even_0.N\[0\]
rlabel metal1 14168 15606 14168 15606 0 divider2.even_0.N\[1\]
rlabel metal1 15778 16422 15778 16422 0 divider2.even_0.N\[2\]
rlabel metal1 17526 1394 17526 1394 0 divider2.even_0.counter\[0\]
rlabel via1 17342 2499 17342 2499 0 divider2.even_0.counter\[1\]
rlabel metal1 17388 2550 17388 2550 0 divider2.even_0.counter\[2\]
rlabel metal1 17825 8602 17825 8602 0 divider2.even_0.out_counter
rlabel metal2 14306 16609 14306 16609 0 divider2.odd_0.counter2\[0\]
rlabel metal1 16997 17782 16997 17782 0 divider2.odd_0.counter2\[1\]
rlabel metal1 12374 17612 12374 17612 0 divider2.odd_0.counter2\[2\]
rlabel metal1 14766 1394 14766 1394 0 divider2.odd_0.counter\[0\]
rlabel metal1 12650 1836 12650 1836 0 divider2.odd_0.counter\[1\]
rlabel metal1 11178 1326 11178 1326 0 divider2.odd_0.counter\[2\]
rlabel metal1 11914 9588 11914 9588 0 divider2.odd_0.initial_begin\[0\]
rlabel metal1 11914 10064 11914 10064 0 divider2.odd_0.initial_begin\[1\]
rlabel metal2 11546 10778 11546 10778 0 divider2.odd_0.initial_begin\[2\]
rlabel metal2 17986 9860 17986 9860 0 divider2.odd_0.old_N\[0\]
rlabel metal2 17802 11356 17802 11356 0 divider2.odd_0.old_N\[1\]
rlabel metal1 15088 6834 15088 6834 0 divider2.odd_0.old_N\[2\]
rlabel metal1 16376 12274 16376 12274 0 divider2.odd_0.out_counter
rlabel metal1 16077 10982 16077 10982 0 divider2.odd_0.out_counter2
rlabel metal1 15686 13838 15686 13838 0 divider2.odd_0.rst_pulse
rlabel metal1 16652 12954 16652 12954 0 divider2.out
rlabel metal2 17986 14212 17986 14212 0 divider2.syncNp\[0\]
rlabel metal2 17802 16796 17802 16796 0 divider2.syncNp\[1\]
rlabel metal1 16146 17306 16146 17306 0 divider2.syncNp\[2\]
rlabel metal1 3588 18394 3588 18394 0 ext_clk
rlabel metal2 18446 1207 18446 1207 0 ext_clk_sel
rlabel metal1 5750 16218 5750 16218 0 ext_clk_syncd
rlabel metal1 3726 17850 3726 17850 0 ext_clk_syncd_pre
rlabel metal2 18446 18479 18446 18479 0 ext_reset
rlabel metal2 17986 1734 17986 1734 0 net1
rlabel via1 12558 12869 12558 12869 0 net10
rlabel metal1 7728 17782 7728 17782 0 net11
rlabel metal2 12926 17952 12926 17952 0 net12
rlabel metal1 10764 17170 10764 17170 0 net13
rlabel metal1 17894 1802 17894 1802 0 net14
rlabel metal1 17434 1462 17434 1462 0 net15
rlabel metal1 15778 2414 15778 2414 0 net16
rlabel metal1 16146 14348 16146 14348 0 net17
rlabel metal2 5842 2142 5842 2142 0 net18
rlabel metal2 3358 2244 3358 2244 0 net19
rlabel metal1 2162 17068 2162 17068 0 net2
rlabel metal1 2484 2958 2484 2958 0 net20
rlabel metal1 2116 16694 2116 16694 0 net21
rlabel metal2 15962 8738 15962 8738 0 net22
rlabel metal2 12834 11152 12834 11152 0 net23
rlabel metal1 2576 2414 2576 2414 0 net24
rlabel metal1 6440 2414 6440 2414 0 net25
rlabel metal2 2484 16660 2484 16660 0 net26
rlabel metal1 3082 16626 3082 16626 0 net27
rlabel metal1 16613 5814 16613 5814 0 net28
rlabel metal2 17618 14382 17618 14382 0 net29
rlabel metal1 1978 17306 1978 17306 0 net3
rlabel metal1 2944 17578 2944 17578 0 net30
rlabel metal1 6348 17170 6348 17170 0 net31
rlabel metal1 14812 17714 14812 17714 0 net32
rlabel metal2 14766 11356 14766 11356 0 net33
rlabel metal2 9982 9180 9982 9180 0 net34
rlabel metal1 1610 6358 1610 6358 0 net35
rlabel metal1 5244 7922 5244 7922 0 net36
rlabel metal1 1610 11798 1610 11798 0 net37
rlabel metal2 12926 17136 12926 17136 0 net38
rlabel metal2 9890 15878 9890 15878 0 net39
rlabel metal2 2530 17510 2530 17510 0 net4
rlabel metal2 5934 16116 5934 16116 0 net40
rlabel metal1 4416 15946 4416 15946 0 net41
rlabel metal1 15594 16558 15594 16558 0 net42
rlabel metal1 16974 14586 16974 14586 0 net43
rlabel metal1 16652 16082 16652 16082 0 net44
rlabel metal1 6992 14042 6992 14042 0 net45
rlabel metal1 9200 16626 9200 16626 0 net46
rlabel metal1 17388 13906 17388 13906 0 net5
rlabel metal2 18262 16422 18262 16422 0 net6
rlabel metal1 16192 16762 16192 16762 0 net7
rlabel metal1 13662 13872 13662 13872 0 net8
rlabel metal2 15318 6494 15318 6494 0 net9
rlabel metal2 15502 19244 15502 19244 0 pll_clk
rlabel metal1 17112 12410 17112 12410 0 pll_clk90
rlabel metal1 18400 2550 18400 2550 0 pll_clk_sel
rlabel metal1 782 10098 782 10098 0 porb
rlabel metal2 13018 17782 13018 17782 0 reset_delay\[0\]
rlabel metal1 9591 16762 9591 16762 0 reset_delay\[1\]
rlabel metal1 8533 17306 8533 17306 0 reset_delay\[2\]
rlabel metal1 1518 18190 1518 18190 0 resetb
rlabel metal1 13110 17646 13110 17646 0 resetb_sync
rlabel metal2 18446 11373 18446 11373 0 sel2[0]
rlabel metal1 18768 15538 18768 15538 0 sel2[1]
rlabel via2 18446 16133 18446 16133 0 sel2[2]
rlabel metal1 18768 3570 18768 3570 0 sel[0]
rlabel metal2 18446 6579 18446 6579 0 sel[1]
rlabel metal2 18446 8891 18446 8891 0 sel[2]
rlabel metal1 5520 13498 5520 13498 0 use_pll_first
rlabel metal2 8234 17527 8234 17527 0 use_pll_second
rlabel metal1 10672 16490 10672 16490 0 user_clk
rlabel metal2 9982 17340 9982 17340 0 user_clk_buffered
<< properties >>
string FIXED_BBOX 0 0 20000 20000
<< end >>
