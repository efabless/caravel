magic
tech sky130A
timestamp 1636515711
<< error_p >>
rect 18080 2240 18090 2560
rect 3040 1770 3041 2170
rect 3200 1920 3201 2170
<< metal4 >>
tri 4160 5280 4320 5440 se
rect 4320 5280 4480 5440
rect 3360 4160 4000 4320
rect 3200 2880 4000 4160
tri 1600 2560 1920 2880 se
rect 1920 2720 2720 2880
tri 2720 2720 2880 2880 sw
tri 3520 2720 3680 2880 ne
rect 3680 2720 4000 2880
rect 4160 3520 4320 5280
tri 4320 5120 4480 5280 nw
rect 5440 4800 18080 5120
rect 4480 3680 4800 4320
rect 1920 2560 3360 2720
rect 1600 2400 3360 2560
tri 3360 2400 3680 2720 sw
rect 4160 2560 4480 3520
rect 5440 3360 6880 4480
rect 7040 3360 15520 4480
rect 15680 3360 18080 4480
rect 5440 2880 18080 3200
rect 6560 2720 7040 2880
tri 4800 2400 5120 2720 se
rect 5120 2400 8000 2720
rect 8800 2560 18080 2880
rect 1600 2080 8000 2400
rect 1600 1760 2080 2080
rect 3840 1920 4960 2080
rect 16000 1920 17920 2560
<< metal5 >>
tri 4000 4960 4160 5120 se
rect 4160 4960 4960 5120
tri 4960 4960 5120 5120 sw
tri 3040 4800 3200 4960 se
tri 3040 4640 3200 4800 ne
rect 3200 4320 5120 4960
tri 3040 4160 3200 4320 se
rect 3200 4160 3360 4320
tri 2880 3680 3040 3840 se
rect 3040 3680 3200 4160
tri 3200 4000 3360 4160 nw
rect 4000 3680 4480 4320
rect 4800 3680 5120 4320
tri 2240 3520 2400 3680 se
rect 2400 3520 5120 3680
tri 1600 3360 1760 3520 se
rect 1760 3360 5120 3520
rect 1600 2720 5120 3360
rect 5440 4480 18080 5120
rect 5440 3360 7200 4480
rect 7840 4320 8160 4480
rect 8800 4320 9120 4480
rect 7360 4000 8160 4320
rect 8320 4000 9120 4320
tri 9120 4160 9440 4480 nw
tri 9440 4160 9600 4320 se
tri 9600 4160 9760 4320 sw
tri 9760 4160 10080 4480 ne
rect 7840 3840 8160 4000
rect 8800 3840 9120 4000
tri 9280 4000 9440 4160 se
rect 9440 4000 9760 4160
tri 9760 4000 9920 4160 sw
rect 9280 3840 9920 4000
rect 7360 3520 8160 3840
rect 7840 3360 8160 3520
rect 8320 3360 9120 3840
rect 9280 3360 9920 3680
rect 10080 3360 10400 4480
tri 11040 4320 11200 4480 ne
rect 10560 4000 10880 4320
tri 10880 4160 11040 4320 sw
tri 10880 4000 11040 4160 nw
tri 11120 3920 11200 4000 se
tri 11120 3840 11200 3920 ne
rect 10560 3520 10880 3840
tri 10880 3680 11040 3840 sw
tri 10880 3520 11040 3680 nw
tri 11040 3360 11200 3520 se
rect 11200 3360 11520 4480
rect 11680 3520 12480 4480
rect 13120 4320 13440 4480
tri 13440 4320 13600 4480 nw
rect 14240 4320 14560 4480
tri 14560 4320 14720 4480 nw
rect 15360 4320 18080 4480
rect 12640 4000 13440 4320
tri 13600 4160 13760 4320 se
tri 13600 4000 13760 4160 ne
rect 13760 4000 14560 4320
tri 14720 4160 14880 4320 se
tri 14720 4000 14880 4160 ne
rect 14880 4000 18080 4320
rect 13120 3840 13440 4000
tri 13440 3840 13600 4000 sw
tri 14080 3840 14240 4000 ne
rect 14240 3840 14560 4000
tri 14560 3840 14720 4000 sw
tri 15200 3840 15360 4000 ne
rect 12640 3520 13920 3840
tri 13920 3680 14080 3840 sw
tri 13920 3520 14080 3680 nw
rect 14240 3520 15040 3840
tri 15040 3680 15200 3840 sw
tri 15040 3520 15200 3680 nw
rect 12160 3360 12480 3520
rect 13120 3360 13440 3520
tri 14080 3360 14240 3520 se
rect 14240 3360 14560 3520
tri 15200 3360 15360 3520 se
rect 15360 3360 18080 4000
rect 5440 2880 18080 3360
rect 6560 2720 7040 2880
tri 8640 2720 8800 2880 ne
rect 1600 2560 8160 2720
rect 8800 2560 18080 2880
tri 1440 2400 1600 2560 se
rect 1600 2400 2080 2560
tri 2080 2400 2240 2560 nw
tri 3040 2400 3200 2560 ne
rect 1440 1920 2080 2400
tri 1440 1760 1600 1920 ne
rect 1600 1760 2080 1920
tri 2241 2170 2441 2370 se
rect 2441 2170 2841 2370
tri 2841 2170 3041 2370 sw
rect 2241 1770 3041 2170
rect 3200 1920 5760 2560
tri 5760 2400 5920 2560 nw
tri 6720 2400 6880 2560 ne
tri 6880 2400 7040 2560 nw
tri 7680 2400 7840 2560 ne
rect 7840 2400 8160 2560
rect 8960 2400 11680 2560
rect 15615 2400 15935 2560
tri 15935 2400 16095 2560 nw
tri 16640 2400 16800 2560 ne
rect 16800 2400 16960 2560
tri 16960 2400 17120 2560 nw
tri 17695 2400 17855 2560 ne
rect 17855 2400 18080 2560
tri 5996 2170 6196 2370 se
rect 6196 2170 6596 2370
tri 6596 2170 6796 2370 sw
tri 2241 1570 2441 1770 ne
rect 2441 1570 2841 1770
tri 2841 1570 3041 1770 nw
rect 5996 1770 6796 2170
tri 5996 1570 6196 1770 ne
rect 6196 1570 6596 1770
tri 6596 1570 6796 1770 nw
tri 6996 2170 7196 2370 se
rect 7196 2170 7596 2370
tri 7596 2170 7796 2370 sw
rect 6996 1770 7796 2170
rect 8960 2080 9120 2400
tri 15996 2170 16196 2370 se
rect 16196 2170 16596 2370
tri 16596 2170 16796 2370 sw
rect 8800 1920 9280 2080
tri 6996 1570 7196 1770 ne
rect 7196 1570 7596 1770
tri 7596 1570 7796 1770 nw
rect 15996 1770 16796 2170
tri 15996 1570 16196 1770 ne
rect 16196 1570 16596 1770
tri 16596 1570 16796 1770 nw
tri 16961 2170 17161 2370 se
rect 17161 2170 17561 2370
tri 17561 2170 17761 2370 sw
rect 16961 1770 17761 2170
rect 17930 2240 18080 2400
rect 17930 1920 18240 2240
tri 16961 1570 17161 1770 ne
rect 17161 1570 17561 1770
tri 17561 1570 17761 1770 nw
<< fillblock >>
rect 1120 1280 18500 5760
<< end >>
