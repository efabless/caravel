module sky130_ef_sc_hd__decap_12(
    input VPWR,
    input VGND,
    input VPB,
    input VNB
  );

endmodule
