* NGSPICE file created from caravel_clocking.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtn_1 abstract view
.subckt sky130_fd_sc_hd__dfrtn_1 CLK_N D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_4 abstract view
.subckt sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd1_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd1_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

.subckt caravel_clocking VGND VPWR core_clk ext_clk ext_clk_sel ext_reset pll_clk
+ pll_clk90 resetb resetb_sync sel2[0] sel2[1] sel2[2] sel[0] sel[1] sel[2] user_clk
XTAP_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_432_ _417_/A1 hold1/X _349_/S VGND VGND VPWR VPWR _432_/Q sky130_fd_sc_hd__dfrtp_1
X_294_ _294_/A _457_/Q _319_/C VGND VGND VPWR VPWR _294_/Y sky130_fd_sc_hd__nand3_1
X_363_ _448_/Q _363_/B VGND VGND VPWR VPWR _363_/X sky130_fd_sc_hd__xor2_1
XFILLER_12_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_415_ _414_/X _443_/Q _473_/Q VGND VGND VPWR VPWR _415_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_277_ _459_/Q VGND VGND VPWR VPWR _279_/A sky130_fd_sc_hd__inv_2
XFILLER_5_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_1_0_pll_clk clkbuf_0_pll_clk/X VGND VGND VPWR VPWR _417_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_9_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_329_ _438_/Q _422_/Q VGND VGND VPWR VPWR _329_/Y sky130_fd_sc_hd__nor2_1
XFILLER_19_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_431_ _417_/A1 _431_/D _349_/S VGND VGND VPWR VPWR _431_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_13_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_293_ _408_/X _289_/Y _292_/Y VGND VGND VPWR VPWR _458_/D sky130_fd_sc_hd__a21bo_1
X_362_ _447_/Q _446_/Q VGND VGND VPWR VPWR _363_/B sky130_fd_sc_hd__nor2_1
XFILLER_12_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__468__RESET_B _349_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_276_ _276_/A _276_/B VGND VGND VPWR VPWR _461_/D sky130_fd_sc_hd__nand2_1
X_414_ _371_/Y _443_/Q _414_/S VGND VGND VPWR VPWR _414_/X sky130_fd_sc_hd__mux2_1
X_345_ _445_/Q _345_/B VGND VGND VPWR VPWR _445_/D sky130_fd_sc_hd__xnor2_1
X_259_ _256_/Y _261_/A _253_/B VGND VGND VPWR VPWR _260_/B sky130_fd_sc_hd__o21bai_1
XFILLER_0_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_328_ _328_/A _328_/B _420_/Q VGND VGND VPWR VPWR _328_/Y sky130_fd_sc_hd__nand3_1
XFILLER_18_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput10 _399_/X VGND VGND VPWR VPWR core_clk sky130_fd_sc_hd__clkbuf_1
XTAP_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_292_ _294_/A _458_/Q _319_/C VGND VGND VPWR VPWR _292_/Y sky130_fd_sc_hd__nand3_1
X_361_ _447_/Q _446_/Q VGND VGND VPWR VPWR _361_/Y sky130_fd_sc_hd__xnor2_1
X_430_ _417_/A1 _430_/D _349_/S VGND VGND VPWR VPWR _431_/D sky130_fd_sc_hd__dfrtp_1
XFILLER_10_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_275_ _352_/A _275_/B _275_/C VGND VGND VPWR VPWR _276_/B sky130_fd_sc_hd__nand3_1
X_413_ _412_/X _438_/Q _449_/Q VGND VGND VPWR VPWR _413_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_344_ _436_/Q _370_/A _450_/Q VGND VGND VPWR VPWR _345_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_258_ _443_/Q _444_/Q _442_/Q _257_/Y VGND VGND VPWR VPWR _261_/A sky130_fd_sc_hd__o211ai_1
XFILLER_9_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_327_ _421_/Q _437_/Q VGND VGND VPWR VPWR _328_/B sky130_fd_sc_hd__or2b_1
XFILLER_18_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__452__RESET_B _349_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_337__6 _459_/CLK VGND VGND VPWR VPWR _447_/CLK sky130_fd_sc_hd__inv_2
XFILLER_6_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput11 _381_/Y VGND VGND VPWR VPWR resetb_sync sky130_fd_sc_hd__buf_2
XFILLER_16_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_360_ _275_/B _419_/X _235_/A _359_/Y VGND VGND VPWR VPWR _360_/Y sky130_fd_sc_hd__o2bb2ai_2
X_291_ _405_/X _289_/Y _290_/Y VGND VGND VPWR VPWR _459_/D sky130_fd_sc_hd__a21bo_1
XFILLER_12_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_274_ _352_/A _275_/B _275_/C VGND VGND VPWR VPWR _276_/A sky130_fd_sc_hd__a21o_1
X_412_ _363_/X _438_/Q _412_/S VGND VGND VPWR VPWR _412_/X sky130_fd_sc_hd__mux2_1
X_343_ _452_/Q _451_/Q VGND VGND VPWR VPWR _370_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_257_ _468_/Q _467_/Q VGND VGND VPWR VPWR _257_/Y sky130_fd_sc_hd__nor2_1
X_326_ _421_/D _421_/Q VGND VGND VPWR VPWR _328_/A sky130_fd_sc_hd__or2b_1
XFILLER_11_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_309_ _309_/A _309_/B VGND VGND VPWR VPWR _403_/S sky130_fd_sc_hd__nor2_1
XFILLER_6_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__445__SET_B _349_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput12 _400_/X VGND VGND VPWR VPWR user_clk sky130_fd_sc_hd__clkbuf_1
XTAP_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input8_A sel[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_290_ _294_/A _459_/Q _319_/C VGND VGND VPWR VPWR _290_/Y sky130_fd_sc_hd__nand3_1
XFILLER_12_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_0_pll_clk pll_clk VGND VGND VPWR VPWR clkbuf_0_pll_clk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_8_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_273_ _461_/Q VGND VGND VPWR VPWR _275_/C sky130_fd_sc_hd__inv_2
X_411_ _410_/X _436_/Q _449_/Q VGND VGND VPWR VPWR _411_/X sky130_fd_sc_hd__mux2_1
X_342_ _340_/Y _338_/A _341_/Y VGND VGND VPWR VPWR _446_/D sky130_fd_sc_hd__o21ai_1
XFILLER_5_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__446__RESET_B _349_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_256_ _256_/A _256_/B _462_/Q VGND VGND VPWR VPWR _256_/Y sky130_fd_sc_hd__nand3_1
XFILLER_1_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_325_ _325_/A VGND VGND VPWR VPWR _450_/D sky130_fd_sc_hd__clkbuf_1
X_239_ _473_/Q _237_/Y _238_/Y VGND VGND VPWR VPWR _239_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_15_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_348__7 _399_/X VGND VGND VPWR VPWR _427_/CLK sky130_fd_sc_hd__inv_2
XTAP_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_272_ _442_/Q VGND VGND VPWR VPWR _275_/B sky130_fd_sc_hd__inv_2
X_410_ _364_/Y _436_/Q _410_/S VGND VGND VPWR VPWR _410_/X sky130_fd_sc_hd__mux2_1
X_341_ _341_/A _392_/X VGND VGND VPWR VPWR _341_/Y sky130_fd_sc_hd__nand2_1
X_255_ _463_/Q VGND VGND VPWR VPWR _256_/B sky130_fd_sc_hd__inv_2
XFILLER_9_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_324_ _406_/X _450_/Q _436_/Q VGND VGND VPWR VPWR _325_/A sky130_fd_sc_hd__mux2_1
XANTENNA__428__SET_B _349_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_238_ _396_/X VGND VGND VPWR VPWR _238_/Y sky130_fd_sc_hd__inv_2
X_307_ _297_/Y _454_/Q _299_/Y VGND VGND VPWR VPWR _454_/D sky130_fd_sc_hd__a21bo_1
XANTENNA__430__RESET_B _349_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__474__SET_B _349_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_271_ _475_/Q _476_/Q _474_/Q VGND VGND VPWR VPWR _352_/A sky130_fd_sc_hd__nor3b_1
X_340_ _446_/Q VGND VGND VPWR VPWR _340_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_469_ _471_/CLK _469_/D _349_/S VGND VGND VPWR VPWR _469_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_254_ _464_/Q VGND VGND VPWR VPWR _256_/A sky130_fd_sc_hd__inv_2
X_323_ _323_/A VGND VGND VPWR VPWR _451_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__434__SET_B _349_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_237_ _467_/Q _466_/Q VGND VGND VPWR VPWR _237_/Y sky130_fd_sc_hd__nor2_1
X_306_ _302_/B _305_/X _298_/Y VGND VGND VPWR VPWR _455_/D sky130_fd_sc_hd__o21ai_1
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input6_A sel2[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_270_ _268_/Y _266_/A _269_/Y VGND VGND VPWR VPWR _462_/D sky130_fd_sc_hd__o21ai_1
X_468_ _471_/CLK _468_/D _349_/S VGND VGND VPWR VPWR _468_/Q sky130_fd_sc_hd__dfrtn_1
X_399_ _418_/X _357_/Y _431_/Q VGND VGND VPWR VPWR _399_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_322_ _409_/X _451_/Q _436_/Q VGND VGND VPWR VPWR _323_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_253_ _396_/S _253_/B _414_/S VGND VGND VPWR VPWR _260_/A sky130_fd_sc_hd__nand3_1
X_236_ _386_/X _220_/Y _235_/Y VGND VGND VPWR VPWR _469_/D sky130_fd_sc_hd__a21bo_1
X_305_ _454_/Q _305_/B VGND VGND VPWR VPWR _305_/X sky130_fd_sc_hd__and2b_1
XANTENNA__440__SET_B _349_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_1_1_0_pll_clk90 clkbuf_0_pll_clk90/X VGND VGND VPWR VPWR _419_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_219_ _473_/Q VGND VGND VPWR VPWR _261_/B sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_0_pll_clk_A pll_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__449__RESET_B _349_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_398_ _397_/X _443_/Q _473_/Q VGND VGND VPWR VPWR _398_/X sky130_fd_sc_hd__mux2_1
X_467_ _467_/CLK _467_/D _349_/S VGND VGND VPWR VPWR _467_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__464__RESET_B _349_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_252_ _464_/Q _463_/Q _462_/Q VGND VGND VPWR VPWR _414_/S sky130_fd_sc_hd__nor3b_2
X_321_ _452_/Q _321_/B VGND VGND VPWR VPWR _452_/D sky130_fd_sc_hd__xor2_1
Xclkbuf_1_0_0_pll_clk90 clkbuf_0_pll_clk90/X VGND VGND VPWR VPWR _471_/CLK sky130_fd_sc_hd__clkbuf_2
XANTENNA__463__SET_B _349_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_235_ _235_/A _260_/C _469_/Q VGND VGND VPWR VPWR _235_/Y sky130_fd_sc_hd__nand3_1
XFILLER_1_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_218_ _443_/Q _444_/Q _442_/Q VGND VGND VPWR VPWR _250_/A sky130_fd_sc_hd__o21ai_1
Xclkbuf_1_1_0_ext_clk clkbuf_0_ext_clk/X VGND VGND VPWR VPWR _418_/A0 sky130_fd_sc_hd__clkbuf_2
XTAP_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0_pll_clk clkbuf_0_pll_clk/X VGND VGND VPWR VPWR _459_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_8_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_466_ _471_/CLK _466_/D _349_/S VGND VGND VPWR VPWR _466_/Q sky130_fd_sc_hd__dfrtn_1
X_397_ _375_/Y _443_/Q _397_/S VGND VGND VPWR VPWR _397_/X sky130_fd_sc_hd__mux2_1
X_245__1 _471_/CLK VGND VGND VPWR VPWR _467_/CLK sky130_fd_sc_hd__inv_2
XANTENNA__433__RESET_B _349_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_251_ _465_/Q VGND VGND VPWR VPWR _253_/B sky130_fd_sc_hd__inv_2
X_320_ _436_/Q _451_/Q _450_/Q VGND VGND VPWR VPWR _321_/B sky130_fd_sc_hd__nor3_1
X_449_ _417_/A1 _449_/D _349_/S VGND VGND VPWR VPWR _449_/Q sky130_fd_sc_hd__dfrtp_4
X_234_ _398_/X _220_/Y _233_/Y VGND VGND VPWR VPWR _470_/D sky130_fd_sc_hd__a21bo_1
X_303_ _456_/Q _298_/Y _299_/Y _309_/B VGND VGND VPWR VPWR _456_/D sky130_fd_sc_hd__o2bb2ai_1
XFILLER_6_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_217_ _214_/Y _215_/X _226_/C VGND VGND VPWR VPWR _217_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_18_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_396_ _220_/Y _473_/Q _396_/S VGND VGND VPWR VPWR _396_/X sky130_fd_sc_hd__mux2_1
X_465_ _465_/CLK _465_/D _349_/S VGND VGND VPWR VPWR _465_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__473__RESET_B _349_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_250_ _250_/A _250_/B VGND VGND VPWR VPWR _396_/S sky130_fd_sc_hd__nor2_1
XANTENNA_input4_A sel2[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_379_ _475_/Q _474_/Q VGND VGND VPWR VPWR _379_/Y sky130_fd_sc_hd__xnor2_1
X_448_ _459_/CLK _448_/D _349_/S VGND VGND VPWR VPWR _448_/Q sky130_fd_sc_hd__dfrtn_1
X_233_ _235_/A _260_/C _470_/Q VGND VGND VPWR VPWR _233_/Y sky130_fd_sc_hd__nand3_1
X_302_ _302_/A _302_/B VGND VGND VPWR VPWR _309_/B sky130_fd_sc_hd__nand2_1
XFILLER_19_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_216_ _443_/Q _444_/Q _442_/Q VGND VGND VPWR VPWR _226_/C sky130_fd_sc_hd__o21a_1
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_308__5 _459_/CLK VGND VGND VPWR VPWR _453_/CLK sky130_fd_sc_hd__inv_2
X_464_ _471_/CLK _464_/D _349_/S VGND VGND VPWR VPWR _464_/Q sky130_fd_sc_hd__dfrtn_1
X_395_ _394_/X _444_/Q _473_/Q VGND VGND VPWR VPWR _395_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__442__RESET_B _349_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_378_ _474_/Q VGND VGND VPWR VPWR _378_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_1_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_447_ _447_/CLK _447_/D _349_/S VGND VGND VPWR VPWR _447_/Q sky130_fd_sc_hd__dfstp_1
X_232_ _395_/X _220_/Y _231_/Y VGND VGND VPWR VPWR _471_/D sky130_fd_sc_hd__a21bo_1
XFILLER_1_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_301_ _455_/Q VGND VGND VPWR VPWR _302_/B sky130_fd_sc_hd__inv_2
XFILLER_19_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_215_ _425_/Q _444_/Q VGND VGND VPWR VPWR _215_/X sky130_fd_sc_hd__and2_1
XANTENNA__429__SET_B _349_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_394_ _377_/X _444_/Q _397_/S VGND VGND VPWR VPWR _394_/X sky130_fd_sc_hd__mux2_1
X_463_ _463_/CLK _463_/D _349_/S VGND VGND VPWR VPWR _463_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_4_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_377_ _471_/Q _377_/B VGND VGND VPWR VPWR _377_/X sky130_fd_sc_hd__xor2_1
XFILLER_13_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_446_ _459_/CLK _446_/D _349_/S VGND VGND VPWR VPWR _446_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0_ext_clk ext_clk VGND VGND VPWR VPWR clkbuf_0_ext_clk/X sky130_fd_sc_hd__clkbuf_16
X_231_ _235_/A _260_/C _471_/Q VGND VGND VPWR VPWR _231_/Y sky130_fd_sc_hd__nand3_1
X_300_ _456_/Q VGND VGND VPWR VPWR _302_/A sky130_fd_sc_hd__inv_2
X_429_ _429_/CLK _429_/D _349_/S VGND VGND VPWR VPWR _429_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_1_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput1 ext_clk_sel VGND VGND VPWR VPWR _380_/A sky130_fd_sc_hd__clkbuf_1
XTAP_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_214_ _425_/Q _444_/Q VGND VGND VPWR VPWR _214_/Y sky130_fd_sc_hd__nor2_1
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__436__RESET_B _349_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_462_ _471_/CLK _462_/D _349_/S VGND VGND VPWR VPWR _462_/Q sky130_fd_sc_hd__dfrtn_1
X_393_ _443_/Q _378_/Y _416_/S VGND VGND VPWR VPWR _393_/X sky130_fd_sc_hd__mux2_1
XANTENNA__451__RESET_B _349_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_376_ _470_/Q _469_/Q VGND VGND VPWR VPWR _377_/B sky130_fd_sc_hd__nor2_1
X_445_ _417_/A1 _445_/D _349_/S VGND VGND VPWR VPWR _445_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA_input2_A ext_reset VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_230_ _230_/A _260_/C _230_/C VGND VGND VPWR VPWR _472_/D sky130_fd_sc_hd__nand3_1
X_428_ _428_/CLK _429_/Q _349_/S VGND VGND VPWR VPWR _428_/Q sky130_fd_sc_hd__dfstp_1
X_359_ _472_/Q _465_/Q VGND VGND VPWR VPWR _359_/Y sky130_fd_sc_hd__xnor2_1
Xinput2 ext_reset VGND VGND VPWR VPWR _381_/A sky130_fd_sc_hd__clkbuf_1
XTAP_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_213_ _213_/A _213_/B _423_/Q VGND VGND VPWR VPWR _213_/Y sky130_fd_sc_hd__nand3_1
XFILLER_18_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__458__SET_B _349_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__476__RESET_B _349_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_461_ _419_/A1 _461_/D _349_/S VGND VGND VPWR VPWR _461_/Q sky130_fd_sc_hd__dfstp_1
X_392_ _391_/X _436_/Q _449_/Q VGND VGND VPWR VPWR _392_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_444_ _360_/Y _444_/D _349_/S VGND VGND VPWR VPWR _444_/Q sky130_fd_sc_hd__dfrtp_4
X_375_ _470_/Q _469_/Q VGND VGND VPWR VPWR _375_/Y sky130_fd_sc_hd__xnor2_1
X_427_ _427_/CLK _428_/Q _349_/S VGND VGND VPWR VPWR _427_/Q sky130_fd_sc_hd__dfstp_1
X_358_ _443_/Q _444_/Q VGND VGND VPWR VPWR _419_/S sky130_fd_sc_hd__nor2_1
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput3 resetb VGND VGND VPWR VPWR _349_/S sky130_fd_sc_hd__buf_12
XTAP_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_289_ _309_/A _333_/B VGND VGND VPWR VPWR _289_/Y sky130_fd_sc_hd__nand2_2
XTAP_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_212_ _443_/Q _424_/Q VGND VGND VPWR VPWR _213_/B sky130_fd_sc_hd__or2b_1
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_391_ _340_/Y _436_/Q _412_/S VGND VGND VPWR VPWR _391_/X sky130_fd_sc_hd__mux2_1
X_460_ _417_/A1 _460_/D _349_/S VGND VGND VPWR VPWR _460_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_4_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_374_ _469_/Q VGND VGND VPWR VPWR _374_/Y sky130_fd_sc_hd__clkinv_2
X_443_ _360_/Y _443_/D _349_/S VGND VGND VPWR VPWR _443_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_426_ _417_/A1 _426_/D VGND VGND VPWR VPWR hold1/A sky130_fd_sc_hd__dfxtp_1
Xinput4 sel2[0] VGND VGND VPWR VPWR _439_/D sky130_fd_sc_hd__clkbuf_1
XTAP_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_288_ _288_/A _319_/C _288_/C VGND VGND VPWR VPWR _460_/D sky130_fd_sc_hd__nand3_1
X_357_ _294_/A _355_/Y _356_/X VGND VGND VPWR VPWR _357_/Y sky130_fd_sc_hd__o21bai_2
XTAP_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_211_ _424_/Q _443_/Q VGND VGND VPWR VPWR _213_/A sky130_fd_sc_hd__or2b_1
XFILLER_10_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_409_ _438_/Q _369_/Y _409_/S VGND VGND VPWR VPWR _409_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__470__SET_B _349_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_390_ _389_/X _442_/Q _473_/Q VGND VGND VPWR VPWR _390_/X sky130_fd_sc_hd__mux2_1
XTAP_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_442_ _360_/Y _442_/D _349_/S VGND VGND VPWR VPWR _442_/Q sky130_fd_sc_hd__dfrtp_4
X_373_ _464_/Q _373_/B VGND VGND VPWR VPWR _373_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__447__SET_B _349_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput5 sel2[1] VGND VGND VPWR VPWR _440_/D sky130_fd_sc_hd__clkbuf_1
X_425_ _419_/A1 _444_/Q VGND VGND VPWR VPWR _425_/Q sky130_fd_sc_hd__dfxtp_1
X_287_ _294_/A _351_/A _282_/B VGND VGND VPWR VPWR _288_/C sky130_fd_sc_hd__o21bai_1
X_356_ _436_/Q _417_/X VGND VGND VPWR VPWR _356_/X sky130_fd_sc_hd__and2b_2
XANTENNA__439__RESET_B _349_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_210_ _210_/A VGND VGND VPWR VPWR _474_/D sky130_fd_sc_hd__clkbuf_1
X_408_ _407_/X _421_/D _449_/Q VGND VGND VPWR VPWR _408_/X sky130_fd_sc_hd__mux2_1
X_339_ _315_/B _338_/A _338_/Y VGND VGND VPWR VPWR _447_/D sky130_fd_sc_hd__o21ai_1
XFILLER_15_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__454__RESET_B _349_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_441_ _360_/Y _441_/D _349_/S VGND VGND VPWR VPWR _444_/D sky130_fd_sc_hd__dfrtp_1
X_372_ _463_/Q _462_/Q VGND VGND VPWR VPWR _373_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_0_ext_clk clkbuf_0_ext_clk/X VGND VGND VPWR VPWR _349_/A1 sky130_fd_sc_hd__clkbuf_2
X_424_ _471_/CLK _443_/Q VGND VGND VPWR VPWR _424_/Q sky130_fd_sc_hd__dfxtp_1
X_286_ _309_/A VGND VGND VPWR VPWR _294_/A sky130_fd_sc_hd__clkbuf_2
X_355_ _460_/Q _453_/Q VGND VGND VPWR VPWR _355_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_19_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput6 sel2[2] VGND VGND VPWR VPWR _441_/D sky130_fd_sc_hd__clkbuf_1
XTAP_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__453__SET_B _349_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_269_ _269_/A _390_/X VGND VGND VPWR VPWR _269_/Y sky130_fd_sc_hd__nand2_1
X_407_ _365_/Y _437_/Q _410_/S VGND VGND VPWR VPWR _407_/X sky130_fd_sc_hd__mux2_1
X_338_ _338_/A _388_/X VGND VGND VPWR VPWR _338_/Y sky130_fd_sc_hd__nand2_1
XFILLER_15_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_384__13 VGND VGND VPWR VPWR _384__13/HI _429_/D sky130_fd_sc_hd__conb_1
X_346__9 _399_/X VGND VGND VPWR VPWR _429_/CLK sky130_fd_sc_hd__inv_2
X_440_ _360_/Y _440_/D _349_/S VGND VGND VPWR VPWR _443_/D sky130_fd_sc_hd__dfstp_1
XFILLER_13_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_371_ _463_/Q _462_/Q VGND VGND VPWR VPWR _371_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_8_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_423_ _471_/CLK _442_/Q VGND VGND VPWR VPWR _423_/Q sky130_fd_sc_hd__dfxtp_1
X_354_ _438_/Q _421_/D VGND VGND VPWR VPWR _417_/S sky130_fd_sc_hd__nor2_1
X_285_ _438_/Q _437_/Q _436_/Q VGND VGND VPWR VPWR _309_/A sky130_fd_sc_hd__o21ai_2
XFILLER_10_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__448__RESET_B _349_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput7 sel[0] VGND VGND VPWR VPWR _433_/D sky130_fd_sc_hd__clkbuf_1
XTAP_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_268_ _462_/Q VGND VGND VPWR VPWR _268_/Y sky130_fd_sc_hd__inv_2
X_406_ _421_/D _368_/Y _409_/S VGND VGND VPWR VPWR _406_/X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_0_pll_clk90_A pll_clk90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_370_ _370_/A _450_/Q VGND VGND VPWR VPWR _409_/S sky130_fd_sc_hd__nand2_1
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_353_ _353_/A VGND VGND VPWR VPWR _397_/S sky130_fd_sc_hd__inv_2
X_422_ _417_/A1 _438_/Q VGND VGND VPWR VPWR _422_/Q sky130_fd_sc_hd__dfxtp_1
X_284_ _333_/B VGND VGND VPWR VPWR _319_/C sky130_fd_sc_hd__clkbuf_2
XTAP_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput8 sel[1] VGND VGND VPWR VPWR _434_/D sky130_fd_sc_hd__clkbuf_1
X_267_ _256_/B _266_/A _266_/Y VGND VGND VPWR VPWR _463_/D sky130_fd_sc_hd__o21ai_1
X_336_ _315_/A _338_/A _335_/Y VGND VGND VPWR VPWR _448_/D sky130_fd_sc_hd__o21ai_1
X_405_ _404_/X _438_/Q _449_/Q VGND VGND VPWR VPWR _405_/X sky130_fd_sc_hd__mux2_1
X_319_ _319_/A _319_/B _319_/C VGND VGND VPWR VPWR _453_/D sky130_fd_sc_hd__nand3_1
XANTENNA__432__RESET_B _349_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input9_A sel[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_421_ _417_/A1 _421_/D VGND VGND VPWR VPWR _421_/Q sky130_fd_sc_hd__dfxtp_1
X_352_ _352_/A VGND VGND VPWR VPWR _416_/S sky130_fd_sc_hd__inv_2
Xinput9 sel[2] VGND VGND VPWR VPWR _435_/D sky130_fd_sc_hd__clkbuf_1
XTAP_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_283_ _449_/Q VGND VGND VPWR VPWR _333_/B sky130_fd_sc_hd__inv_2
XTAP_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__457__RESET_B _349_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_266_ _266_/A _415_/X VGND VGND VPWR VPWR _266_/Y sky130_fd_sc_hd__nand2_1
X_335_ _338_/A _413_/X VGND VGND VPWR VPWR _335_/Y sky130_fd_sc_hd__nand2_1
X_404_ _367_/X _438_/Q _410_/S VGND VGND VPWR VPWR _404_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_318_ _315_/Y _333_/A _312_/B VGND VGND VPWR VPWR _319_/B sky130_fd_sc_hd__o21bai_1
XFILLER_16_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1 hold1/A VGND VGND VPWR VPWR hold1/X sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA__465__SET_B _349_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_420_ _417_/A1 _436_/Q VGND VGND VPWR VPWR _420_/Q sky130_fd_sc_hd__dfxtp_1
X_351_ _351_/A VGND VGND VPWR VPWR _410_/S sky130_fd_sc_hd__inv_2
X_282_ _351_/A _282_/B _282_/C VGND VGND VPWR VPWR _288_/A sky130_fd_sc_hd__nand3b_1
XFILLER_5_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_334_ _341_/A VGND VGND VPWR VPWR _338_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_403_ _289_/Y _449_/Q _403_/S VGND VGND VPWR VPWR _403_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_248_ _238_/Y _466_/Q _240_/Y VGND VGND VPWR VPWR _466_/D sky130_fd_sc_hd__a21bo_1
XFILLER_14_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_317_ _438_/Q _437_/Q _436_/Q _316_/Y VGND VGND VPWR VPWR _333_/A sky130_fd_sc_hd__o211ai_1
XANTENNA__441__RESET_B _349_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_350_ _350_/A VGND VGND VPWR VPWR _426_/D sky130_fd_sc_hd__buf_1
XFILLER_14_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_281_ _438_/Q _421_/D _436_/Q VGND VGND VPWR VPWR _282_/C sky130_fd_sc_hd__o21a_1
XTAP_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__466__RESET_B _349_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_402_ _401_/X _444_/Q _473_/Q VGND VGND VPWR VPWR _402_/X sky130_fd_sc_hd__mux2_1
X_264_ _256_/A _266_/A _263_/Y VGND VGND VPWR VPWR _464_/D sky130_fd_sc_hd__o21ai_1
XFILLER_2_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_333_ _333_/A _333_/B VGND VGND VPWR VPWR _341_/A sky130_fd_sc_hd__nand2_1
X_247_ _243_/B _246_/X _239_/Y VGND VGND VPWR VPWR _467_/D sky130_fd_sc_hd__o21ai_1
XFILLER_14_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_316_ _456_/Q _455_/Q VGND VGND VPWR VPWR _316_/Y sky130_fd_sc_hd__nor2_1
X_249__2 _471_/CLK VGND VGND VPWR VPWR _465_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_280_ _460_/Q VGND VGND VPWR VPWR _282_/B sky130_fd_sc_hd__inv_2
XANTENNA_input7_A sel[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__435__RESET_B _349_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_263_ _266_/A _402_/X VGND VGND VPWR VPWR _263_/Y sky130_fd_sc_hd__nand2_1
X_401_ _373_/X _444_/Q _414_/S VGND VGND VPWR VPWR _401_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_332_ _328_/Y _331_/Y _289_/Y VGND VGND VPWR VPWR _449_/D sky130_fd_sc_hd__o21a_1
XFILLER_17_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_246_ _466_/Q _396_/X VGND VGND VPWR VPWR _246_/X sky130_fd_sc_hd__and2b_1
XFILLER_14_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_315_ _315_/A _315_/B _446_/Q VGND VGND VPWR VPWR _315_/Y sky130_fd_sc_hd__nand3_1
X_229_ _235_/A _353_/A _226_/B VGND VGND VPWR VPWR _230_/C sky130_fd_sc_hd__o21bai_1
XFILLER_6_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_400_ _418_/X _360_/Y _431_/Q VGND VGND VPWR VPWR _400_/X sky130_fd_sc_hd__mux2_1
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_262_ _269_/A VGND VGND VPWR VPWR _266_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__475__RESET_B _349_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_331_ _329_/Y _330_/X _282_/C VGND VGND VPWR VPWR _331_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_2_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_314_ _447_/Q VGND VGND VPWR VPWR _315_/B sky130_fd_sc_hd__inv_2
XFILLER_11_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_228_ _250_/A VGND VGND VPWR VPWR _235_/A sky130_fd_sc_hd__clkbuf_2
X_265__3 _471_/CLK VGND VGND VPWR VPWR _463_/CLK sky130_fd_sc_hd__inv_2
XANTENNA__460__SET_B _349_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_476_ _419_/A1 _476_/D _349_/S VGND VGND VPWR VPWR _476_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__444__RESET_B _349_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_261_ _261_/A _261_/B VGND VGND VPWR VPWR _269_/A sky130_fd_sc_hd__nand2_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_330_ _438_/Q _422_/Q VGND VGND VPWR VPWR _330_/X sky130_fd_sc_hd__and2_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__437__SET_B _349_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_459_ _459_/CLK _459_/D _349_/S VGND VGND VPWR VPWR _459_/Q sky130_fd_sc_hd__dfrtp_1
X_244_ _468_/Q _239_/Y _240_/Y _250_/B VGND VGND VPWR VPWR _468_/D sky130_fd_sc_hd__o2bb2ai_1
X_313_ _448_/Q VGND VGND VPWR VPWR _315_/A sky130_fd_sc_hd__inv_2
X_227_ _261_/B VGND VGND VPWR VPWR _260_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_10_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__469__RESET_B _349_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_475_ _419_/A1 _475_/D _349_/S VGND VGND VPWR VPWR _475_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input5_A sel2[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_260_ _260_/A _260_/B _260_/C VGND VGND VPWR VPWR _465_/D sky130_fd_sc_hd__nand3_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_389_ _268_/Y _442_/Q _414_/S VGND VGND VPWR VPWR _389_/X sky130_fd_sc_hd__mux2_1
X_458_ _459_/CLK _458_/D _349_/S VGND VGND VPWR VPWR _458_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__443__SET_B _349_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_243_ _243_/A _243_/B VGND VGND VPWR VPWR _250_/B sky130_fd_sc_hd__nand2_1
XFILLER_11_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_312_ _312_/A _312_/B _412_/S VGND VGND VPWR VPWR _319_/A sky130_fd_sc_hd__nand3_1
XFILLER_9_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_226_ _353_/A _226_/B _226_/C VGND VGND VPWR VPWR _230_/A sky130_fd_sc_hd__nand3b_1
XFILLER_6_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_209_ _393_/X _474_/Q _442_/Q VGND VGND VPWR VPWR _210_/A sky130_fd_sc_hd__mux2_1
XANTENNA__438__RESET_B _349_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_474_ _419_/A1 _474_/D _349_/S VGND VGND VPWR VPWR _474_/Q sky130_fd_sc_hd__dfstp_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_457_ _417_/A1 _457_/D _349_/S VGND VGND VPWR VPWR _457_/Q sky130_fd_sc_hd__dfrtp_2
X_388_ _387_/X _437_/Q _449_/Q VGND VGND VPWR VPWR _388_/X sky130_fd_sc_hd__mux2_1
XTAP_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_242_ _467_/Q VGND VGND VPWR VPWR _243_/B sky130_fd_sc_hd__inv_2
X_311_ _448_/Q _447_/Q _446_/Q VGND VGND VPWR VPWR _412_/S sky130_fd_sc_hd__nor3b_2
XFILLER_9_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_225_ _472_/Q VGND VGND VPWR VPWR _226_/B sky130_fd_sc_hd__inv_2
XFILLER_17_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_208_ _208_/A VGND VGND VPWR VPWR _475_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_473_ _419_/A1 _473_/D _349_/S VGND VGND VPWR VPWR _473_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__472__SET_B _349_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_387_ _361_/Y _437_/Q _412_/S VGND VGND VPWR VPWR _387_/X sky130_fd_sc_hd__mux2_1
X_456_ _459_/CLK _456_/D _349_/S VGND VGND VPWR VPWR _456_/Q sky130_fd_sc_hd__dfrtn_1
XTAP_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_310_ _453_/Q VGND VGND VPWR VPWR _312_/B sky130_fd_sc_hd__inv_2
X_241_ _468_/Q VGND VGND VPWR VPWR _243_/A sky130_fd_sc_hd__inv_2
X_439_ _360_/Y _439_/D _349_/S VGND VGND VPWR VPWR _442_/D sky130_fd_sc_hd__dfrtp_1
X_224_ _224_/A _224_/B _469_/Q VGND VGND VPWR VPWR _353_/A sky130_fd_sc_hd__nand3_1
XFILLER_10_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_207_ _416_/X _475_/Q _442_/Q VGND VGND VPWR VPWR _208_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_347__8 _399_/X VGND VGND VPWR VPWR _428_/CLK sky130_fd_sc_hd__inv_2
X_472_ _419_/A1 _472_/D _349_/S VGND VGND VPWR VPWR _472_/Q sky130_fd_sc_hd__dfstp_1
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_386_ _385_/X _442_/Q _473_/Q VGND VGND VPWR VPWR _386_/X sky130_fd_sc_hd__mux2_1
XANTENNA__462__RESET_B _349_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_455_ _455_/CLK _455_/D _349_/S VGND VGND VPWR VPWR _455_/Q sky130_fd_sc_hd__dfstp_1
XTAP_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input3_A resetb VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_240_ _466_/Q _261_/B _396_/X VGND VGND VPWR VPWR _240_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_14_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_369_ _451_/Q _450_/Q VGND VGND VPWR VPWR _369_/Y sky130_fd_sc_hd__xnor2_1
X_438_ _357_/Y _438_/D _349_/S VGND VGND VPWR VPWR _438_/Q sky130_fd_sc_hd__dfrtp_4
X_223_ _470_/Q VGND VGND VPWR VPWR _224_/B sky130_fd_sc_hd__inv_2
XFILLER_8_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__455__SET_B _349_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_471_ _471_/CLK _471_/D _349_/S VGND VGND VPWR VPWR _471_/Q sky130_fd_sc_hd__dfrtp_1
Xsplit2 _437_/Q VGND VGND VPWR VPWR _421_/D sky130_fd_sc_hd__clkbuf_2
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__431__RESET_B _349_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_385_ _374_/Y _442_/Q _397_/S VGND VGND VPWR VPWR _385_/X sky130_fd_sc_hd__mux2_1
X_454_ _459_/CLK _454_/D _349_/S VGND VGND VPWR VPWR _454_/Q sky130_fd_sc_hd__dfrtn_1
XTAP_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_299_ _454_/Q _333_/B _403_/X VGND VGND VPWR VPWR _299_/Y sky130_fd_sc_hd__nand3b_1
X_437_ _357_/Y _437_/D _349_/S VGND VGND VPWR VPWR _437_/Q sky130_fd_sc_hd__dfstp_4
X_368_ _450_/Q VGND VGND VPWR VPWR _368_/Y sky130_fd_sc_hd__clkinv_2
X_222_ _471_/Q VGND VGND VPWR VPWR _224_/A sky130_fd_sc_hd__inv_2
XFILLER_10_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_pll_clk90 pll_clk90 VGND VGND VPWR VPWR clkbuf_0_pll_clk90/X sky130_fd_sc_hd__clkbuf_16
XANTENNA__456__RESET_B _349_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__461__SET_B _349_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_470_ _471_/CLK _470_/D _349_/S VGND VGND VPWR VPWR _470_/Q sky130_fd_sc_hd__dfstp_1
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_453_ _453_/CLK _453_/D _349_/S VGND VGND VPWR VPWR _453_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__471__RESET_B _349_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_0_ext_clk_A ext_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_367_ _459_/Q _367_/B VGND VGND VPWR VPWR _367_/X sky130_fd_sc_hd__xor2_1
X_436_ _357_/Y _436_/D _349_/S VGND VGND VPWR VPWR _436_/Q sky130_fd_sc_hd__dfrtp_4
X_298_ _449_/Q _296_/Y _297_/Y VGND VGND VPWR VPWR _298_/Y sky130_fd_sc_hd__o21bai_1
Xrebuffer3 _403_/X VGND VGND VPWR VPWR _305_/B sky130_fd_sc_hd__buf_2
X_221_ _213_/Y _217_/Y _220_/Y VGND VGND VPWR VPWR _473_/D sky130_fd_sc_hd__o21a_1
XFILLER_12_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_419_ _461_/Q _419_/A1 _419_/S VGND VGND VPWR VPWR _419_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_383_ _476_/Q _383_/B VGND VGND VPWR VPWR _476_/D sky130_fd_sc_hd__xor2_1
X_452_ _417_/A1 _452_/D _349_/S VGND VGND VPWR VPWR _452_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_15_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_435_ _357_/Y _435_/D _349_/S VGND VGND VPWR VPWR _438_/D sky130_fd_sc_hd__dfrtp_1
X_366_ _458_/Q _457_/Q VGND VGND VPWR VPWR _367_/B sky130_fd_sc_hd__nor2_1
X_297_ _305_/B VGND VGND VPWR VPWR _297_/Y sky130_fd_sc_hd__inv_2
Xrebuffer4 _403_/S VGND VGND VPWR VPWR _312_/A sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_3_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_220_ _250_/A _261_/B VGND VGND VPWR VPWR _220_/Y sky130_fd_sc_hd__nand2_2
XFILLER_10_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input1_A ext_clk_sel VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_304__4 _459_/CLK VGND VGND VPWR VPWR _455_/CLK sky130_fd_sc_hd__inv_2
X_418_ _418_/A0 _432_/Q _431_/D VGND VGND VPWR VPWR _418_/X sky130_fd_sc_hd__mux2_1
X_349_ hold1/A _349_/A1 _349_/S VGND VGND VPWR VPWR _350_/A sky130_fd_sc_hd__mux2_2
XFILLER_0_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_382_ _475_/Q _442_/Q _474_/Q VGND VGND VPWR VPWR _383_/B sky130_fd_sc_hd__nor3_1
X_451_ _417_/A1 _451_/D _349_/S VGND VGND VPWR VPWR _451_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_365_ _458_/Q _457_/Q VGND VGND VPWR VPWR _365_/Y sky130_fd_sc_hd__xnor2_1
X_296_ _455_/Q _454_/Q VGND VGND VPWR VPWR _296_/Y sky130_fd_sc_hd__nor2_1
X_434_ _357_/Y _434_/D _349_/S VGND VGND VPWR VPWR _437_/D sky130_fd_sc_hd__dfstp_1
XFILLER_3_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__467__SET_B _349_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_279_ _279_/A _279_/B _457_/Q VGND VGND VPWR VPWR _351_/A sky130_fd_sc_hd__nand3_1
X_417_ _445_/Q _417_/A1 _417_/S VGND VGND VPWR VPWR _417_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__450__SET_B _349_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_381_ _381_/A _427_/Q VGND VGND VPWR VPWR _381_/Y sky130_fd_sc_hd__nor2_1
XFILLER_17_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_450_ _459_/CLK _450_/D _349_/S VGND VGND VPWR VPWR _450_/Q sky130_fd_sc_hd__dfstp_2
XTAP_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__427__SET_B _349_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__349__S _349_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_433_ _357_/Y _433_/D _349_/S VGND VGND VPWR VPWR _436_/D sky130_fd_sc_hd__dfrtp_1
XFILLER_13_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_364_ _457_/Q VGND VGND VPWR VPWR _364_/Y sky130_fd_sc_hd__clkinv_2
X_295_ _411_/X _289_/Y _294_/Y VGND VGND VPWR VPWR _457_/D sky130_fd_sc_hd__a21bo_1
XFILLER_12_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_416_ _444_/Q _379_/Y _416_/S VGND VGND VPWR VPWR _416_/X sky130_fd_sc_hd__mux2_1
X_278_ _458_/Q VGND VGND VPWR VPWR _279_/B sky130_fd_sc_hd__inv_2
XANTENNA__459__RESET_B _349_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_380_ _380_/A VGND VGND VPWR VPWR _430_/D sky130_fd_sc_hd__inv_2
XFILLER_16_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

