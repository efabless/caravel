magic
tech sky130A
magscale 1 2
timestamp 1637274818
<< nwell >>
rect -38 8965 18898 9531
rect -38 7877 18898 8443
rect -38 6789 18898 7355
rect -38 5701 18898 6267
rect -38 4613 18898 5179
rect -38 3525 18898 4091
rect -38 2437 18898 3003
rect -38 1349 18898 1915
rect -38 261 18898 827
<< pwell >>
rect 29 -17 63 17
rect 305 -17 339 17
rect 1409 -17 1443 17
rect 2512 -11 2536 11
rect 2697 -17 2731 17
rect 3801 -17 3835 17
rect 4905 -17 4939 17
rect 5273 -17 5307 17
rect 6377 -17 6411 17
rect 7115 -10 7147 12
rect 7481 -17 7515 17
rect 7575 -10 7607 12
rect 7849 -17 7883 17
rect 8401 -17 8435 17
rect 10240 -11 10264 11
rect 10425 -17 10459 17
rect 11070 -17 11104 17
rect 11345 -17 11379 17
rect 12449 -17 12483 17
rect 12816 -11 12840 11
rect 13001 -17 13035 17
rect 14105 -17 14139 17
rect 15209 -17 15243 17
rect 15577 -17 15611 17
rect 16681 -17 16715 17
rect 16957 -17 16991 17
rect 17601 -17 17635 17
rect 17968 -11 17992 11
rect 18155 -10 18187 12
rect 18521 -17 18555 17
rect 18797 -17 18831 17
<< obsli1 >>
rect 0 0 19015 9809
rect 0 -17 18860 0
<< obsm1 >>
rect 0 0 19027 9840
rect 0 -48 18860 0
<< metal2 >>
rect 1398 11200 1454 12000
rect 4250 11200 4306 12000
rect 7102 11200 7158 12000
rect 9954 11200 10010 12000
rect 12806 11200 12862 12000
rect 15658 11200 15714 12000
rect 18510 11200 18566 12000
<< obsm2 >>
rect 388 11144 1342 11257
rect 1510 11144 4194 11257
rect 4362 11144 7046 11257
rect 7214 11144 9898 11257
rect 10066 11144 12750 11257
rect 12918 11144 15602 11257
rect 15770 11144 18454 11257
rect 18622 11144 18658 11257
rect 388 0 18658 11144
rect 6144 -48 6452 0
rect 12443 -48 12751 0
<< metal3 >>
rect 19200 11160 20000 11280
rect 19200 9664 20000 9784
rect 19200 8168 20000 8288
rect 19200 6672 20000 6792
rect 19200 5176 20000 5296
rect 19200 3680 20000 3800
rect 19200 2184 20000 2304
rect 19200 688 20000 808
<< obsm3 >>
rect 2989 11080 19120 11253
rect 2989 9864 19200 11080
rect 2989 9584 19120 9864
rect 2989 8368 19200 9584
rect 2989 8088 19120 8368
rect 2989 6872 19200 8088
rect 2989 6592 19120 6872
rect 2989 5376 19200 6592
rect 2989 5096 19120 5376
rect 2989 3880 19200 5096
rect 2989 3600 19120 3880
rect 2989 2384 19200 3600
rect 2989 2104 19120 2384
rect 2989 888 19200 2104
rect 2989 608 19120 888
rect 2989 0 19200 608
rect 6138 -33 6458 0
rect 12437 -33 12757 0
<< metal4 >>
rect 2989 -48 3309 9840
rect 6138 -48 6458 9840
rect 9287 -48 9607 9840
rect 12437 -48 12757 9840
rect 15586 -48 15906 9840
<< obsm4 >>
rect 9607 -48 9608 9840
<< metal5 >>
rect 0 7978 18860 8298
rect 0 6341 18860 6661
rect 0 4704 18860 5024
rect 0 3066 18860 3386
rect 0 1429 18860 1749
<< labels >>
rlabel metal5 s 0 3066 18860 3386 6 VGND
port 1 nsew ground input
rlabel metal5 s 0 6341 18860 6661 6 VGND
port 1 nsew ground input
rlabel metal4 s 6138 -48 6458 9840 6 VGND
port 1 nsew ground input
rlabel metal4 s 12437 -48 12757 9840 6 VGND
port 1 nsew ground input
rlabel metal5 s 0 1429 18860 1749 6 VPWR
port 2 nsew power input
rlabel metal5 s 0 4704 18860 5024 6 VPWR
port 2 nsew power input
rlabel metal5 s 0 7978 18860 8298 6 VPWR
port 2 nsew power input
rlabel metal4 s 2989 -48 3309 9840 6 VPWR
port 2 nsew power input
rlabel metal4 s 9287 -48 9607 9840 6 VPWR
port 2 nsew power input
rlabel metal4 s 15586 -48 15906 9840 6 VPWR
port 2 nsew power input
rlabel metal2 s 7102 11200 7158 12000 6 core_clk
port 3 nsew signal output
rlabel metal2 s 4250 11200 4306 12000 6 ext_clk
port 4 nsew signal input
rlabel metal3 s 19200 688 20000 808 6 ext_clk_sel
port 5 nsew signal input
rlabel metal3 s 19200 11160 20000 11280 6 ext_reset
port 6 nsew signal input
rlabel metal2 s 15658 11200 15714 12000 6 pll_clk
port 7 nsew signal input
rlabel metal2 s 18510 11200 18566 12000 6 pll_clk90
port 8 nsew signal input
rlabel metal2 s 1398 11200 1454 12000 6 resetb
port 9 nsew signal input
rlabel metal2 s 12806 11200 12862 12000 6 resetb_sync
port 10 nsew signal output
rlabel metal3 s 19200 6672 20000 6792 6 sel2[0]
port 11 nsew signal input
rlabel metal3 s 19200 8168 20000 8288 6 sel2[1]
port 12 nsew signal input
rlabel metal3 s 19200 9664 20000 9784 6 sel2[2]
port 13 nsew signal input
rlabel metal3 s 19200 2184 20000 2304 6 sel[0]
port 14 nsew signal input
rlabel metal3 s 19200 3680 20000 3800 6 sel[1]
port 15 nsew signal input
rlabel metal3 s 19200 5176 20000 5296 6 sel[2]
port 16 nsew signal input
rlabel metal2 s 9954 11200 10010 12000 6 user_clk
port 17 nsew signal output
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 20000 12000
string LEFview TRUE
string GDS_FILE /home/ma/ef/caravel_openframe/openlane/caravel_clocking/runs/caravel_clocking/results/magic/caravel_clocking.gds
string GDS_END 1020802
string GDS_START 357236
<< end >>

