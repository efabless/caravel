magic
tech sky130A
magscale 1 2
timestamp 1695675344
<< checkpaint >>
rect 674054 99659 678702 116976
<< metal1 >>
rect 675778 116066 675830 116072
rect 675778 115848 675830 115854
rect 675682 113513 675734 115709
rect 675586 112736 675638 112742
rect 675586 112558 675638 112564
rect 675588 108330 675636 112558
rect 675682 108981 675734 113341
rect 675586 108324 675638 108330
rect 675586 108146 675638 108152
rect 675588 100462 675636 108146
rect 675586 100456 675638 100462
rect 675586 100278 675638 100284
rect 675682 99896 675734 108797
rect 675780 102343 675828 115848
rect 675874 109636 675926 109642
rect 675874 109458 675926 109464
rect 675778 102337 675830 102343
rect 675778 102119 675830 102125
rect 675876 101791 675924 109458
rect 677378 103462 677384 103674
rect 677436 103514 677442 103674
rect 677436 103462 677658 103514
rect 675874 101785 675926 101791
rect 675874 101567 675926 101573
rect 675876 101554 675924 101567
<< via1 >>
rect 675778 115854 675830 116066
rect 675682 113341 675734 113513
rect 675586 112564 675638 112736
rect 675682 108797 675734 108981
rect 675586 108152 675638 108324
rect 675586 100284 675638 100456
rect 675874 109464 675926 109636
rect 675778 102125 675830 102337
rect 677384 103462 677436 103674
rect 675874 101573 675926 101785
<< metal2 >>
rect 675772 115854 675778 116066
rect 675830 116064 675836 116066
rect 676699 116064 676708 116230
rect 675830 116016 676708 116064
rect 675830 115854 675836 116016
rect 676699 116010 676708 116016
rect 676768 116010 676777 116230
rect 677187 115272 677196 115332
rect 677416 115325 677425 115332
rect 677416 115279 677607 115325
rect 677416 115272 677425 115279
rect 677189 114863 677198 114923
rect 677418 114916 677427 114923
rect 677418 114870 677607 114916
rect 677418 114863 677427 114870
rect 677186 114718 677195 114778
rect 677415 114774 677424 114778
rect 677415 114722 677607 114774
rect 677415 114718 677424 114722
rect 675676 113341 675682 113513
rect 675734 113453 675740 113513
rect 675734 113449 676020 113453
rect 675734 113397 677607 113449
rect 675734 113341 675740 113397
rect 675580 112736 677607 112738
rect 675580 112564 675586 112736
rect 675638 112686 677607 112736
rect 675638 112682 677262 112686
rect 675638 112564 675644 112682
rect 677220 111689 677290 111694
rect 677216 111469 677225 111689
rect 677285 111529 677295 111689
rect 677285 111477 677607 111529
rect 677285 111469 677294 111477
rect 677220 111464 677290 111469
rect 676980 110620 676989 110840
rect 677049 110680 677058 110840
rect 677049 110628 677607 110680
rect 677049 110620 677058 110628
rect 676758 110243 676767 110463
rect 676827 110302 676836 110463
rect 676827 110250 677607 110302
rect 676827 110243 676836 110250
rect 676543 109796 676552 110016
rect 676612 109850 676621 110016
rect 676612 109798 677607 109850
rect 676612 109796 676621 109798
rect 675868 109636 677607 109637
rect 675868 109464 675874 109636
rect 675926 109585 677607 109636
rect 675926 109581 677286 109585
rect 675926 109464 675932 109581
rect 675676 108797 675682 108981
rect 675734 108912 675740 108981
rect 675734 108908 677272 108912
rect 675734 108856 677607 108908
rect 675734 108797 675740 108856
rect 675580 108324 677286 108326
rect 675580 108152 675586 108324
rect 675638 108322 677286 108324
rect 675638 108270 677607 108322
rect 675638 108152 675644 108270
rect 677373 106895 677382 107115
rect 677442 106951 677451 107115
rect 677442 106899 677616 106951
rect 677442 106895 677451 106899
rect 677379 106510 677439 106514
rect 677374 106505 677444 106510
rect 677374 106285 677379 106505
rect 677439 106285 677444 106505
rect 677374 106275 677444 106285
rect 677384 106029 677436 106275
rect 677384 105977 677607 106029
rect 677380 105865 677440 105874
rect 677380 105636 677440 105645
rect 677384 103674 677436 105636
rect 677384 103456 677436 103462
rect 676885 102577 676894 102797
rect 676954 102633 676963 102797
rect 676954 102581 677607 102633
rect 676954 102577 676963 102581
rect 675773 102337 675835 102343
rect 675773 102125 675778 102337
rect 675830 102179 675835 102337
rect 676285 102179 676363 102189
rect 675830 102125 676291 102179
rect 675773 102123 676291 102125
rect 675773 102118 675835 102123
rect 676285 101963 676291 102123
rect 676357 101963 676363 102179
rect 676285 101954 676363 101963
rect 675870 101785 675931 101792
rect 675870 101573 675874 101785
rect 675926 101627 675931 101785
rect 675926 101573 676249 101627
rect 675870 101571 676249 101573
rect 675870 101566 675931 101571
rect 675580 100284 675586 100456
rect 675638 100339 675644 100456
rect 675638 100284 676031 100339
rect 675580 100283 676031 100284
rect 675991 100057 676031 100283
rect 676209 100259 676249 101571
rect 676473 100422 676482 100642
rect 676542 100478 676551 100642
rect 676653 100616 676662 100904
rect 676790 100744 676800 100904
rect 676790 100616 677607 100744
rect 676542 100426 677607 100478
rect 676542 100422 676551 100426
rect 676209 100219 677607 100259
rect 675991 100017 677607 100057
<< via2 >>
rect 676708 116010 676768 116230
rect 677196 115272 677416 115332
rect 677198 114863 677418 114923
rect 677195 114718 677415 114778
rect 677225 111469 677285 111689
rect 676989 110620 677049 110840
rect 676767 110243 676827 110463
rect 676552 109796 676612 110016
rect 677382 106895 677442 107115
rect 677379 106285 677439 106505
rect 677380 105645 677440 105865
rect 676894 102577 676954 102797
rect 676291 101963 676357 102179
rect 676482 100422 676542 100642
rect 676662 100616 676790 100904
<< metal3 >>
rect 676708 116235 676768 117452
rect 676703 116230 676773 116235
rect 676703 116010 676708 116230
rect 676768 116010 676773 116230
rect 676703 116005 676773 116010
rect 677177 115796 677607 115920
rect 677177 115711 677247 115796
rect 675407 115641 677247 115711
rect 677191 115332 677421 115337
rect 675942 115272 677196 115332
rect 677416 115272 677421 115332
rect 675942 115159 676002 115272
rect 677191 115267 677421 115272
rect 675407 115089 676002 115159
rect 677193 114923 677423 114928
rect 676200 114863 677198 114923
rect 677418 114863 677423 114923
rect 676200 114515 676260 114863
rect 677193 114858 677423 114863
rect 677190 114778 677420 114783
rect 675407 114445 676260 114515
rect 676326 114718 677195 114778
rect 677415 114718 677420 114778
rect 676326 113871 676386 114718
rect 677190 114713 677420 114718
rect 675407 113801 676386 113871
rect 675407 111961 677290 112031
rect 677220 111689 677290 111961
rect 675407 111409 677054 111479
rect 677220 111469 677225 111689
rect 677285 111469 677290 111689
rect 677220 111464 677290 111469
rect 676984 110840 677054 111409
rect 675407 110765 676832 110835
rect 676762 110463 676832 110765
rect 676984 110620 676989 110840
rect 677049 110620 677054 110840
rect 676984 110615 677054 110620
rect 676762 110243 676767 110463
rect 676827 110243 676832 110463
rect 676762 110238 676832 110243
rect 675407 110121 676617 110191
rect 676547 110016 676617 110121
rect 676547 109796 676552 110016
rect 676612 109796 676617 110016
rect 676547 109790 676617 109796
rect 675407 107637 677442 107707
rect 675407 107085 677250 107155
rect 677382 107120 677442 107637
rect 677180 106827 677250 107085
rect 677377 107115 677447 107120
rect 677377 106895 677382 107115
rect 677442 106895 677447 107115
rect 677377 106890 677447 106895
rect 677180 106761 677616 106827
rect 675407 106510 677379 106511
rect 675407 106505 677444 106510
rect 675407 106441 677379 106505
rect 677374 106285 677379 106441
rect 677439 106285 677444 106505
rect 677374 106280 677444 106285
rect 677375 105866 677445 105870
rect 675407 105865 677445 105866
rect 675407 105806 677380 105865
rect 675407 105796 675887 105806
rect 677375 105645 677380 105806
rect 677440 105645 677445 105865
rect 677375 105640 677445 105645
rect 675407 105172 677260 105386
rect 675407 104601 676955 104671
rect 675407 103375 676790 103503
rect 675407 102761 676542 102831
rect 676286 102179 676362 102187
rect 676286 101963 676291 102179
rect 676357 101963 676362 102179
rect 676286 101958 676362 101963
rect 675407 100921 676153 100991
rect 676087 100152 676153 100921
rect 676291 100284 676357 101958
rect 676482 100647 676542 102761
rect 676662 100909 676790 103375
rect 676894 102802 676954 104601
rect 677046 103436 677260 105172
rect 677046 103222 677607 103436
rect 676889 102797 676959 102802
rect 676889 102577 676894 102797
rect 676954 102577 676959 102797
rect 676889 102572 676959 102577
rect 676657 100904 676795 100909
rect 676477 100642 676547 100647
rect 676477 100422 676482 100642
rect 676542 100422 676547 100642
rect 676657 100616 676662 100904
rect 676790 100616 676795 100904
rect 676657 100611 676795 100616
rect 676477 100417 676547 100422
rect 676291 100218 677607 100284
rect 676087 100086 677607 100152
<< properties >>
string flatten true
<< end >>
