magic
tech sky130A
magscale 1 2
timestamp 1665749831
<< obsli1 >>
rect 184 527 18860 10897
<< obsm1 >>
rect 184 76 19214 11416
<< metal2 >>
rect 1398 11200 1454 12000
rect 4250 11200 4306 12000
rect 7102 11200 7158 12000
rect 9954 11200 10010 12000
rect 12806 11200 12862 12000
rect 15658 11200 15714 12000
rect 18510 11200 18566 12000
<< obsm2 >>
rect 480 11144 1342 11422
rect 1510 11144 4194 11422
rect 4362 11144 7046 11422
rect 7214 11144 9898 11422
rect 10066 11144 12750 11422
rect 12918 11144 15602 11422
rect 15770 11144 18454 11422
rect 18622 11144 19208 11422
rect 480 70 19208 11144
<< metal3 >>
rect 19200 11160 20000 11280
rect 19200 9664 20000 9784
rect 19200 8168 20000 8288
rect 19200 6672 20000 6792
rect 19200 5176 20000 5296
rect 19200 3680 20000 3800
rect 19200 2184 20000 2304
rect 19200 688 20000 808
<< obsm3 >>
rect 565 11080 19120 11250
rect 565 9864 19200 11080
rect 565 9584 19120 9864
rect 565 8368 19200 9584
rect 565 8088 19120 8368
rect 565 6872 19200 8088
rect 565 6592 19120 6872
rect 565 5376 19200 6592
rect 565 5096 19120 5376
rect 565 3880 19200 5096
rect 565 3600 19120 3880
rect 565 2384 19200 3600
rect 565 2104 19120 2384
rect 565 888 19200 2104
rect 565 608 19120 888
rect 565 511 19200 608
<< metal4 >>
rect 3104 496 3424 10928
rect 4654 496 4974 10928
rect 6204 496 6524 10928
rect 7754 496 8074 10928
rect 9304 496 9624 10928
rect 10854 496 11174 10928
rect 12404 496 12724 10928
rect 13954 496 14274 10928
rect 15504 496 15824 10928
rect 17054 496 17374 10928
rect 18604 496 18924 10928
<< obsm4 >>
rect 14411 987 15424 8533
rect 15904 987 16974 8533
rect 17454 987 17605 8533
<< metal5 >>
rect 136 9882 18924 10202
rect 136 8192 18908 8512
rect 136 6502 18924 6822
rect 136 4812 18908 5132
rect 136 3122 18924 3442
<< labels >>
rlabel metal4 s 4654 496 4974 10928 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 7754 496 8074 10928 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 10854 496 11174 10928 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 13954 496 14274 10928 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 17054 496 17374 10928 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 136 4812 18908 5132 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 136 8192 18908 8512 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 3104 496 3424 10928 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 6204 496 6524 10928 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 9304 496 9624 10928 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 12404 496 12724 10928 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 15504 496 15824 10928 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 18604 496 18924 10928 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 136 3122 18924 3442 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 136 6502 18924 6822 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 136 9882 18924 10202 6 VPWR
port 2 nsew power bidirectional
rlabel metal2 s 7102 11200 7158 12000 6 core_clk
port 3 nsew signal output
rlabel metal2 s 4250 11200 4306 12000 6 ext_clk
port 4 nsew signal input
rlabel metal3 s 19200 688 20000 808 6 ext_clk_sel
port 5 nsew signal input
rlabel metal3 s 19200 11160 20000 11280 6 ext_reset
port 6 nsew signal input
rlabel metal2 s 15658 11200 15714 12000 6 pll_clk
port 7 nsew signal input
rlabel metal2 s 18510 11200 18566 12000 6 pll_clk90
port 8 nsew signal input
rlabel metal2 s 1398 11200 1454 12000 6 resetb
port 9 nsew signal input
rlabel metal2 s 12806 11200 12862 12000 6 resetb_sync
port 10 nsew signal output
rlabel metal3 s 19200 6672 20000 6792 6 sel2[0]
port 11 nsew signal input
rlabel metal3 s 19200 8168 20000 8288 6 sel2[1]
port 12 nsew signal input
rlabel metal3 s 19200 9664 20000 9784 6 sel2[2]
port 13 nsew signal input
rlabel metal3 s 19200 2184 20000 2304 6 sel[0]
port 14 nsew signal input
rlabel metal3 s 19200 3680 20000 3800 6 sel[1]
port 15 nsew signal input
rlabel metal3 s 19200 5176 20000 5296 6 sel[2]
port 16 nsew signal input
rlabel metal2 s 9954 11200 10010 12000 6 user_clk
port 17 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 20000 12000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1397874
string GDS_FILE ../gds/caravel_clocking.gds
string GDS_START 391844
<< end >>

