* NGSPICE file created from caravel.ext - technology: sky130A

.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VPWR X VNB VPB
X0 VPWR a_75_212# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1 a_75_212# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2 a_75_212# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3 VGND a_75_212# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_1 A VGND VPWR X VNB VPB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
.ends

.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VPB VPWR VNB
D0 VNB DIODE sky130_fd_pr__diode_pw2nd_05v5 pj=5.36e+06u area=4.347e+11p
.ends

.subckt sky130_fd_sc_hd__buf_2 A VGND VPWR X VNB VPB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VPWR X VNB VPB
X0 a_219_297# a_27_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VGND B_N a_27_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VPWR A a_301_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 X a_219_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_301_297# a_27_53# a_219_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 X a_219_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_27_53# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VGND A a_219_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
.ends

.subckt sky130_fd_sc_hd__or2_1 A B VGND VPWR X VNB VPB
X0 VGND A a_68_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_68_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 X a_68_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A a_150_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 X a_68_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_150_297# B a_68_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VPWR X VNB VPB
X0 a_558_47# a_381_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND X a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_841_47# a_664_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR A a_62_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VGND A a_62_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_558_47# a_381_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 X a_62_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR X a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_841_47# a_664_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 X a_62_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VPWR a_558_47# a_664_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VGND a_558_47# a_664_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VPWR X VNB VPB
X0 a_244_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=820000u l=250000u
X1 VPWR a_244_47# a_355_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=820000u l=250000u
X2 X a_355_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND a_244_47# a_355_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=250000u
X6 X a_355_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_244_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=250000u
.ends

.subckt sky130_fd_sc_hd__decap_3 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
.ends

.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
R0 HI VPWR sky130_fd_pr__res_generic_po w=480000u l=45000u
R1 VGND LO sky130_fd_pr__res_generic_po w=480000u l=45000u
.ends

.subckt sky130_fd_sc_hd__dfbbn_1 CLK_N D RESET_B SET_B VGND VPWR Q Q_N VNB VPB
X0 a_791_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_1555_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VPWR RESET_B a_941_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 a_1415_315# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_791_47# a_941_21# a_647_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5 VGND a_1415_315# a_1363_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_1340_413# a_27_47# a_1256_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR CLK_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X8 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_473_413# a_193_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X10 a_1555_47# a_941_21# a_1415_315# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X11 VPWR a_1415_315# a_2136_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X12 a_1256_413# a_193_47# a_1112_329# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 a_581_47# a_27_47# a_473_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X14 a_647_21# a_473_413# a_791_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X15 a_647_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 VPWR a_941_21# a_891_329# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X17 a_557_413# a_193_47# a_473_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 Q a_2136_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_473_413# a_27_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 a_891_329# a_473_413# a_647_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X22 Q_N a_1415_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VGND RESET_B a_941_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 Q a_2136_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 VPWR a_647_21# a_557_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 a_1112_329# a_647_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X27 VGND a_647_21# a_581_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 VGND a_1415_315# a_2136_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X30 VPWR a_941_21# a_1672_329# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X31 VPWR a_1415_315# a_1340_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X32 a_1363_47# a_193_47# a_1256_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X33 Q_N a_1415_315# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X34 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X35 a_1159_47# a_647_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X36 a_1672_329# a_1256_413# a_1415_315# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X37 VGND CLK_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X38 a_1256_413# a_27_47# a_1159_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X39 a_1415_315# a_1256_413# a_1555_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
.ends

.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VPWR Q VNB VPB
X0 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X3 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X8 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X10 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X13 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X20 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X24 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
.ends

.subckt sky130_fd_sc_hd__einvp_8 A TE VGND VPWR Z VNB VPB
X0 VPWR a_27_47# a_215_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X1 a_215_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_193_47# A Z VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_215_309# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X4 Z A a_215_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND TE a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_215_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR a_27_47# a_215_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X8 a_215_309# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X9 Z A a_215_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_193_47# TE VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 Z A a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_193_47# TE VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_193_47# TE VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_193_47# TE VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_193_47# A Z VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_193_47# A Z VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_193_47# A Z VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_215_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND TE a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 VPWR a_27_47# a_215_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X21 VGND TE a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 VGND TE a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 Z A a_215_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 Z A a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 a_215_309# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X26 Z A a_215_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_215_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 Z A a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 VPWR a_27_47# a_215_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X30 Z A a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 a_215_309# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X32 VPWR TE a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 VGND TE a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VPWR X VNB VPB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__inv_2 A VGND VPWR Y VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__and2_1 A B VGND VPWR X VNB VPB
X0 VPWR B a_59_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 X a_59_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND B a_145_75# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_59_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 X a_59_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_145_75# A a_59_75# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__decap_6 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
.ends

.subckt sky130_fd_sc_hd__decap_8 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
.ends

.subckt gpio_logic_high gpio_logic1 vccd1 vssd1
XFILLER_3_3 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_3 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_0 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_5 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_6 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_7 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_8 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_9 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_3 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_3 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_4
Xgpio_logic_high vssd1 vssd1 vccd1 vccd1 gpio_logic1 gpio_logic_high/LO sky130_fd_sc_hd__conb_1
XFILLER_4_9 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_9 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
.ends

.subckt sky130_fd_sc_hd__buf_6 A VGND VPWR X VNB VPB
X0 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_161_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A a_161_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VPWR A a_161_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_161_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VPWR X VNB VPB
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X33 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X36 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X37 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X38 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X39 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__ebufn_8 A TE_B VGND VPWR Z VNB VPB
X0 VPWR TE_B a_407_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X1 a_455_47# a_301_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Z a_116_47# a_407_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Z a_116_47# a_455_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_116_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_407_309# a_116_47# Z VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR TE_B a_407_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X7 a_407_309# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X8 VGND a_301_47# a_455_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VGND a_301_47# a_455_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Z a_116_47# a_407_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_116_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND a_301_47# a_455_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_407_309# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X14 VGND a_301_47# a_455_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_455_47# a_116_47# Z VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VPWR TE_B a_407_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X17 a_455_47# a_116_47# Z VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_455_47# a_116_47# Z VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_301_47# TE_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_455_47# a_301_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 a_301_47# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_455_47# a_301_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_455_47# a_301_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 a_407_309# a_116_47# Z VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 Z a_116_47# a_455_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 Z a_116_47# a_455_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 VPWR A a_116_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 Z a_116_47# a_407_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 Z a_116_47# a_455_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 a_407_309# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X31 VGND A a_116_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X32 VPWR TE_B a_407_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X33 a_407_309# a_116_47# Z VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 Z a_116_47# a_407_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 a_407_309# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X36 a_455_47# a_116_47# Z VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X37 a_407_309# a_116_47# Z VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VPWR X VNB VPB
X0 VPWR a_505_21# a_535_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_505_21# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_218_374# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VGND a_505_21# a_439_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_76_199# A0 a_218_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_505_21# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_439_47# A0 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_535_374# A1 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_76_199# A1 a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_218_47# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt gpio_control_block gpio_defaults[0] gpio_defaults[10] gpio_defaults[11] gpio_defaults[12]
+ gpio_defaults[1] gpio_defaults[2] gpio_defaults[3] gpio_defaults[4] gpio_defaults[5]
+ gpio_defaults[6] gpio_defaults[7] gpio_defaults[8] gpio_defaults[9] mgmt_gpio_in
+ mgmt_gpio_oeb mgmt_gpio_out one pad_gpio_ana_en pad_gpio_ana_pol pad_gpio_ana_sel
+ pad_gpio_dm[0] pad_gpio_dm[1] pad_gpio_dm[2] pad_gpio_holdover pad_gpio_ib_mode_sel
+ pad_gpio_in pad_gpio_inenb pad_gpio_out pad_gpio_outenb pad_gpio_slow_sel pad_gpio_vtrip_sel
+ resetn resetn_out serial_clock serial_clock_out serial_data_in serial_data_out serial_load
+ serial_load_out user_gpio_in user_gpio_oeb user_gpio_out vccd1 vssd zero dw_1110_1538#
+ vccd vssd1
X_131_ _131_/A vssd vccd _131_/X vssd vccd sky130_fd_sc_hd__clkbuf_1
X_200_ _200_/A vssd vccd _201_/A vssd vccd sky130_fd_sc_hd__buf_1
X_114_ _114_/A vssd vccd _114_/X vssd vccd sky130_fd_sc_hd__clkbuf_1
XANTENNA_5 user_gpio_oeb vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput31 _205_/X vssd vccd pad_gpio_outenb vssd vccd sky130_fd_sc_hd__buf_2
X_130_ _136_/A _132_/B vssd vccd _131_/A vssd vccd sky130_fd_sc_hd__or2b_1
XFILLER_0_58 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_113_ _187_/A _113_/B vssd vccd _114_/A vssd vccd sky130_fd_sc_hd__or2_1
XANTENNA_6 user_gpio_out vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput32 _212_/Q vssd vccd pad_gpio_slow_sel vssd vccd sky130_fd_sc_hd__buf_2
Xoutput21 _220_/Q vssd vccd pad_gpio_ana_en vssd vccd sky130_fd_sc_hd__buf_2
X_189_ _189_/A _189_/B vssd vccd _190_/A vssd vccd sky130_fd_sc_hd__or2_1
XANTENNA_7 serial_data_in vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_112_ _202_/A vssd vccd _187_/A vssd vccd sky130_fd_sc_hd__dlymetal6s2s_1
Xhold10 _226_/D vssd vccd _211_/D vssd vccd sky130_fd_sc_hd__clkdlybuf4s25_1
Xoutput33 _213_/Q vssd vccd pad_gpio_vtrip_sel vssd vccd sky130_fd_sc_hd__buf_2
Xoutput22 _222_/Q vssd vccd pad_gpio_ana_pol vssd vccd sky130_fd_sc_hd__buf_2
X_188_ _188_/A vssd vccd _188_/X vssd vccd sky130_fd_sc_hd__clkbuf_1
X_111_ _111_/A vssd vccd _111_/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xoutput34 _202_/X vssd vccd resetn_out vssd vccd sky130_fd_sc_hd__buf_2
Xoutput23 _221_/Q vssd vccd pad_gpio_ana_sel vssd vccd sky130_fd_sc_hd__buf_2
Xhold11 _224_/D vssd vccd _210_/D vssd vccd sky130_fd_sc_hd__clkdlybuf4s25_1
X_187_ _187_/A _189_/A vssd vccd _188_/A vssd vccd sky130_fd_sc_hd__or2b_1
X_110_ _136_/A _113_/B vssd vccd _111_/A vssd vccd sky130_fd_sc_hd__or2b_1
Xhold12 _230_/D vssd vccd _221_/D vssd vccd sky130_fd_sc_hd__clkdlybuf4s25_1
Xoutput35 _203_/X vssd vccd serial_clock_out vssd vccd sky130_fd_sc_hd__clkbuf_1
Xoutput24 _217_/Q vssd vccd pad_gpio_dm[0] vssd vccd sky130_fd_sc_hd__buf_2
X_186_ _186_/A vssd vccd _186_/X vssd vccd sky130_fd_sc_hd__buf_1
X_169_ _169_/A _171_/B vssd vccd _170_/A vssd vccd sky130_fd_sc_hd__or2b_1
Xhold13 _233_/D vssd vccd hold1/A vssd vccd sky130_fd_sc_hd__clkdlybuf4s25_1
XPHY_0 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xoutput36 _199_/X vssd vccd serial_data_out vssd vccd sky130_fd_sc_hd__buf_2
Xoutput25 _218_/Q vssd vccd pad_gpio_dm[1] vssd vccd sky130_fd_sc_hd__buf_2
X_185_ _185_/A vssd vccd _186_/A vssd vccd sky130_fd_sc_hd__buf_1
X_168_ _168_/A vssd vccd _168_/X vssd vccd sky130_fd_sc_hd__buf_1
Xhold14 _231_/D vssd vccd _222_/D vssd vccd sky130_fd_sc_hd__clkdlybuf4s25_1
XPHY_1 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xoutput37 _204_/X vssd vccd serial_load_out vssd vccd sky130_fd_sc_hd__clkbuf_1
Xoutput26 _219_/Q vssd vccd pad_gpio_dm[2] vssd vccd sky130_fd_sc_hd__buf_2
Xconst_source vssd vssd vccd vccd one zero sky130_fd_sc_hd__conb_1
X_184_ _184_/A vssd vccd _184_/X vssd vccd sky130_fd_sc_hd__clkbuf_1
X_167_ _173_/A vssd vccd _168_/A vssd vccd sky130_fd_sc_hd__buf_1
Xhold15 _232_/D vssd vccd hold4/A vssd vccd sky130_fd_sc_hd__clkdlybuf4s25_1
X_219_ _129_/X hold8/X _133_/X _131_/X vssd vccd _219_/Q _219_/Q_N vssd vccd sky130_fd_sc_hd__dfbbn_1
XPHY_2 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xoutput27 _211_/Q vssd vccd pad_gpio_holdover vssd vccd sky130_fd_sc_hd__buf_2
X_166_ _166_/A vssd vccd _166_/X vssd vccd sky130_fd_sc_hd__clkbuf_1
X_235_ _203_/A _235_/D _202_/A vssd vccd hold8/A vssd vccd sky130_fd_sc_hd__dfrtp_1
X_183_ _183_/A _183_/B vssd vccd _184_/A vssd vccd sky130_fd_sc_hd__or2_1
Xoutput28 _215_/Q vssd vccd pad_gpio_ib_mode_sel vssd vccd sky130_fd_sc_hd__buf_2
X_149_ _149_/A vssd vccd _149_/X vssd vccd sky130_fd_sc_hd__buf_1
Xhold16 _228_/D vssd vccd hold2/A vssd vccd sky130_fd_sc_hd__clkdlybuf4s25_1
X_218_ _135_/X hold5/X _139_/X _137_/X vssd vccd _218_/Q _218_/Q_N vssd vccd sky130_fd_sc_hd__dfbbn_1
XPHY_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_182_ _182_/A vssd vccd _182_/X vssd vccd sky130_fd_sc_hd__clkbuf_1
X_217_ _141_/X hold6/X _146_/X _144_/X vssd vccd _217_/Q _206_/A0 vssd vccd sky130_fd_sc_hd__dfbbn_1
X_234_ _203_/A _234_/D _202_/A vssd vccd _235_/D vssd vccd sky130_fd_sc_hd__dfrtp_1
X_148_ _173_/A vssd vccd _149_/A vssd vccd sky130_fd_sc_hd__buf_1
X_165_ _183_/A _165_/B vssd vccd _166_/A vssd vccd sky130_fd_sc_hd__or2_1
Xhold17 _234_/D vssd vccd hold6/A vssd vccd sky130_fd_sc_hd__clkdlybuf4s25_1
XPHY_4 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xoutput29 _214_/Q vssd vccd pad_gpio_inenb vssd vccd sky130_fd_sc_hd__buf_2
X_164_ _164_/A vssd vccd _164_/X vssd vccd sky130_fd_sc_hd__clkbuf_1
X_233_ _203_/A _233_/D _202_/A vssd vccd _234_/D vssd vccd sky130_fd_sc_hd__dfrtp_1
X_181_ _187_/A _183_/B vssd vccd _182_/A vssd vccd sky130_fd_sc_hd__or2b_1
X_216_ _149_/X hold3/X _153_/X _151_/X vssd vccd _216_/Q _216_/Q_N vssd vccd sky130_fd_sc_hd__dfbbn_1
X_147_ _147_/A vssd vccd _173_/A vssd vccd sky130_fd_sc_hd__buf_1
Xhold18 _225_/D vssd vccd hold3/A vssd vccd sky130_fd_sc_hd__clkdlybuf4s25_1
XPHY_5 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_180_ _180_/A vssd vccd _180_/X vssd vccd sky130_fd_sc_hd__buf_1
X_232_ _203_/A _232_/D _202_/A vssd vccd _233_/D vssd vccd sky130_fd_sc_hd__dfrtp_1
X_163_ _169_/A _165_/B vssd vccd _164_/A vssd vccd sky130_fd_sc_hd__or2b_1
Xhold19 _235_/D vssd vccd hold5/A vssd vccd sky130_fd_sc_hd__clkdlybuf4s25_1
XPHY_6 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_146_ _146_/A vssd vccd _146_/X vssd vccd sky130_fd_sc_hd__clkbuf_1
X_129_ _129_/A vssd vccd _129_/X vssd vccd sky130_fd_sc_hd__buf_1
X_215_ _155_/X hold2/X _160_/X _157_/X vssd vccd _215_/Q _215_/Q_N vssd vccd sky130_fd_sc_hd__dfbbn_1
X_231_ _231_/CLK _231_/D _202_/A vssd vccd _232_/D vssd vccd sky130_fd_sc_hd__dfrtp_1
X_162_ _162_/A vssd vccd _162_/X vssd vccd sky130_fd_sc_hd__buf_1
Xinput1 gpio_defaults[0] vssd vccd _189_/A vssd vccd sky130_fd_sc_hd__clkbuf_1
X_214_ _162_/X hold7/X _166_/X _164_/X vssd vccd _214_/Q _214_/Q_N vssd vccd sky130_fd_sc_hd__dfbbn_1
X_145_ _152_/A _145_/B vssd vccd _146_/A vssd vccd sky130_fd_sc_hd__or2_1
XPHY_7 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_128_ _140_/A vssd vccd _129_/A vssd vccd sky130_fd_sc_hd__buf_1
Xinput2 gpio_defaults[10] vssd vccd _145_/B vssd vccd sky130_fd_sc_hd__clkbuf_1
Xgpio_in_buf _197_/Y gpio_in_buf/TE vssd vccd user_gpio_in vssd vccd sky130_fd_sc_hd__einvp_8
X_230_ _231_/CLK _230_/D _202_/A vssd vccd _231_/D vssd vccd sky130_fd_sc_hd__dfrtp_1
X_161_ _173_/A vssd vccd _162_/A vssd vccd sky130_fd_sc_hd__buf_1
XPHY_8 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_144_ _144_/A vssd vccd _144_/X vssd vccd sky130_fd_sc_hd__clkbuf_1
X_127_ _127_/A vssd vccd _127_/X vssd vccd sky130_fd_sc_hd__clkbuf_1
X_213_ _168_/X hold1/X _172_/X _170_/X vssd vccd _213_/Q _213_/Q_N vssd vccd sky130_fd_sc_hd__dfbbn_1
X_160_ _160_/A vssd vccd _160_/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput3 gpio_defaults[11] vssd vccd _138_/B vssd vccd sky130_fd_sc_hd__clkbuf_1
X_212_ _174_/X hold4/X _178_/X _176_/X vssd vccd _212_/Q _212_/Q_N vssd vccd sky130_fd_sc_hd__dfbbn_1
X_143_ _169_/A _145_/B vssd vccd _144_/A vssd vccd sky130_fd_sc_hd__or2b_1
XPHY_9 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_126_ _152_/A _126_/B vssd vccd _127_/A vssd vccd sky130_fd_sc_hd__or2_1
X_109_ _189_/B vssd vccd _136_/A vssd vccd sky130_fd_sc_hd__dlymetal6s2s_1
Xinput4 gpio_defaults[12] vssd vccd _132_/B vssd vccd sky130_fd_sc_hd__clkbuf_1
X_125_ _189_/B vssd vccd _152_/A vssd vccd sky130_fd_sc_hd__dlymetal6s2s_1
X_142_ _189_/B vssd vccd _169_/A vssd vccd sky130_fd_sc_hd__dlymetal6s2s_1
X_211_ _180_/X _211_/D _184_/X _182_/X vssd vccd _211_/Q _211_/Q_N vssd vccd sky130_fd_sc_hd__dfbbn_1
X_108_ _202_/A vssd vccd _189_/B vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput5 gpio_defaults[1] vssd vccd _152_/B vssd vccd sky130_fd_sc_hd__clkbuf_1
X_210_ _186_/X _210_/D _190_/X _188_/X vssd vccd _210_/Q _210_/Q_N vssd vccd sky130_fd_sc_hd__dfbbn_1
X_141_ _141_/A vssd vccd _141_/X vssd vccd sky130_fd_sc_hd__buf_1
X_124_ _124_/A vssd vccd _124_/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0_serial_clock clkbuf_0_serial_clock/X vssd vccd _203_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
X_115__1 serial_load vssd vccd _200_/A vssd vccd sky130_fd_sc_hd__inv_2
Xinput6 gpio_defaults[2] vssd vccd _183_/B vssd vccd sky130_fd_sc_hd__clkbuf_1
X_140_ _140_/A vssd vccd _141_/A vssd vccd sky130_fd_sc_hd__buf_1
Xinput20 user_gpio_out vssd vccd _208_/A0 vssd vccd sky130_fd_sc_hd__clkbuf_1
X_123_ _136_/A _126_/B vssd vccd _124_/A vssd vccd sky130_fd_sc_hd__or2b_1
X_115__2 serial_load vssd vccd _185_/A vssd vccd sky130_fd_sc_hd__inv_2
Xinput7 gpio_defaults[3] vssd vccd _165_/B vssd vccd sky130_fd_sc_hd__clkbuf_1
X_199_ _199_/A vssd vccd _199_/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput10 gpio_defaults[6] vssd vccd _119_/B vssd vccd sky130_fd_sc_hd__clkbuf_1
X_122_ _122_/A vssd vccd _122_/X vssd vccd sky130_fd_sc_hd__buf_1
X_115__3 serial_load vssd vccd _179_/A vssd vccd sky130_fd_sc_hd__inv_2
Xinput8 gpio_defaults[4] vssd vccd _159_/B vssd vccd sky130_fd_sc_hd__clkbuf_1
X_198_ one hold8/A vssd vccd _199_/A vssd vccd sky130_fd_sc_hd__and2_1
Xinput11 gpio_defaults[7] vssd vccd _113_/B vssd vccd sky130_fd_sc_hd__clkbuf_1
X_121_ _140_/A vssd vccd _122_/A vssd vccd sky130_fd_sc_hd__buf_1
X_115__4 serial_load vssd vccd _147_/A vssd vccd sky130_fd_sc_hd__inv_2
Xinput9 gpio_defaults[5] vssd vccd _126_/B vssd vccd sky130_fd_sc_hd__clkbuf_1
X_197_ _209_/A vssd vccd _197_/Y vssd vccd sky130_fd_sc_hd__inv_2
X_120_ _120_/A vssd vccd _120_/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput12 gpio_defaults[8] vssd vccd _177_/B vssd vccd sky130_fd_sc_hd__clkbuf_1
X_115__5 serial_load vssd vccd _116_/A vssd vccd sky130_fd_sc_hd__inv_2
Xhold1 hold1/A vssd vccd hold1/X vssd vccd sky130_fd_sc_hd__clkdlybuf4s25_1
X_196_ _196_/A vssd vccd _206_/S vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput13 gpio_defaults[9] vssd vccd _171_/B vssd vccd sky130_fd_sc_hd__clkbuf_1
X_179_ _179_/A vssd vccd _180_/A vssd vccd sky130_fd_sc_hd__buf_1
Xhold2 hold2/A vssd vccd hold2/X vssd vccd sky130_fd_sc_hd__clkdlybuf4s25_1
Xgpio_logic_high gpio_in_buf/TE vccd1 vssd1 gpio_logic_high
Xinput14 mgmt_gpio_oeb vssd vccd _207_/S vssd vccd sky130_fd_sc_hd__clkbuf_1
X_195_ _219_/Q _218_/Q vssd vccd _196_/A vssd vccd sky130_fd_sc_hd__or2b_1
X_178_ _178_/A vssd vccd _178_/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xhold3 hold3/A vssd vccd hold3/X vssd vccd sky130_fd_sc_hd__clkdlybuf4s25_1
XPHY_30 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_194_ _194_/A vssd vccd _194_/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput15 mgmt_gpio_out vssd vccd _207_/A0 vssd vccd sky130_fd_sc_hd__clkbuf_1
X_177_ _183_/A _177_/B vssd vccd _178_/A vssd vccd sky130_fd_sc_hd__or2_1
X_229_ _231_/CLK hold9/A _202_/A vssd vccd _230_/D vssd vccd sky130_fd_sc_hd__dfrtp_1
Xhold4 hold4/A vssd vccd hold4/X vssd vccd sky130_fd_sc_hd__clkdlybuf4s25_1
XPHY_31 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_20 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_193_ _216_/Q _207_/S vssd vccd _194_/A vssd vccd sky130_fd_sc_hd__and2_1
X_176_ _176_/A vssd vccd _176_/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput16 pad_gpio_in vssd vccd _209_/A vssd vccd sky130_fd_sc_hd__clkbuf_1
X_228_ _231_/CLK _228_/D _202_/A vssd vccd hold9/A vssd vccd sky130_fd_sc_hd__dfrtp_1
X_159_ _183_/A _159_/B vssd vccd _160_/A vssd vccd sky130_fd_sc_hd__or2_1
Xhold5 hold5/A vssd vccd hold5/X vssd vccd sky130_fd_sc_hd__clkdlybuf4s25_1
XPHY_32 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_21 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_10 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_192_ _192_/A vssd vccd _192_/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput17 resetn vssd vccd _202_/A vssd vccd sky130_fd_sc_hd__buf_6
X_175_ _187_/A _177_/B vssd vccd _176_/A vssd vccd sky130_fd_sc_hd__or2b_1
X_158_ _189_/B vssd vccd _183_/A vssd vccd sky130_fd_sc_hd__clkbuf_1
X_227_ _231_/CLK hold7/A _202_/A vssd vccd _228_/D vssd vccd sky130_fd_sc_hd__dfrtp_1
Xhold6 hold6/A vssd vccd hold6/X vssd vccd sky130_fd_sc_hd__clkdlybuf4s25_1
Xclkbuf_1_0_0_serial_clock clkbuf_0_serial_clock/X vssd vccd _231_/CLK vssd vccd sky130_fd_sc_hd__clkbuf_2
XPHY_33 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_22 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_11 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xclkbuf_0_serial_clock serial_clock vssd vccd clkbuf_0_serial_clock/X vssd vccd sky130_fd_sc_hd__clkbuf_16
X_191_ _214_/Q _216_/Q vssd vccd _192_/A vssd vccd sky130_fd_sc_hd__or2b_1
X_157_ _157_/A vssd vccd _157_/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput18 serial_data_in vssd vccd _223_/D vssd vccd sky130_fd_sc_hd__clkbuf_1
X_226_ _231_/CLK _226_/D _202_/A vssd vccd hold7/A vssd vccd sky130_fd_sc_hd__dfrtp_1
X_174_ _174_/A vssd vccd _174_/X vssd vccd sky130_fd_sc_hd__buf_1
X_209_ _209_/A _192_/X vssd vccd mgmt_gpio_in vssd vccd sky130_fd_sc_hd__ebufn_8
Xhold7 hold7/A vssd vccd hold7/X vssd vccd sky130_fd_sc_hd__clkdlybuf4s25_1
XPHY_12 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_34 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_23 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_190_ _190_/A vssd vccd _190_/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput19 user_gpio_oeb vssd vccd _205_/A0 vssd vccd sky130_fd_sc_hd__clkbuf_1
X_173_ _173_/A vssd vccd _174_/A vssd vccd sky130_fd_sc_hd__buf_1
X_225_ _231_/CLK _225_/D _202_/A vssd vccd _226_/D vssd vccd sky130_fd_sc_hd__dfrtp_1
X_156_ _169_/A _159_/B vssd vccd _157_/A vssd vccd sky130_fd_sc_hd__or2b_1
Xhold8 hold8/A vssd vccd hold8/X vssd vccd sky130_fd_sc_hd__clkdlybuf4s25_1
X_139_ _139_/A vssd vccd _139_/X vssd vccd sky130_fd_sc_hd__clkbuf_1
X_208_ _208_/A0 _207_/X _210_/Q vssd vccd _208_/X vssd vccd sky130_fd_sc_hd__mux2_1
XPHY_35 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_24 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_13 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_172_ _172_/A vssd vccd _172_/X vssd vccd sky130_fd_sc_hd__clkbuf_1
X_224_ _231_/CLK _224_/D _202_/A vssd vccd _225_/D vssd vccd sky130_fd_sc_hd__dfrtp_1
X_155_ _155_/A vssd vccd _155_/X vssd vccd sky130_fd_sc_hd__buf_1
X_207_ _207_/A0 _206_/X _207_/S vssd vccd _207_/X vssd vccd sky130_fd_sc_hd__mux2_1
X_138_ _152_/A _138_/B vssd vccd _139_/A vssd vccd sky130_fd_sc_hd__or2_1
Xhold9 hold9/A vssd vccd hold9/X vssd vccd sky130_fd_sc_hd__clkdlybuf4s25_1
XPHY_36 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_25 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_14 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_171_ _183_/A _171_/B vssd vccd _172_/A vssd vccd sky130_fd_sc_hd__or2_1
X_223_ _203_/A _223_/D _202_/A vssd vccd _224_/D vssd vccd sky130_fd_sc_hd__dfrtp_1
X_154_ _173_/A vssd vccd _155_/A vssd vccd sky130_fd_sc_hd__buf_1
X_137_ _137_/A vssd vccd _137_/X vssd vccd sky130_fd_sc_hd__clkbuf_1
X_206_ _206_/A0 _207_/A0 _206_/S vssd vccd _206_/X vssd vccd sky130_fd_sc_hd__mux2_1
XPHY_37 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_26 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_170_ _170_/A vssd vccd _170_/X vssd vccd sky130_fd_sc_hd__clkbuf_1
X_153_ _153_/A vssd vccd _153_/X vssd vccd sky130_fd_sc_hd__clkbuf_1
X_222_ _201_/X _222_/D _114_/X _111_/X vssd vccd _222_/Q _222_/Q_N vssd vccd sky130_fd_sc_hd__dfbbn_1
X_205_ _205_/A0 _194_/X _210_/Q vssd vccd _205_/X vssd vccd sky130_fd_sc_hd__mux2_1
X_136_ _136_/A _138_/B vssd vccd _137_/A vssd vccd sky130_fd_sc_hd__or2b_1
X_119_ _187_/A _119_/B vssd vccd _120_/A vssd vccd sky130_fd_sc_hd__or2_1
XPHY_27 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_16 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_0 mgmt_gpio_oeb vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_152_ _152_/A _152_/B vssd vccd _153_/A vssd vccd sky130_fd_sc_hd__or2_1
X_221_ _140_/A _221_/D _120_/X _118_/X vssd vccd _221_/Q _221_/Q_N vssd vccd sky130_fd_sc_hd__dfbbn_1
X_118_ _118_/A vssd vccd _118_/X vssd vccd sky130_fd_sc_hd__clkbuf_1
X_204_ serial_load vssd vccd _204_/X vssd vccd sky130_fd_sc_hd__buf_2
X_135_ _135_/A vssd vccd _135_/X vssd vccd sky130_fd_sc_hd__buf_1
XPHY_28 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_17 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_1 mgmt_gpio_out vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_151_ _151_/A vssd vccd _151_/X vssd vccd sky130_fd_sc_hd__clkbuf_1
X_203_ _203_/A vssd vccd _203_/X vssd vccd sky130_fd_sc_hd__buf_2
X_134_ _140_/A vssd vccd _135_/A vssd vccd sky130_fd_sc_hd__buf_1
X_220_ _122_/X hold9/X _127_/X _124_/X vssd vccd _220_/Q _220_/Q_N vssd vccd sky130_fd_sc_hd__dfbbn_1
X_117_ _136_/A _119_/B vssd vccd _118_/A vssd vccd sky130_fd_sc_hd__or2b_1
XPHY_29 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_18 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_2 one vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_150_ _169_/A _152_/B vssd vccd _151_/A vssd vccd sky130_fd_sc_hd__or2b_1
X_133_ _133_/A vssd vccd _133_/X vssd vccd sky130_fd_sc_hd__clkbuf_1
X_202_ _202_/A vssd vccd _202_/X vssd vccd sky130_fd_sc_hd__clkbuf_1
XPHY_19 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_3 one vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_116_ _116_/A vssd vccd _140_/A vssd vccd sky130_fd_sc_hd__buf_1
X_201_ _201_/A vssd vccd _201_/X vssd vccd sky130_fd_sc_hd__buf_1
X_132_ _152_/A _132_/B vssd vccd _133_/A vssd vccd sky130_fd_sc_hd__or2_1
XANTENNA_4 pad_gpio_in vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput30 _208_/X vssd vccd pad_gpio_out vssd vccd sky130_fd_sc_hd__buf_2
.ends

.subckt sky130_fd_sc_hd__decap_12 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
.ends

.subckt gpio_defaults_block VGND gpio_defaults[0] gpio_defaults[10] gpio_defaults[11]
+ gpio_defaults[12] gpio_defaults[1] gpio_defaults[2] gpio_defaults[3] gpio_defaults[4]
+ gpio_defaults[5] gpio_defaults[6] gpio_defaults[7] gpio_defaults[8] gpio_defaults[9]
+ VPWR
Xgpio_default_value\[8\] VGND VGND VPWR VPWR gpio_default_value\[8\]/HI gpio_defaults[8]
+ sky130_fd_sc_hd__conb_1
Xgpio_default_value\[6\] VGND VGND VPWR VPWR gpio_default_value\[6\]/HI gpio_defaults[6]
+ sky130_fd_sc_hd__conb_1
XFILLER_1_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_0 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xgpio_default_value\[4\] VGND VGND VPWR VPWR gpio_default_value\[4\]/HI gpio_defaults[4]
+ sky130_fd_sc_hd__conb_1
XPHY_2 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_4 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_5 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xgpio_default_value\[2\] VGND VGND VPWR VPWR gpio_default_value\[2\]/HI gpio_defaults[2]
+ sky130_fd_sc_hd__conb_1
XFILLER_1_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xgpio_default_value\[12\] VGND VGND VPWR VPWR gpio_default_value\[12\]/HI gpio_defaults[12]
+ sky130_fd_sc_hd__conb_1
Xgpio_default_value\[0\] VGND VGND VPWR VPWR gpio_default_value\[0\]/HI gpio_defaults[0]
+ sky130_fd_sc_hd__conb_1
XFILLER_1_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xgpio_default_value\[10\] VGND VGND VPWR VPWR gpio_defaults[10] gpio_default_value\[10\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xgpio_default_value\[9\] VGND VGND VPWR VPWR gpio_default_value\[9\]/HI gpio_defaults[9]
+ sky130_fd_sc_hd__conb_1
XFILLER_2_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xgpio_default_value\[7\] VGND VGND VPWR VPWR gpio_default_value\[7\]/HI gpio_defaults[7]
+ sky130_fd_sc_hd__conb_1
XFILLER_2_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xgpio_default_value\[5\] VGND VGND VPWR VPWR gpio_default_value\[5\]/HI gpio_defaults[5]
+ sky130_fd_sc_hd__conb_1
XFILLER_2_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xgpio_default_value\[3\] VGND VGND VPWR VPWR gpio_default_value\[3\]/HI gpio_defaults[3]
+ sky130_fd_sc_hd__conb_1
XFILLER_2_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xgpio_default_value\[1\] VGND VGND VPWR VPWR gpio_defaults[1] gpio_default_value\[1\]/LO
+ sky130_fd_sc_hd__conb_1
Xgpio_default_value\[11\] VGND VGND VPWR VPWR gpio_default_value\[11\]/HI gpio_defaults[11]
+ sky130_fd_sc_hd__conb_1
.ends

.subckt sky130_fd_sc_hd__or3_2 A B C VGND VPWR X VNB VPB
X0 VPWR a_30_53# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND a_30_53# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X a_30_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_112_297# C a_30_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 X a_30_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND A a_30_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_30_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VGND C a_30_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_184_297# B a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VPWR A a_184_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VPWR Q VNB VPB
X0 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X4 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X10 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X12 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X15 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X22 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X26 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkinv_1 A VGND VPWR Y VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VPWR X VNB VPB
X0 a_79_21# C1 a_635_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR A2 a_319_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_417_47# A2 a_319_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_79_21# A1 a_417_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_319_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_319_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_319_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_79_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_635_297# B1 a_319_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VPWR X VNB VPB
X0 VPWR a_82_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_646_47# B2 a_82_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_574_369# a_313_47# a_82_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 a_574_369# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 VGND a_82_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR B2 a_574_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X6 X a_82_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 X a_82_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_313_47# A2_N a_313_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X9 a_313_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_313_297# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X11 VGND A2_N a_313_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_82_21# a_313_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VGND B1 a_646_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__einvp_2 A TE VGND VPWR Z VNB VPB
X0 VPWR a_27_47# a_215_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X1 a_204_47# A Z VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR TE a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 Z A a_204_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_215_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Z A a_215_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_204_47# TE VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND TE a_204_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_215_309# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X9 VGND TE a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__einvn_8 A TE_B VGND VPWR Z VNB VPB
X0 a_204_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_215_47# A Z VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Z A a_204_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_204_309# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X7 a_204_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR TE_B a_204_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X10 Z A a_204_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_204_309# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X12 a_215_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 Z A a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_215_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_215_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VPWR TE_B a_204_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X17 a_215_47# A Z VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_204_309# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X19 a_215_47# A Z VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_215_47# A Z VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 a_204_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 VPWR TE_B a_204_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X23 a_204_309# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X24 Z A a_204_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 Z A a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 Z A a_204_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_204_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 Z A a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 VPWR TE_B a_204_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X30 Z A a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 a_215_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X32 VPWR TE_B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 VGND TE_B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VPWR X VNB VPB
X0 X a_91_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_91_21# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_360_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR B1 a_91_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_360_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND A2 a_360_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_360_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR a_91_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND a_91_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 X a_91_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_677_47# B1 a_360_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_460_297# A2 a_360_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_91_21# C1 a_677_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_91_21# A3 a_460_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__or2_2 A B VGND VPWR X VNB VPB
X0 a_121_297# B a_39_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 X a_39_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR a_39_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_39_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND a_39_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR A a_121_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VGND A a_39_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_39_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__einvn_4 A TE_B VGND VPWR Z VNB VPB
X0 VGND a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_204_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR TE_B a_204_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X4 Z A a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_204_309# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X6 a_215_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Z A a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Z A a_204_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR TE_B a_204_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X10 a_204_309# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X11 a_215_47# A Z VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_215_47# A Z VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_215_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_204_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VPWR TE_B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 Z A a_204_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VGND TE_B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand2_2 A B VGND VPWR Y VNB VPB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VPWR X VNB VPB
X0 VPWR a_38_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR A1 a_497_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 X a_38_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_141_47# B2 a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_497_297# A2 a_38_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND A1 a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR C1 a_38_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_237_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_38_47# B2 a_237_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_225_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 X a_38_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_141_47# C1 a_38_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND a_38_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_225_47# B1 a_141_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VPWR X VNB VPB
X0 VPWR A2 a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_277_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_79_21# B1 a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_277_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_361_47# A2 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_277_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VGND B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_79_21# A1 a_361_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VPWR X VNB VPB
X0 VPWR A3 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_299_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_352_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_549_47# A1 a_21_199# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 X a_21_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND a_21_199# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_665_47# A2 a_549_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR A1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_299_297# B1 a_21_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_21_199# B2 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VGND A3 a_665_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR a_21_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 X a_21_199# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_21_199# B1 a_352_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VPWR X VNB VPB
X0 VPWR a_27_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND A2 a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_27_297# B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_27_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND a_27_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_381_47# A1 a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_109_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_109_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VPWR Y VNB VPB
X0 VGND A2 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Y B1 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR A1 a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_29_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y A2 a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND A1 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_112_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_112_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_29_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_29_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor2_2 A B VGND VPWR Y VNB VPB
X0 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VPWR X VNB VPB
X0 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VGND D a_304_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_198_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_27_47# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_304_47# C a_198_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VPWR D a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VPWR X VNB VPB
X0 a_301_47# B2 a_81_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VGND A2 a_301_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_383_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_301_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 X a_81_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 X a_81_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR A1 a_579_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_81_21# B1 a_301_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_579_297# A2 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_81_21# B2 a_383_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VPWR X VNB VPB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_465_47# A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_109_297# B1 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_205_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR A2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_193_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_27_47# B1 a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_109_297# C1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND A2 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VPWR Y VNB VPB
X0 VGND A2 a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y A1 a_114_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_114_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_285_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VPWR X VNB VPB
X0 a_108_21# B1 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_346_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X a_108_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_108_21# A3 a_430_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_430_297# A2 a_346_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR a_108_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_346_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND A2 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 X a_108_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR B1 a_108_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VGND a_108_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_346_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VPWR Y VNB VPB
X0 Y A2 a_734_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_300_47# B2 a_28_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_300_47# B1 a_28_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_300_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_300_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_734_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_28_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y C1 a_28_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR B1 a_382_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_382_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_28_47# B1 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_28_47# B2 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VGND A1 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 Y B2 a_382_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VPWR A1 a_734_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VGND A2 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_382_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_734_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__einvp_1 A TE VGND VPWR Z VNB VPB
X0 a_276_297# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Z A a_204_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR TE a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 Z A a_276_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_204_47# TE VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND TE a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and3_2 A B C VGND VPWR X VNB VPB
X0 VPWR a_29_311# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X a_29_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A a_29_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VGND a_29_311# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_184_53# B a_112_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR C a_29_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 X a_29_311# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_112_53# A a_29_311# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_29_311# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VGND C a_184_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VPWR X VNB VPB
X0 VPWR A1 a_485_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_485_297# a_297_93# a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_297_93# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_581_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_79_21# a_297_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND A2 a_581_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_297_93# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_485_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VPWR X VNB VPB
X0 VGND A2 a_393_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_496_297# A4 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_393_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A1 a_697_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND A4 a_393_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_697_297# A2 a_597_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_393_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_393_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_597_297# A3 a_496_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VPWR X VNB VPB
X0 a_294_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VPWR A2_N a_295_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 VPWR B1 a_665_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 VGND a_84_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 X a_84_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_581_47# a_295_369# a_84_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR a_84_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_665_369# B2 a_84_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X8 VGND B2 a_581_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_295_369# A2_N a_294_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 X a_84_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_84_21# a_295_369# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X12 a_295_369# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X13 a_581_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VPWR X VNB VPB
X0 VPWR A1 a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_470_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_384_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_384_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VPWR Y VNB VPB
X0 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_27_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_475_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR A1 a_475_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_27_47# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_475_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 Y A2 a_475_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkinv_2 A VGND VPWR Y VNB VPB
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VPWR X VNB VPB
X0 a_429_297# A2 a_345_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND A2 a_345_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_345_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_345_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_629_297# B2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR B1 a_629_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_79_21# B2 a_345_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_345_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_79_21# A3 a_429_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_345_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkinv_8 A VGND VPWR Y VNB VPB
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VPWR X VNB VPB
X0 a_27_47# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR C1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR A1 a_373_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_182_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_182_47# B1 a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_373_297# A2 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_110_47# C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND A1 a_182_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VPWR X VNB VPB
X0 VPWR a_80_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X a_80_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND a_80_199# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_386_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_80_199# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_80_199# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_386_297# B1 a_80_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_458_47# A1 a_80_199# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR A1 a_386_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND A2 a_458_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VPWR Y VNB VPB
X0 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_298_47# C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VGND A1 a_497_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_664_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A2 a_497_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_298_47# B1 a_497_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_497_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y D1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_497_47# B1 a_298_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 Y A2 a_664_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_27_47# C1 a_298_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VPWR D1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_27_47# D1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_497_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 Y D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 VPWR A1 a_664_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_664_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__o2bb2ai_2 A1_N A2_N B1 B2 VGND VPWR Y VNB VPB
X0 a_113_297# A2_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_113_47# A2_N a_113_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR B1 a_730_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR A2_N a_113_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_730_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_471_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_471_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y B2 a_730_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_113_297# A2_N a_113_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_113_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND A1_N a_113_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND B2 a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VPWR a_113_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_113_297# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y a_113_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_730_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 Y a_113_297# a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_471_47# a_113_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VPWR A1_N a_113_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND B1 a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and2_2 A B VGND VPWR X VNB VPB
X0 X a_61_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR a_61_75# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR B a_61_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VGND B a_147_75# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 X a_61_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND a_61_75# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_61_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_147_75# A a_61_75# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VPWR X VNB VPB
X0 a_27_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_27_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_277_297# B a_205_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR A a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_205_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR a_27_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND a_27_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND C a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_109_297# D a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VGND A a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VPWR Y VNB VPB
X0 a_109_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_467_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_467_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y A1 a_467_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_109_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND A2 a_467_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_27_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VPWR A1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_109_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt digital_pll clockp[0] clockp[1] dco div[0] div[1] div[2] div[3] div[4] enable
+ ext_trim[0] ext_trim[10] ext_trim[11] ext_trim[12] ext_trim[13] ext_trim[14] ext_trim[15]
+ ext_trim[16] ext_trim[17] ext_trim[18] ext_trim[19] ext_trim[1] ext_trim[20] ext_trim[21]
+ ext_trim[22] ext_trim[23] ext_trim[24] ext_trim[25] ext_trim[2] ext_trim[3] ext_trim[4]
+ ext_trim[5] ext_trim[6] ext_trim[7] ext_trim[8] ext_trim[9] osc resetb VPWR VGND
XFILLER_22_133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__338__A1 ext_trim[7] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_294_ _297_/C _302_/C _301_/A VGND VPWR _294_/X VGND VPWR sky130_fd_sc_hd__or3_2
X_363_ _328_/A _363_/D _318_/X VGND VPWR _363_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
Xringosc.dstage\[1\].id.delayint0 ringosc.dstage\[1\].id.delayen1/Z VGND VPWR ringosc.dstage\[1\].id.delayen0/A
+ VGND VPWR sky130_fd_sc_hd__clkinv_1
X_346_ _288_/B ext_trim[3] dco VGND VPWR _346_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_277_ _362_/Q _272_/B _363_/Q _267_/B _226_/B VGND VPWR _359_/D VGND VPWR sky130_fd_sc_hd__a311o_2
X_200_ _196_/A _199_/Y _196_/A _199_/Y VGND VPWR _200_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_2
Xringosc.dstage\[11\].id.delayen1 ringosc.dstage\[11\].id.delayen1/A _331_/X VGND
+ VPWR ringosc.dstage\[11\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvp_2
X_329_ _292_/B _232_/B _370_/Q VGND VPWR _329_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xringosc.dstage\[10\].id.delayenb0 ringosc.dstage\[10\].id.delayenb1/A _332_/X VGND
+ VPWR ringosc.dstage\[10\].id.delayen0/Z VGND VPWR sky130_fd_sc_hd__einvn_8
Xringosc.dstage\[9\].id.delayenb0 ringosc.dstage\[9\].id.delayenb1/A _334_/X VGND
+ VPWR ringosc.dstage\[9\].id.delayen0/Z VGND VPWR sky130_fd_sc_hd__einvn_8
X_293_ _367_/Q _221_/B _302_/B _370_/Q _232_/B VGND VPWR _293_/X VGND VPWR sky130_fd_sc_hd__o311a_2
X_362_ _328_/A _362_/D _319_/X VGND VPWR _362_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_276_ _276_/A _276_/B VGND VPWR _360_/D VGND VPWR sky130_fd_sc_hd__or2_2
X_345_ _300_/X ext_trim[17] dco VGND VPWR _345_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_259_ _366_/Q _220_/Y _262_/A VGND VPWR _259_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_328_ _328_/A VGND VPWR clockp[0] VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_20_5 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xringosc.dstage\[10\].id.delayenb1 ringosc.dstage\[10\].id.delayenb1/A _333_/X VGND
+ VPWR ringosc.dstage\[10\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvn_4
Xringosc.dstage\[9\].id.delayenb1 ringosc.dstage\[9\].id.delayenb1/A _335_/X VGND
+ VPWR ringosc.dstage\[9\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvn_4
X_361_ _328_/A _361_/D _320_/X VGND VPWR _361_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_292_ _301_/A _292_/B VGND VPWR _299_/B VGND VPWR sky130_fd_sc_hd__nand2_2
X_275_ _267_/A _267_/B _360_/Q _359_/Q _272_/D VGND VPWR _276_/B VGND VPWR sky130_fd_sc_hd__o221a_2
X_344_ _286_/X ext_trim[4] dco VGND VPWR _344_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xringosc.dstage\[4\].id.delayen0 ringosc.dstage\[4\].id.delayen0/A _344_/X VGND VPWR
+ ringosc.dstage\[4\].id.delayen0/Z VGND VPWR sky130_fd_sc_hd__einvp_2
XFILLER_0_37 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_258_ _262_/A _262_/B VGND VPWR _258_/X VGND VPWR sky130_fd_sc_hd__or2_2
X_189_ _371_/Q _226_/B VGND VPWR _371_/D VGND VPWR sky130_fd_sc_hd__or2_2
X_327_ _327_/A VGND VPWR _327_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_15_67 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__210__B1 div[0] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xringosc.dstage\[5\].id.delayenb0 ringosc.dstage\[5\].id.delayenb1/A _342_/X VGND
+ VPWR ringosc.ibufp10/A VGND VPWR sky130_fd_sc_hd__einvn_8
Xringosc.dstage\[10\].id.delaybuf0 ringosc.dstage\[9\].id.delayen0/Z VGND VPWR ringosc.dstage\[10\].id.delayenb1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_2
Xringosc.dstage\[9\].id.delaybuf0 ringosc.dstage\[8\].id.delayen0/Z VGND VPWR ringosc.dstage\[9\].id.delayenb1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_2
XANTENNA__201__B1 div[2] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_7_90 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_360_ _328_/A _360_/D _321_/X VGND VPWR _360_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_291_ _369_/Q _368_/Q _367_/Q _370_/Q VGND VPWR _291_/X VGND VPWR sky130_fd_sc_hd__a31o_2
X_274_ _272_/D _268_/A _273_/Y _276_/A VGND VPWR _361_/D VGND VPWR sky130_fd_sc_hd__a31o_2
X_343_ _301_/Y ext_trim[18] dco VGND VPWR _343_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xringosc.dstage\[4\].id.delayen1 ringosc.dstage\[4\].id.delayen1/A _345_/X VGND VPWR
+ ringosc.dstage\[4\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvp_2
X_257_ _236_/A _251_/X _256_/Y _368_/Q _236_/Y VGND VPWR _368_/D VGND VPWR sky130_fd_sc_hd__a32o_2
X_188_ _372_/Q _272_/D _371_/Q _226_/B VGND VPWR _372_/D VGND VPWR sky130_fd_sc_hd__a22o_2
X_326_ _370_/Q VGND VPWR _326_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_309_ _327_/A VGND VPWR _309_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__210__A1 div[1] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xringosc.dstage\[5\].id.delayenb1 ringosc.dstage\[5\].id.delayenb1/A _343_/X VGND
+ VPWR ringosc.dstage\[5\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvn_4
XANTENNA__201__A1 div[3] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xringosc.dstage\[10\].id.delaybuf1 ringosc.dstage\[10\].id.delayenb1/A VGND VPWR ringosc.dstage\[10\].id.delayen1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xringosc.dstage\[9\].id.delaybuf1 ringosc.dstage\[9\].id.delayenb1/A VGND VPWR ringosc.dstage\[9\].id.delayen1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_290_ _369_/Q _368_/Q _297_/C _370_/Q VGND VPWR _290_/X VGND VPWR sky130_fd_sc_hd__a31o_2
X_273_ _267_/A _267_/B _267_/C VGND VPWR _273_/Y VGND VPWR sky130_fd_sc_hd__o21ai_2
X_342_ _283_/X ext_trim[5] dco VGND VPWR _342_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_4_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_187_ _372_/Q _226_/B _373_/Q _272_/D VGND VPWR _373_/D VGND VPWR sky130_fd_sc_hd__a22o_2
X_325_ _327_/A VGND VPWR _325_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_256_ _256_/A _256_/B VGND VPWR _256_/Y VGND VPWR sky130_fd_sc_hd__nand2_2
X_308_ _327_/A VGND VPWR _308_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_239_ _288_/A _239_/B VGND VPWR _239_/Y VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_6_38 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xringosc.dstage\[5\].id.delaybuf0 ringosc.dstage\[4\].id.delayen0/Z VGND VPWR ringosc.dstage\[5\].id.delayenb1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_2
X_272_ _362_/Q _272_/B _363_/Q _272_/D VGND VPWR _276_/A VGND VPWR sky130_fd_sc_hd__and4_2
Xringosc.dstage\[1\].id.delayenb0 ringosc.dstage\[1\].id.delayenb1/A _350_/X VGND
+ VPWR ringosc.dstage\[1\].id.delayen0/Z VGND VPWR sky130_fd_sc_hd__einvn_8
X_341_ _299_/B ext_trim[19] dco VGND VPWR _341_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xringosc.dstage\[8\].id.delayint0 ringosc.dstage\[8\].id.delayen1/Z VGND VPWR ringosc.dstage\[8\].id.delayen0/A
+ VGND VPWR sky130_fd_sc_hd__clkinv_1
XANTENNA__340__A1 ext_trim[6] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA__181__A enable VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA__331__A1 ext_trim[24] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_255_ _297_/A _236_/A _254_/X VGND VPWR _369_/D VGND VPWR sky130_fd_sc_hd__o21ai_2
X_186_ _374_/Q _272_/D _359_/Q _226_/B VGND VPWR _374_/D VGND VPWR sky130_fd_sc_hd__a22o_2
X_324_ _327_/A VGND VPWR _324_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_238_ _224_/A _220_/A _224_/B _237_/X VGND VPWR _262_/A VGND VPWR sky130_fd_sc_hd__o22a_2
X_307_ _327_/A VGND VPWR _307_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_169_ _374_/Q VGND VPWR _193_/B VGND VPWR sky130_fd_sc_hd__inv_2
XPHY_0 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xringosc.dstage\[1\].id.delayenb1 ringosc.dstage\[1\].id.delayenb1/A _351_/X VGND
+ VPWR ringosc.dstage\[1\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvn_4
Xringosc.dstage\[5\].id.delaybuf1 ringosc.dstage\[5\].id.delayenb1/A VGND VPWR ringosc.dstage\[5\].id.delayen1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_271_ _362_/Q _272_/B _363_/Q _269_/Y _272_/D VGND VPWR _362_/D VGND VPWR sky130_fd_sc_hd__o221a_2
X_340_ _279_/X ext_trim[6] dco VGND VPWR _340_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xringosc.dstage\[1\].id.delayen0 ringosc.dstage\[1\].id.delayen0/A _350_/X VGND VPWR
+ ringosc.dstage\[1\].id.delayen0/Z VGND VPWR sky130_fd_sc_hd__einvp_2
XANTENNA__181__B resetb VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_0_19 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_185_ _375_/Q _272_/D _360_/Q _226_/B VGND VPWR _375_/D VGND VPWR sky130_fd_sc_hd__a22o_2
X_254_ _244_/Y _253_/A _244_/A _253_/Y _236_/Y VGND VPWR _254_/X VGND VPWR sky130_fd_sc_hd__a221o_2
X_323_ _327_/A VGND VPWR _323_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_237_ _365_/Q _220_/Y _224_/A _220_/A VGND VPWR _237_/X VGND VPWR sky130_fd_sc_hd__a22o_2
X_306_ _327_/A VGND VPWR _306_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_168_ _359_/Q VGND VPWR _267_/B VGND VPWR sky130_fd_sc_hd__inv_2
XANTENNA__204__A1 div[2] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_16_115 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_270_ _164_/Y _269_/Y _226_/B VGND VPWR _363_/D VGND VPWR sky130_fd_sc_hd__a21oi_2
Xringosc.dstage\[1\].id.delayen1 ringosc.dstage\[1\].id.delayen1/A _351_/X VGND VPWR
+ ringosc.dstage\[1\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvp_2
X_322_ _327_/A VGND VPWR _322_/X VGND VPWR sky130_fd_sc_hd__buf_1
Xringosc.dstage\[1\].id.delaybuf0 ringosc.dstage\[0\].id.delayen0/Z VGND VPWR ringosc.dstage\[1\].id.delayenb1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_2
X_184_ _376_/Q _272_/D _361_/Q _226_/B VGND VPWR _376_/D VGND VPWR sky130_fd_sc_hd__a22o_2
Xringosc.dstage\[4\].id.delayint0 ringosc.dstage\[4\].id.delayen1/Z VGND VPWR ringosc.dstage\[4\].id.delayen0/A
+ VGND VPWR sky130_fd_sc_hd__clkinv_1
X_253_ _253_/A VGND VPWR _253_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_305_ _327_/A VGND VPWR _305_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_167_ _360_/Q VGND VPWR _267_/A VGND VPWR sky130_fd_sc_hd__inv_2
X_236_ _236_/A VGND VPWR _236_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_219_ _219_/A _219_/B VGND VPWR _220_/A VGND VPWR sky130_fd_sc_hd__or2_2
Xringosc.dstage\[9\].id.delayen0 ringosc.dstage\[9\].id.delayen0/A _334_/X VGND VPWR
+ ringosc.dstage\[9\].id.delayen0/Z VGND VPWR sky130_fd_sc_hd__einvp_2
XPHY_2 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__352__A1 ext_trim[0] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA__330__S dco VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA__343__A1 ext_trim[18] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA__334__A1 ext_trim[9] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA__356__D osc VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xringosc.dstage\[1\].id.delaybuf1 ringosc.dstage\[1\].id.delayenb1/A VGND VPWR ringosc.dstage\[1\].id.delayen1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_252_ _280_/B _220_/A _251_/X VGND VPWR _253_/A VGND VPWR sky130_fd_sc_hd__o21ai_2
X_183_ _377_/Q _272_/D _362_/Q _226_/B VGND VPWR _377_/D VGND VPWR sky130_fd_sc_hd__a22o_2
X_321_ _327_/A VGND VPWR _321_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_304_ _288_/A _239_/B _302_/B _370_/Q _232_/B VGND VPWR _304_/X VGND VPWR sky130_fd_sc_hd__o311a_2
X_235_ _301_/A _220_/Y _224_/X _234_/X VGND VPWR _236_/A VGND VPWR sky130_fd_sc_hd__o31a_2
X_166_ _361_/Q VGND VPWR _267_/C VGND VPWR sky130_fd_sc_hd__inv_2
XANTENNA__333__S dco VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_218_ _164_/Y _165_/Y div[4] _216_/B _214_/X VGND VPWR _219_/B VGND VPWR sky130_fd_sc_hd__o221ai_2
Xringosc.dstage\[9\].id.delayen1 ringosc.dstage\[9\].id.delayen1/A _335_/X VGND VPWR
+ ringosc.dstage\[9\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvp_2
XPHY_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_94 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__341__S dco VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_251_ _256_/A _256_/B VGND VPWR _251_/X VGND VPWR sky130_fd_sc_hd__or2_2
X_320_ _327_/A VGND VPWR _320_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__336__S dco VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_182_ dco _182_/B VGND VPWR _327_/A VGND VPWR sky130_fd_sc_hd__nor2_2
X_234_ _219_/B _225_/Y _220_/A _233_/X _226_/X VGND VPWR _234_/X VGND VPWR sky130_fd_sc_hd__o221a_2
X_303_ _297_/A _368_/Q _367_/Q _302_/X VGND VPWR _303_/X VGND VPWR sky130_fd_sc_hd__o31a_2
X_165_ _378_/Q VGND VPWR _165_/Y VGND VPWR sky130_fd_sc_hd__inv_2
Xringosc.dstage\[0\].id.delayint0 ringosc.dstage\[0\].id.delayen1/Z VGND VPWR ringosc.dstage\[0\].id.delayen0/A
+ VGND VPWR sky130_fd_sc_hd__clkinv_1
Xringosc.iss.reseten0 ringosc.iss.const1/HI _182_/B VGND VPWR ringosc.ibufp00/A VGND
+ VPWR sky130_fd_sc_hd__einvp_1
X_217_ _201_/Y _203_/Y _205_/Y _211_/Y _216_/Y VGND VPWR _219_/A VGND VPWR sky130_fd_sc_hd__o221a_2
XANTENNA__344__S dco VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XPHY_4 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__339__S dco VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xringosc.dstage\[8\].id.delayenb0 ringosc.dstage\[8\].id.delayenb1/A _336_/X VGND
+ VPWR ringosc.dstage\[8\].id.delayen0/Z VGND VPWR sky130_fd_sc_hd__einvn_8
X_250_ _301_/A _236_/A _249_/X VGND VPWR _370_/D VGND VPWR sky130_fd_sc_hd__o21ai_2
XANTENNA__352__S dco VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_181_ enable resetb VGND VPWR _182_/B VGND VPWR sky130_fd_sc_hd__nand2_2
X_233_ _365_/Q _364_/Q _233_/C VGND VPWR _233_/X VGND VPWR sky130_fd_sc_hd__or3_2
X_302_ _370_/Q _302_/B _302_/C VGND VPWR _302_/X VGND VPWR sky130_fd_sc_hd__and3_2
XANTENNA__347__S dco VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_164_ _363_/Q VGND VPWR _164_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_216_ div[4] _216_/B VGND VPWR _216_/Y VGND VPWR sky130_fd_sc_hd__nand2_2
Xringosc.iss.delayint0 ringosc.iss.delayen1/Z VGND VPWR ringosc.iss.delayen0/A VGND
+ VPWR sky130_fd_sc_hd__clkinv_1
XANTENNA__355__A1 ext_trim[25] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XPHY_5 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__346__A1 ext_trim[3] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA__337__A1 ext_trim[21] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA__355__S dco VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xringosc.dstage\[8\].id.delayenb1 ringosc.dstage\[8\].id.delayenb1/A _337_/X VGND
+ VPWR ringosc.dstage\[8\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvn_4
X_180_ _378_/Q _272_/D _363_/Q _226_/B VGND VPWR _378_/D VGND VPWR sky130_fd_sc_hd__a22o_2
X_378_ _328_/A _378_/D _327_/X VGND VPWR _378_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_232_ _370_/Q _232_/B VGND VPWR _233_/C VGND VPWR sky130_fd_sc_hd__or2_2
X_301_ _301_/A _301_/B VGND VPWR _301_/Y VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_10_10 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_215_ _214_/A _214_/B _214_/X VGND VPWR _216_/B VGND VPWR sky130_fd_sc_hd__a21bo_2
Xringosc.dstage\[6\].id.delayen0 ringosc.dstage\[6\].id.delayen0/A _340_/X VGND VPWR
+ ringosc.dstage\[6\].id.delayen0/Z VGND VPWR sky130_fd_sc_hd__einvp_2
XANTENNA__207__A div[1] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XPHY_6 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_377_ _328_/A _377_/D _327_/A VGND VPWR _377_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
Xringosc.dstage\[4\].id.delayenb0 ringosc.dstage\[4\].id.delayenb1/A _344_/X VGND
+ VPWR ringosc.dstage\[4\].id.delayen0/Z VGND VPWR sky130_fd_sc_hd__einvn_8
Xringosc.dstage\[8\].id.delaybuf0 ringosc.dstage\[7\].id.delayen0/Z VGND VPWR ringosc.dstage\[8\].id.delayenb1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_2
X_231_ _297_/C _302_/B VGND VPWR _232_/B VGND VPWR sky130_fd_sc_hd__or2_2
X_300_ _221_/A _366_/Q _301_/A _302_/C _296_/X VGND VPWR _300_/X VGND VPWR sky130_fd_sc_hd__o41a_2
Xringosc.dstage\[10\].id.delayen0 ringosc.dstage\[10\].id.delayen0/A _332_/X VGND
+ VPWR ringosc.dstage\[10\].id.delayen0/Z VGND VPWR sky130_fd_sc_hd__einvp_2
X_214_ _214_/A _214_/B VGND VPWR _214_/X VGND VPWR sky130_fd_sc_hd__or2_2
Xringosc.dstage\[6\].id.delayen1 ringosc.dstage\[6\].id.delayen1/A _341_/X VGND VPWR
+ ringosc.dstage\[6\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvp_2
XPHY_7 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_32 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_120 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_376_ _328_/A _376_/D _305_/X VGND VPWR _376_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
Xringosc.dstage\[4\].id.delayenb1 ringosc.dstage\[4\].id.delayenb1/A _345_/X VGND
+ VPWR ringosc.dstage\[4\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvn_4
Xringosc.dstage\[8\].id.delaybuf1 ringosc.dstage\[8\].id.delayenb1/A VGND VPWR ringosc.dstage\[8\].id.delayen1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_230_ _302_/B VGND VPWR _301_/B VGND VPWR sky130_fd_sc_hd__inv_2
X_359_ _328_/A _359_/D _322_/X VGND VPWR _359_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
Xringosc.dstage\[10\].id.delayen1 ringosc.dstage\[10\].id.delayen1/A _333_/X VGND
+ VPWR ringosc.dstage\[10\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvp_2
X_213_ _362_/Q _377_/Q _190_/Y _197_/X VGND VPWR _214_/B VGND VPWR sky130_fd_sc_hd__o2bb2a_2
XANTENNA__349__A1 ext_trim[15] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XPHY_8 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_375_ _328_/A _375_/D _306_/X VGND VPWR _375_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_358_ _328_/A _358_/D _323_/X VGND VPWR _358_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_289_ _297_/A _368_/Q _370_/Q _284_/X VGND VPWR _289_/X VGND VPWR sky130_fd_sc_hd__o31a_2
Xringosc.dstage\[4\].id.delaybuf0 ringosc.dstage\[3\].id.delayen0/Z VGND VPWR ringosc.dstage\[4\].id.delayenb1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_2
X_212_ _363_/Q _378_/Q _164_/Y _165_/Y VGND VPWR _214_/A VGND VPWR sky130_fd_sc_hd__a22o_2
Xringosc.dstage\[7\].id.delayint0 ringosc.dstage\[7\].id.delayen1/Z VGND VPWR ringosc.dstage\[7\].id.delayen0/A
+ VGND VPWR sky130_fd_sc_hd__clkinv_1
Xringosc.dstage\[0\].id.delayenb0 ringosc.dstage\[0\].id.delayenb1/A _352_/X VGND
+ VPWR ringosc.dstage\[0\].id.delayen0/Z VGND VPWR sky130_fd_sc_hd__einvn_8
XPHY_9 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_23 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_374_ _328_/A _374_/D _307_/X VGND VPWR _374_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_288_ _288_/A _288_/B VGND VPWR _288_/X VGND VPWR sky130_fd_sc_hd__or2_2
X_357_ _328_/A _357_/D _324_/X VGND VPWR _358_/D VGND VPWR sky130_fd_sc_hd__dfrtp_2
Xringosc.dstage\[3\].id.delayen0 ringosc.dstage\[3\].id.delayen0/A _346_/X VGND VPWR
+ ringosc.dstage\[3\].id.delayen0/Z VGND VPWR sky130_fd_sc_hd__einvp_2
XFILLER_10_36 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xringosc.dstage\[0\].id.delayenb1 ringosc.dstage\[0\].id.delayenb1/A _353_/X VGND
+ VPWR ringosc.dstage\[0\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvn_4
X_211_ div[1] _207_/B _210_/X VGND VPWR _211_/Y VGND VPWR sky130_fd_sc_hd__a21oi_2
Xringosc.dstage\[4\].id.delaybuf1 ringosc.dstage\[4\].id.delayenb1/A VGND VPWR ringosc.dstage\[4\].id.delayen1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xringosc.iss.delayenb0 ringosc.iss.delayenb1/A ringosc.iss.ctrlen0/X VGND VPWR ringosc.ibufp00/A
+ VGND VPWR sky130_fd_sc_hd__einvn_8
XANTENNA__330__A1 ext_trim[11] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_373_ _328_/A _373_/D _308_/X VGND VPWR _373_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_356_ _328_/A osc _325_/X VGND VPWR _357_/D VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_287_ _297_/A _368_/Q _370_/Q _288_/A _284_/X VGND VPWR _287_/X VGND VPWR sky130_fd_sc_hd__o41a_2
Xringosc.dstage\[3\].id.delayen1 ringosc.dstage\[3\].id.delayen1/A _347_/X VGND VPWR
+ ringosc.dstage\[3\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvp_2
X_210_ div[1] _207_/B div[0] _209_/Y _207_/Y VGND VPWR _210_/X VGND VPWR sky130_fd_sc_hd__o221a_2
X_339_ _303_/X ext_trim[20] dco VGND VPWR _339_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xringosc.iss.delayenb1 ringosc.iss.delayenb1/A _355_/X VGND VPWR ringosc.iss.delayen1/Z
+ VGND VPWR sky130_fd_sc_hd__einvn_4
Xringosc.dstage\[0\].id.delaybuf0 ringosc.ibufp00/A VGND VPWR ringosc.dstage\[0\].id.delayenb1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_2
Xringosc.dstage\[3\].id.delayint0 ringosc.dstage\[3\].id.delayen1/Z VGND VPWR ringosc.dstage\[3\].id.delayen0/A
+ VGND VPWR sky130_fd_sc_hd__clkinv_1
X_372_ _328_/A _372_/D _309_/X VGND VPWR _372_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XANTENNA__182__A dco VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_286_ _297_/A _368_/Q _370_/Q _367_/Q _284_/X VGND VPWR _286_/X VGND VPWR sky130_fd_sc_hd__o41a_2
X_355_ _304_/X ext_trim[25] dco VGND VPWR _355_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XANTENNA__177__A div[0] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_338_ _290_/X ext_trim[7] dco VGND VPWR _338_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_269_ _362_/Q _272_/B VGND VPWR _269_/Y VGND VPWR sky130_fd_sc_hd__nand2_2
Xringosc.dstage\[0\].id.delaybuf1 ringosc.dstage\[0\].id.delayenb1/A VGND VPWR ringosc.dstage\[0\].id.delayen1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_7_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_7 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_59 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xringosc.iss.delaybuf0 ringosc.iss.delayenb1/A VGND VPWR ringosc.iss.delayen1/A VGND
+ VPWR sky130_fd_sc_hd__clkbuf_1
X_371_ _328_/A _371_/D _310_/X VGND VPWR _371_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_14_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_285_ _297_/A _368_/Q _370_/Q _297_/C _284_/X VGND VPWR _285_/X VGND VPWR sky130_fd_sc_hd__o41a_2
X_354_ _282_/X ext_trim[12] dco VGND VPWR _354_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_199_ _361_/Q _376_/Q _192_/Y VGND VPWR _199_/Y VGND VPWR sky130_fd_sc_hd__a21oi_2
X_337_ _293_/X ext_trim[21] dco VGND VPWR _337_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_268_ _268_/A VGND VPWR _272_/B VGND VPWR sky130_fd_sc_hd__inv_2
XANTENNA__351__A1 ext_trim[14] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA__333__A1 ext_trim[23] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA__342__A1 ext_trim[5] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_370_ _328_/A _370_/D _311_/X VGND VPWR _370_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
Xringosc.dstage\[0\].id.delayen0 ringosc.dstage\[0\].id.delayen0/A _352_/X VGND VPWR
+ ringosc.dstage\[0\].id.delayen0/Z VGND VPWR sky130_fd_sc_hd__einvp_2
X_284_ _370_/Q _302_/C _288_/B VGND VPWR _284_/X VGND VPWR sky130_fd_sc_hd__o21a_2
X_353_ _291_/X ext_trim[13] dco VGND VPWR _353_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_267_ _267_/A _267_/B _267_/C VGND VPWR _268_/A VGND VPWR sky130_fd_sc_hd__or3_2
Xringosc.dstage\[7\].id.delayenb0 ringosc.dstage\[7\].id.delayenb1/A _338_/X VGND
+ VPWR ringosc.dstage\[7\].id.delayen0/Z VGND VPWR sky130_fd_sc_hd__einvn_8
X_198_ _191_/X _197_/X _191_/X _197_/X VGND VPWR _202_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_2
X_336_ _281_/X ext_trim[8] dco VGND VPWR _336_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_11_50 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_319_ _327_/A VGND VPWR _319_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_8_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__331__S dco VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xringosc.dstage\[0\].id.delayen1 ringosc.dstage\[0\].id.delayen1/A _353_/X VGND VPWR
+ ringosc.dstage\[0\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvp_2
X_283_ _370_/Q _302_/C _288_/A _288_/B VGND VPWR _283_/X VGND VPWR sky130_fd_sc_hd__o31a_2
X_352_ _233_/C ext_trim[0] dco VGND VPWR _352_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_10_19 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_197_ _361_/Q _376_/Q _192_/Y _196_/Y VGND VPWR _197_/X VGND VPWR sky130_fd_sc_hd__o2bb2a_2
X_266_ _364_/Q _236_/A _224_/B _236_/Y VGND VPWR _364_/D VGND VPWR sky130_fd_sc_hd__o22a_2
Xringosc.dstage\[7\].id.delayenb1 ringosc.dstage\[7\].id.delayenb1/A _339_/X VGND
+ VPWR ringosc.dstage\[7\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvn_4
X_335_ _296_/X ext_trim[22] dco VGND VPWR _335_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XANTENNA__334__S dco VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_249_ _246_/Y _248_/A _246_/A _248_/Y _236_/Y VGND VPWR _249_/X VGND VPWR sky130_fd_sc_hd__a221o_2
X_318_ _327_/A VGND VPWR _318_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_22_72 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xringosc.dstage\[8\].id.delayen0 ringosc.dstage\[8\].id.delayen0/A _336_/X VGND VPWR
+ ringosc.dstage\[8\].id.delayen0/Z VGND VPWR sky130_fd_sc_hd__einvp_2
XFILLER_8_63 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__342__S dco VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_282_ _370_/Q _302_/C _367_/Q _288_/B VGND VPWR _282_/X VGND VPWR sky130_fd_sc_hd__o31a_2
X_351_ _298_/X ext_trim[14] dco VGND VPWR _351_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XANTENNA__337__S dco VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_334_ _285_/X ext_trim[9] dco VGND VPWR _334_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_265_ _224_/A _236_/A _236_/Y _264_/X VGND VPWR _365_/D VGND VPWR sky130_fd_sc_hd__o22ai_2
X_196_ _196_/A VGND VPWR _196_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XANTENNA__354__A1 ext_trim[12] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_317_ _327_/A VGND VPWR _317_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__350__S dco VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA__345__A1 ext_trim[17] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_179_ _272_/D VGND VPWR _226_/B VGND VPWR sky130_fd_sc_hd__inv_2
X_248_ _248_/A VGND VPWR _248_/Y VGND VPWR sky130_fd_sc_hd__inv_2
Xringosc.dstage\[3\].id.delayenb0 ringosc.dstage\[3\].id.delayenb1/A _346_/X VGND
+ VPWR ringosc.dstage\[3\].id.delayen0/Z VGND VPWR sky130_fd_sc_hd__einvn_8
Xringosc.dstage\[7\].id.delaybuf0 ringosc.dstage\[6\].id.delayen0/Z VGND VPWR ringosc.dstage\[7\].id.delayenb1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_2
XANTENNA__336__A1 ext_trim[8] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xringosc.dstage\[11\].id.delayint0 ringosc.dstage\[11\].id.delayen1/Z VGND VPWR ringosc.dstage\[11\].id.delayen0/A
+ VGND VPWR sky130_fd_sc_hd__clkinv_1
XANTENNA__345__S dco VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xringosc.dstage\[8\].id.delayen1 ringosc.dstage\[8\].id.delayen1/A _337_/X VGND VPWR
+ ringosc.dstage\[8\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvp_2
XFILLER_4_129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__218__B1 div[4] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_5_32 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_63 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_281_ _297_/C _302_/C _370_/Q _288_/B VGND VPWR _281_/X VGND VPWR sky130_fd_sc_hd__o31a_2
X_350_ _289_/X ext_trim[1] dco VGND VPWR _350_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XANTENNA__353__S dco VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA__202__A div[3] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA__348__S dco VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XPHY_40 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_195_ _360_/Q _375_/Q _193_/Y _194_/X VGND VPWR _196_/A VGND VPWR sky130_fd_sc_hd__a22o_2
X_264_ _224_/B _237_/X _224_/B _237_/X VGND VPWR _264_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_2
X_333_ _326_/X ext_trim[23] dco VGND VPWR _333_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_15_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_247_ _370_/Q _220_/Y _301_/A _220_/A VGND VPWR _248_/A VGND VPWR sky130_fd_sc_hd__o22a_2
X_316_ _327_/A VGND VPWR _316_/X VGND VPWR sky130_fd_sc_hd__buf_1
Xringosc.dstage\[3\].id.delayenb1 ringosc.dstage\[3\].id.delayenb1/A _347_/X VGND
+ VPWR ringosc.dstage\[3\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvn_4
X_178_ _358_/D _358_/Q _358_/D _358_/Q VGND VPWR _272_/D VGND VPWR sky130_fd_sc_hd__a2bb2o_2
Xringosc.dstage\[7\].id.delaybuf1 ringosc.dstage\[7\].id.delayenb1/A VGND VPWR ringosc.dstage\[7\].id.delayen1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_7_116 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_127 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_30 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_280_ _369_/Q _280_/B VGND VPWR _302_/C VGND VPWR sky130_fd_sc_hd__or2_2
XPHY_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_30 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_78 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_263_ _236_/A _258_/X _262_/Y _366_/Q _236_/Y VGND VPWR _366_/D VGND VPWR sky130_fd_sc_hd__a32o_2
X_194_ _360_/Q _375_/Q _360_/Q _375_/Q VGND VPWR _194_/X VGND VPWR sky130_fd_sc_hd__o2bb2a_2
X_332_ _288_/X ext_trim[10] dco VGND VPWR _332_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_315_ _327_/A VGND VPWR _315_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_177_ div[0] VGND VPWR _177_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_246_ _246_/A VGND VPWR _246_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_22_31 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_229_ _369_/Q _368_/Q VGND VPWR _302_/B VGND VPWR sky130_fd_sc_hd__or2_2
Xringosc.dstage\[3\].id.delaybuf0 ringosc.dstage\[2\].id.delayen0/Z VGND VPWR ringosc.dstage\[3\].id.delayenb1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_2
Xringosc.dstage\[6\].id.delayint0 ringosc.dstage\[6\].id.delayen1/Z VGND VPWR ringosc.dstage\[6\].id.delayen0/A
+ VGND VPWR sky130_fd_sc_hd__clkinv_1
XFILLER_14_43 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xringosc.ibufp10 ringosc.ibufp10/A VGND VPWR ringosc.ibufp11/A VGND VPWR sky130_fd_sc_hd__clkinv_2
XANTENNA__216__A div[4] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XPHY_42 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_331_ _302_/X ext_trim[24] dco VGND VPWR _331_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_193_ _267_/B _193_/B VGND VPWR _193_/Y VGND VPWR sky130_fd_sc_hd__nor2_2
X_262_ _262_/A _262_/B VGND VPWR _262_/Y VGND VPWR sky130_fd_sc_hd__nand2_2
XANTENNA__348__A1 ext_trim[2] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA__339__A1 ext_trim[20] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_245_ _256_/B _244_/A _256_/A _220_/A _301_/B VGND VPWR _246_/A VGND VPWR sky130_fd_sc_hd__o32a_2
X_314_ _327_/A VGND VPWR _314_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_176_ _364_/Q VGND VPWR _224_/B VGND VPWR sky130_fd_sc_hd__inv_2
Xringosc.dstage\[5\].id.delayen0 ringosc.dstage\[5\].id.delayen0/A _342_/X VGND VPWR
+ ringosc.ibufp10/A VGND VPWR sky130_fd_sc_hd__einvp_2
Xringosc.dstage\[3\].id.delaybuf1 ringosc.dstage\[3\].id.delayenb1/A VGND VPWR ringosc.dstage\[3\].id.delayen1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_228_ _297_/C VGND VPWR _239_/B VGND VPWR sky130_fd_sc_hd__inv_2
Xringosc.ibufp00 ringosc.ibufp00/A VGND VPWR ringosc.ibufp01/A VGND VPWR sky130_fd_sc_hd__clkinv_2
Xringosc.ibufp11 ringosc.ibufp11/A VGND VPWR clockp[1] VGND VPWR sky130_fd_sc_hd__clkinv_8
XPHY_43 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_261_ _367_/Q _260_/X _367_/Q _260_/X VGND VPWR _367_/D VGND VPWR sky130_fd_sc_hd__o2bb2a_2
X_330_ _287_/X ext_trim[11] dco VGND VPWR _330_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_192_ _361_/Q _376_/Q VGND VPWR _192_/Y VGND VPWR sky130_fd_sc_hd__nor2_2
X_313_ _327_/A VGND VPWR _313_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_175_ _365_/Q VGND VPWR _224_/A VGND VPWR sky130_fd_sc_hd__inv_2
X_244_ _244_/A VGND VPWR _244_/Y VGND VPWR sky130_fd_sc_hd__inv_2
Xringosc.dstage\[5\].id.delayen1 ringosc.dstage\[5\].id.delayen1/A _343_/X VGND VPWR
+ ringosc.dstage\[5\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvp_2
X_227_ _367_/Q _366_/Q VGND VPWR _297_/C VGND VPWR sky130_fd_sc_hd__or2_2
Xringosc.dstage\[2\].id.delayint0 ringosc.dstage\[2\].id.delayen1/Z VGND VPWR ringosc.dstage\[2\].id.delayen0/A
+ VGND VPWR sky130_fd_sc_hd__clkinv_1
Xringosc.ibufp01 ringosc.ibufp01/A VGND VPWR _328_/A VGND VPWR sky130_fd_sc_hd__clkinv_8
XPHY_44 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_260_ _221_/B _220_/A _236_/A _259_/X VGND VPWR _260_/X VGND VPWR sky130_fd_sc_hd__o211a_2
X_191_ _362_/Q _377_/Q _190_/Y VGND VPWR _191_/X VGND VPWR sky130_fd_sc_hd__a21o_2
X_243_ _297_/A _220_/Y _369_/Q _220_/A VGND VPWR _244_/A VGND VPWR sky130_fd_sc_hd__o22a_2
X_312_ _327_/A VGND VPWR _312_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_174_ _366_/Q VGND VPWR _221_/B VGND VPWR sky130_fd_sc_hd__inv_2
X_226_ _372_/Q _226_/B _373_/Q _371_/Q VGND VPWR _226_/X VGND VPWR sky130_fd_sc_hd__and4_2
Xringosc.dstage\[11\].id.delayenb0 ringosc.dstage\[11\].id.delayenb1/A _330_/X VGND
+ VPWR ringosc.iss.delayenb1/A VGND VPWR sky130_fd_sc_hd__einvn_8
XFILLER_17_12 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_209_ _209_/A VGND VPWR _209_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XPHY_12 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_190_ _362_/Q _377_/Q VGND VPWR _190_/Y VGND VPWR sky130_fd_sc_hd__nor2_2
X_242_ _368_/Q _220_/Y _280_/B _220_/A VGND VPWR _256_/B VGND VPWR sky130_fd_sc_hd__a22o_2
X_311_ _327_/A VGND VPWR _311_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_173_ _367_/Q VGND VPWR _221_/A VGND VPWR sky130_fd_sc_hd__inv_2
X_225_ _177_/Y _209_/A _210_/X _205_/A _216_/Y VGND VPWR _225_/Y VGND VPWR sky130_fd_sc_hd__o2111ai_2
Xringosc.dstage\[11\].id.delayenb1 ringosc.dstage\[11\].id.delayenb1/A _331_/X VGND
+ VPWR ringosc.dstage\[11\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvn_4
XFILLER_0_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_208_ _267_/B _193_/B _193_/Y VGND VPWR _209_/A VGND VPWR sky130_fd_sc_hd__a21oi_2
XFILLER_0_105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_35 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_13 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__211__A1 div[1] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_310_ _327_/A VGND VPWR _310_/X VGND VPWR sky130_fd_sc_hd__buf_1
Xringosc.iss.const1 VGND VGND VPWR VPWR ringosc.iss.const1/HI ringosc.iss.const1/LO
+ sky130_fd_sc_hd__conb_1
X_241_ _239_/Y _262_/B _262_/A _220_/A _239_/B VGND VPWR _256_/A VGND VPWR sky130_fd_sc_hd__o32a_2
Xringosc.dstage\[2\].id.delayen0 ringosc.dstage\[2\].id.delayen0/A _348_/X VGND VPWR
+ ringosc.dstage\[2\].id.delayen0/Z VGND VPWR sky130_fd_sc_hd__einvp_2
X_172_ _368_/Q VGND VPWR _280_/B VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_6_100 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_122 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_224_ _224_/A _224_/B _292_/B VGND VPWR _224_/X VGND VPWR sky130_fd_sc_hd__or3_2
Xringosc.dstage\[6\].id.delayenb0 ringosc.dstage\[6\].id.delayenb1/A _340_/X VGND
+ VPWR ringosc.dstage\[6\].id.delayen0/Z VGND VPWR sky130_fd_sc_hd__einvn_8
Xringosc.dstage\[11\].id.delaybuf0 ringosc.dstage\[10\].id.delayen0/Z VGND VPWR ringosc.dstage\[11\].id.delayenb1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_2
X_207_ div[1] _207_/B VGND VPWR _207_/Y VGND VPWR sky130_fd_sc_hd__nand2_2
XFILLER_6_71 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_36 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_38 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_240_ _366_/Q _220_/Y _221_/B _220_/A VGND VPWR _262_/B VGND VPWR sky130_fd_sc_hd__a22o_2
Xringosc.dstage\[2\].id.delayen1 ringosc.dstage\[2\].id.delayen1/A _349_/X VGND VPWR
+ ringosc.dstage\[2\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvp_2
X_171_ _369_/Q VGND VPWR _297_/A VGND VPWR sky130_fd_sc_hd__inv_2
X_369_ _328_/A _369_/D _312_/X VGND VPWR _369_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_223_ _297_/A _280_/B _223_/C VGND VPWR _292_/B VGND VPWR sky130_fd_sc_hd__or3_2
XANTENNA__350__A1 ext_trim[1] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA__341__A1 ext_trim[19] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA__332__A1 ext_trim[10] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_206_ _193_/Y _194_/X _193_/Y _194_/X VGND VPWR _207_/B VGND VPWR sky130_fd_sc_hd__o2bb2ai_2
Xringosc.dstage\[6\].id.delayenb1 ringosc.dstage\[6\].id.delayenb1/A _341_/X VGND
+ VPWR ringosc.dstage\[6\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvn_4
Xringosc.dstage\[11\].id.delaybuf1 ringosc.dstage\[11\].id.delayenb1/A VGND VPWR ringosc.dstage\[11\].id.delayen1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_37 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xringosc.iss.delayen0 ringosc.iss.delayen0/A _354_/X VGND VPWR ringosc.ibufp00/A VGND
+ VPWR sky130_fd_sc_hd__einvp_2
X_170_ _370_/Q VGND VPWR _301_/A VGND VPWR sky130_fd_sc_hd__inv_2
X_368_ _328_/A _368_/D _313_/X VGND VPWR _368_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_299_ _329_/X _299_/B VGND VPWR _299_/X VGND VPWR sky130_fd_sc_hd__and2_2
X_222_ _223_/C VGND VPWR _288_/A VGND VPWR sky130_fd_sc_hd__inv_2
X_205_ _205_/A VGND VPWR _205_/Y VGND VPWR sky130_fd_sc_hd__inv_2
Xringosc.dstage\[2\].id.delayenb0 ringosc.dstage\[2\].id.delayenb1/A _348_/X VGND
+ VPWR ringosc.dstage\[2\].id.delayen0/Z VGND VPWR sky130_fd_sc_hd__einvn_8
Xringosc.dstage\[6\].id.delaybuf0 ringosc.ibufp10/A VGND VPWR ringosc.dstage\[6\].id.delayenb1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_2
Xringosc.dstage\[10\].id.delayint0 ringosc.dstage\[10\].id.delayen1/Z VGND VPWR ringosc.dstage\[10\].id.delayen0/A
+ VGND VPWR sky130_fd_sc_hd__clkinv_1
Xringosc.dstage\[9\].id.delayint0 ringosc.dstage\[9\].id.delayen1/Z VGND VPWR ringosc.dstage\[9\].id.delayen0/A
+ VGND VPWR sky130_fd_sc_hd__clkinv_1
XFILLER_6_62 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_38 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xringosc.iss.delayen1 ringosc.iss.delayen1/A _355_/X VGND VPWR ringosc.iss.delayen1/Z
+ VGND VPWR sky130_fd_sc_hd__einvp_2
XFILLER_15_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_298_ _301_/A _302_/C _221_/A _297_/X _296_/X VGND VPWR _298_/X VGND VPWR sky130_fd_sc_hd__o311a_2
X_367_ _328_/A _367_/D _314_/X VGND VPWR _367_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_221_ _221_/A _221_/B VGND VPWR _223_/C VGND VPWR sky130_fd_sc_hd__or2_2
X_204_ div[2] _200_/X _203_/A _201_/Y VGND VPWR _205_/A VGND VPWR sky130_fd_sc_hd__o211a_2
XANTENNA__332__S dco VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_22_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xringosc.dstage\[2\].id.delayenb1 ringosc.dstage\[2\].id.delayenb1/A _349_/X VGND
+ VPWR ringosc.dstage\[2\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvn_4
Xringosc.dstage\[6\].id.delaybuf1 ringosc.dstage\[6\].id.delayenb1/A VGND VPWR ringosc.dstage\[6\].id.delayen1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_1
XPHY_28 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__353__A1 ext_trim[13] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_297_ _297_/A _368_/Q _297_/C _301_/A VGND VPWR _297_/X VGND VPWR sky130_fd_sc_hd__or4_2
X_366_ _328_/A _366_/D _315_/X VGND VPWR _366_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XANTENNA__344__A1 ext_trim[4] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA__340__S dco VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA__335__A1 ext_trim[22] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA__335__S dco VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_220_ _220_/A VGND VPWR _220_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_349_ _295_/X ext_trim[15] dco VGND VPWR _349_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_203_ _203_/A VGND VPWR _203_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_10 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xringosc.iss.ctrlen0 _182_/B _354_/X VGND VPWR ringosc.iss.ctrlen0/X VGND VPWR sky130_fd_sc_hd__or2_2
XANTENNA__343__S dco VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_6_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xringosc.dstage\[2\].id.delaybuf0 ringosc.dstage\[1\].id.delayen0/Z VGND VPWR ringosc.dstage\[2\].id.delayenb1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_2
Xringosc.dstage\[5\].id.delayint0 ringosc.dstage\[5\].id.delayen1/Z VGND VPWR ringosc.dstage\[5\].id.delayen0/A
+ VGND VPWR sky130_fd_sc_hd__clkinv_1
XANTENNA__338__S dco VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_365_ _328_/A _365_/D _316_/X VGND VPWR _365_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_296_ _367_/Q _221_/B _302_/C _301_/A _295_/X VGND VPWR _296_/X VGND VPWR sky130_fd_sc_hd__o41a_2
XANTENNA__351__S dco VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_279_ _367_/Q _288_/B VGND VPWR _279_/X VGND VPWR sky130_fd_sc_hd__or2_2
X_348_ _284_/X ext_trim[2] dco VGND VPWR _348_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_202_ div[3] _202_/B VGND VPWR _203_/A VGND VPWR sky130_fd_sc_hd__or2_2
XANTENNA__346__S dco VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xringosc.dstage\[7\].id.delayen0 ringosc.dstage\[7\].id.delayen0/A _338_/X VGND VPWR
+ ringosc.dstage\[7\].id.delayen0/Z VGND VPWR sky130_fd_sc_hd__einvp_2
XPHY_19 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xringosc.dstage\[2\].id.delaybuf1 ringosc.dstage\[2\].id.delayenb1/A VGND VPWR ringosc.dstage\[2\].id.delayen1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__354__S dco VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA__349__S dco VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_3_33 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_295_ _301_/A _302_/B _221_/A _294_/X _293_/X VGND VPWR _295_/X VGND VPWR sky130_fd_sc_hd__o311a_2
X_364_ _328_/A _364_/D _317_/X VGND VPWR _364_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_278_ _370_/Q _302_/B VGND VPWR _288_/B VGND VPWR sky130_fd_sc_hd__or2_2
X_347_ _299_/X ext_trim[16] dco VGND VPWR _347_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_201_ div[3] _202_/B div[2] _200_/X VGND VPWR _201_/Y VGND VPWR sky130_fd_sc_hd__a22oi_2
XFILLER_9_87 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xringosc.dstage\[11\].id.delayen0 ringosc.dstage\[11\].id.delayen0/A _330_/X VGND
+ VPWR ringosc.iss.delayenb1/A VGND VPWR sky130_fd_sc_hd__einvp_2
Xringosc.dstage\[7\].id.delayen1 ringosc.dstage\[7\].id.delayen1/A _339_/X VGND VPWR
+ ringosc.dstage\[7\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvp_2
XFILLER_15_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__347__A1 ext_trim[16] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
.ends

* Black-box entry subcircuit for sky130_ef_io__com_bus_slice_5um abstract view
.subckt sky130_ef_io__com_bus_slice_5um AMUXBUS_A AMUXBUS_B VSSA VDDA VSWITCH VDDIO_Q
+ VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
.ends

* Black-box entry subcircuit for sky130_ef_io__com_bus_slice_10um abstract view
.subckt sky130_ef_io__com_bus_slice_10um AMUXBUS_A AMUXBUS_B VSSA VDDA VSWITCH VDDIO_Q
+ VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
.ends

* Black-box entry subcircuit for sky130_ef_io__com_bus_slice_20um abstract view
.subckt sky130_ef_io__com_bus_slice_20um AMUXBUS_A AMUXBUS_B VSSA VDDA VSWITCH VDDIO_Q
+ VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
.ends

* Black-box entry subcircuit for sky130_ef_io__gpiov2_pad_wrapped abstract view
.subckt sky130_ef_io__gpiov2_pad_wrapped IN_H PAD_A_NOESD_H PAD_A_ESD_0_H PAD_A_ESD_1_H
+ PAD DM[2] DM[1] DM[0] HLD_H_N IN INP_DIS IB_MODE_SEL ENABLE_H ENABLE_VDDA_H ENABLE_INP_H
+ OE_N TIE_HI_ESD TIE_LO_ESD SLOW VTRIP_SEL HLD_OVR ANALOG_EN ANALOG_SEL ENABLE_VDDIO
+ ENABLE_VSWITCH_H ANALOG_POL OUT AMUXBUS_A AMUXBUS_B VSSA VDDA VSWITCH VDDIO_Q VCCHIB
+ VDDIO VCCD VSSIO VSSD VSSIO_Q
.ends

* Black-box entry subcircuit for sky130_ef_io__com_bus_slice_1um abstract view
.subckt sky130_ef_io__com_bus_slice_1um AMUXBUS_A AMUXBUS_B VSSA VDDA VSWITCH VDDIO_Q
+ VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
.ends

* Black-box entry subcircuit for sky130_ef_io__vccd_lvc_clamped_pad abstract view
.subckt sky130_ef_io__vccd_lvc_clamped_pad AMUXBUS_A AMUXBUS_B VCCD_PAD VSSA VDDA
+ VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
.ends

* Black-box entry subcircuit for sky130_ef_io__disconnect_vdda_slice_5um abstract view
.subckt sky130_ef_io__disconnect_vdda_slice_5um AMUXBUS_A AMUXBUS_B VSWITCH VDDIO_Q
+ VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
.ends

* Black-box entry subcircuit for sky130_ef_io__corner_pad abstract view
.subckt sky130_ef_io__corner_pad AMUXBUS_A AMUXBUS_B VSSA VDDA VSWITCH VDDIO_Q VCCHIB
+ VDDIO VCCD VSSIO VSSD VSSIO_Q
.ends

* Black-box entry subcircuit for sky130_ef_io__vddio_hvc_clamped_pad abstract view
.subckt sky130_ef_io__vddio_hvc_clamped_pad AMUXBUS_A AMUXBUS_B VDDIO_PAD VSSA VDDA
+ VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
.ends

* Black-box entry subcircuit for sky130_ef_io__vssio_hvc_clamped_pad abstract view
.subckt sky130_ef_io__vssio_hvc_clamped_pad AMUXBUS_A AMUXBUS_B VSSIO_PAD VSSA VDDA
+ VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
.ends

* Black-box entry subcircuit for sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um abstract view
.subckt sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um AMUXBUS_A AMUXBUS_B
+ VSSA VDDA VDDIO_Q VDDIO VCCD VSSIO VSSD VSSIO_Q VSWITCH VCCHIB
.ends

* Black-box entry subcircuit for sky130_ef_io__vdda_hvc_clamped_pad abstract view
.subckt sky130_ef_io__vdda_hvc_clamped_pad AMUXBUS_A AMUXBUS_B VDDA_PAD VSSA VDDA
+ VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
.ends

* Black-box entry subcircuit for sky130_ef_io__vssd_lvc_clamped3_pad abstract view
.subckt sky130_ef_io__vssd_lvc_clamped3_pad AMUXBUS_A AMUXBUS_B VSSD_PAD VSSA VDDA
+ VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q VCCD1 VSSD1
.ends

* Black-box entry subcircuit for sky130_ef_io__vssd_lvc_clamped_pad abstract view
.subckt sky130_ef_io__vssd_lvc_clamped_pad AMUXBUS_A AMUXBUS_B VSSD_PAD VSSA VDDA
+ VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
.ends

* Black-box entry subcircuit for sky130_ef_io__vccd_lvc_clamped3_pad abstract view
.subckt sky130_ef_io__vccd_lvc_clamped3_pad AMUXBUS_A AMUXBUS_B VCCD_PAD VSSA VDDA
+ VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q VCCD1 VSSD1
.ends

* Black-box entry subcircuit for sky130_ef_io__vssa_hvc_clamped_pad abstract view
.subckt sky130_ef_io__vssa_hvc_clamped_pad AMUXBUS_A AMUXBUS_B VSSA_PAD VSSA VDDA
+ VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
.ends

* Black-box entry subcircuit for sky130_fd_io__top_xres4v2 abstract view
.subckt sky130_fd_io__top_xres4v2 PAD_A_ESD_H XRES_H_N FILT_IN_H ENABLE_VDDIO TIE_WEAK_HI_H
+ ENABLE_H PULLUP_H EN_VDDIO_SIG_H TIE_LO_ESD TIE_HI_ESD DISABLE_PULLUP_H INP_SEL_H
+ VSSIO VSSA VSSD AMUXBUS_B AMUXBUS_A VDDIO_Q VDDIO VSWITCH VDDA VCCD VCCHIB VSSIO_Q
+ PAD
.ends

.subckt chip_io clock clock_core por flash_clk flash_clk_core flash_clk_ieb_core flash_clk_oeb_core
+ flash_csb flash_csb_core flash_csb_ieb_core flash_csb_oeb_core flash_io0 flash_io0_di_core
+ flash_io0_do_core flash_io0_oeb_core flash_io1 flash_io1_di_core flash_io1_do_core
+ flash_io1_oeb_core gpio gpio_in_core gpio_inenb_core gpio_mode0_core gpio_mode1_core
+ gpio_out_core gpio_outenb_core vccd_pad vdda_pad vddio_pad vddio_pad2 vssa_pad vssd_pad
+ vssio_pad vssio_pad2 mprj_io[0] mprj_io_analog_en[0] mprj_io_analog_pol[0] mprj_io_analog_sel[0]
+ mprj_io_dm[0] mprj_io_dm[1] mprj_io_dm[2] mprj_io_holdover[0] mprj_io_ib_mode_sel[0]
+ mprj_io_inp_dis[0] mprj_io_oeb[0] mprj_io_out[0] mprj_io_slow_sel[0] mprj_io_vtrip_sel[0]
+ mprj_io_in[0] mprj_analog_io[3] mprj_io[10] mprj_io_analog_en[10] mprj_io_analog_pol[10]
+ mprj_io_analog_sel[10] mprj_io_dm[30] mprj_io_dm[31] mprj_io_dm[32] mprj_io_holdover[10]
+ mprj_io_ib_mode_sel[10] mprj_io_inp_dis[10] mprj_io_oeb[10] mprj_io_out[10] mprj_io_slow_sel[10]
+ mprj_io_vtrip_sel[10] mprj_io_in[10] mprj_analog_io[4] mprj_io[11] mprj_io_analog_en[11]
+ mprj_io_analog_pol[11] mprj_io_analog_sel[11] mprj_io_dm[33] mprj_io_dm[34] mprj_io_dm[35]
+ mprj_io_holdover[11] mprj_io_ib_mode_sel[11] mprj_io_inp_dis[11] mprj_io_oeb[11]
+ mprj_io_out[11] mprj_io_slow_sel[11] mprj_io_vtrip_sel[11] mprj_io_in[11] mprj_analog_io[5]
+ mprj_io[12] mprj_io_analog_en[12] mprj_io_analog_pol[12] mprj_io_analog_sel[12]
+ mprj_io_dm[36] mprj_io_dm[37] mprj_io_dm[38] mprj_io_holdover[12] mprj_io_ib_mode_sel[12]
+ mprj_io_inp_dis[12] mprj_io_oeb[12] mprj_io_out[12] mprj_io_slow_sel[12] mprj_io_vtrip_sel[12]
+ mprj_io_in[12] mprj_analog_io[6] mprj_io[13] mprj_io_analog_en[13] mprj_io_analog_pol[13]
+ mprj_io_analog_sel[13] mprj_io_dm[39] mprj_io_dm[40] mprj_io_dm[41] mprj_io_holdover[13]
+ mprj_io_ib_mode_sel[13] mprj_io_inp_dis[13] mprj_io_oeb[13] mprj_io_out[13] mprj_io_slow_sel[13]
+ mprj_io_vtrip_sel[13] mprj_io_in[13] mprj_analog_io[7] mprj_io[14] mprj_io_analog_en[14]
+ mprj_io_analog_pol[14] mprj_io_analog_sel[14] mprj_io_dm[42] mprj_io_dm[43] mprj_io_dm[44]
+ mprj_io_holdover[14] mprj_io_ib_mode_sel[14] mprj_io_inp_dis[14] mprj_io_oeb[14]
+ mprj_io_out[14] mprj_io_slow_sel[14] mprj_io_vtrip_sel[14] mprj_io_in[14] mprj_analog_io[8]
+ mprj_io[15] mprj_io_analog_en[15] mprj_io_analog_pol[15] mprj_io_analog_sel[15]
+ mprj_io_dm[45] mprj_io_dm[46] mprj_io_dm[47] mprj_io_holdover[15] mprj_io_ib_mode_sel[15]
+ mprj_io_inp_dis[15] mprj_io_oeb[15] mprj_io_out[15] mprj_io_slow_sel[15] mprj_io_vtrip_sel[15]
+ mprj_io_in[15] mprj_analog_io[9] mprj_io[16] mprj_io_analog_en[16] mprj_io_analog_pol[16]
+ mprj_io_analog_sel[16] mprj_io_dm[48] mprj_io_dm[49] mprj_io_dm[50] mprj_io_holdover[16]
+ mprj_io_ib_mode_sel[16] mprj_io_inp_dis[16] mprj_io_oeb[16] mprj_io_out[16] mprj_io_slow_sel[16]
+ mprj_io_vtrip_sel[16] mprj_io_in[16] mprj_analog_io[10] mprj_io[17] mprj_io_analog_en[17]
+ mprj_io_analog_pol[17] mprj_io_analog_sel[17] mprj_io_dm[51] mprj_io_dm[52] mprj_io_dm[53]
+ mprj_io_holdover[17] mprj_io_ib_mode_sel[17] mprj_io_inp_dis[17] mprj_io_oeb[17]
+ mprj_io_out[17] mprj_io_slow_sel[17] mprj_io_vtrip_sel[17] mprj_io_in[17] mprj_analog_io[11]
+ mprj_io[18] mprj_io_analog_en[18] mprj_io_analog_pol[18] mprj_io_analog_sel[18]
+ mprj_io_dm[54] mprj_io_dm[55] mprj_io_dm[56] mprj_io_holdover[18] mprj_io_ib_mode_sel[18]
+ mprj_io_inp_dis[18] mprj_io_oeb[18] mprj_io_out[18] mprj_io_slow_sel[18] mprj_io_vtrip_sel[18]
+ mprj_io_in[18] mprj_io[1] mprj_io_analog_en[1] mprj_io_analog_pol[1] mprj_io_analog_sel[1]
+ mprj_io_dm[3] mprj_io_dm[4] mprj_io_dm[5] mprj_io_holdover[1] mprj_io_ib_mode_sel[1]
+ mprj_io_inp_dis[1] mprj_io_oeb[1] mprj_io_out[1] mprj_io_slow_sel[1] mprj_io_vtrip_sel[1]
+ mprj_io_in[1] mprj_io[2] mprj_io_analog_en[2] mprj_io_analog_pol[2] mprj_io_analog_sel[2]
+ mprj_io_dm[6] mprj_io_dm[7] mprj_io_dm[8] mprj_io_holdover[2] mprj_io_ib_mode_sel[2]
+ mprj_io_inp_dis[2] mprj_io_oeb[2] mprj_io_out[2] mprj_io_slow_sel[2] mprj_io_vtrip_sel[2]
+ mprj_io_in[2] mprj_io[3] mprj_io_analog_en[3] mprj_io_analog_pol[3] mprj_io_analog_sel[3]
+ mprj_io_dm[10] mprj_io_dm[11] mprj_io_dm[9] mprj_io_holdover[3] mprj_io_ib_mode_sel[3]
+ mprj_io_inp_dis[3] mprj_io_oeb[3] mprj_io_out[3] mprj_io_slow_sel[3] mprj_io_vtrip_sel[3]
+ mprj_io_in[3] mprj_io[4] mprj_io_analog_en[4] mprj_io_analog_pol[4] mprj_io_analog_sel[4]
+ mprj_io_dm[12] mprj_io_dm[13] mprj_io_dm[14] mprj_io_holdover[4] mprj_io_ib_mode_sel[4]
+ mprj_io_inp_dis[4] mprj_io_oeb[4] mprj_io_out[4] mprj_io_slow_sel[4] mprj_io_vtrip_sel[4]
+ mprj_io_in[4] mprj_io[5] mprj_io_analog_en[5] mprj_io_analog_pol[5] mprj_io_analog_sel[5]
+ mprj_io_dm[15] mprj_io_dm[16] mprj_io_dm[17] mprj_io_holdover[5] mprj_io_ib_mode_sel[5]
+ mprj_io_inp_dis[5] mprj_io_oeb[5] mprj_io_out[5] mprj_io_slow_sel[5] mprj_io_vtrip_sel[5]
+ mprj_io_in[5] mprj_io[6] mprj_io_analog_en[6] mprj_io_analog_pol[6] mprj_io_analog_sel[6]
+ mprj_io_dm[18] mprj_io_dm[19] mprj_io_dm[20] mprj_io_holdover[6] mprj_io_ib_mode_sel[6]
+ mprj_io_inp_dis[6] mprj_io_oeb[6] mprj_io_out[6] mprj_io_slow_sel[6] mprj_io_vtrip_sel[6]
+ mprj_io_in[6] mprj_analog_io[0] mprj_io[7] mprj_io_analog_en[7] mprj_io_analog_pol[7]
+ mprj_io_analog_sel[7] mprj_io_dm[21] mprj_io_dm[22] mprj_io_dm[23] mprj_io_holdover[7]
+ mprj_io_ib_mode_sel[7] mprj_io_inp_dis[7] mprj_io_oeb[7] mprj_io_out[7] mprj_io_slow_sel[7]
+ mprj_io_vtrip_sel[7] mprj_io_in[7] mprj_analog_io[1] mprj_io[8] mprj_io_analog_en[8]
+ mprj_io_analog_pol[8] mprj_io_analog_sel[8] mprj_io_dm[24] mprj_io_dm[25] mprj_io_dm[26]
+ mprj_io_holdover[8] mprj_io_ib_mode_sel[8] mprj_io_inp_dis[8] mprj_io_oeb[8] mprj_io_out[8]
+ mprj_io_slow_sel[8] mprj_io_vtrip_sel[8] mprj_io_in[8] mprj_analog_io[2] mprj_io[9]
+ mprj_io_analog_en[9] mprj_io_analog_pol[9] mprj_io_analog_sel[9] mprj_io_dm[27]
+ mprj_io_dm[28] mprj_io_dm[29] mprj_io_holdover[9] mprj_io_ib_mode_sel[9] mprj_io_inp_dis[9]
+ mprj_io_oeb[9] mprj_io_out[9] mprj_io_slow_sel[9] mprj_io_vtrip_sel[9] mprj_io_in[9]
+ mprj_analog_io[12] mprj_io[19] mprj_io_analog_en[19] mprj_io_analog_pol[19] mprj_io_analog_sel[19]
+ mprj_io_dm[57] mprj_io_dm[58] mprj_io_dm[59] mprj_io_holdover[19] mprj_io_ib_mode_sel[19]
+ mprj_io_inp_dis[19] mprj_io_oeb[19] mprj_io_out[19] mprj_io_slow_sel[19] mprj_io_vtrip_sel[19]
+ mprj_io_in[19] mprj_analog_io[22] mprj_io[29] mprj_io_analog_en[29] mprj_io_analog_pol[29]
+ mprj_io_analog_sel[29] mprj_io_dm[87] mprj_io_dm[88] mprj_io_dm[89] mprj_io_holdover[29]
+ mprj_io_ib_mode_sel[29] mprj_io_inp_dis[29] mprj_io_oeb[29] mprj_io_out[29] mprj_io_slow_sel[29]
+ mprj_io_vtrip_sel[29] mprj_io_in[29] mprj_analog_io[23] mprj_io[30] mprj_io_analog_en[30]
+ mprj_io_analog_pol[30] mprj_io_analog_sel[30] mprj_io_dm[90] mprj_io_dm[91] mprj_io_dm[92]
+ mprj_io_holdover[30] mprj_io_ib_mode_sel[30] mprj_io_inp_dis[30] mprj_io_oeb[30]
+ mprj_io_out[30] mprj_io_slow_sel[30] mprj_io_vtrip_sel[30] mprj_io_in[30] mprj_analog_io[24]
+ mprj_io[31] mprj_io_analog_en[31] mprj_io_analog_pol[31] mprj_io_analog_sel[31]
+ mprj_io_dm[93] mprj_io_dm[94] mprj_io_dm[95] mprj_io_holdover[31] mprj_io_ib_mode_sel[31]
+ mprj_io_inp_dis[31] mprj_io_oeb[31] mprj_io_out[31] mprj_io_slow_sel[31] mprj_io_vtrip_sel[31]
+ mprj_io_in[31] mprj_analog_io[25] mprj_io[32] mprj_io_analog_en[32] mprj_io_analog_pol[32]
+ mprj_io_analog_sel[32] mprj_io_dm[96] mprj_io_dm[97] mprj_io_dm[98] mprj_io_holdover[32]
+ mprj_io_ib_mode_sel[32] mprj_io_inp_dis[32] mprj_io_oeb[32] mprj_io_out[32] mprj_io_slow_sel[32]
+ mprj_io_vtrip_sel[32] mprj_io_in[32] mprj_analog_io[26] mprj_io[33] mprj_io_analog_en[33]
+ mprj_io_analog_pol[33] mprj_io_analog_sel[33] mprj_io_dm[100] mprj_io_dm[101] mprj_io_dm[99]
+ mprj_io_holdover[33] mprj_io_ib_mode_sel[33] mprj_io_inp_dis[33] mprj_io_oeb[33]
+ mprj_io_out[33] mprj_io_slow_sel[33] mprj_io_vtrip_sel[33] mprj_io_in[33] mprj_analog_io[27]
+ mprj_io[34] mprj_io_analog_en[34] mprj_io_analog_pol[34] mprj_io_analog_sel[34]
+ mprj_io_dm[102] mprj_io_dm[103] mprj_io_dm[104] mprj_io_holdover[34] mprj_io_ib_mode_sel[34]
+ mprj_io_inp_dis[34] mprj_io_oeb[34] mprj_io_out[34] mprj_io_slow_sel[34] mprj_io_vtrip_sel[34]
+ mprj_io_in[34] mprj_analog_io[28] mprj_io[35] mprj_io_analog_en[35] mprj_io_analog_pol[35]
+ mprj_io_analog_sel[35] mprj_io_dm[105] mprj_io_dm[106] mprj_io_dm[107] mprj_io_holdover[35]
+ mprj_io_ib_mode_sel[35] mprj_io_inp_dis[35] mprj_io_oeb[35] mprj_io_out[35] mprj_io_slow_sel[35]
+ mprj_io_vtrip_sel[35] mprj_io_in[35] mprj_io[36] mprj_io_analog_en[36] mprj_io_analog_pol[36]
+ mprj_io_analog_sel[36] mprj_io_dm[108] mprj_io_dm[109] mprj_io_dm[110] mprj_io_holdover[36]
+ mprj_io_ib_mode_sel[36] mprj_io_inp_dis[36] mprj_io_oeb[36] mprj_io_out[36] mprj_io_slow_sel[36]
+ mprj_io_vtrip_sel[36] mprj_io_in[36] mprj_io[37] mprj_io_analog_en[37] mprj_io_analog_pol[37]
+ mprj_io_analog_sel[37] mprj_io_dm[111] mprj_io_dm[112] mprj_io_dm[113] mprj_io_holdover[37]
+ mprj_io_ib_mode_sel[37] mprj_io_inp_dis[37] mprj_io_oeb[37] mprj_io_out[37] mprj_io_slow_sel[37]
+ mprj_io_vtrip_sel[37] mprj_io_in[37] mprj_analog_io[13] mprj_io[20] mprj_io_analog_en[20]
+ mprj_io_analog_pol[20] mprj_io_analog_sel[20] mprj_io_dm[60] mprj_io_dm[61] mprj_io_dm[62]
+ mprj_io_holdover[20] mprj_io_ib_mode_sel[20] mprj_io_inp_dis[20] mprj_io_oeb[20]
+ mprj_io_out[20] mprj_io_slow_sel[20] mprj_io_vtrip_sel[20] mprj_io_in[20] mprj_analog_io[14]
+ mprj_io[21] mprj_io_analog_en[21] mprj_io_analog_pol[21] mprj_io_analog_sel[21]
+ mprj_io_dm[63] mprj_io_dm[64] mprj_io_dm[65] mprj_io_holdover[21] mprj_io_ib_mode_sel[21]
+ mprj_io_inp_dis[21] mprj_io_oeb[21] mprj_io_out[21] mprj_io_slow_sel[21] mprj_io_vtrip_sel[21]
+ mprj_io_in[21] mprj_analog_io[15] mprj_io[22] mprj_io_analog_en[22] mprj_io_analog_pol[22]
+ mprj_io_analog_sel[22] mprj_io_dm[66] mprj_io_dm[67] mprj_io_dm[68] mprj_io_holdover[22]
+ mprj_io_ib_mode_sel[22] mprj_io_inp_dis[22] mprj_io_oeb[22] mprj_io_out[22] mprj_io_slow_sel[22]
+ mprj_io_vtrip_sel[22] mprj_io_in[22] mprj_analog_io[16] mprj_io[23] mprj_io_analog_en[23]
+ mprj_io_analog_pol[23] mprj_io_analog_sel[23] mprj_io_dm[69] mprj_io_dm[70] mprj_io_dm[71]
+ mprj_io_holdover[23] mprj_io_ib_mode_sel[23] mprj_io_inp_dis[23] mprj_io_oeb[23]
+ mprj_io_out[23] mprj_io_slow_sel[23] mprj_io_vtrip_sel[23] mprj_io_in[23] mprj_analog_io[17]
+ mprj_io[24] mprj_io_analog_en[24] mprj_io_analog_pol[24] mprj_io_analog_sel[24]
+ mprj_io_dm[72] mprj_io_dm[73] mprj_io_dm[74] mprj_io_holdover[24] mprj_io_ib_mode_sel[24]
+ mprj_io_inp_dis[24] mprj_io_oeb[24] mprj_io_out[24] mprj_io_slow_sel[24] mprj_io_vtrip_sel[24]
+ mprj_io_in[24] mprj_analog_io[18] mprj_io[25] mprj_io_analog_en[25] mprj_io_analog_pol[25]
+ mprj_io_analog_sel[25] mprj_io_dm[75] mprj_io_dm[76] mprj_io_dm[77] mprj_io_holdover[25]
+ mprj_io_ib_mode_sel[25] mprj_io_inp_dis[25] mprj_io_oeb[25] mprj_io_out[25] mprj_io_slow_sel[25]
+ mprj_io_vtrip_sel[25] mprj_io_in[25] mprj_analog_io[19] mprj_io[26] mprj_io_analog_en[26]
+ mprj_io_analog_pol[26] mprj_io_analog_sel[26] mprj_io_dm[78] mprj_io_dm[79] mprj_io_dm[80]
+ mprj_io_holdover[26] mprj_io_ib_mode_sel[26] mprj_io_inp_dis[26] mprj_io_oeb[26]
+ mprj_io_out[26] mprj_io_slow_sel[26] mprj_io_vtrip_sel[26] mprj_io_in[26] mprj_analog_io[20]
+ mprj_io[27] mprj_io_analog_en[27] mprj_io_analog_pol[27] mprj_io_analog_sel[27]
+ mprj_io_dm[81] mprj_io_dm[82] mprj_io_dm[83] mprj_io_holdover[27] mprj_io_ib_mode_sel[27]
+ mprj_io_inp_dis[27] mprj_io_oeb[27] mprj_io_out[27] mprj_io_slow_sel[27] mprj_io_vtrip_sel[27]
+ mprj_io_in[27] mprj_analog_io[21] mprj_io[28] mprj_io_analog_en[28] mprj_io_analog_pol[28]
+ mprj_io_analog_sel[28] mprj_io_dm[84] mprj_io_dm[85] mprj_io_dm[86] mprj_io_holdover[28]
+ mprj_io_ib_mode_sel[28] mprj_io_inp_dis[28] mprj_io_oeb[28] mprj_io_out[28] mprj_io_slow_sel[28]
+ mprj_io_vtrip_sel[28] mprj_io_in[28] porb_h resetb resetb_core_h vdda vssa vccd1_pad
+ vdda1_pad vdda1_pad2 vssa1_pad vssa1_pad2 vccd1 vdda1 vssd1 vssd1_pad vccd2_pad
+ vdda2_pad vssa2_pad vccd2 vdda2 vddio vssd2 vssd2_pad vssa2 flash_io0_ieb_core vssio
+ vssa1 flash_io1_ieb_core vccd vssd
XFILLER_592 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_581 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_570 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xclock_pad clock_pad/IN_H clock_pad/PAD_A_NOESD_H clock_pad/PAD_A_ESD_0_H clock_pad/PAD_A_ESD_1_H
+ clock vssd vssd vccd vddio clock_core por vssd porb_h porb_h clock_pad/TIE_LO_ESD
+ vccd clock_pad/TIE_HI_ESD clock_pad/TIE_LO_ESD vssd vssd vssd vssd vssd vccd vssa
+ vssd vssd gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
Xmprj_pads.area2_io_pad\[17\] mprj_pads.area2_io_pad\[17\]/IN_H mprj_pads.area2_io_pad\[17\]/PAD_A_NOESD_H
+ mprj_pads.area2_io_pad\[17\]/PAD_A_ESD_0_H mprj_pads.area2_io_pad\[17\]/PAD_A_ESD_1_H
+ mprj_io[36] mprj_io_dm[110] mprj_io_dm[109] mprj_io_dm[108] vddio mprj_io_in[36]
+ mprj_io_inp_dis[36] mprj_io_ib_mode_sel[36] porb_h porb_h mprj_pads.area2_io_pad\[17\]/TIE_LO_ESD
+ mprj_io_oeb[36] mprj_pads.area2_io_pad\[17\]/TIE_HI_ESD mprj_pads.area2_io_pad\[17\]/TIE_LO_ESD
+ mprj_io_slow_sel[36] mprj_io_vtrip_sel[36] mprj_io_holdover[36] mprj_io_analog_en[36]
+ mprj_io_analog_sel[36] vccd vssio mprj_io_analog_pol[36] mprj_io_out[36] gpio_pad/AMUXBUS_A
+ gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd
+ gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_25 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_14 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_69 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_58 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_47 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_36 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xmgmt_vccd_lvclamp_pad gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vccd_pad vssa vdda vddio
+ gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__vccd_lvc_clamped_pad
Xmprj_pads.area2_io_pad\[7\] mprj_pads.area2_io_pad\[7\]/IN_H mprj_pads.area2_io_pad\[7\]/PAD_A_NOESD_H
+ mprj_analog_io[19] mprj_pads.area2_io_pad\[7\]/PAD_A_ESD_1_H mprj_io[26] mprj_io_dm[80]
+ mprj_io_dm[79] mprj_io_dm[78] vddio mprj_io_in[26] mprj_io_inp_dis[26] mprj_io_ib_mode_sel[26]
+ porb_h porb_h mprj_pads.area2_io_pad\[7\]/TIE_LO_ESD mprj_io_oeb[26] mprj_pads.area2_io_pad\[7\]/TIE_HI_ESD
+ mprj_pads.area2_io_pad\[7\]/TIE_LO_ESD mprj_io_slow_sel[26] mprj_io_vtrip_sel[26]
+ mprj_io_holdover[26] mprj_io_analog_en[26] mprj_io_analog_sel[26] vccd vssio mprj_io_analog_pol[26]
+ mprj_io_out[26] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_218 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_207 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_796 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_785 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_763 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_752 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_741 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_730 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_593 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_582 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_571 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_560 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_390 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
Xmprj_pads.area1_io_pad\[7\] mprj_pads.area1_io_pad\[7\]/IN_H mprj_pads.area1_io_pad\[7\]/PAD_A_NOESD_H
+ mprj_analog_io[0] mprj_pads.area1_io_pad\[7\]/PAD_A_ESD_1_H mprj_io[7] mprj_io_dm[23]
+ mprj_io_dm[22] mprj_io_dm[21] vddio mprj_io_in[7] mprj_io_inp_dis[7] mprj_io_ib_mode_sel[7]
+ porb_h porb_h mprj_pads.area1_io_pad\[7\]/TIE_LO_ESD mprj_io_oeb[7] mprj_pads.area1_io_pad\[7\]/TIE_HI_ESD
+ mprj_pads.area1_io_pad\[7\]/TIE_LO_ESD mprj_io_slow_sel[7] mprj_io_vtrip_sel[7]
+ mprj_io_holdover[7] mprj_io_analog_en[7] mprj_io_analog_sel[7] vccd vssio mprj_io_analog_pol[7]
+ mprj_io_out[7] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_59 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_48 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_37 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_26 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_15 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_219 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_208 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_797 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_786 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_775 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_753 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_742 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_731 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_720 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_583 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_572 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_561 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_550 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_380 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_391 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
Xmprj_pads.area1_io_pad\[11\] mprj_pads.area1_io_pad\[11\]/IN_H mprj_pads.area1_io_pad\[11\]/PAD_A_NOESD_H
+ mprj_analog_io[4] mprj_pads.area1_io_pad\[11\]/PAD_A_ESD_1_H mprj_io[11] mprj_io_dm[35]
+ mprj_io_dm[34] mprj_io_dm[33] vddio mprj_io_in[11] mprj_io_inp_dis[11] mprj_io_ib_mode_sel[11]
+ porb_h porb_h mprj_pads.area1_io_pad\[11\]/TIE_LO_ESD mprj_io_oeb[11] mprj_pads.area1_io_pad\[11\]/TIE_HI_ESD
+ mprj_pads.area1_io_pad\[11\]/TIE_LO_ESD mprj_io_slow_sel[11] mprj_io_vtrip_sel[11]
+ mprj_io_holdover[11] mprj_io_analog_en[11] mprj_io_analog_sel[11] vccd vssio mprj_io_analog_pol[11]
+ mprj_io_out[11] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_49 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_38 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_27 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_16 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_798 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_787 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_776 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_765 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_754 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_743 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_732 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_721 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_710 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_595 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_573 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_562 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_551 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_540 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_370 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_381 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_392 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
Xmprj_pads.area2_io_pad\[15\] mprj_pads.area2_io_pad\[15\]/IN_H mprj_pads.area2_io_pad\[15\]/PAD_A_NOESD_H
+ mprj_analog_io[27] mprj_pads.area2_io_pad\[15\]/PAD_A_ESD_1_H mprj_io[34] mprj_io_dm[104]
+ mprj_io_dm[103] mprj_io_dm[102] vddio mprj_io_in[34] mprj_io_inp_dis[34] mprj_io_ib_mode_sel[34]
+ porb_h porb_h mprj_pads.area2_io_pad\[15\]/TIE_LO_ESD mprj_io_oeb[34] mprj_pads.area2_io_pad\[15\]/TIE_HI_ESD
+ mprj_pads.area2_io_pad\[15\]/TIE_LO_ESD mprj_io_slow_sel[34] mprj_io_vtrip_sel[34]
+ mprj_io_holdover[34] mprj_io_analog_en[34] mprj_io_analog_sel[34] vccd vssio mprj_io_analog_pol[34]
+ mprj_io_out[34] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_39 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_28 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
Xmprj_pads.area2_io_pad\[5\] mprj_pads.area2_io_pad\[5\]/IN_H mprj_pads.area2_io_pad\[5\]/PAD_A_NOESD_H
+ mprj_analog_io[17] mprj_pads.area2_io_pad\[5\]/PAD_A_ESD_1_H mprj_io[24] mprj_io_dm[74]
+ mprj_io_dm[73] mprj_io_dm[72] vddio mprj_io_in[24] mprj_io_inp_dis[24] mprj_io_ib_mode_sel[24]
+ porb_h porb_h mprj_pads.area2_io_pad\[5\]/TIE_LO_ESD mprj_io_oeb[24] mprj_pads.area2_io_pad\[5\]/TIE_HI_ESD
+ mprj_pads.area2_io_pad\[5\]/TIE_LO_ESD mprj_io_slow_sel[24] mprj_io_vtrip_sel[24]
+ mprj_io_holdover[24] mprj_io_analog_en[24] mprj_io_analog_sel[24] vccd vssio mprj_io_analog_pol[24]
+ mprj_io_out[24] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_799 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_788 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_777 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_766 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_744 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_733 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_722 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_711 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_700 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_596 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_585 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_563 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_552 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_541 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_530 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_360 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_371 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_382 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_190 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_29 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_18 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xmprj_pads.area1_io_pad\[5\] mprj_pads.area1_io_pad\[5\]/IN_H mprj_pads.area1_io_pad\[5\]/PAD_A_NOESD_H
+ mprj_pads.area1_io_pad\[5\]/PAD_A_ESD_0_H mprj_pads.area1_io_pad\[5\]/PAD_A_ESD_1_H
+ mprj_io[5] mprj_io_dm[17] mprj_io_dm[16] mprj_io_dm[15] vddio mprj_io_in[5] mprj_io_inp_dis[5]
+ mprj_io_ib_mode_sel[5] porb_h porb_h mprj_pads.area1_io_pad\[5\]/TIE_LO_ESD mprj_io_oeb[5]
+ mprj_pads.area1_io_pad\[5\]/TIE_HI_ESD mprj_pads.area1_io_pad\[5\]/TIE_LO_ESD mprj_io_slow_sel[5]
+ mprj_io_vtrip_sel[5] mprj_io_holdover[5] mprj_io_analog_en[5] mprj_io_analog_sel[5]
+ vccd vssio mprj_io_analog_pol[5] mprj_io_out[5] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B
+ vssa1 vdda1 vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
Xdisconnect_vdda_0 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vddio gpio_pad/VDDIO_Q vccd
+ vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__disconnect_vdda_slice_5um
XFILLER_734 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_723 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_712 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_701 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_789 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_778 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_767 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_756 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_745 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_597 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_586 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_575 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_553 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_542 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_531 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_520 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_361 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_372 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_394 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_19 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_191 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
Xdisconnect_vdda_1 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vddio gpio_pad/VDDIO_Q vccd
+ vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__disconnect_vdda_slice_5um
XFILLER_779 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_768 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_757 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_735 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_724 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_713 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_702 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_598 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_587 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_576 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_565 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_543 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_532 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_521 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_510 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xuser2_corner gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__corner_pad
Xmgmt_vddio_hvclamp_pad\[0\] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vddio_pad vssa
+ vdda vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__vddio_hvc_clamped_pad
XFILLER_340 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_351 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_373 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_384 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_395 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_181 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_170 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xdisconnect_vdda_2 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vddio gpio_pad/VDDIO_Q vccd
+ vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__disconnect_vdda_slice_5um
Xmprj_pads.area2_io_pad\[13\] mprj_pads.area2_io_pad\[13\]/IN_H mprj_pads.area2_io_pad\[13\]/PAD_A_NOESD_H
+ mprj_analog_io[25] mprj_pads.area2_io_pad\[13\]/PAD_A_ESD_1_H mprj_io[32] mprj_io_dm[98]
+ mprj_io_dm[97] mprj_io_dm[96] vddio mprj_io_in[32] mprj_io_inp_dis[32] mprj_io_ib_mode_sel[32]
+ porb_h porb_h mprj_pads.area2_io_pad\[13\]/TIE_LO_ESD mprj_io_oeb[32] mprj_pads.area2_io_pad\[13\]/TIE_HI_ESD
+ mprj_pads.area2_io_pad\[13\]/TIE_LO_ESD mprj_io_slow_sel[32] mprj_io_vtrip_sel[32]
+ mprj_io_holdover[32] mprj_io_analog_en[32] mprj_io_analog_sel[32] vccd vssio mprj_io_analog_pol[32]
+ mprj_io_out[32] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
Xmgmt_vssio_hvclamp_pad\[1\] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssio_pad2 vssa2
+ vdda2 vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__vssio_hvc_clamped_pad
XFILLER_769 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_758 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_747 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_725 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_714 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_703 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xmprj_pads.area2_io_pad\[3\] mprj_pads.area2_io_pad\[3\]/IN_H mprj_pads.area2_io_pad\[3\]/PAD_A_NOESD_H
+ mprj_analog_io[15] mprj_pads.area2_io_pad\[3\]/PAD_A_ESD_1_H mprj_io[22] mprj_io_dm[68]
+ mprj_io_dm[67] mprj_io_dm[66] vddio mprj_io_in[22] mprj_io_inp_dis[22] mprj_io_ib_mode_sel[22]
+ porb_h porb_h mprj_pads.area2_io_pad\[3\]/TIE_LO_ESD mprj_io_oeb[22] mprj_pads.area2_io_pad\[3\]/TIE_HI_ESD
+ mprj_pads.area2_io_pad\[3\]/TIE_LO_ESD mprj_io_slow_sel[22] mprj_io_vtrip_sel[22]
+ mprj_io_holdover[22] mprj_io_analog_en[22] mprj_io_analog_sel[22] vccd vssio mprj_io_analog_pol[22]
+ mprj_io_out[22] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_500 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_599 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_588 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_577 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_566 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_555 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_533 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_522 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_511 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_374 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_341 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_352 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_385 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_396 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_160 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_182 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_171 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
Xbus_tie_1 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xmprj_pads.area1_io_pad\[3\] mprj_pads.area1_io_pad\[3\]/IN_H mprj_pads.area1_io_pad\[3\]/PAD_A_NOESD_H
+ mprj_pads.area1_io_pad\[3\]/PAD_A_ESD_0_H mprj_pads.area1_io_pad\[3\]/PAD_A_ESD_1_H
+ mprj_io[3] mprj_io_dm[11] mprj_io_dm[10] mprj_io_dm[9] vddio mprj_io_in[3] mprj_io_inp_dis[3]
+ mprj_io_ib_mode_sel[3] porb_h porb_h mprj_pads.area1_io_pad\[3\]/TIE_LO_ESD mprj_io_oeb[3]
+ mprj_pads.area1_io_pad\[3\]/TIE_HI_ESD mprj_pads.area1_io_pad\[3\]/TIE_LO_ESD mprj_io_slow_sel[3]
+ mprj_io_vtrip_sel[3] mprj_io_holdover[3] mprj_io_analog_en[3] mprj_io_analog_sel[3]
+ vccd vssio mprj_io_analog_pol[3] mprj_io_out[3] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B
+ vssa1 vdda1 vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_759 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_748 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_737 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_726 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_715 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_704 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_589 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_578 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_567 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_556 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_545 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_523 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_512 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_501 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_320 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_342 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_353 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_375 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_386 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_397 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_161 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_150 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_183 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_172 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
Xbus_tie_2 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
XFILLER_749 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_738 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_716 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_705 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xuser2_vdda_hvclamp_pad gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vdda2_pad vssa2 vdda2
+ vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__vdda_hvc_clamped_pad
XFILLER_579 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_568 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_557 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_546 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_535 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_513 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_502 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
Xmprj_pads.area1_io_pad\[18\] mprj_pads.area1_io_pad\[18\]/IN_H mprj_pads.area1_io_pad\[18\]/PAD_A_NOESD_H
+ mprj_analog_io[11] mprj_pads.area1_io_pad\[18\]/PAD_A_ESD_1_H mprj_io[18] mprj_io_dm[56]
+ mprj_io_dm[55] mprj_io_dm[54] vddio mprj_io_in[18] mprj_io_inp_dis[18] mprj_io_ib_mode_sel[18]
+ porb_h porb_h mprj_pads.area1_io_pad\[18\]/TIE_LO_ESD mprj_io_oeb[18] mprj_pads.area1_io_pad\[18\]/TIE_HI_ESD
+ mprj_pads.area1_io_pad\[18\]/TIE_LO_ESD mprj_io_slow_sel[18] mprj_io_vtrip_sel[18]
+ mprj_io_holdover[18] mprj_io_analog_en[18] mprj_io_analog_sel[18] vccd vssio mprj_io_analog_pol[18]
+ mprj_io_out[18] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_310 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_321 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_343 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_354 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_376 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_387 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_398 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_162 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_151 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_140 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_184 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_173 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
Xbus_tie_70 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xmprj_pads.area2_io_pad\[11\] mprj_pads.area2_io_pad\[11\]/IN_H mprj_pads.area2_io_pad\[11\]/PAD_A_NOESD_H
+ mprj_analog_io[23] mprj_pads.area2_io_pad\[11\]/PAD_A_ESD_1_H mprj_io[30] mprj_io_dm[92]
+ mprj_io_dm[91] mprj_io_dm[90] vddio mprj_io_in[30] mprj_io_inp_dis[30] mprj_io_ib_mode_sel[30]
+ porb_h porb_h mprj_pads.area2_io_pad\[11\]/TIE_LO_ESD mprj_io_oeb[30] mprj_pads.area2_io_pad\[11\]/TIE_HI_ESD
+ mprj_pads.area2_io_pad\[11\]/TIE_LO_ESD mprj_io_slow_sel[30] mprj_io_vtrip_sel[30]
+ mprj_io_holdover[30] mprj_io_analog_en[30] mprj_io_analog_sel[30] vccd vssio mprj_io_analog_pol[30]
+ mprj_io_out[30] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
Xbus_tie_3 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
XFILLER_739 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_728 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_706 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_569 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_558 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_547 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_536 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_525 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_503 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
Xmprj_pads.area2_io_pad\[1\] mprj_pads.area2_io_pad\[1\]/IN_H mprj_pads.area2_io_pad\[1\]/PAD_A_NOESD_H
+ mprj_analog_io[13] mprj_pads.area2_io_pad\[1\]/PAD_A_ESD_1_H mprj_io[20] mprj_io_dm[62]
+ mprj_io_dm[61] mprj_io_dm[60] vddio mprj_io_in[20] mprj_io_inp_dis[20] mprj_io_ib_mode_sel[20]
+ porb_h porb_h mprj_pads.area2_io_pad\[1\]/TIE_LO_ESD mprj_io_oeb[20] mprj_pads.area2_io_pad\[1\]/TIE_HI_ESD
+ mprj_pads.area2_io_pad\[1\]/TIE_LO_ESD mprj_io_slow_sel[20] mprj_io_vtrip_sel[20]
+ mprj_io_holdover[20] mprj_io_analog_en[20] mprj_io_analog_sel[20] vccd vssio mprj_io_analog_pol[20]
+ mprj_io_out[20] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_300 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_344 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_355 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_377 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_388 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_399 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_141 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_163 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_152 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_185 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_174 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
Xbus_tie_4 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_60 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_71 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
XFILLER_729 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_718 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_707 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
Xmprj_pads.area1_io_pad\[1\] mprj_pads.area1_io_pad\[1\]/IN_H mprj_pads.area1_io_pad\[1\]/PAD_A_NOESD_H
+ mprj_pads.area1_io_pad\[1\]/PAD_A_ESD_0_H mprj_pads.area1_io_pad\[1\]/PAD_A_ESD_1_H
+ mprj_io[1] mprj_io_dm[5] mprj_io_dm[4] mprj_io_dm[3] vddio mprj_io_in[1] mprj_io_inp_dis[1]
+ mprj_io_ib_mode_sel[1] porb_h porb_h mprj_pads.area1_io_pad\[1\]/TIE_LO_ESD mprj_io_oeb[1]
+ mprj_pads.area1_io_pad\[1\]/TIE_HI_ESD mprj_pads.area1_io_pad\[1\]/TIE_LO_ESD mprj_io_slow_sel[1]
+ mprj_io_vtrip_sel[1] mprj_io_holdover[1] mprj_io_analog_en[1] mprj_io_analog_sel[1]
+ vccd vssio mprj_io_analog_pol[1] mprj_io_out[1] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B
+ vssa1 vdda1 vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_559 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_548 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_537 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_526 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_515 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_301 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_323 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_334 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_378 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_389 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_164 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_153 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_142 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_131 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_120 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xuser1_vssd_lvclamp_pad gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssd1_pad vssa1 vdda1
+ vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q vccd1 vssd1 sky130_ef_io__vssd_lvc_clamped3_pad
Xgpio_pad gpio_pad/IN_H gpio_pad/PAD_A_NOESD_H gpio_pad/PAD_A_ESD_0_H gpio_pad/PAD_A_ESD_1_H
+ gpio gpio_mode1_core gpio_mode1_core gpio_mode0_core vddio gpio_in_core gpio_inenb_core
+ vssd porb_h porb_h gpio_pad/TIE_LO_ESD gpio_outenb_core gpio_pad/TIE_HI_ESD gpio_pad/TIE_LO_ESD
+ vssd vssd vssd vssd vssd vccd vssa vssd gpio_out_core gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B
+ vssa vdda vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
Xbus_tie_5 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_50 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_61 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_72 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
XFILLER_719 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_516 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_505 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_549 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_538 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_527 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_302 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_324 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_335 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_357 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_368 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_379 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_165 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_154 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_132 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xmprj_pads.area1_io_pad\[16\] mprj_pads.area1_io_pad\[16\]/IN_H mprj_pads.area1_io_pad\[16\]/PAD_A_NOESD_H
+ mprj_analog_io[9] mprj_pads.area1_io_pad\[16\]/PAD_A_ESD_1_H mprj_io[16] mprj_io_dm[50]
+ mprj_io_dm[49] mprj_io_dm[48] vddio mprj_io_in[16] mprj_io_inp_dis[16] mprj_io_ib_mode_sel[16]
+ porb_h porb_h mprj_pads.area1_io_pad\[16\]/TIE_LO_ESD mprj_io_oeb[16] mprj_pads.area1_io_pad\[16\]/TIE_HI_ESD
+ mprj_pads.area1_io_pad\[16\]/TIE_LO_ESD mprj_io_slow_sel[16] mprj_io_vtrip_sel[16]
+ mprj_io_holdover[16] mprj_io_analog_en[16] mprj_io_analog_sel[16] vccd vssio mprj_io_analog_pol[16]
+ mprj_io_out[16] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_121 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_110 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_198 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_187 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xuser1_vdda_hvclamp_pad\[0\] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vdda1_pad vssa1
+ vdda1 vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__vdda_hvc_clamped_pad
Xbus_tie_6 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_40 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_51 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_62 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
XFILLER_709 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xmgmt_vssd_lvclamp_pad gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssd_pad vssa vdda vddio
+ gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__vssd_lvc_clamped_pad
XFILLER_539 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_528 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_517 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_506 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_303 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_325 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_336 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_358 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_369 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_166 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_155 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_144 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_133 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_122 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_111 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_100 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_199 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_188 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
Xuser2_vccd_lvclamp_pad gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vccd2_pad vssa2 vdda2
+ vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q vccd2 vssd2 sky130_ef_io__vccd_lvc_clamped3_pad
Xbus_tie_30 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_41 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_52 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_63 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_7 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
XFILLER_529 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_518 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_507 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_304 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_326 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_337 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_359 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
Xmgmt_vssa_hvclamp_pad gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa_pad vssa vdda vddio
+ gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__vssa_hvc_clamped_pad
XFILLER_167 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_145 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_134 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_123 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_112 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_101 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_189 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_SB1 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_690 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xmgmt_corner\[1\] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__corner_pad
Xuser1_vssa_hvclamp_pad\[1\] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1_pad2 vssa1
+ vdda1 vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__vssa_hvc_clamped_pad
Xbus_tie_31 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_20 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_42 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_53 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_64 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_8 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
XFILLER_519 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_508 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_327 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_338 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_157 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_146 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_135 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_124 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_113 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_102 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_SB2 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_168 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_691 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xmprj_pads.area1_io_pad\[14\] mprj_pads.area1_io_pad\[14\]/IN_H mprj_pads.area1_io_pad\[14\]/PAD_A_NOESD_H
+ mprj_analog_io[7] mprj_pads.area1_io_pad\[14\]/PAD_A_ESD_1_H mprj_io[14] mprj_io_dm[44]
+ mprj_io_dm[43] mprj_io_dm[42] vddio mprj_io_in[14] mprj_io_inp_dis[14] mprj_io_ib_mode_sel[14]
+ porb_h porb_h mprj_pads.area1_io_pad\[14\]/TIE_LO_ESD mprj_io_oeb[14] mprj_pads.area1_io_pad\[14\]/TIE_HI_ESD
+ mprj_pads.area1_io_pad\[14\]/TIE_LO_ESD mprj_io_slow_sel[14] mprj_io_vtrip_sel[14]
+ mprj_io_holdover[14] mprj_io_analog_en[14] mprj_io_analog_sel[14] vccd vssio mprj_io_analog_pol[14]
+ mprj_io_out[14] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
Xbus_tie_32 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_21 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_10 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_9 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_43 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_54 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_65 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
XFILLER_509 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_306 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_317 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_SB3 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_169 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_158 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_147 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_136 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_125 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_114 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_103 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_692 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_681 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xmprj_pads.area2_io_pad\[18\] mprj_pads.area2_io_pad\[18\]/IN_H mprj_pads.area2_io_pad\[18\]/PAD_A_NOESD_H
+ mprj_pads.area2_io_pad\[18\]/PAD_A_ESD_0_H mprj_pads.area2_io_pad\[18\]/PAD_A_ESD_1_H
+ mprj_io[37] mprj_io_dm[113] mprj_io_dm[112] mprj_io_dm[111] vddio mprj_io_in[37]
+ mprj_io_inp_dis[37] mprj_io_ib_mode_sel[37] porb_h porb_h mprj_pads.area2_io_pad\[18\]/TIE_LO_ESD
+ mprj_io_oeb[37] mprj_pads.area2_io_pad\[18\]/TIE_HI_ESD mprj_pads.area2_io_pad\[18\]/TIE_LO_ESD
+ mprj_io_slow_sel[37] mprj_io_vtrip_sel[37] mprj_io_holdover[37] mprj_io_analog_en[37]
+ mprj_io_analog_sel[37] vccd vssio mprj_io_analog_pol[37] mprj_io_out[37] gpio_pad/AMUXBUS_A
+ gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd
+ gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
Xbus_tie_33 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_22 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_11 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_44 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_55 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_66 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xmprj_pads.area2_io_pad\[8\] mprj_pads.area2_io_pad\[8\]/IN_H mprj_pads.area2_io_pad\[8\]/PAD_A_NOESD_H
+ mprj_analog_io[20] mprj_pads.area2_io_pad\[8\]/PAD_A_ESD_1_H mprj_io[27] mprj_io_dm[83]
+ mprj_io_dm[82] mprj_io_dm[81] vddio mprj_io_in[27] mprj_io_inp_dis[27] mprj_io_ib_mode_sel[27]
+ porb_h porb_h mprj_pads.area2_io_pad\[8\]/TIE_LO_ESD mprj_io_oeb[27] mprj_pads.area2_io_pad\[8\]/TIE_HI_ESD
+ mprj_pads.area2_io_pad\[8\]/TIE_LO_ESD mprj_io_slow_sel[27] mprj_io_vtrip_sel[27]
+ mprj_io_holdover[27] mprj_io_analog_en[27] mprj_io_analog_sel[27] vccd vssio mprj_io_analog_pol[27]
+ mprj_io_out[27] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_307 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_318 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_159 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_148 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_137 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_126 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_115 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_104 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_693 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_660 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_671 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_682 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_490 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xbus_tie_34 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_23 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_12 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_45 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_56 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_67 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xmprj_pads.area1_io_pad\[8\] mprj_pads.area1_io_pad\[8\]/IN_H mprj_pads.area1_io_pad\[8\]/PAD_A_NOESD_H
+ mprj_analog_io[1] mprj_pads.area1_io_pad\[8\]/PAD_A_ESD_1_H mprj_io[8] mprj_io_dm[26]
+ mprj_io_dm[25] mprj_io_dm[24] vddio mprj_io_in[8] mprj_io_inp_dis[8] mprj_io_ib_mode_sel[8]
+ porb_h porb_h mprj_pads.area1_io_pad\[8\]/TIE_LO_ESD mprj_io_oeb[8] mprj_pads.area1_io_pad\[8\]/TIE_HI_ESD
+ mprj_pads.area1_io_pad\[8\]/TIE_LO_ESD mprj_io_slow_sel[8] mprj_io_vtrip_sel[8]
+ mprj_io_holdover[8] mprj_io_analog_en[8] mprj_io_analog_sel[8] vccd vssio mprj_io_analog_pol[8]
+ mprj_io_out[8] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
Xresetb_pad resetb_pad/PAD_A_ESD_H resetb_core_h vssio vccd resetb_pad/PAD_A_ESD_H
+ porb_h vssio vssio resetb_pad/TIE_LO_ESD resetb_pad/TIE_HI_ESD vssio vssio vssio
+ vssa vssd gpio_pad/AMUXBUS_B gpio_pad/AMUXBUS_A gpio_pad/VDDIO_Q vddio vddio vdda
+ vccd vccd gpio_pad/VSSIO_Q resetb sky130_fd_io__top_xres4v2
XFILLER_308 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_319 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_149 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_138 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_127 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_116 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_105 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_694 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_650 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_672 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_683 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_491 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_480 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xbus_tie_24 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_13 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_35 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_46 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_57 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_68 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xmprj_pads.area1_io_pad\[12\] mprj_pads.area1_io_pad\[12\]/IN_H mprj_pads.area1_io_pad\[12\]/PAD_A_NOESD_H
+ mprj_analog_io[5] mprj_pads.area1_io_pad\[12\]/PAD_A_ESD_1_H mprj_io[12] mprj_io_dm[38]
+ mprj_io_dm[37] mprj_io_dm[36] vddio mprj_io_in[12] mprj_io_inp_dis[12] mprj_io_ib_mode_sel[12]
+ porb_h porb_h mprj_pads.area1_io_pad\[12\]/TIE_LO_ESD mprj_io_oeb[12] mprj_pads.area1_io_pad\[12\]/TIE_HI_ESD
+ mprj_pads.area1_io_pad\[12\]/TIE_LO_ESD mprj_io_slow_sel[12] mprj_io_vtrip_sel[12]
+ mprj_io_holdover[12] mprj_io_analog_en[12] mprj_io_analog_sel[12] vccd vssio mprj_io_analog_pol[12]
+ mprj_io_out[12] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_810 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_309 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_139 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_128 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_106 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_695 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_640 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_651 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_662 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_673 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_684 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_492 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_481 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_470 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xbus_tie_25 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_14 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_36 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_47 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_58 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_69 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xmprj_pads.area2_io_pad\[16\] mprj_pads.area2_io_pad\[16\]/IN_H mprj_pads.area2_io_pad\[16\]/PAD_A_NOESD_H
+ mprj_analog_io[28] mprj_pads.area2_io_pad\[16\]/PAD_A_ESD_1_H mprj_io[35] mprj_io_dm[107]
+ mprj_io_dm[106] mprj_io_dm[105] vddio mprj_io_in[35] mprj_io_inp_dis[35] mprj_io_ib_mode_sel[35]
+ porb_h porb_h mprj_pads.area2_io_pad\[16\]/TIE_LO_ESD mprj_io_oeb[35] mprj_pads.area2_io_pad\[16\]/TIE_HI_ESD
+ mprj_pads.area2_io_pad\[16\]/TIE_LO_ESD mprj_io_slow_sel[35] mprj_io_vtrip_sel[35]
+ mprj_io_holdover[35] mprj_io_analog_en[35] mprj_io_analog_sel[35] vccd vssio mprj_io_analog_pol[35]
+ mprj_io_out[35] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
Xmprj_pads.area2_io_pad\[6\] mprj_pads.area2_io_pad\[6\]/IN_H mprj_pads.area2_io_pad\[6\]/PAD_A_NOESD_H
+ mprj_analog_io[18] mprj_pads.area2_io_pad\[6\]/PAD_A_ESD_1_H mprj_io[25] mprj_io_dm[77]
+ mprj_io_dm[76] mprj_io_dm[75] vddio mprj_io_in[25] mprj_io_inp_dis[25] mprj_io_ib_mode_sel[25]
+ porb_h porb_h mprj_pads.area2_io_pad\[6\]/TIE_LO_ESD mprj_io_oeb[25] mprj_pads.area2_io_pad\[6\]/TIE_HI_ESD
+ mprj_pads.area2_io_pad\[6\]/TIE_LO_ESD mprj_io_slow_sel[25] mprj_io_vtrip_sel[25]
+ mprj_io_holdover[25] mprj_io_analog_en[25] mprj_io_analog_sel[25] vccd vssio mprj_io_analog_pol[25]
+ mprj_io_out[25] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_811 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_800 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xflash_csb_pad flash_csb_pad/IN_H flash_csb_pad/PAD_A_NOESD_H flash_csb_pad/PAD_A_ESD_0_H
+ flash_csb_pad/PAD_A_ESD_1_H flash_csb vccd vccd vssd vddio flash_csb_pad/IN flash_csb_pad/INP_DIS
+ vssd porb_h porb_h flash_csb_pad/INP_DIS flash_csb_oeb_core flash_csb_pad/TIE_HI_ESD
+ flash_csb_pad/INP_DIS vssd vssd vssd vssd vssd vccd vssa vssd flash_csb_core gpio_pad/AMUXBUS_A
+ gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q
+ sky130_ef_io__gpiov2_pad_wrapped
XFILLER_129 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_118 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_107 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_696 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_630 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_641 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_663 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_674 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_685 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_493 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_482 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_471 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_460 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xbus_tie_26 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_15 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_37 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_48 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_59 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
XFILLER_290 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
Xmprj_pads.area1_io_pad\[6\] mprj_pads.area1_io_pad\[6\]/IN_H mprj_pads.area1_io_pad\[6\]/PAD_A_NOESD_H
+ mprj_pads.area1_io_pad\[6\]/PAD_A_ESD_0_H mprj_pads.area1_io_pad\[6\]/PAD_A_ESD_1_H
+ mprj_io[6] mprj_io_dm[20] mprj_io_dm[19] mprj_io_dm[18] vddio mprj_io_in[6] mprj_io_inp_dis[6]
+ mprj_io_ib_mode_sel[6] porb_h porb_h mprj_pads.area1_io_pad\[6\]/TIE_LO_ESD mprj_io_oeb[6]
+ mprj_pads.area1_io_pad\[6\]/TIE_HI_ESD mprj_pads.area1_io_pad\[6\]/TIE_LO_ESD mprj_io_slow_sel[6]
+ mprj_io_vtrip_sel[6] mprj_io_holdover[6] mprj_io_analog_en[6] mprj_io_analog_sel[6]
+ vccd vssio mprj_io_analog_pol[6] mprj_io_out[6] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B
+ vssa1 vdda1 vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_801 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_119 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_108 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_697 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_620 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_631 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_653 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_664 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_675 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_686 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_483 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_472 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_450 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_461 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
Xbus_tie_27 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_16 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_38 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_49 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
XFILLER_291 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
Xmprj_pads.area1_io_pad\[10\] mprj_pads.area1_io_pad\[10\]/IN_H mprj_pads.area1_io_pad\[10\]/PAD_A_NOESD_H
+ mprj_analog_io[3] mprj_pads.area1_io_pad\[10\]/PAD_A_ESD_1_H mprj_io[10] mprj_io_dm[32]
+ mprj_io_dm[31] mprj_io_dm[30] vddio mprj_io_in[10] mprj_io_inp_dis[10] mprj_io_ib_mode_sel[10]
+ porb_h porb_h mprj_pads.area1_io_pad\[10\]/TIE_LO_ESD mprj_io_oeb[10] mprj_pads.area1_io_pad\[10\]/TIE_HI_ESD
+ mprj_pads.area1_io_pad\[10\]/TIE_LO_ESD mprj_io_slow_sel[10] mprj_io_vtrip_sel[10]
+ mprj_io_holdover[10] mprj_io_analog_en[10] mprj_io_analog_sel[10] vccd vssio mprj_io_analog_pol[10]
+ mprj_io_out[10] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
Xflash_io1_pad flash_io1_pad/IN_H flash_io1_pad/PAD_A_NOESD_H flash_io1_pad/PAD_A_ESD_0_H
+ flash_io1_pad/PAD_A_ESD_1_H flash_io1 flash_io1_ieb_core flash_io1_ieb_core flash_io1_oeb_core
+ vddio flash_io1_di_core flash_io1_ieb_core vssd porb_h porb_h flash_io1_pad/TIE_LO_ESD
+ flash_io1_oeb_core flash_io1_pad/TIE_HI_ESD flash_io1_pad/TIE_LO_ESD vssd vssd vssd
+ vssd vssd vccd vssa vssd flash_io1_do_core gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B
+ vssa vdda vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_109 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_698 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_610 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_621 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_632 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_643 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_654 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_665 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_676 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_687 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xmgmt_vddio_hvclamp_pad\[1\] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vddio_pad2 vssa2
+ vdda2 vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__vddio_hvc_clamped_pad
XFILLER_495 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_473 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_440 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_451 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_462 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
Xbus_tie_28 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_17 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_39 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
XFILLER_270 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_292 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
Xmprj_pads.area2_io_pad\[14\] mprj_pads.area2_io_pad\[14\]/IN_H mprj_pads.area2_io_pad\[14\]/PAD_A_NOESD_H
+ mprj_analog_io[26] mprj_pads.area2_io_pad\[14\]/PAD_A_ESD_1_H mprj_io[33] mprj_io_dm[101]
+ mprj_io_dm[100] mprj_io_dm[99] vddio mprj_io_in[33] mprj_io_inp_dis[33] mprj_io_ib_mode_sel[33]
+ porb_h porb_h mprj_pads.area2_io_pad\[14\]/TIE_LO_ESD mprj_io_oeb[33] mprj_pads.area2_io_pad\[14\]/TIE_HI_ESD
+ mprj_pads.area2_io_pad\[14\]/TIE_LO_ESD mprj_io_slow_sel[33] mprj_io_vtrip_sel[33]
+ mprj_io_holdover[33] mprj_io_analog_en[33] mprj_io_analog_sel[33] vccd vssio mprj_io_analog_pol[33]
+ mprj_io_out[33] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_803 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xmprj_pads.area2_io_pad\[4\] mprj_pads.area2_io_pad\[4\]/IN_H mprj_pads.area2_io_pad\[4\]/PAD_A_NOESD_H
+ mprj_analog_io[16] mprj_pads.area2_io_pad\[4\]/PAD_A_ESD_1_H mprj_io[23] mprj_io_dm[71]
+ mprj_io_dm[70] mprj_io_dm[69] vddio mprj_io_in[23] mprj_io_inp_dis[23] mprj_io_ib_mode_sel[23]
+ porb_h porb_h mprj_pads.area2_io_pad\[4\]/TIE_LO_ESD mprj_io_oeb[23] mprj_pads.area2_io_pad\[4\]/TIE_HI_ESD
+ mprj_pads.area2_io_pad\[4\]/TIE_LO_ESD mprj_io_slow_sel[23] mprj_io_vtrip_sel[23]
+ mprj_io_holdover[23] mprj_io_analog_en[23] mprj_io_analog_sel[23] vccd vssio mprj_io_analog_pol[23]
+ mprj_io_out[23] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_600 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_611 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_622 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_644 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_655 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_666 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_677 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_688 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_496 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_485 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xbus_tie_29 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_18 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
XFILLER_430 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_441 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_452 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_463 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_293 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
Xmprj_pads.area1_io_pad\[4\] mprj_pads.area1_io_pad\[4\]/IN_H mprj_pads.area1_io_pad\[4\]/PAD_A_NOESD_H
+ mprj_pads.area1_io_pad\[4\]/PAD_A_ESD_0_H mprj_pads.area1_io_pad\[4\]/PAD_A_ESD_1_H
+ mprj_io[4] mprj_io_dm[14] mprj_io_dm[13] mprj_io_dm[12] vddio mprj_io_in[4] mprj_io_inp_dis[4]
+ mprj_io_ib_mode_sel[4] porb_h porb_h mprj_pads.area1_io_pad\[4\]/TIE_LO_ESD mprj_io_oeb[4]
+ mprj_pads.area1_io_pad\[4\]/TIE_HI_ESD mprj_pads.area1_io_pad\[4\]/TIE_LO_ESD mprj_io_slow_sel[4]
+ mprj_io_vtrip_sel[4] mprj_io_holdover[4] mprj_io_analog_en[4] mprj_io_analog_sel[4]
+ vccd vssio mprj_io_analog_pol[4] mprj_io_out[4] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B
+ vssa1 vdda1 vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_804 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_601 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_612 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_634 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_645 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_656 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_667 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_678 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_90 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_497 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_486 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_475 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xbus_tie_19 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
XFILLER_420 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_431 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_442 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_453 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_250 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_272 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_283 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_805 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_602 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_624 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_635 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_646 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_657 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_668 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_679 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_91 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_80 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_498 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_487 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_476 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_410 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_421 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_432 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_443 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_465 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_251 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_240 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_273 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_284 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
Xuser2_vssd_lvclamp_pad gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssd2_pad vssa2 vdda2
+ vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q vccd2 vssd2 sky130_ef_io__vssd_lvc_clamped3_pad
Xmprj_pads.area2_io_pad\[12\] mprj_pads.area2_io_pad\[12\]/IN_H mprj_pads.area2_io_pad\[12\]/PAD_A_NOESD_H
+ mprj_analog_io[24] mprj_pads.area2_io_pad\[12\]/PAD_A_ESD_1_H mprj_io[31] mprj_io_dm[95]
+ mprj_io_dm[94] mprj_io_dm[93] vddio mprj_io_in[31] mprj_io_inp_dis[31] mprj_io_ib_mode_sel[31]
+ porb_h porb_h mprj_pads.area2_io_pad\[12\]/TIE_LO_ESD mprj_io_oeb[31] mprj_pads.area2_io_pad\[12\]/TIE_HI_ESD
+ mprj_pads.area2_io_pad\[12\]/TIE_LO_ESD mprj_io_slow_sel[31] mprj_io_vtrip_sel[31]
+ mprj_io_holdover[31] mprj_io_analog_en[31] mprj_io_analog_sel[31] vccd vssio mprj_io_analog_pol[31]
+ mprj_io_out[31] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_806 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xmgmt_vssio_hvclamp_pad\[0\] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssio_pad vssa
+ vdda vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__vssio_hvc_clamped_pad
XFILLER_603 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_625 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_636 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_647 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_658 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_669 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_92 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_81 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
Xmprj_pads.area2_io_pad\[2\] mprj_pads.area2_io_pad\[2\]/IN_H mprj_pads.area2_io_pad\[2\]/PAD_A_NOESD_H
+ mprj_analog_io[14] mprj_pads.area2_io_pad\[2\]/PAD_A_ESD_1_H mprj_io[21] mprj_io_dm[65]
+ mprj_io_dm[64] mprj_io_dm[63] vddio mprj_io_in[21] mprj_io_inp_dis[21] mprj_io_ib_mode_sel[21]
+ porb_h porb_h mprj_pads.area2_io_pad\[2\]/TIE_LO_ESD mprj_io_oeb[21] mprj_pads.area2_io_pad\[2\]/TIE_HI_ESD
+ mprj_pads.area2_io_pad\[2\]/TIE_LO_ESD mprj_io_slow_sel[21] mprj_io_vtrip_sel[21]
+ mprj_io_holdover[21] mprj_io_analog_en[21] mprj_io_analog_sel[21] vccd vssio mprj_io_analog_pol[21]
+ mprj_io_out[21] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_499 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_488 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_477 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_400 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_411 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_422 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_433 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_455 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_466 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_252 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_241 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_274 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_285 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_807 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xuser2_vssa_hvclamp_pad gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2_pad vssa2 vdda2
+ vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__vssa_hvc_clamped_pad
Xmprj_pads.area1_io_pad\[2\] mprj_pads.area1_io_pad\[2\]/IN_H mprj_pads.area1_io_pad\[2\]/PAD_A_NOESD_H
+ mprj_pads.area1_io_pad\[2\]/PAD_A_ESD_0_H mprj_pads.area1_io_pad\[2\]/PAD_A_ESD_1_H
+ mprj_io[2] mprj_io_dm[8] mprj_io_dm[7] mprj_io_dm[6] vddio mprj_io_in[2] mprj_io_inp_dis[2]
+ mprj_io_ib_mode_sel[2] porb_h porb_h mprj_pads.area1_io_pad\[2\]/TIE_LO_ESD mprj_io_oeb[2]
+ mprj_pads.area1_io_pad\[2\]/TIE_HI_ESD mprj_pads.area1_io_pad\[2\]/TIE_LO_ESD mprj_io_slow_sel[2]
+ mprj_io_vtrip_sel[2] mprj_io_holdover[2] mprj_io_analog_en[2] mprj_io_analog_sel[2]
+ vccd vssio mprj_io_analog_pol[2] mprj_io_out[2] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B
+ vssa1 vdda1 vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_5 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_604 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_615 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_626 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_637 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_648 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_659 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_93 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_82 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_71 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_60 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_489 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_478 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_401 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_412 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_423 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_445 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_456 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_467 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_253 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_242 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_275 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_286 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_808 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_6 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_605 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_616 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_627 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_638 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_649 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_94 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_72 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_61 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_50 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_479 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_468 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_402 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_413 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_435 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_446 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_457 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_232 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_221 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_276 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_287 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
Xmprj_pads.area1_io_pad\[17\] mprj_pads.area1_io_pad\[17\]/IN_H mprj_pads.area1_io_pad\[17\]/PAD_A_NOESD_H
+ mprj_analog_io[10] mprj_pads.area1_io_pad\[17\]/PAD_A_ESD_1_H mprj_io[17] mprj_io_dm[53]
+ mprj_io_dm[52] mprj_io_dm[51] vddio mprj_io_in[17] mprj_io_inp_dis[17] mprj_io_ib_mode_sel[17]
+ porb_h porb_h mprj_pads.area1_io_pad\[17\]/TIE_LO_ESD mprj_io_oeb[17] mprj_pads.area1_io_pad\[17\]/TIE_HI_ESD
+ mprj_pads.area1_io_pad\[17\]/TIE_LO_ESD mprj_io_slow_sel[17] mprj_io_vtrip_sel[17]
+ mprj_io_holdover[17] mprj_io_analog_en[17] mprj_io_analog_sel[17] vccd vssio mprj_io_analog_pol[17]
+ mprj_io_out[17] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
Xuser1_vdda_hvclamp_pad\[1\] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vdda1_pad2 vssa1
+ vdda1 vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__vdda_hvc_clamped_pad
XFILLER_809 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xmprj_pads.area2_io_pad\[10\] mprj_pads.area2_io_pad\[10\]/IN_H mprj_pads.area2_io_pad\[10\]/PAD_A_NOESD_H
+ mprj_analog_io[22] mprj_pads.area2_io_pad\[10\]/PAD_A_ESD_1_H mprj_io[29] mprj_io_dm[89]
+ mprj_io_dm[88] mprj_io_dm[87] vddio mprj_io_in[29] mprj_io_inp_dis[29] mprj_io_ib_mode_sel[29]
+ porb_h porb_h mprj_pads.area2_io_pad\[10\]/TIE_LO_ESD mprj_io_oeb[29] mprj_pads.area2_io_pad\[10\]/TIE_HI_ESD
+ mprj_pads.area2_io_pad\[10\]/TIE_LO_ESD mprj_io_slow_sel[29] mprj_io_vtrip_sel[29]
+ mprj_io_holdover[29] mprj_io_analog_en[29] mprj_io_analog_sel[29] vccd vssio mprj_io_analog_pol[29]
+ mprj_io_out[29] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_7 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_606 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_617 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_628 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_639 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_95 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_73 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_62 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_51 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_40 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_469 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_425 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_436 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_447 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_458 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xmprj_pads.area2_io_pad\[0\] mprj_pads.area2_io_pad\[0\]/IN_H mprj_pads.area2_io_pad\[0\]/PAD_A_NOESD_H
+ mprj_analog_io[12] mprj_pads.area2_io_pad\[0\]/PAD_A_ESD_1_H mprj_io[19] mprj_io_dm[59]
+ mprj_io_dm[58] mprj_io_dm[57] vddio mprj_io_in[19] mprj_io_inp_dis[19] mprj_io_ib_mode_sel[19]
+ porb_h porb_h mprj_pads.area2_io_pad\[0\]/TIE_LO_ESD mprj_io_oeb[19] mprj_pads.area2_io_pad\[0\]/TIE_HI_ESD
+ mprj_pads.area2_io_pad\[0\]/TIE_LO_ESD mprj_io_slow_sel[19] mprj_io_vtrip_sel[19]
+ mprj_io_holdover[19] mprj_io_analog_en[19] mprj_io_analog_sel[19] vccd vssio mprj_io_analog_pol[19]
+ mprj_io_out[19] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_255 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_233 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_222 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_200 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_266 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_8 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_607 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_618 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_629 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_96 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_74 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_63 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_52 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_41 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
Xmprj_pads.area1_io_pad\[0\] mprj_pads.area1_io_pad\[0\]/IN_H mprj_pads.area1_io_pad\[0\]/PAD_A_NOESD_H
+ mprj_pads.area1_io_pad\[0\]/PAD_A_ESD_0_H mprj_pads.area1_io_pad\[0\]/PAD_A_ESD_1_H
+ mprj_io[0] mprj_io_dm[2] mprj_io_dm[1] mprj_io_dm[0] vddio mprj_io_in[0] mprj_io_inp_dis[0]
+ mprj_io_ib_mode_sel[0] porb_h porb_h mprj_pads.area1_io_pad\[0\]/TIE_LO_ESD mprj_io_oeb[0]
+ mprj_pads.area1_io_pad\[0\]/TIE_HI_ESD mprj_pads.area1_io_pad\[0\]/TIE_LO_ESD mprj_io_slow_sel[0]
+ mprj_io_vtrip_sel[0] mprj_io_holdover[0] mprj_io_analog_en[0] mprj_io_analog_sel[0]
+ vccd vssio mprj_io_analog_pol[0] mprj_io_out[0] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B
+ vssa1 vdda1 vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_415 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_426 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_437 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_448 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_459 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_256 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_234 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_223 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_201 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_267 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_289 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_790 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_9 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_608 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_619 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_86 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_75 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_64 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_53 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_42 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_31 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_20 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_405 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_416 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_427 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_438 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_449 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_257 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_235 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_224 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_202 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_268 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_791 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_780 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xmgmt_vdda_hvclamp_pad gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vdda_pad vssa vdda vddio
+ gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__vdda_hvc_clamped_pad
Xmprj_pads.area1_io_pad\[15\] mprj_pads.area1_io_pad\[15\]/IN_H mprj_pads.area1_io_pad\[15\]/PAD_A_NOESD_H
+ mprj_analog_io[8] mprj_pads.area1_io_pad\[15\]/PAD_A_ESD_1_H mprj_io[15] mprj_io_dm[47]
+ mprj_io_dm[46] mprj_io_dm[45] vddio mprj_io_in[15] mprj_io_inp_dis[15] mprj_io_ib_mode_sel[15]
+ porb_h porb_h mprj_pads.area1_io_pad\[15\]/TIE_LO_ESD mprj_io_oeb[15] mprj_pads.area1_io_pad\[15\]/TIE_HI_ESD
+ mprj_pads.area1_io_pad\[15\]/TIE_LO_ESD mprj_io_slow_sel[15] mprj_io_vtrip_sel[15]
+ mprj_io_holdover[15] mprj_io_analog_en[15] mprj_io_analog_sel[15] vccd vssio mprj_io_analog_pol[15]
+ mprj_io_out[15] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_609 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_98 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_87 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_76 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_65 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_54 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_32 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_21 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_10 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_406 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_417 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_428 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_439 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_258 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_236 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_225 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_269 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_792 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_781 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_770 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xmprj_pads.area2_io_pad\[9\] mprj_pads.area2_io_pad\[9\]/IN_H mprj_pads.area2_io_pad\[9\]/PAD_A_NOESD_H
+ mprj_analog_io[21] mprj_pads.area2_io_pad\[9\]/PAD_A_ESD_1_H mprj_io[28] mprj_io_dm[86]
+ mprj_io_dm[85] mprj_io_dm[84] vddio mprj_io_in[28] mprj_io_inp_dis[28] mprj_io_ib_mode_sel[28]
+ porb_h porb_h mprj_pads.area2_io_pad\[9\]/TIE_LO_ESD mprj_io_oeb[28] mprj_pads.area2_io_pad\[9\]/TIE_HI_ESD
+ mprj_pads.area2_io_pad\[9\]/TIE_LO_ESD mprj_io_slow_sel[28] mprj_io_vtrip_sel[28]
+ mprj_io_holdover[28] mprj_io_analog_en[28] mprj_io_analog_sel[28] vccd vssio mprj_io_analog_pol[28]
+ mprj_io_out[28] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
Xflash_io0_pad flash_io0_pad/IN_H flash_io0_pad/PAD_A_NOESD_H flash_io0_pad/PAD_A_ESD_0_H
+ flash_io0_pad/PAD_A_ESD_1_H flash_io0 flash_io0_ieb_core flash_io0_ieb_core flash_io0_oeb_core
+ vddio flash_io0_di_core flash_io0_ieb_core vssd porb_h porb_h flash_io0_pad/TIE_LO_ESD
+ flash_io0_oeb_core flash_io0_pad/TIE_HI_ESD flash_io0_pad/TIE_LO_ESD vssd vssd vssd
+ vssd vssd vccd vssa vssd flash_io0_do_core gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B
+ vssa vdda vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_99 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_88 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_77 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_66 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_55 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_44 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_33 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_22 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_11 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_407 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_418 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_429 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_259 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_215 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_204 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_782 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_771 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_760 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_590 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xmgmt_corner\[0\] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__corner_pad
Xuser1_vssa_hvclamp_pad\[0\] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1_pad vssa1
+ vdda1 vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__vssa_hvc_clamped_pad
Xmprj_pads.area1_io_pad\[9\] mprj_pads.area1_io_pad\[9\]/IN_H mprj_pads.area1_io_pad\[9\]/PAD_A_NOESD_H
+ mprj_analog_io[2] mprj_pads.area1_io_pad\[9\]/PAD_A_ESD_1_H mprj_io[9] mprj_io_dm[29]
+ mprj_io_dm[28] mprj_io_dm[27] vddio mprj_io_in[9] mprj_io_inp_dis[9] mprj_io_ib_mode_sel[9]
+ porb_h porb_h mprj_pads.area1_io_pad\[9\]/TIE_LO_ESD mprj_io_oeb[9] mprj_pads.area1_io_pad\[9\]/TIE_HI_ESD
+ mprj_pads.area1_io_pad\[9\]/TIE_LO_ESD mprj_io_slow_sel[9] mprj_io_vtrip_sel[9]
+ mprj_io_holdover[9] mprj_io_analog_en[9] mprj_io_analog_sel[9] vccd vssio mprj_io_analog_pol[9]
+ mprj_io_out[9] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_89 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_78 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_67 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_45 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_34 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_23 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_12 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xflash_clk_pad flash_clk_pad/IN_H flash_clk_pad/PAD_A_NOESD_H flash_clk_pad/PAD_A_ESD_0_H
+ flash_clk_pad/PAD_A_ESD_1_H flash_clk vccd vccd vssd vddio flash_clk_pad/IN flash_clk_pad/INP_DIS
+ vssd porb_h porb_h flash_clk_pad/INP_DIS flash_clk_oeb_core flash_clk_pad/TIE_HI_ESD
+ flash_clk_pad/INP_DIS vssd vssd vssd vssd vssd vccd vssa vssd flash_clk_core gpio_pad/AMUXBUS_A
+ gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q
+ sky130_ef_io__gpiov2_pad_wrapped
XFILLER_408 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_419 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_249 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_238 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_216 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_205 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_794 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_772 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_761 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_750 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_591 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
Xuser1_vccd_lvclamp_pad gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vccd1_pad vssa1 vdda1
+ vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q vccd1 vssd1 sky130_ef_io__vccd_lvc_clamped3_pad
XFILLER_580 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xmprj_pads.area1_io_pad\[13\] mprj_pads.area1_io_pad\[13\]/IN_H mprj_pads.area1_io_pad\[13\]/PAD_A_NOESD_H
+ mprj_analog_io[6] mprj_pads.area1_io_pad\[13\]/PAD_A_ESD_1_H mprj_io[13] mprj_io_dm[41]
+ mprj_io_dm[40] mprj_io_dm[39] vddio mprj_io_in[13] mprj_io_inp_dis[13] mprj_io_ib_mode_sel[13]
+ porb_h porb_h mprj_pads.area1_io_pad\[13\]/TIE_LO_ESD mprj_io_oeb[13] mprj_pads.area1_io_pad\[13\]/TIE_HI_ESD
+ mprj_pads.area1_io_pad\[13\]/TIE_LO_ESD mprj_io_slow_sel[13] mprj_io_vtrip_sel[13]
+ mprj_io_holdover[13] mprj_io_analog_en[13] mprj_io_analog_sel[13] vccd vssio mprj_io_analog_pol[13]
+ mprj_io_out[13] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_79 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_68 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_57 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_46 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_35 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_24 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_13 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
Xuser1_corner gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__corner_pad
XFILLER_409 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_239 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_217 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_206 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_795 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_784 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_773 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_762 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_751 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_740 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
.ends

.subckt sky130_fd_sc_hd__dfbbp_1 CLK D RESET_B SET_B VGND VPWR Q Q_N VNB VPB
X0 a_788_47# a_942_21# a_648_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 VPWR RESET_B a_942_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 VGND a_1429_21# a_1364_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR a_942_21# a_1663_329# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X4 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR a_1429_21# a_1341_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_474_413# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X8 a_1545_47# a_942_21# a_1429_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X9 VPWR a_1429_21# a_2136_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X10 a_582_47# a_193_47# a_474_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X11 a_1429_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_648_21# a_474_413# a_788_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X13 a_1341_413# a_193_47# a_1255_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_1663_329# a_1255_47# a_1429_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X15 a_1160_47# a_648_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X16 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_1255_47# a_27_47# a_1113_329# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 Q a_2136_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_648_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 a_788_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 Q_N a_1429_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 VGND RESET_B a_942_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 Q a_2136_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 VPWR a_942_21# a_892_329# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X25 a_558_413# a_27_47# a_474_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 VGND a_648_21# a_582_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 a_892_329# a_474_413# a_648_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X28 VGND a_1429_21# a_2136_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X30 a_474_413# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X31 a_1364_47# a_27_47# a_1255_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X32 a_1255_47# a_193_47# a_1160_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X33 Q_N a_1429_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X34 a_1545_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X35 VPWR a_648_21# a_558_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X36 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X37 a_1113_329# a_648_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X38 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X39 a_1429_21# a_1255_47# a_1545_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
.ends

.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VPWR X VNB VPB
X0 VPWR S a_591_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 a_591_369# A0 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_79_21# A1 a_306_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND S a_578_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_306_369# a_257_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X7 a_79_21# A0 a_288_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_288_47# a_257_199# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_257_199# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_578_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_257_199# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X13 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__inv_8 A VGND VPWR Y VNB VPB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt spare_logic_block spare_xfq[0] spare_xfq[1] spare_xfqn[0] spare_xfqn[1] spare_xi[0]
+ spare_xi[1] spare_xi[2] spare_xi[3] spare_xib spare_xmx[0] spare_xmx[1] spare_xna[0]
+ spare_xna[1] spare_xno[0] spare_xno[1] spare_xz[0] spare_xz[10] spare_xz[11] spare_xz[12]
+ spare_xz[13] spare_xz[14] spare_xz[15] spare_xz[16] spare_xz[17] spare_xz[18] spare_xz[19]
+ spare_xz[1] spare_xz[20] spare_xz[21] spare_xz[22] spare_xz[23] spare_xz[24] spare_xz[25]
+ spare_xz[26] spare_xz[2] spare_xz[3] spare_xz[4] spare_xz[5] spare_xz[6] spare_xz[7]
+ spare_xz[8] spare_xz[9] vssd vccd
XFILLER_0_24 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_57 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_57 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xspare_logic_const\[8\] vssd vssd vccd vccd spare_logic_const\[8\]/HI spare_xz[8]
+ sky130_fd_sc_hd__conb_1
XFILLER_3_35 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xspare_logic_nor\[0\] spare_xz[9] spare_xz[11] vssd vccd spare_xno[0] vssd vccd sky130_fd_sc_hd__nor2_2
XFILLER_0_47 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_47 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xspare_logic_const\[22\] vssd vssd vccd vccd spare_logic_const\[22\]/HI spare_xz[22]
+ sky130_fd_sc_hd__conb_1
XFILLER_9_57 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_24 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_25 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xspare_logic_const\[15\] vssd vssd vccd vccd spare_logic_const\[15\]/HI spare_xz[15]
+ sky130_fd_sc_hd__conb_1
XFILLER_9_36 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_59 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xspare_logic_const\[6\] vssd vssd vccd vccd spare_logic_const\[6\]/HI spare_xz[6]
+ sky130_fd_sc_hd__conb_1
XFILLER_11_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_48 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xspare_logic_const\[20\] vssd vssd vccd vccd spare_logic_const\[20\]/HI spare_xz[20]
+ sky130_fd_sc_hd__conb_1
XFILLER_9_16 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_17 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XPHY_0 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_61 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xspare_logic_const\[13\] vssd vssd vccd vccd spare_logic_const\[13\]/HI spare_xz[13]
+ sky130_fd_sc_hd__conb_1
XFILLER_1_62 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XPHY_1 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_61 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_29 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xspare_logic_const\[4\] vssd vssd vccd vccd spare_logic_const\[4\]/HI spare_xz[4]
+ sky130_fd_sc_hd__conb_1
XFILLER_7_51 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XPHY_2 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_41 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xspare_logic_flop\[0\] spare_xz[21] spare_xz[19] spare_xz[25] spare_xz[23] vssd vccd
+ spare_xfq[0] spare_xfqn[0] vssd vccd sky130_fd_sc_hd__dfbbp_1
XPHY_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xspare_logic_mux\[1\] spare_xz[14] spare_xz[16] spare_xz[18] vssd vccd spare_xmx[1]
+ vssd vccd sky130_fd_sc_hd__mux2_2
XFILLER_4_53 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_20 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xspare_logic_const\[11\] vssd vssd vccd vccd spare_logic_const\[11\]/HI spare_xz[11]
+ sky130_fd_sc_hd__conb_1
XFILLER_10_52 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XPHY_4 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_8 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xspare_logic_const\[2\] vssd vssd vccd vccd spare_logic_const\[2\]/HI spare_xz[2]
+ sky130_fd_sc_hd__conb_1
XPHY_5 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xspare_logic_inv\[3\] spare_xz[3] vssd vccd spare_xi[3] vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_10_21 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XPHY_6 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_66 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XPHY_7 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xspare_logic_const\[0\] vssd vssd vccd vccd spare_logic_const\[0\]/HI spare_xz[0]
+ sky130_fd_sc_hd__conb_1
XFILLER_10_34 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_8 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xspare_logic_inv\[1\] spare_xz[1] vssd vccd spare_xi[1] vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_10_46 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_48 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XPHY_9 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xspare_logic_const\[25\] vssd vssd vccd vccd spare_logic_const\[25\]/HI spare_xz[25]
+ sky130_fd_sc_hd__conb_1
XFILLER_6_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xspare_logic_nand\[1\] spare_xz[6] spare_xz[8] vssd vccd spare_xna[1] vssd vccd sky130_fd_sc_hd__nand2_2
XFILLER_1_38 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_14 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xspare_logic_const\[18\] vssd vssd vccd vccd spare_logic_const\[18\]/HI spare_xz[18]
+ sky130_fd_sc_hd__conb_1
XFILLER_10_59 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_27 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xspare_logic_const\[9\] vssd vssd vccd vccd spare_logic_const\[9\]/HI spare_xz[9]
+ sky130_fd_sc_hd__conb_1
XFILLER_8_8 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xspare_logic_nor\[1\] spare_xz[10] spare_xz[12] vssd vccd spare_xno[1] vssd vccd sky130_fd_sc_hd__nor2_2
XFILLER_7_39 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xspare_logic_const\[23\] vssd vssd vccd vccd spare_logic_const\[23\]/HI spare_xz[23]
+ sky130_fd_sc_hd__conb_1
XFILLER_4_29 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xspare_logic_const\[16\] vssd vssd vccd vccd spare_logic_const\[16\]/HI spare_xz[16]
+ sky130_fd_sc_hd__conb_1
XFILLER_2_41 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_52 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xspare_logic_const\[7\] vssd vssd vccd vccd spare_logic_const\[7\]/HI spare_xz[7]
+ sky130_fd_sc_hd__conb_1
Xspare_logic_biginv spare_xz[4] vssd vccd spare_xib vssd vccd sky130_fd_sc_hd__inv_8
XFILLER_8_41 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xspare_logic_const\[21\] vssd vssd vccd vccd spare_logic_const\[21\]/HI spare_xz[21]
+ sky130_fd_sc_hd__conb_1
XFILLER_5_31 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_54 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_41 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_53 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_20 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_43 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xspare_logic_const\[14\] vssd vssd vccd vccd spare_logic_const\[14\]/HI spare_xz[14]
+ sky130_fd_sc_hd__conb_1
XFILLER_2_66 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_53 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_22 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_66 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xspare_logic_const\[5\] vssd vssd vccd vccd spare_logic_const\[5\]/HI spare_xz[5]
+ sky130_fd_sc_hd__conb_1
XFILLER_4_8 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_66 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_12 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_66 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XPHY_20 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xspare_logic_flop\[1\] spare_xz[22] spare_xz[20] spare_xz[26] spare_xz[24] vssd vccd
+ spare_xfq[1] spare_xfqn[1] vssd vccd sky130_fd_sc_hd__dfbbp_1
XFILLER_0_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_57 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XPHY_21 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_10 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xspare_logic_const\[12\] vssd vssd vccd vccd spare_logic_const\[12\]/HI spare_xz[12]
+ sky130_fd_sc_hd__conb_1
XFILLER_2_47 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XPHY_22 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_11 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_57 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xspare_logic_const\[3\] vssd vssd vccd vccd spare_logic_const\[3\]/HI spare_xz[3]
+ sky130_fd_sc_hd__conb_1
XFILLER_2_8 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XPHY_12 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_23 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_13 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xspare_logic_mux\[0\] spare_xz[13] spare_xz[15] spare_xz[17] vssd vccd spare_xmx[0]
+ vssd vccd sky130_fd_sc_hd__mux2_2
Xspare_logic_const\[10\] vssd vssd vccd vccd spare_logic_const\[10\]/HI spare_xz[10]
+ sky130_fd_sc_hd__conb_1
XFILLER_11_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_14 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_29 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xspare_logic_const\[1\] vssd vssd vccd vccd spare_logic_const\[1\]/HI spare_xz[1]
+ sky130_fd_sc_hd__conb_1
XPHY_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xspare_logic_inv\[2\] spare_xz[2] vssd vccd spare_xi[2] vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_8_29 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xspare_logic_const\[26\] vssd vssd vccd vccd spare_logic_const\[26\]/HI spare_xz[26]
+ sky130_fd_sc_hd__conb_1
XFILLER_5_19 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_16 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_29 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_17 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xspare_logic_const\[19\] vssd vssd vccd vccd spare_logic_const\[19\]/HI spare_xz[19]
+ sky130_fd_sc_hd__conb_1
XFILLER_6_41 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_63 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XPHY_18 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_53 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xspare_logic_inv\[0\] spare_xz[0] vssd vccd spare_xi[0] vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_0_66 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_9 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_10 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XPHY_19 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xspare_logic_const\[24\] vssd vssd vccd vccd spare_logic_const\[24\]/HI spare_xz[24]
+ sky130_fd_sc_hd__conb_1
XFILLER_3_66 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xspare_logic_nand\[0\] spare_xz[5] spare_xz[7] vssd vccd spare_xna[0] vssd vccd sky130_fd_sc_hd__nand2_2
XFILLER_0_34 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_66 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xspare_logic_const\[17\] vssd vssd vccd vccd spare_logic_const\[17\]/HI spare_xz[17]
+ sky130_fd_sc_hd__conb_1
.ends

* Black-box entry subcircuit for mgmt_core_wrapper abstract view
.subckt mgmt_core_wrapper VGND VPWR core_clk core_rstn debug_in debug_mode debug_oeb
+ debug_out flash_clk flash_csb flash_io0_di flash_io0_do flash_io0_oeb flash_io1_di
+ flash_io1_do flash_io1_oeb flash_io2_di flash_io2_do flash_io2_oeb flash_io3_di
+ flash_io3_do flash_io3_oeb gpio_in_pad gpio_inenb_pad gpio_mode0_pad gpio_mode1_pad
+ gpio_out_pad gpio_outenb_pad hk_ack_i hk_cyc_o hk_dat_i[0] hk_dat_i[10] hk_dat_i[11]
+ hk_dat_i[12] hk_dat_i[13] hk_dat_i[14] hk_dat_i[15] hk_dat_i[16] hk_dat_i[17] hk_dat_i[18]
+ hk_dat_i[19] hk_dat_i[1] hk_dat_i[20] hk_dat_i[21] hk_dat_i[22] hk_dat_i[23] hk_dat_i[24]
+ hk_dat_i[25] hk_dat_i[26] hk_dat_i[27] hk_dat_i[28] hk_dat_i[29] hk_dat_i[2] hk_dat_i[30]
+ hk_dat_i[31] hk_dat_i[3] hk_dat_i[4] hk_dat_i[5] hk_dat_i[6] hk_dat_i[7] hk_dat_i[8]
+ hk_dat_i[9] hk_stb_o irq[0] irq[1] irq[2] irq[3] irq[4] irq[5] la_iena[0] la_iena[100]
+ la_iena[101] la_iena[102] la_iena[103] la_iena[104] la_iena[105] la_iena[106] la_iena[107]
+ la_iena[108] la_iena[109] la_iena[10] la_iena[110] la_iena[111] la_iena[112] la_iena[113]
+ la_iena[114] la_iena[115] la_iena[116] la_iena[117] la_iena[118] la_iena[119] la_iena[11]
+ la_iena[120] la_iena[121] la_iena[122] la_iena[123] la_iena[124] la_iena[125] la_iena[126]
+ la_iena[127] la_iena[12] la_iena[13] la_iena[14] la_iena[15] la_iena[16] la_iena[17]
+ la_iena[18] la_iena[19] la_iena[1] la_iena[20] la_iena[21] la_iena[22] la_iena[23]
+ la_iena[24] la_iena[25] la_iena[26] la_iena[27] la_iena[28] la_iena[29] la_iena[2]
+ la_iena[30] la_iena[31] la_iena[32] la_iena[33] la_iena[34] la_iena[35] la_iena[36]
+ la_iena[37] la_iena[38] la_iena[39] la_iena[3] la_iena[40] la_iena[41] la_iena[42]
+ la_iena[43] la_iena[44] la_iena[45] la_iena[46] la_iena[47] la_iena[48] la_iena[49]
+ la_iena[4] la_iena[50] la_iena[51] la_iena[52] la_iena[53] la_iena[54] la_iena[55]
+ la_iena[56] la_iena[57] la_iena[58] la_iena[59] la_iena[5] la_iena[60] la_iena[61]
+ la_iena[62] la_iena[63] la_iena[64] la_iena[65] la_iena[66] la_iena[67] la_iena[68]
+ la_iena[69] la_iena[6] la_iena[70] la_iena[71] la_iena[72] la_iena[73] la_iena[74]
+ la_iena[75] la_iena[76] la_iena[77] la_iena[78] la_iena[79] la_iena[7] la_iena[80]
+ la_iena[81] la_iena[82] la_iena[83] la_iena[84] la_iena[85] la_iena[86] la_iena[87]
+ la_iena[88] la_iena[89] la_iena[8] la_iena[90] la_iena[91] la_iena[92] la_iena[93]
+ la_iena[94] la_iena[95] la_iena[96] la_iena[97] la_iena[98] la_iena[99] la_iena[9]
+ la_input[0] la_input[100] la_input[101] la_input[102] la_input[103] la_input[104]
+ la_input[105] la_input[106] la_input[107] la_input[108] la_input[109] la_input[10]
+ la_input[110] la_input[111] la_input[112] la_input[113] la_input[114] la_input[115]
+ la_input[116] la_input[117] la_input[118] la_input[119] la_input[11] la_input[120]
+ la_input[121] la_input[122] la_input[123] la_input[124] la_input[125] la_input[126]
+ la_input[127] la_input[12] la_input[13] la_input[14] la_input[15] la_input[16] la_input[17]
+ la_input[18] la_input[19] la_input[1] la_input[20] la_input[21] la_input[22] la_input[23]
+ la_input[24] la_input[25] la_input[26] la_input[27] la_input[28] la_input[29] la_input[2]
+ la_input[30] la_input[31] la_input[32] la_input[33] la_input[34] la_input[35] la_input[36]
+ la_input[37] la_input[38] la_input[39] la_input[3] la_input[40] la_input[41] la_input[42]
+ la_input[43] la_input[44] la_input[45] la_input[46] la_input[47] la_input[48] la_input[49]
+ la_input[4] la_input[50] la_input[51] la_input[52] la_input[53] la_input[54] la_input[55]
+ la_input[56] la_input[57] la_input[58] la_input[59] la_input[5] la_input[60] la_input[61]
+ la_input[62] la_input[63] la_input[64] la_input[65] la_input[66] la_input[67] la_input[68]
+ la_input[69] la_input[6] la_input[70] la_input[71] la_input[72] la_input[73] la_input[74]
+ la_input[75] la_input[76] la_input[77] la_input[78] la_input[79] la_input[7] la_input[80]
+ la_input[81] la_input[82] la_input[83] la_input[84] la_input[85] la_input[86] la_input[87]
+ la_input[88] la_input[89] la_input[8] la_input[90] la_input[91] la_input[92] la_input[93]
+ la_input[94] la_input[95] la_input[96] la_input[97] la_input[98] la_input[99] la_input[9]
+ la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104] la_oenb[105]
+ la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109] la_oenb[10] la_oenb[110] la_oenb[111]
+ la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117] la_oenb[118]
+ la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121] la_oenb[122] la_oenb[123] la_oenb[124]
+ la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12] la_oenb[13] la_oenb[14] la_oenb[15]
+ la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20] la_oenb[21]
+ la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27] la_oenb[28]
+ la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33] la_oenb[34]
+ la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3] la_oenb[40]
+ la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46] la_oenb[47]
+ la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52] la_oenb[53]
+ la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59] la_oenb[5]
+ la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65] la_oenb[66]
+ la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6] la_oenb[70] la_oenb[71] la_oenb[72]
+ la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76] la_oenb[77] la_oenb[78] la_oenb[79]
+ la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84] la_oenb[85]
+ la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89] la_oenb[8] la_oenb[90] la_oenb[91]
+ la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97] la_oenb[98]
+ la_oenb[99] la_oenb[9] la_output[0] la_output[100] la_output[101] la_output[102]
+ la_output[103] la_output[104] la_output[105] la_output[106] la_output[107] la_output[108]
+ la_output[109] la_output[10] la_output[110] la_output[111] la_output[112] la_output[113]
+ la_output[114] la_output[115] la_output[116] la_output[117] la_output[118] la_output[119]
+ la_output[11] la_output[120] la_output[121] la_output[122] la_output[123] la_output[124]
+ la_output[125] la_output[126] la_output[127] la_output[12] la_output[13] la_output[14]
+ la_output[15] la_output[16] la_output[17] la_output[18] la_output[19] la_output[1]
+ la_output[20] la_output[21] la_output[22] la_output[23] la_output[24] la_output[25]
+ la_output[26] la_output[27] la_output[28] la_output[29] la_output[2] la_output[30]
+ la_output[31] la_output[32] la_output[33] la_output[34] la_output[35] la_output[36]
+ la_output[37] la_output[38] la_output[39] la_output[3] la_output[40] la_output[41]
+ la_output[42] la_output[43] la_output[44] la_output[45] la_output[46] la_output[47]
+ la_output[48] la_output[49] la_output[4] la_output[50] la_output[51] la_output[52]
+ la_output[53] la_output[54] la_output[55] la_output[56] la_output[57] la_output[58]
+ la_output[59] la_output[5] la_output[60] la_output[61] la_output[62] la_output[63]
+ la_output[64] la_output[65] la_output[66] la_output[67] la_output[68] la_output[69]
+ la_output[6] la_output[70] la_output[71] la_output[72] la_output[73] la_output[74]
+ la_output[75] la_output[76] la_output[77] la_output[78] la_output[79] la_output[7]
+ la_output[80] la_output[81] la_output[82] la_output[83] la_output[84] la_output[85]
+ la_output[86] la_output[87] la_output[88] la_output[89] la_output[8] la_output[90]
+ la_output[91] la_output[92] la_output[93] la_output[94] la_output[95] la_output[96]
+ la_output[97] la_output[98] la_output[99] la_output[9] mprj_ack_i mprj_adr_o[0]
+ mprj_adr_o[10] mprj_adr_o[11] mprj_adr_o[12] mprj_adr_o[13] mprj_adr_o[14] mprj_adr_o[15]
+ mprj_adr_o[16] mprj_adr_o[17] mprj_adr_o[18] mprj_adr_o[19] mprj_adr_o[1] mprj_adr_o[20]
+ mprj_adr_o[21] mprj_adr_o[22] mprj_adr_o[23] mprj_adr_o[24] mprj_adr_o[25] mprj_adr_o[26]
+ mprj_adr_o[27] mprj_adr_o[28] mprj_adr_o[29] mprj_adr_o[2] mprj_adr_o[30] mprj_adr_o[31]
+ mprj_adr_o[3] mprj_adr_o[4] mprj_adr_o[5] mprj_adr_o[6] mprj_adr_o[7] mprj_adr_o[8]
+ mprj_adr_o[9] mprj_cyc_o mprj_dat_i[0] mprj_dat_i[10] mprj_dat_i[11] mprj_dat_i[12]
+ mprj_dat_i[13] mprj_dat_i[14] mprj_dat_i[15] mprj_dat_i[16] mprj_dat_i[17] mprj_dat_i[18]
+ mprj_dat_i[19] mprj_dat_i[1] mprj_dat_i[20] mprj_dat_i[21] mprj_dat_i[22] mprj_dat_i[23]
+ mprj_dat_i[24] mprj_dat_i[25] mprj_dat_i[26] mprj_dat_i[27] mprj_dat_i[28] mprj_dat_i[29]
+ mprj_dat_i[2] mprj_dat_i[30] mprj_dat_i[31] mprj_dat_i[3] mprj_dat_i[4] mprj_dat_i[5]
+ mprj_dat_i[6] mprj_dat_i[7] mprj_dat_i[8] mprj_dat_i[9] mprj_dat_o[0] mprj_dat_o[10]
+ mprj_dat_o[11] mprj_dat_o[12] mprj_dat_o[13] mprj_dat_o[14] mprj_dat_o[15] mprj_dat_o[16]
+ mprj_dat_o[17] mprj_dat_o[18] mprj_dat_o[19] mprj_dat_o[1] mprj_dat_o[20] mprj_dat_o[21]
+ mprj_dat_o[22] mprj_dat_o[23] mprj_dat_o[24] mprj_dat_o[25] mprj_dat_o[26] mprj_dat_o[27]
+ mprj_dat_o[28] mprj_dat_o[29] mprj_dat_o[2] mprj_dat_o[30] mprj_dat_o[31] mprj_dat_o[3]
+ mprj_dat_o[4] mprj_dat_o[5] mprj_dat_o[6] mprj_dat_o[7] mprj_dat_o[8] mprj_dat_o[9]
+ mprj_sel_o[0] mprj_sel_o[1] mprj_sel_o[2] mprj_sel_o[3] mprj_stb_o mprj_wb_iena
+ mprj_we_o qspi_enabled ser_rx ser_tx spi_csb spi_enabled spi_sck spi_sdi spi_sdo
+ spi_sdoenb sram_ro_addr[0] sram_ro_addr[1] sram_ro_addr[2] sram_ro_addr[3] sram_ro_addr[4]
+ sram_ro_addr[5] sram_ro_addr[6] sram_ro_addr[7] sram_ro_clk sram_ro_csb sram_ro_data[0]
+ sram_ro_data[10] sram_ro_data[11] sram_ro_data[12] sram_ro_data[13] sram_ro_data[14]
+ sram_ro_data[15] sram_ro_data[16] sram_ro_data[17] sram_ro_data[18] sram_ro_data[19]
+ sram_ro_data[1] sram_ro_data[20] sram_ro_data[21] sram_ro_data[22] sram_ro_data[23]
+ sram_ro_data[24] sram_ro_data[25] sram_ro_data[26] sram_ro_data[27] sram_ro_data[28]
+ sram_ro_data[29] sram_ro_data[2] sram_ro_data[30] sram_ro_data[31] sram_ro_data[3]
+ sram_ro_data[4] sram_ro_data[5] sram_ro_data[6] sram_ro_data[7] sram_ro_data[8]
+ sram_ro_data[9] trap uart_enabled user_irq_ena[0] user_irq_ena[1] user_irq_ena[2]
.ends

* Black-box entry subcircuit for simple_por abstract view
.subckt simple_por vdd1v8 vdd3v3 vss3v3 porb_h por_l porb_l vss1v8
.ends

.subckt sky130_fd_sc_hd__nor2_1 A B VGND VPWR Y VNB VPB
X0 VPWR A a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_109_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VPWR Y VNB VPB
X0 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_193_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y A a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_109_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VPWR X VNB VPB
X0 a_81_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_299_297# B1 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR A1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_299_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_384_47# A1 a_81_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand2_1 A B VGND VPWR Y VNB VPB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A a_113_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_113_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VPWR X VNB VPB
X0 a_298_297# a_27_413# a_215_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_215_297# a_27_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_298_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR B1_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_382_47# A1 a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND B1_N a_27_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VPWR A1 a_298_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND A2 a_382_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VPWR X VNB VPB
X0 VPWR A1 a_382_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_297_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_297_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND A2 a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_382_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkinv_4 A VGND VPWR Y VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VPWR Y VNB VPB
X0 VPWR A a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_193_297# B a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_109_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VPWR Y VNB VPB
X0 Y A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X2 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VPWR Y VNB VPB
X0 a_377_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_47_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_129_47# B a_47_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_285_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y a_47_47# a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND A a_129_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR A a_47_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR a_47_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Y B a_377_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VPWR Y VNB VPB
X0 a_281_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND a_531_21# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR C_N a_531_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_281_297# a_531_21# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 Y a_531_21# a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND C_N a_531_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_27_297# B a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 Y a_531_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VPWR Q VNB VPB
X0 VGND a_652_21# a_586_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_956_413# a_476_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VPWR a_476_47# a_652_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_586_47# a_193_47# a_476_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X4 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5 a_476_47# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X6 a_1056_47# a_476_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X8 a_652_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_1224_47# a_27_47# a_1032_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_562_413# a_27_47# a_476_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VGND a_1032_413# a_1602_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 VPWR a_1182_261# a_1140_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 Q a_1602_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_1032_413# a_193_47# a_1056_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_476_47# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 a_1296_47# a_1182_261# a_1224_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 VPWR a_652_21# a_562_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 VPWR SET_B a_1032_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 a_1032_413# a_27_47# a_956_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 a_1182_261# a_1032_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X22 Q a_1602_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X24 a_1140_413# a_193_47# a_1032_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 VPWR a_1032_413# a_1602_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X26 a_796_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X28 a_1182_261# a_1032_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=540000u l=150000u
X29 a_652_21# a_476_47# a_796_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X31 VGND SET_B a_1296_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__inv_4 A VGND VPWR Y VNB VPB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VPWR X VNB VPB
X0 VGND A1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_510_47# B1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_79_21# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_79_21# A2 a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_297_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_79_21# C1 a_510_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_215_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__dfrtn_1 CLK_N D RESET_B VGND VPWR Q VNB VPB
X0 a_1217_47# a_193_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_1108_47# a_27_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X3 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_651_413# a_193_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR CLK_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X8 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X10 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_1108_47# a_193_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_543_47# a_193_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X13 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_543_47# a_27_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 a_1270_413# a_27_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X20 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_639_47# a_27_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X24 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 VGND CLK_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VPWR Y VNB VPB
X0 a_388_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_105_352# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_297_47# a_105_352# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_297_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR A1 a_388_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND A2 a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR B1_N a_105_352# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 Y a_105_352# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VPWR Q VNB VPB
X0 VGND a_652_21# a_586_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_956_413# a_476_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_1136_413# a_193_47# a_1028_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR a_476_47# a_652_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_586_47# a_193_47# a_476_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X5 a_1228_47# a_27_47# a_1028_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X7 a_476_47# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X8 a_1056_47# a_476_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X10 a_652_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VPWR a_1602_47# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_562_413# a_27_47# a_476_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VGND a_1028_413# a_1602_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VGND a_1602_47# Q VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 Q a_1602_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_1028_413# a_193_47# a_1056_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_476_47# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 VPWR a_1028_413# a_1602_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VPWR a_652_21# a_562_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 Q a_1602_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 a_1028_413# a_27_47# a_956_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 VPWR a_1178_261# a_1136_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X25 a_1178_261# a_1028_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X26 a_796_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 a_1300_47# a_1178_261# a_1228_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X29 a_1178_261# a_1028_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=540000u l=150000u
X30 a_652_21# a_476_47# a_796_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X31 VPWR SET_B a_1028_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X32 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X33 VGND SET_B a_1300_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VPWR Q VNB VPB
X0 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X3 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X8 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X12 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X16 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X24 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X29 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X31 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X32 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X33 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VPWR Y VNB VPB
X0 Y a_53_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_232_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR A_N a_53_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VGND A_N a_53_93# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_316_47# B a_232_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 Y a_53_93# a_316_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__xor2_1 A B VGND VPWR X VNB VPB
X0 X a_35_297# a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X B a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_35_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_117_297# B a_35_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR B a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND A a_35_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_285_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR A a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VPWR Q VNB VPB
X0 a_1178_261# a_1028_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1 VGND a_652_21# a_586_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VPWR a_1028_413# a_1598_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 a_1178_261# a_1028_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=540000u l=150000u
X4 VGND a_1598_47# Q VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_956_413# a_476_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_1136_413# a_193_47# a_1028_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR a_1598_47# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR a_476_47# a_652_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_586_47# a_193_47# a_476_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X10 VGND a_1598_47# Q VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X12 Q a_1598_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_476_47# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X14 a_1056_47# a_476_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X16 a_652_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_1224_47# a_27_47# a_1028_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 a_562_413# a_27_47# a_476_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 a_1028_413# a_193_47# a_1056_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 a_476_47# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 Q a_1598_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_1296_47# a_1178_261# a_1224_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 VGND a_1028_413# a_1598_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 VPWR a_652_21# a_562_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 VPWR a_1598_47# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 VGND SET_B a_1296_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 Q a_1598_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 a_1028_413# a_27_47# a_956_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 VPWR a_1178_261# a_1136_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X31 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X32 Q a_1598_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 a_796_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X34 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X35 Q a_1598_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X36 Q a_1598_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X37 a_652_21# a_476_47# a_796_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X38 VPWR SET_B a_1028_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X39 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VPWR Q VNB VPB
X0 Q a_1059_315# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_891_413# a_193_47# a_634_159# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2 a_561_413# a_27_47# a_466_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 Q a_1059_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VGND a_634_159# a_592_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR a_891_413# a_1059_315# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_466_413# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VPWR a_634_159# a_561_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_634_159# a_466_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X11 a_634_159# a_466_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X12 a_975_413# a_193_47# a_891_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VGND a_1059_315# a_1017_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_891_413# a_27_47# a_634_159# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 a_592_47# a_193_47# a_466_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X17 a_1017_47# a_27_47# a_891_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X18 VPWR a_1059_315# a_975_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 a_466_413# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X20 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X21 VGND a_891_413# a_1059_315# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_12 A VGND VPWR X VNB VPB
X0 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR A a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_109_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VPWR A a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND A a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VGND A a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_109_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_109_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 a_109_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VPWR Y VNB VPB
X0 VGND a_91_199# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR A a_245_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_91_199# C_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_245_297# B a_161_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_91_199# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_161_297# a_91_199# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VPWR Y VNB VPB
X0 VPWR A1 a_110_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A2 a_110_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_806_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_110_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_110_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_110_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR A1 a_110_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_27_47# B1 a_1314_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 Y A2 a_110_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 Y C1 a_978_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 Y C1 a_806_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 a_27_47# B1 a_806_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_110_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 a_806_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 a_978_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X28 a_1314_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__dlygate4sd1_1 A VGND VPWR X VNB VPB
X0 X a_299_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VPWR a_193_47# a_299_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND a_193_47# a_299_93# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 X a_299_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VPWR X VNB VPB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt caravel_clocking core_clk ext_clk ext_clk_sel ext_reset pll_clk pll_clk90
+ resetb resetb_sync sel2[0] sel2[1] sel2[2] sel[0] sel[1] sel[2] user_clk VPWR VGND
X_432_ _386_/Y _460_/Q _432_/S VGND VPWR _432_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_3_12 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xrebuffer7 _455_/Q VGND VPWR _361_/C VGND VPWR sky130_fd_sc_hd__clkbuf_2
X_363_ _363_/A _363_/B VGND VPWR _363_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
X_294_ _296_/A _476_/Q _329_/B VGND VPWR _294_/Y VGND VPWR sky130_fd_sc_hd__nand3_1
X_415_ _366_/Y _455_/Q _417_/S VGND VPWR _415_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_277_ _434_/S _278_/B _278_/C VGND VPWR _279_/A VGND VPWR sky130_fd_sc_hd__a21o_1
Xclkbuf_1_1_0_pll_clk clkbuf_0_pll_clk/X VGND VPWR _435_/A1 VGND VPWR sky130_fd_sc_hd__clkbuf_2
X_329_ _335_/A _329_/B VGND VPWR _338_/A VGND VPWR sky130_fd_sc_hd__nand2_1
Xsplit8 split8/A VGND VPWR _440_/D VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_13_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_78 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_431_ _430_/X _462_/Q _491_/Q VGND VPWR _431_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_13_101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_293_ _424_/X _291_/Y _292_/Y VGND VPWR _477_/D VGND VPWR sky130_fd_sc_hd__a21bo_1
X_362_ _361_/A _361_/C _456_/Q VGND VPWR _363_/B VGND VPWR sky130_fd_sc_hd__o21a_1
X_276_ _479_/Q VGND VPWR _278_/C VGND VPWR sky130_fd_sc_hd__clkinv_4
X_414_ _413_/X _454_/Q _467_/Q VGND VPWR _414_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_259_ _259_/A _480_/Q VGND VPWR _259_/Y VGND VPWR sky130_fd_sc_hd__nand2_1
X_328_ _324_/Y _327_/Y _291_/Y VGND VPWR _467_/D VGND VPWR sky130_fd_sc_hd__o21a_1
XFILLER_18_87 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_140 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__479__SET_B _347_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xoutput10 _399_/X VGND VPWR core_clk VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__283__A2 _439_/D VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_430_ _385_/X _462_/Q _430_/S VGND VPWR _430_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_361_ _361_/A _456_/Q _361_/C VGND VPWR _363_/A VGND VPWR sky130_fd_sc_hd__nor3_1
Xrebuffer9 _454_/Q VGND VPWR _341_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_292_ _296_/A _477_/Q _335_/B VGND VPWR _292_/Y VGND VPWR sky130_fd_sc_hd__nand3_1
X_275_ _460_/Q VGND VPWR _278_/B VGND VPWR sky130_fd_sc_hd__clkinv_4
X_413_ _337_/Y _454_/Q _417_/S VGND VPWR _413_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_120 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_258_ _482_/Q _481_/Q VGND VPWR _259_/A VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_9_79 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_68 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_327_ _325_/Y _326_/X _284_/C VGND VPWR _327_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
Xoutput11 _393_/Y VGND VPWR resetb_sync VGND VPWR sky130_fd_sc_hd__buf_2
XANTENNA__485__SET_B _347_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_291_ _291_/A _329_/B VGND VPWR _291_/Y VGND VPWR sky130_fd_sc_hd__nand2_2
X_360_ _473_/Q _472_/Q VGND VPWR _360_/Y VGND VPWR sky130_fd_sc_hd__xnor2_1
X_489_ _489_/CLK _489_/D _347_/S VGND VPWR _489_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_274_ _493_/Q _494_/Q _492_/Q VGND VPWR _434_/S VGND VPWR sky130_fd_sc_hd__nor3b_2
X_343_ _463_/Q _343_/B VGND VPWR _463_/D VGND VPWR sky130_fd_sc_hd__xnor2_1
X_412_ _365_/X _363_/B _467_/Q VGND VPWR _412_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XANTENNA__477__RESET_B _347_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_257_ _397_/S _257_/B _430_/S VGND VPWR _262_/A VGND VPWR sky130_fd_sc_hd__nand3_1
XFILLER_9_14 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_326_ _440_/D _440_/Q VGND VPWR _326_/X VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_18_45 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_309_ _466_/Q _465_/Q _464_/Q VGND VPWR _417_/S VGND VPWR sky130_fd_sc_hd__nor3b_2
XFILLER_19_120 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__445__SET_B _347_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xoutput12 _400_/X VGND VPWR user_clk VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA_input8_A sel[1] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_13_126 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_488_ _489_/CLK _488_/D _347_/S VGND VPWR _488_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XANTENNA__422__A1 _439_/D VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_290_ _290_/A _335_/B _290_/C VGND VPWR _478_/D VGND VPWR sky130_fd_sc_hd__nand3_1
XFILLER_12_14 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0_pll_clk pll_clk VGND VPWR clkbuf_0_pll_clk/X VGND VPWR sky130_fd_sc_hd__clkbuf_16
X_273_ _271_/Y _272_/A _272_/Y VGND VPWR _480_/D VGND VPWR sky130_fd_sc_hd__o21ai_1
X_411_ _360_/Y _363_/Y _467_/Q VGND VPWR _411_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_342_ _342_/A _342_/B _468_/Q VGND VPWR _343_/B VGND VPWR sky130_fd_sc_hd__nand3_1
XFILLER_2_147 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_256_ _482_/Q _481_/Q _480_/Q VGND VPWR _430_/S VGND VPWR sky130_fd_sc_hd__nor3b_2
XFILLER_0_17 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_325_ _440_/D _440_/Q VGND VPWR _325_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_18_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_239_ _243_/A _269_/B _489_/Q VGND VPWR _239_/Y VGND VPWR sky130_fd_sc_hd__nand3_1
X_308_ _471_/Q VGND VPWR _310_/B VGND VPWR sky130_fd_sc_hd__inv_2
XANTENNA__468__SET_B _347_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_13_138 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_487_ _437_/A1 _487_/D _347_/S VGND VPWR _487_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_8_131 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_345__8 _399_/X VGND VPWR _446_/CLK VGND VPWR sky130_fd_sc_hd__inv_4
X_272_ _272_/A _402_/X VGND VPWR _272_/Y VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_12_59 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_410_ _358_/Y _359_/Y _467_/Q VGND VPWR _410_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_341_ _341_/A VGND VPWR _342_/B VGND VPWR sky130_fd_sc_hd__clkinv_4
XANTENNA__486__RESET_B _347_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_255_ _483_/Q VGND VPWR _257_/B VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_324_ _324_/A _324_/B _438_/Q VGND VPWR _324_/Y VGND VPWR sky130_fd_sc_hd__nand3_1
X_238_ _238_/A _269_/B _238_/C VGND VPWR _490_/D VGND VPWR sky130_fd_sc_hd__nand3_1
X_307_ _456_/Q _455_/Q _454_/Q _306_/Y VGND VPWR _398_/S VGND VPWR sky130_fd_sc_hd__o211a_1
XFILLER_19_188 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_166 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_17 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_28 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_59 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_0 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_82 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_486_ _489_/CLK _486_/D _347_/S VGND VPWR _486_/Q VGND VPWR sky130_fd_sc_hd__dfrtn_1
X_271_ _480_/Q VGND VPWR _271_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_340_ _470_/Q _469_/Q VGND VPWR _342_/A VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_4_83 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_469_ _478_/CLK _469_/D _347_/S VGND VPWR _469_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_254_ _462_/Q _461_/Q _460_/Q _253_/Y VGND VPWR _397_/S VGND VPWR sky130_fd_sc_hd__o211a_1
X_323_ _439_/Q _439_/D VGND VPWR _324_/B VGND VPWR sky130_fd_sc_hd__or2b_1
X_237_ _243_/A _353_/A _234_/B VGND VPWR _238_/C VGND VPWR sky130_fd_sc_hd__o21bai_1
X_306_ _474_/Q _473_/Q VGND VPWR _306_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
XANTENNA__470__RESET_B _347_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_19_178 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_112 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_192 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__425__A1 _439_/D VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_485_ _485_/CLK _485_/D _347_/S VGND VPWR _485_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XANTENNA_input6_A sel2[2] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_270_ _270_/A _270_/B VGND VPWR _481_/D VGND VPWR sky130_fd_sc_hd__nand2_1
X_399_ _436_/X _355_/Y _449_/Q VGND VPWR _399_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_468_ _478_/CLK _468_/D _347_/S VGND VPWR _468_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
X_322_ _439_/D _439_/Q VGND VPWR _324_/A VGND VPWR sky130_fd_sc_hd__or2b_1
X_253_ _486_/Q _485_/Q VGND VPWR _253_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
X_236_ _236_/A VGND VPWR _243_/A VGND VPWR sky130_fd_sc_hd__clkbuf_2
Xclkbuf_1_1_0_pll_clk90 clkbuf_0_pll_clk90/X VGND VPWR _437_/A1 VGND VPWR sky130_fd_sc_hd__clkbuf_2
X_219_ _219_/A VGND VPWR _492_/D VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_0_pll_clk_A pll_clk VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA__449__RESET_B _347_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XPHY_2 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_484_ _489_/CLK _484_/D _347_/S VGND VPWR _484_/Q VGND VPWR sky130_fd_sc_hd__dfrtn_1
X_398_ _291_/Y _467_/Q _398_/S VGND VPWR _398_/X VGND VPWR sky130_fd_sc_hd__mux2_2
XANTENNA__464__RESET_B _347_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_467_ _435_/A1 _467_/D _347_/S VGND VPWR _467_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_321_ _321_/A VGND VPWR _468_/D VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0_0_pll_clk90 clkbuf_0_pll_clk90/X VGND VPWR _489_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_2
XANTENNA__463__SET_B _347_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_235_ _263_/B VGND VPWR _269_/B VGND VPWR sky130_fd_sc_hd__clkbuf_2
X_304_ _304_/A VGND VPWR _472_/D VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_10_40 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_218_ _409_/X _492_/Q _460_/Q VGND VPWR _219_/A VGND VPWR sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0_ext_clk clkbuf_0_ext_clk/X VGND VPWR _436_/A0 VGND VPWR sky130_fd_sc_hd__clkbuf_2
XANTENNA__489__RESET_B _347_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XPHY_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_483_ _483_/CLK _483_/D _347_/S VGND VPWR _483_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_16_50 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0_pll_clk clkbuf_0_pll_clk/X VGND VPWR _478_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_2
X_397_ _229_/Y _491_/Q _397_/S VGND VPWR _397_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_466_ _435_/A1 _466_/D _347_/S VGND VPWR _466_/Q VGND VPWR sky130_fd_sc_hd__dfrtn_1
X_251_ _251_/A VGND VPWR _484_/D VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_320_ _425_/X _468_/Q _320_/S VGND VPWR _321_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_449_ _435_/A1 _449_/D _347_/S VGND VPWR _449_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_234_ _353_/A _234_/B _234_/C VGND VPWR _238_/A VGND VPWR sky130_fd_sc_hd__nand3b_1
X_303_ _472_/Q _410_/X _398_/X VGND VPWR _304_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_19_72 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_217_ _217_/A VGND VPWR _493_/D VGND VPWR sky130_fd_sc_hd__clkbuf_1
XPHY_4 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_75 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_482_ _489_/CLK _482_/D _347_/S VGND VPWR _482_/Q VGND VPWR sky130_fd_sc_hd__dfrtn_1
XFILLER_16_62 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__446__SET_B _347_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_465_ _465_/CLK _465_/D _347_/S VGND VPWR _465_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XANTENNA_input4_A sel2[0] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_250_ _484_/Q _427_/X _397_/X VGND VPWR _251_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_305__5 _435_/A1 VGND VPWR _471_/CLK VGND VPWR sky130_fd_sc_hd__inv_4
X_379_ _460_/Q _461_/Q _462_/Q VGND VPWR _380_/B VGND VPWR sky130_fd_sc_hd__o21a_1
XANTENNA__492__SET_B _347_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_448_ _435_/A1 _448_/D _347_/S VGND VPWR _449_/D VGND VPWR sky130_fd_sc_hd__dfrtp_1
XANTENNA__347__S _347_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_233_ _490_/Q VGND VPWR _234_/B VGND VPWR sky130_fd_sc_hd__inv_2
X_302_ _302_/A VGND VPWR _473_/D VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_19_105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_216_ _434_/X _493_/Q _460_/Q VGND VPWR _217_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XPHY_5 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_98 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_481_ _481_/CLK _481_/D _347_/S VGND VPWR _481_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_12_144 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_464_ _435_/A1 _464_/D _347_/S VGND VPWR _464_/Q VGND VPWR sky130_fd_sc_hd__dfrtn_1
X_395_ _494_/Q _395_/B VGND VPWR _494_/D VGND VPWR sky130_fd_sc_hd__xor2_1
XANTENNA__452__SET_B _347_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_447_ _447_/CLK _447_/D _347_/S VGND VPWR hold2/A VGND VPWR sky130_fd_sc_hd__dfstp_1
X_378_ _460_/Q _462_/Q _461_/Q VGND VPWR _380_/A VGND VPWR sky130_fd_sc_hd__nor3_1
X_232_ _232_/A _487_/Q VGND VPWR _353_/A VGND VPWR sky130_fd_sc_hd__nand2_1
X_301_ _473_/Q _411_/X _398_/X VGND VPWR _302_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_1_45 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_6 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__467__RESET_B _347_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_480_ _489_/CLK _480_/D _347_/S VGND VPWR _480_/Q VGND VPWR sky130_fd_sc_hd__dfrtn_1
XFILLER_5_108 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_394_ _493_/Q _460_/Q _492_/Q VGND VPWR _395_/B VGND VPWR sky130_fd_sc_hd__nor3_1
X_463_ _435_/A1 _463_/D _347_/S VGND VPWR _463_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XANTENNA__482__RESET_B _347_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_446_ _446_/CLK hold2/X _347_/S VGND VPWR hold3/A VGND VPWR sky130_fd_sc_hd__dfstp_1
X_377_ _485_/Q _484_/Q VGND VPWR _377_/Y VGND VPWR sky130_fd_sc_hd__xnor2_1
XFILLER_8_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_0_ext_clk ext_clk VGND VPWR clkbuf_0_ext_clk/X VGND VPWR sky130_fd_sc_hd__clkbuf_16
X_231_ _489_/Q _488_/Q VGND VPWR _232_/A VGND VPWR sky130_fd_sc_hd__nor2_1
X_429_ _382_/X _380_/B _491_/Q VGND VPWR _429_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_19_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput1 ext_clk_sel VGND VPWR _392_/A VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_7 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_67 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__481__SET_B _347_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_393_ _393_/A _445_/Q VGND VPWR _393_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
X_462_ _357_/Y _462_/D _347_/S VGND VPWR _462_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_4_131 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__451__RESET_B _347_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_445_ _445_/CLK hold3/X _347_/S VGND VPWR _445_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_376_ _460_/Q _461_/Q VGND VPWR _376_/Y VGND VPWR sky130_fd_sc_hd__xnor2_1
XANTENNA_input2_A ext_reset VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_230_ _222_/Y _226_/Y _229_/Y VGND VPWR _491_/D VGND VPWR sky130_fd_sc_hd__o21a_1
X_428_ _377_/Y _380_/Y _491_/Q VGND VPWR _428_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_359_ _361_/A _361_/C VGND VPWR _359_/Y VGND VPWR sky130_fd_sc_hd__xnor2_1
Xinput2 ext_reset VGND VPWR _393_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_267__3 _489_/CLK VGND VPWR _481_/CLK VGND VPWR sky130_fd_sc_hd__inv_4
XANTENNA__458__SET_B _347_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_16_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_8 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_88 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_66 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_461_ _357_/Y _461_/D _347_/S VGND VPWR _461_/Q VGND VPWR sky130_fd_sc_hd__dfstp_4
XFILLER_4_14 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_392_ _392_/A VGND VPWR _448_/D VGND VPWR sky130_fd_sc_hd__clkinv_4
XFILLER_13_34 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__491__RESET_B _347_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_444_ _478_/CLK _444_/D VGND VPWR hold1/A VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_375_ _484_/Q VGND VPWR _375_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_427_ _375_/Y _376_/Y _491_/Q VGND VPWR _427_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_358_ _472_/Q VGND VPWR _358_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
Xinput3 resetb VGND VPWR _347_/S VGND VPWR sky130_fd_sc_hd__buf_12
X_289_ _296_/A _352_/A _284_/B VGND VPWR _290_/C VGND VPWR sky130_fd_sc_hd__o21bai_1
XPHY_9 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_34 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__421__A1 _439_/D VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_460_ _357_/Y _460_/D _347_/S VGND VPWR _460_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_391_ _493_/Q _492_/Q VGND VPWR _391_/Y VGND VPWR sky130_fd_sc_hd__xnor2_1
XFILLER_4_100 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__460__RESET_B _347_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_443_ _437_/A1 _462_/Q VGND VPWR _443_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_374_ _469_/Q _468_/Q VGND VPWR _374_/Y VGND VPWR sky130_fd_sc_hd__xnor2_1
XFILLER_6_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_357_ _278_/B _437_/X _243_/A _356_/Y VGND VPWR _357_/Y VGND VPWR sky130_fd_sc_hd__o2bb2ai_2
Xinput4 sel2[0] VGND VPWR _457_/D VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_288_ _291_/A VGND VPWR _296_/A VGND VPWR sky130_fd_sc_hd__clkbuf_2
X_426_ _374_/Y _440_/D _426_/S VGND VPWR _426_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_18_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_409_ _390_/Y _461_/Q _434_/S VGND VPWR _409_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_11_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_390_ _492_/Q VGND VPWR _390_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_346__7 _399_/X VGND VPWR _445_/CLK VGND VPWR sky130_fd_sc_hd__inv_4
X_442_ _489_/CLK _461_/Q VGND VPWR _442_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_373_ _468_/Q VGND VPWR _373_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_0_170 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__447__SET_B _347_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xinput5 sel2[1] VGND VPWR _458_/D VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_356_ _490_/Q _483_/Q VGND VPWR _356_/Y VGND VPWR sky130_fd_sc_hd__xnor2_1
X_287_ _456_/Q _455_/Q _454_/Q VGND VPWR _291_/A VGND VPWR sky130_fd_sc_hd__o21ai_1
X_425_ _373_/Y _439_/D _426_/S VGND VPWR _425_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_408_ _407_/X _462_/Q _491_/Q VGND VPWR _408_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_339_ _337_/Y _338_/A _338_/Y VGND VPWR _464_/D VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_12_139 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__454__RESET_B _347_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_14_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_187 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_441_ _437_/A1 _460_/Q VGND VPWR _441_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_1_127 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_372_ _477_/Q _372_/B VGND VPWR _372_/X VGND VPWR sky130_fd_sc_hd__xor2_1
Xclkbuf_1_0_0_ext_clk clkbuf_0_ext_clk/X VGND VPWR _347_/A1 VGND VPWR sky130_fd_sc_hd__clkbuf_2
X_286_ _329_/B VGND VPWR _335_/B VGND VPWR sky130_fd_sc_hd__clkbuf_2
X_424_ _423_/X _440_/D _467_/Q VGND VPWR _424_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_355_ _342_/B _435_/X _296_/A _354_/Y VGND VPWR _355_/Y VGND VPWR sky130_fd_sc_hd__o2bb2ai_2
XFILLER_19_47 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_14 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xinput6 sel2[2] VGND VPWR _459_/D VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_269_ _269_/A _269_/B _481_/Q VGND VPWR _270_/B VGND VPWR sky130_fd_sc_hd__nand3_1
X_407_ _389_/X _462_/Q _432_/S VGND VPWR _407_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_338_ _338_/A _414_/X VGND VPWR _338_/Y VGND VPWR sky130_fd_sc_hd__nand2_1
XANTENNA__494__RESET_B _347_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA__349__B _439_/D VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_13_49 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_371_ _476_/Q _475_/Q VGND VPWR _372_/B VGND VPWR sky130_fd_sc_hd__nor2_1
X_440_ _435_/A1 _440_/D VGND VPWR _440_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA__476__SET_B _347_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_5_83 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_92 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_285_ _467_/Q VGND VPWR _329_/B VGND VPWR sky130_fd_sc_hd__clkinv_4
X_423_ _372_/X split8/A _423_/S VGND VPWR _423_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_354_ _478_/Q _471_/Q VGND VPWR _354_/Y VGND VPWR sky130_fd_sc_hd__xnor2_1
Xinput7 sel[0] VGND VPWR _451_/D VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__448__RESET_B _347_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_4_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_268_ _272_/A _404_/X VGND VPWR _270_/A VGND VPWR sky130_fd_sc_hd__nand2_1
X_406_ _405_/X _461_/Q _491_/Q VGND VPWR _406_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_337_ _464_/Q VGND VPWR _337_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_0_pll_clk90_A pll_clk90 VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_370_ _476_/Q _475_/Q VGND VPWR _370_/Y VGND VPWR sky130_fd_sc_hd__xnor2_1
X_353_ _353_/A VGND VPWR _432_/S VGND VPWR sky130_fd_sc_hd__clkinv_4
X_422_ _421_/X _439_/D _467_/Q VGND VPWR _422_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_284_ _352_/A _284_/B _284_/C VGND VPWR _290_/A VGND VPWR sky130_fd_sc_hd__nand3b_1
Xinput8 sel[1] VGND VPWR _452_/D VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_19_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_405_ _387_/Y _461_/Q _432_/S VGND VPWR _405_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_336_ _336_/A _336_/B VGND VPWR _465_/D VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_17_191 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__439__D _439_/D VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_319_ _319_/A VGND VPWR _469_/D VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_11_131 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_300__4 _478_/CLK VGND VPWR _473_/CLK VGND VPWR sky130_fd_sc_hd__inv_4
XFILLER_12_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input9_A sel[2] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_0_196 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_421_ _370_/Y _439_/D _423_/S VGND VPWR _421_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xinput9 sel[2] VGND VPWR _453_/D VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_352_ _352_/A VGND VPWR _423_/S VGND VPWR sky130_fd_sc_hd__clkinv_4
X_283_ _440_/D _439_/D _454_/Q VGND VPWR _284_/C VGND VPWR sky130_fd_sc_hd__o21a_1
XANTENNA__457__RESET_B _347_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_266_ _266_/A _266_/B VGND VPWR _482_/D VGND VPWR sky130_fd_sc_hd__nand2_1
X_404_ _403_/X _461_/Q _491_/Q VGND VPWR _404_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_335_ _335_/A _335_/B _465_/Q VGND VPWR _336_/B VGND VPWR sky130_fd_sc_hd__nand3_1
XFILLER_2_42 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_249_ _249_/A VGND VPWR _485_/D VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_318_ _426_/X _469_/Q _320_/S VGND VPWR _319_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XANTENNA__472__RESET_B _347_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_11_143 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_396__13 VGND VGND VPWR VPWR _396__13/HI _447_/D sky130_fd_sc_hd__conb_1
Xhold1 hold1/A VGND VPWR hold1/X VGND VPWR sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA__465__SET_B _347_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_14_40 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_420_ _419_/X _420_/A1 _467_/Q VGND VPWR _420_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_282_ _478_/Q VGND VPWR _284_/B VGND VPWR sky130_fd_sc_hd__inv_2
X_351_ _470_/Q _469_/Q _468_/Q VGND VPWR _426_/S VGND VPWR sky130_fd_sc_hd__nor3b_1
XFILLER_18_138 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_403_ _383_/Y _461_/Q _430_/S VGND VPWR _403_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_334_ _338_/A _416_/X VGND VPWR _336_/A VGND VPWR sky130_fd_sc_hd__nand2_1
XANTENNA__323__B_N _439_/D VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_265_ _269_/A _269_/B _482_/Q VGND VPWR _266_/B VGND VPWR sky130_fd_sc_hd__nand3_1
XFILLER_2_10 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_30 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_196 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_248_ _485_/Q _428_/X _397_/X VGND VPWR _249_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_317_ _470_/Q _317_/B VGND VPWR _470_/D VGND VPWR sky130_fd_sc_hd__xor2_1
XANTENNA__488__SET_B _347_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_4_107 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold2 hold2/A VGND VPWR hold2/X VGND VPWR sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA__471__SET_B _347_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_0_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_350_ _462_/Q _461_/Q VGND VPWR _437_/S VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_14_52 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_281_ _281_/A _475_/Q VGND VPWR _352_/A VGND VPWR sky130_fd_sc_hd__nand2_1
X_479_ _437_/A1 _479_/D _347_/S VGND VPWR _479_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XANTENNA__466__RESET_B _347_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_264_ _272_/A _431_/X VGND VPWR _266_/A VGND VPWR sky130_fd_sc_hd__nand2_1
X_402_ _401_/X _460_/Q _491_/Q VGND VPWR _402_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_11_75 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_316_ _454_/Q _469_/Q _468_/Q VGND VPWR _317_/B VGND VPWR sky130_fd_sc_hd__nor3_1
XFILLER_9_190 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold3 hold3/A VGND VPWR hold3/X VGND VPWR sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_144 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_122 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_99 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_280_ _477_/Q _476_/Q VGND VPWR _281_/A VGND VPWR sky130_fd_sc_hd__nor2_1
XANTENNA_input7_A sel[0] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_478_ _478_/CLK _478_/D _347_/S VGND VPWR _478_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_263_ _269_/A _263_/B VGND VPWR _272_/A VGND VPWR sky130_fd_sc_hd__nand2_1
XPHY_30 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_401_ _271_/Y _460_/Q _430_/S VGND VPWR _401_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_332_ _332_/A _332_/B VGND VPWR _466_/D VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_14_132 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_246_ _246_/A VGND VPWR _486_/D VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_315_ _315_/A _315_/B _335_/B VGND VPWR _471_/D VGND VPWR sky130_fd_sc_hd__nand3_1
XANTENNA__450__RESET_B _347_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_229_ _236_/A _263_/B VGND VPWR _229_/Y VGND VPWR sky130_fd_sc_hd__nand2_2
XFILLER_8_55 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_75 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_131 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_494_ _437_/A1 _494_/D _347_/S VGND VPWR _494_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_477_ _478_/CLK _477_/D _347_/S VGND VPWR _477_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_262_ _262_/A _262_/B _269_/B VGND VPWR _483_/D VGND VPWR sky130_fd_sc_hd__nand3_1
X_400_ _436_/X _357_/Y _449_/Q VGND VPWR _400_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XPHY_31 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_331_ _335_/A _335_/B _466_/Q VGND VPWR _332_/B VGND VPWR sky130_fd_sc_hd__nand3_1
XANTENNA__475__RESET_B _347_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_245_ _486_/Q _429_/X _397_/X VGND VPWR _246_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_314_ _312_/Y _335_/A _310_/B VGND VPWR _315_/B VGND VPWR sky130_fd_sc_hd__o21bai_1
XFILLER_0_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_228_ _491_/Q VGND VPWR _263_/B VGND VPWR sky130_fd_sc_hd__clkinv_4
X_493_ _437_/A1 _493_/D _347_/S VGND VPWR _493_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XANTENNA__322__A _439_/D VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_476_ _478_/CLK _476_/D _347_/S VGND VPWR _476_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_261_ _259_/Y _269_/A _257_/B VGND VPWR _262_/B VGND VPWR sky130_fd_sc_hd__o21bai_1
XPHY_32 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_330_ _338_/A _418_/X VGND VPWR _332_/A VGND VPWR sky130_fd_sc_hd__nand2_1
X_333__6 _435_/A1 VGND VPWR _465_/CLK VGND VPWR sky130_fd_sc_hd__inv_4
XPHY_10 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_459_ _357_/Y _459_/D _347_/S VGND VPWR _462_/D VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_244_ _433_/X _229_/Y _243_/Y VGND VPWR _487_/D VGND VPWR sky130_fd_sc_hd__a21bo_1
X_313_ _313_/A1 _313_/A2 _313_/B1 _306_/Y VGND VPWR _335_/A VGND VPWR sky130_fd_sc_hd__o211ai_4
XANTENNA__483__SET_B _347_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_227_ _462_/Q _461_/Q _460_/Q VGND VPWR _236_/A VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_3_166 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_199 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__469__RESET_B _347_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_492_ _437_/A1 _492_/D _347_/S VGND VPWR _492_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_475_ _435_/A1 _475_/D _347_/S VGND VPWR _475_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XPHY_33 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input5_A sel2[1] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_260_ _462_/Q _461_/Q _460_/Q _253_/Y VGND VPWR _269_/A VGND VPWR sky130_fd_sc_hd__o211ai_4
XPHY_22 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_458_ _357_/Y _458_/D _347_/S VGND VPWR _461_/D VGND VPWR sky130_fd_sc_hd__dfstp_1
X_389_ _489_/Q _389_/B VGND VPWR _389_/X VGND VPWR sky130_fd_sc_hd__xor2_1
XANTENNA__484__RESET_B _347_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_14_146 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_243_ _243_/A _263_/B _487_/Q VGND VPWR _243_/Y VGND VPWR sky130_fd_sc_hd__nand3_1
X_312_ _312_/A _464_/Q VGND VPWR _312_/Y VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_13_190 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_226_ _223_/Y _224_/X _234_/C VGND VPWR _226_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
X_491_ _437_/A1 _491_/D _347_/S VGND VPWR _491_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_474_ _478_/CLK _474_/D _347_/S VGND VPWR _474_/Q VGND VPWR sky130_fd_sc_hd__dfrtn_1
XPHY_12 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_199 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__453__RESET_B _347_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_388_ _488_/Q _487_/Q VGND VPWR _389_/B VGND VPWR sky130_fd_sc_hd__nor2_1
X_457_ _357_/Y _457_/D _347_/S VGND VPWR _460_/D VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_242_ _406_/X _229_/Y _241_/Y VGND VPWR _488_/D VGND VPWR sky130_fd_sc_hd__a21bo_1
X_311_ _466_/Q _465_/Q VGND VPWR _312_/A VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_9_151 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_225_ _462_/Q _461_/Q _460_/Q VGND VPWR _234_/C VGND VPWR sky130_fd_sc_hd__o21a_1
X_490_ _437_/A1 _490_/D _347_/S VGND VPWR _490_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_0_105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_36 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_473_ _473_/CLK _473_/D _347_/S VGND VPWR _473_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XPHY_35 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__493__RESET_B _347_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_9_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_13 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_387_ _488_/Q _487_/Q VGND VPWR _387_/Y VGND VPWR sky130_fd_sc_hd__xnor2_1
X_456_ _355_/Y _456_/D _347_/S VGND VPWR _456_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_310_ _310_/A _310_/B _417_/S VGND VPWR _315_/A VGND VPWR sky130_fd_sc_hd__nand3_1
X_241_ _243_/A _263_/B _488_/Q VGND VPWR _241_/Y VGND VPWR sky130_fd_sc_hd__nand3_1
X_439_ _435_/A1 _439_/D VGND VPWR _439_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_224_ _462_/Q _443_/Q VGND VPWR _224_/X VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_17_47 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_147 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_472_ _478_/CLK _472_/D _347_/S VGND VPWR _472_/Q VGND VPWR sky130_fd_sc_hd__dfrtn_1
XPHY_36 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xrebuffer10 _454_/Q VGND VPWR _313_/B1 VGND VPWR sky130_fd_sc_hd__clkbuf_1
XPHY_14 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__462__RESET_B _347_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_386_ _487_/Q VGND VPWR _386_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_455_ _355_/Y _455_/D _347_/S VGND VPWR _455_/Q VGND VPWR sky130_fd_sc_hd__dfstp_4
XANTENNA_input3_A resetb VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_11_49 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_344__9 _399_/X VGND VPWR _447_/CLK VGND VPWR sky130_fd_sc_hd__inv_4
X_240_ _408_/X _229_/Y _239_/Y VGND VPWR _489_/D VGND VPWR sky130_fd_sc_hd__a21bo_1
X_369_ _475_/Q VGND VPWR _369_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_438_ _435_/A1 _454_/Q VGND VPWR _438_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_223_ _462_/Q _443_/Q VGND VPWR _223_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_2_170 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__487__RESET_B _347_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xsplit15 _456_/Q VGND VPWR split8/A VGND VPWR sky130_fd_sc_hd__clkbuf_2
XANTENNA__455__SET_B _347_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_471_ _471_/CLK _471_/D _347_/S VGND VPWR _471_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XPHY_37 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xrebuffer11 _454_/Q VGND VPWR _361_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XPHY_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_385_ _482_/Q _385_/B VGND VPWR _385_/X VGND VPWR sky130_fd_sc_hd__xor2_1
X_454_ _355_/Y _454_/D _347_/S VGND VPWR _454_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_437_ _479_/Q _437_/A1 _437_/S VGND VPWR _437_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_368_ _466_/Q _368_/B VGND VPWR _368_/X VGND VPWR sky130_fd_sc_hd__xor2_1
XFILLER_3_95 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_299_ _299_/A VGND VPWR _474_/D VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_222_ _222_/A _222_/B _441_/Q VGND VPWR _222_/Y VGND VPWR sky130_fd_sc_hd__nand3_1
XFILLER_6_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_pll_clk90 pll_clk90 VGND VPWR clkbuf_0_pll_clk90/X VGND VPWR sky130_fd_sc_hd__clkbuf_16
XANTENNA__478__SET_B _347_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA__456__RESET_B _347_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA__461__SET_B _347_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_470_ _478_/CLK _470_/D _347_/S VGND VPWR _470_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XPHY_38 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xrebuffer12 _361_/A VGND VPWR _320_/S VGND VPWR sky130_fd_sc_hd__dlygate4sd1_1
XPHY_16 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_384_ _481_/Q _480_/Q VGND VPWR _385_/B VGND VPWR sky130_fd_sc_hd__nor2_1
X_453_ _355_/Y _453_/D _347_/S VGND VPWR _456_/D VGND VPWR sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_0_ext_clk_A ext_clk VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_436_ _436_/A0 _450_/Q _449_/D VGND VPWR _436_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_367_ _465_/Q _464_/Q VGND VPWR _368_/B VGND VPWR sky130_fd_sc_hd__nor2_1
X_298_ _474_/Q _412_/X _398_/X VGND VPWR _299_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_221_ _442_/Q _461_/Q VGND VPWR _222_/B VGND VPWR sky130_fd_sc_hd__or2b_1
XFILLER_6_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_419_ _369_/Y _419_/A1 _423_/S VGND VPWR _419_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xsplit4 _455_/Q VGND VPWR _439_/D VGND VPWR sky130_fd_sc_hd__clkbuf_4
XPHY_28 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xrebuffer13 _454_/Q VGND VPWR _419_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd1_1
XPHY_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_383_ _481_/Q _480_/Q VGND VPWR _383_/Y VGND VPWR sky130_fd_sc_hd__xnor2_1
X_452_ _355_/Y _452_/D _347_/S VGND VPWR _455_/D VGND VPWR sky130_fd_sc_hd__dfstp_1
X_366_ _465_/Q _464_/Q VGND VPWR _366_/Y VGND VPWR sky130_fd_sc_hd__xnor2_1
X_297_ _420_/X _291_/Y _296_/Y VGND VPWR _475_/D VGND VPWR sky130_fd_sc_hd__a21bo_1
X_435_ _463_/Q _435_/A1 _435_/S VGND VPWR _435_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_3_20 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_220_ _461_/Q _442_/Q VGND VPWR _222_/A VGND VPWR sky130_fd_sc_hd__or2b_1
XANTENNA_input1_A ext_clk_sel VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_6_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_349_ _440_/D _439_/D VGND VPWR _435_/S VGND VPWR sky130_fd_sc_hd__nor2_1
X_418_ _417_/X split8/A _467_/Q VGND VPWR _418_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XANTENNA__490__SET_B _347_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XPHY_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_247__1 _489_/CLK VGND VPWR _485_/CLK VGND VPWR sky130_fd_sc_hd__inv_4
XPHY_18 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xrebuffer14 _419_/A1 VGND VPWR _420_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd1_1
XANTENNA__480__RESET_B _347_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_382_ _486_/Q _382_/B VGND VPWR _382_/X VGND VPWR sky130_fd_sc_hd__xor2_1
X_451_ _355_/Y _451_/D _347_/S VGND VPWR _454_/D VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_434_ _391_/Y _462_/Q _434_/S VGND VPWR _434_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_296_ _296_/A _475_/Q _329_/B VGND VPWR _296_/Y VGND VPWR sky130_fd_sc_hd__nand3_1
X_365_ _474_/Q _365_/B VGND VPWR _365_/X VGND VPWR sky130_fd_sc_hd__xor2_1
Xrebuffer5 split8/A VGND VPWR _313_/A1 VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_348_ _348_/A VGND VPWR _444_/D VGND VPWR sky130_fd_sc_hd__buf_1
X_279_ _279_/A _279_/B VGND VPWR _479_/D VGND VPWR sky130_fd_sc_hd__nand2_1
X_417_ _368_/X _456_/Q _417_/S VGND VPWR _417_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_2_196 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_252__2 _489_/CLK VGND VPWR _483_/CLK VGND VPWR sky130_fd_sc_hd__inv_4
XPHY_19 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_450_ _435_/A1 hold1/X _347_/S VGND VPWR _450_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_381_ _485_/Q _484_/Q VGND VPWR _382_/B VGND VPWR sky130_fd_sc_hd__nor2_1
X_433_ _432_/X _460_/Q _491_/Q VGND VPWR _433_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_295_ _422_/X _291_/Y _294_/Y VGND VPWR _476_/D VGND VPWR sky130_fd_sc_hd__a21bo_1
X_364_ _473_/Q _472_/Q VGND VPWR _365_/B VGND VPWR sky130_fd_sc_hd__nor2_1
Xrebuffer6 _455_/Q VGND VPWR _313_/A2 VGND VPWR sky130_fd_sc_hd__dlygate4sd1_1
X_347_ hold1/A _347_/A1 _347_/S VGND VPWR _348_/A VGND VPWR sky130_fd_sc_hd__mux2_2
XANTENNA__459__RESET_B _347_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_278_ _434_/S _278_/B _278_/C VGND VPWR _279_/B VGND VPWR sky130_fd_sc_hd__nand3_1
X_416_ _415_/X _455_/Q _467_/Q VGND VPWR _416_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XANTENNA__473__SET_B _347_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_9_87 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_43 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__474__RESET_B _347_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xrebuffer16 _398_/S VGND VPWR _310_/A VGND VPWR sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_6_66 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_380_ _380_/A _380_/B VGND VPWR _380_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_16_196 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
.ends

.subckt gpio_defaults_block_1803 VGND VPWR gpio_defaults[0] gpio_defaults[10] gpio_defaults[11]
+ gpio_defaults[12] gpio_defaults[1] gpio_defaults[2] gpio_defaults[3] gpio_defaults[4]
+ gpio_defaults[5] gpio_defaults[6] gpio_defaults[7] gpio_defaults[8] gpio_defaults[9]
Xgpio_default_value\[8\] VGND VGND VPWR VPWR gpio_default_value\[8\]/HI gpio_defaults[8]
+ sky130_fd_sc_hd__conb_1
Xgpio_default_value\[6\] VGND VGND VPWR VPWR gpio_default_value\[6\]/HI gpio_defaults[6]
+ sky130_fd_sc_hd__conb_1
XFILLER_1_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_0 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xgpio_default_value\[4\] VGND VGND VPWR VPWR gpio_default_value\[4\]/HI gpio_defaults[4]
+ sky130_fd_sc_hd__conb_1
XPHY_2 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_4 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_5 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xgpio_default_value\[2\] VGND VGND VPWR VPWR gpio_default_value\[2\]/HI gpio_defaults[2]
+ sky130_fd_sc_hd__conb_1
XFILLER_1_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xgpio_default_value\[12\] VGND VGND VPWR VPWR gpio_defaults[12] gpio_default_value\[12\]/LO
+ sky130_fd_sc_hd__conb_1
Xgpio_default_value\[0\] VGND VGND VPWR VPWR gpio_defaults[0] gpio_default_value\[0\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xgpio_default_value\[10\] VGND VGND VPWR VPWR gpio_default_value\[10\]/HI gpio_defaults[10]
+ sky130_fd_sc_hd__conb_1
XFILLER_1_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xgpio_default_value\[9\] VGND VGND VPWR VPWR gpio_default_value\[9\]/HI gpio_defaults[9]
+ sky130_fd_sc_hd__conb_1
XFILLER_2_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xgpio_default_value\[7\] VGND VGND VPWR VPWR gpio_default_value\[7\]/HI gpio_defaults[7]
+ sky130_fd_sc_hd__conb_1
XFILLER_2_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xgpio_default_value\[5\] VGND VGND VPWR VPWR gpio_default_value\[5\]/HI gpio_defaults[5]
+ sky130_fd_sc_hd__conb_1
XFILLER_2_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xgpio_default_value\[3\] VGND VGND VPWR VPWR gpio_default_value\[3\]/HI gpio_defaults[3]
+ sky130_fd_sc_hd__conb_1
XFILLER_2_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xgpio_default_value\[1\] VGND VGND VPWR VPWR gpio_defaults[1] gpio_default_value\[1\]/LO
+ sky130_fd_sc_hd__conb_1
Xgpio_default_value\[11\] VGND VGND VPWR VPWR gpio_defaults[11] gpio_default_value\[11\]/LO
+ sky130_fd_sc_hd__conb_1
.ends

.subckt user_id_programming mask_rev[0] mask_rev[10] mask_rev[11] mask_rev[12] mask_rev[13]
+ mask_rev[14] mask_rev[15] mask_rev[16] mask_rev[17] mask_rev[18] mask_rev[19] mask_rev[1]
+ mask_rev[20] mask_rev[21] mask_rev[22] mask_rev[23] mask_rev[24] mask_rev[25] mask_rev[26]
+ mask_rev[27] mask_rev[28] mask_rev[29] mask_rev[2] mask_rev[30] mask_rev[31] mask_rev[3]
+ mask_rev[4] mask_rev[5] mask_rev[6] mask_rev[7] mask_rev[8] mask_rev[9] VGND VPWR
Xmask_rev_value\[1\] VGND VGND VPWR VPWR mask_rev_value\[1\]/HI mask_rev[1] sky130_fd_sc_hd__conb_1
XFILLER_6_12 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xmask_rev_value\[30\] VGND VGND VPWR VPWR mask_rev_value\[30\]/HI mask_rev[30] sky130_fd_sc_hd__conb_1
XFILLER_0_47 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xmask_rev_value\[23\] VGND VGND VPWR VPWR mask_rev_value\[23\]/HI mask_rev[23] sky130_fd_sc_hd__conb_1
XFILLER_0_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xmask_rev_value\[16\] VGND VGND VPWR VPWR mask_rev_value\[16\]/HI mask_rev[16] sky130_fd_sc_hd__conb_1
XFILLER_0_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xmask_rev_value\[21\] VGND VGND VPWR VPWR mask_rev_value\[21\]/HI mask_rev[21] sky130_fd_sc_hd__conb_1
XFILLER_3_6 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_28 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_18 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_0 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xmask_rev_value\[14\] VGND VGND VPWR VPWR mask_rev_value\[14\]/HI mask_rev[14] sky130_fd_sc_hd__conb_1
XPHY_1 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xmask_rev_value\[8\] VGND VGND VPWR VPWR mask_rev_value\[8\]/HI mask_rev[8] sky130_fd_sc_hd__conb_1
XPHY_2 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_6 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xmask_rev_value\[12\] VGND VGND VPWR VPWR mask_rev_value\[12\]/HI mask_rev[12] sky130_fd_sc_hd__conb_1
XPHY_4 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_10 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xmask_rev_value\[6\] VGND VGND VPWR VPWR mask_rev_value\[6\]/HI mask_rev[6] sky130_fd_sc_hd__conb_1
XFILLER_1_33 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_5 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_6 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xmask_rev_value\[28\] VGND VGND VPWR VPWR mask_rev_value\[28\]/HI mask_rev[28] sky130_fd_sc_hd__conb_1
XFILLER_8_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_24 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xmask_rev_value\[10\] VGND VGND VPWR VPWR mask_rev_value\[10\]/HI mask_rev[10] sky130_fd_sc_hd__conb_1
XPHY_7 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_46 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_35 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xmask_rev_value\[4\] VGND VGND VPWR VPWR mask_rev_value\[4\]/HI mask_rev[4] sky130_fd_sc_hd__conb_1
XFILLER_7_46 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_8 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_36 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_9 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_26 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xmask_rev_value\[26\] VGND VGND VPWR VPWR mask_rev_value\[26\]/HI mask_rev[26] sky130_fd_sc_hd__conb_1
XFILLER_6_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xmask_rev_value\[19\] VGND VGND VPWR VPWR mask_rev_value\[19\]/HI mask_rev[19] sky130_fd_sc_hd__conb_1
XFILLER_7_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xmask_rev_value\[2\] VGND VGND VPWR VPWR mask_rev_value\[2\]/HI mask_rev[2] sky130_fd_sc_hd__conb_1
Xmask_rev_value\[31\] VGND VGND VPWR VPWR mask_rev_value\[31\]/HI mask_rev[31] sky130_fd_sc_hd__conb_1
Xmask_rev_value\[24\] VGND VGND VPWR VPWR mask_rev_value\[24\]/HI mask_rev[24] sky130_fd_sc_hd__conb_1
XFILLER_5_40 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xmask_rev_value\[17\] VGND VGND VPWR VPWR mask_rev_value\[17\]/HI mask_rev[17] sky130_fd_sc_hd__conb_1
Xmask_rev_value\[0\] VGND VGND VPWR VPWR mask_rev_value\[0\]/HI mask_rev[11] sky130_fd_sc_hd__conb_1
XFILLER_5_31 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_32 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xmask_rev_value\[22\] VGND VGND VPWR VPWR mask_rev_value\[22\]/HI mask_rev[22] sky130_fd_sc_hd__conb_1
XFILLER_2_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xmask_rev_value\[15\] VGND VGND VPWR VPWR mask_rev_value\[15\]/HI mask_rev[15] sky130_fd_sc_hd__conb_1
XFILLER_2_44 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_32 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_11 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xmask_rev_value\[9\] VGND VGND VPWR VPWR mask_rev_value\[9\]/HI mask_rev[9] sky130_fd_sc_hd__conb_1
XFILLER_8_44 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_23 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xmask_rev_value\[20\] VGND VGND VPWR VPWR mask_rev_value\[20\]/HI mask_rev[20] sky130_fd_sc_hd__conb_1
XPHY_10 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xmask_rev_value\[13\] VGND VGND VPWR VPWR mask_rev_value\[13\]/HI mask_rev[13] sky130_fd_sc_hd__conb_1
Xmask_rev_value\[7\] VGND VGND VPWR VPWR mask_rev_value\[7\]/HI mask_rev[7] sky130_fd_sc_hd__conb_1
XFILLER_2_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_11 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_12 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xmask_rev_value\[29\] VGND VGND VPWR VPWR mask_rev_value\[29\]/HI mask_rev[29] sky130_fd_sc_hd__conb_1
XPHY_13 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xmask_rev_value\[11\] VGND VGND VPWR VPWR mask_rev_value\[11\]/HI mask_rev[0] sky130_fd_sc_hd__conb_1
XPHY_14 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xmask_rev_value\[5\] VGND VGND VPWR VPWR mask_rev_value\[5\]/HI mask_rev[5] sky130_fd_sc_hd__conb_1
XPHY_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xmask_rev_value\[27\] VGND VGND VPWR VPWR mask_rev_value\[27\]/HI mask_rev[27] sky130_fd_sc_hd__conb_1
XPHY_16 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_40 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_30 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_17 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_42 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xmask_rev_value\[3\] VGND VGND VPWR VPWR mask_rev_value\[3\]/HI mask_rev[3] sky130_fd_sc_hd__conb_1
XFILLER_6_32 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xmask_rev_value\[25\] VGND VGND VPWR VPWR mask_rev_value\[25\]/HI mask_rev[25] sky130_fd_sc_hd__conb_1
Xmask_rev_value\[18\] VGND VGND VPWR VPWR mask_rev_value\[18\]/HI mask_rev[18] sky130_fd_sc_hd__conb_1
.ends

.subckt gpio_defaults_block_0403 VGND VPWR gpio_defaults[0] gpio_defaults[10] gpio_defaults[11]
+ gpio_defaults[12] gpio_defaults[1] gpio_defaults[2] gpio_defaults[3] gpio_defaults[4]
+ gpio_defaults[5] gpio_defaults[6] gpio_defaults[7] gpio_defaults[8] gpio_defaults[9]
Xgpio_default_value\[8\] VGND VGND VPWR VPWR gpio_default_value\[8\]/HI gpio_defaults[8]
+ sky130_fd_sc_hd__conb_1
Xgpio_default_value\[6\] VGND VGND VPWR VPWR gpio_default_value\[6\]/HI gpio_defaults[6]
+ sky130_fd_sc_hd__conb_1
XFILLER_1_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_0 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xgpio_default_value\[4\] VGND VGND VPWR VPWR gpio_default_value\[4\]/HI gpio_defaults[4]
+ sky130_fd_sc_hd__conb_1
XPHY_2 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_4 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_5 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xgpio_default_value\[2\] VGND VGND VPWR VPWR gpio_default_value\[2\]/HI gpio_defaults[2]
+ sky130_fd_sc_hd__conb_1
XFILLER_1_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xgpio_default_value\[12\] VGND VGND VPWR VPWR gpio_default_value\[12\]/HI gpio_defaults[12]
+ sky130_fd_sc_hd__conb_1
Xgpio_default_value\[0\] VGND VGND VPWR VPWR gpio_defaults[0] gpio_default_value\[0\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xgpio_default_value\[10\] VGND VGND VPWR VPWR gpio_defaults[10] gpio_default_value\[10\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xgpio_default_value\[9\] VGND VGND VPWR VPWR gpio_default_value\[9\]/HI gpio_defaults[9]
+ sky130_fd_sc_hd__conb_1
XFILLER_2_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xgpio_default_value\[7\] VGND VGND VPWR VPWR gpio_default_value\[7\]/HI gpio_defaults[7]
+ sky130_fd_sc_hd__conb_1
XFILLER_2_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xgpio_default_value\[5\] VGND VGND VPWR VPWR gpio_default_value\[5\]/HI gpio_defaults[5]
+ sky130_fd_sc_hd__conb_1
XFILLER_2_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xgpio_default_value\[3\] VGND VGND VPWR VPWR gpio_default_value\[3\]/HI gpio_defaults[3]
+ sky130_fd_sc_hd__conb_1
XFILLER_2_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xgpio_default_value\[1\] VGND VGND VPWR VPWR gpio_defaults[1] gpio_default_value\[1\]/LO
+ sky130_fd_sc_hd__conb_1
Xgpio_default_value\[11\] VGND VGND VPWR VPWR gpio_default_value\[11\]/HI gpio_defaults[11]
+ sky130_fd_sc_hd__conb_1
.ends

.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VPWR X VNB VPB
X0 VPWR B a_207_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 X a_207_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_297_47# a_27_413# a_207_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 X a_207_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_207_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VGND B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand2_4 A B VGND VPWR Y VNB VPB
X0 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__inv_12 A VGND VPWR Y VNB VPB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_8 A VGND VPWR X VNB VPB
X0 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_4 A VGND VPWR X VNB VPB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__inv_6 A VGND VPWR Y VNB VPB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand2_8 A B VGND VPWR Y VNB VPB
X0 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VPWR X VNB VPB
X0 VPWR a_212_413# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_297_47# a_27_413# a_212_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 X a_212_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_212_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_212_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR B a_212_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VGND B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VGND a_212_413# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkinv_16 A VGND VPWR Y VNB VPB
X0 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X32 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X33 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X35 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X37 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X39 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt mprj2_logic_high HI vccd2 vssd2
XFILLER_0_57 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_209 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_69 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_15 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_81 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_1_181 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_29 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_3 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_193 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_1_95 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XPHY_0 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_1 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_1_85 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_1_41 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_53 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_2 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_3 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_1_141 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_197 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_153 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_165 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_209 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_1_57 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_113 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_69 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_169 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_125 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_15 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_181 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_137 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_193 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_1_29 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_107 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_141 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_197 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_153 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_165 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_113 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_3 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_169 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_125 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_137 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_81 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_3
Xinst vssd2 vssd2 vccd2 vccd2 HI inst/LO sky130_fd_sc_hd__conb_1
XFILLER_0_85 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_41 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_109 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_97 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_53 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_3
.ends

.subckt mprj_logic_high HI[0] HI[100] HI[101] HI[102] HI[103] HI[104] HI[105] HI[106]
+ HI[107] HI[108] HI[109] HI[10] HI[110] HI[111] HI[112] HI[113] HI[114] HI[115] HI[116]
+ HI[117] HI[118] HI[119] HI[11] HI[120] HI[121] HI[122] HI[123] HI[124] HI[125] HI[126]
+ HI[127] HI[128] HI[129] HI[12] HI[130] HI[131] HI[132] HI[133] HI[134] HI[135] HI[136]
+ HI[137] HI[138] HI[139] HI[13] HI[140] HI[141] HI[142] HI[143] HI[144] HI[145] HI[146]
+ HI[147] HI[148] HI[149] HI[14] HI[150] HI[151] HI[152] HI[153] HI[154] HI[155] HI[156]
+ HI[157] HI[158] HI[159] HI[15] HI[160] HI[161] HI[162] HI[163] HI[164] HI[165] HI[166]
+ HI[167] HI[168] HI[169] HI[16] HI[170] HI[171] HI[172] HI[173] HI[174] HI[175] HI[176]
+ HI[177] HI[178] HI[179] HI[17] HI[180] HI[181] HI[182] HI[183] HI[184] HI[185] HI[186]
+ HI[187] HI[188] HI[189] HI[18] HI[190] HI[191] HI[192] HI[193] HI[194] HI[195] HI[196]
+ HI[197] HI[198] HI[199] HI[19] HI[1] HI[200] HI[201] HI[202] HI[203] HI[204] HI[205]
+ HI[206] HI[207] HI[208] HI[209] HI[20] HI[210] HI[211] HI[212] HI[213] HI[214] HI[215]
+ HI[216] HI[217] HI[218] HI[219] HI[21] HI[220] HI[221] HI[222] HI[223] HI[224] HI[225]
+ HI[226] HI[227] HI[228] HI[229] HI[22] HI[230] HI[231] HI[232] HI[233] HI[234] HI[235]
+ HI[236] HI[237] HI[238] HI[239] HI[23] HI[240] HI[241] HI[242] HI[243] HI[244] HI[245]
+ HI[246] HI[247] HI[248] HI[249] HI[24] HI[250] HI[251] HI[252] HI[253] HI[254] HI[255]
+ HI[256] HI[257] HI[258] HI[259] HI[25] HI[260] HI[261] HI[262] HI[263] HI[264] HI[265]
+ HI[266] HI[267] HI[268] HI[269] HI[26] HI[270] HI[271] HI[272] HI[273] HI[274] HI[275]
+ HI[276] HI[277] HI[278] HI[279] HI[27] HI[280] HI[281] HI[282] HI[283] HI[284] HI[285]
+ HI[286] HI[288] HI[289] HI[28] HI[290] HI[291] HI[292] HI[293] HI[294] HI[295] HI[296]
+ HI[297] HI[298] HI[299] HI[29] HI[2] HI[300] HI[301] HI[302] HI[303] HI[304] HI[305]
+ HI[306] HI[307] HI[308] HI[309] HI[30] HI[310] HI[311] HI[312] HI[313] HI[314] HI[315]
+ HI[316] HI[317] HI[318] HI[319] HI[31] HI[320] HI[321] HI[322] HI[323] HI[324] HI[325]
+ HI[326] HI[327] HI[328] HI[329] HI[32] HI[330] HI[331] HI[332] HI[333] HI[334] HI[335]
+ HI[336] HI[337] HI[338] HI[339] HI[33] HI[340] HI[341] HI[342] HI[343] HI[344] HI[345]
+ HI[346] HI[347] HI[348] HI[349] HI[34] HI[350] HI[351] HI[352] HI[353] HI[354] HI[355]
+ HI[356] HI[357] HI[358] HI[359] HI[35] HI[360] HI[361] HI[362] HI[363] HI[364] HI[365]
+ HI[366] HI[367] HI[368] HI[369] HI[36] HI[370] HI[371] HI[372] HI[373] HI[374] HI[375]
+ HI[376] HI[377] HI[378] HI[379] HI[37] HI[380] HI[381] HI[382] HI[383] HI[384] HI[385]
+ HI[386] HI[387] HI[388] HI[389] HI[38] HI[390] HI[391] HI[392] HI[393] HI[394] HI[395]
+ HI[396] HI[397] HI[398] HI[399] HI[39] HI[3] HI[400] HI[401] HI[402] HI[403] HI[404]
+ HI[405] HI[406] HI[407] HI[408] HI[409] HI[40] HI[410] HI[411] HI[412] HI[413] HI[414]
+ HI[415] HI[416] HI[417] HI[418] HI[419] HI[41] HI[420] HI[421] HI[422] HI[423] HI[424]
+ HI[425] HI[426] HI[427] HI[428] HI[42] HI[430] HI[431] HI[432] HI[433] HI[434] HI[435]
+ HI[436] HI[437] HI[438] HI[439] HI[43] HI[440] HI[441] HI[442] HI[443] HI[444] HI[445]
+ HI[446] HI[447] HI[448] HI[449] HI[44] HI[450] HI[451] HI[452] HI[453] HI[454] HI[455]
+ HI[456] HI[457] HI[458] HI[459] HI[45] HI[460] HI[461] HI[462] HI[46] HI[47] HI[48]
+ HI[49] HI[4] HI[50] HI[51] HI[52] HI[53] HI[54] HI[55] HI[56] HI[57] HI[58] HI[59]
+ HI[5] HI[60] HI[61] HI[62] HI[63] HI[64] HI[65] HI[66] HI[67] HI[68] HI[69] HI[6]
+ HI[70] HI[71] HI[72] HI[73] HI[74] HI[75] HI[76] HI[77] HI[78] HI[79] HI[7] HI[80]
+ HI[81] HI[82] HI[83] HI[84] HI[85] HI[86] HI[87] HI[88] HI[89] HI[8] HI[90] HI[91]
+ HI[92] HI[93] HI[94] HI[95] HI[96] HI[97] HI[98] HI[99] HI[9] vccd1 HI[287] HI[429]
+ vssd1
Xinsts\[210\] vssd1 vssd1 vccd1 vccd1 HI[210] insts\[210\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[308\] vssd1 vssd1 vccd1 vccd1 HI[308] insts\[308\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[425\] vssd1 vssd1 vccd1 vccd1 HI[425] insts\[425\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[160\] vssd1 vssd1 vccd1 vccd1 HI[160] insts\[160\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_357 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_302 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[258\] vssd1 vssd1 vccd1 vccd1 HI[258] insts\[258\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[40\] vssd1 vssd1 vccd1 vccd1 HI[40] insts\[40\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[375\] vssd1 vssd1 vccd1 vccd1 HI[375] insts\[375\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[88\] vssd1 vssd1 vccd1 vccd1 HI[88] insts\[88\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_165 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[123\] vssd1 vssd1 vccd1 vccd1 HI[123] insts\[123\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_669 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[338\] vssd1 vssd1 vccd1 vccd1 HI[338] insts\[338\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[240\] vssd1 vssd1 vccd1 vccd1 HI[240] insts\[240\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[9\] vssd1 vssd1 vccd1 vccd1 HI[9] insts\[9\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[455\] vssd1 vssd1 vccd1 vccd1 HI[455] insts\[455\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[288\] vssd1 vssd1 vccd1 vccd1 HI[288] insts\[288\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[190\] vssd1 vssd1 vccd1 vccd1 HI[190] insts\[190\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[70\] vssd1 vssd1 vccd1 vccd1 HI[70] insts\[70\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[203\] vssd1 vssd1 vccd1 vccd1 HI[203] insts\[203\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_561 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[418\] vssd1 vssd1 vccd1 vccd1 HI[418] insts\[418\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[153\] vssd1 vssd1 vccd1 vccd1 HI[153] insts\[153\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[320\] vssd1 vssd1 vccd1 vccd1 HI[320] insts\[320\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[33\] vssd1 vssd1 vccd1 vccd1 HI[33] insts\[33\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[368\] vssd1 vssd1 vccd1 vccd1 HI[368] insts\[368\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[270\] vssd1 vssd1 vccd1 vccd1 HI[270] insts\[270\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_177 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_486 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[116\] vssd1 vssd1 vccd1 vccd1 HI[116] insts\[116\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[400\] vssd1 vssd1 vccd1 vccd1 HI[400] insts\[400\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[233\] vssd1 vssd1 vccd1 vccd1 HI[233] insts\[233\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_209 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[183\] vssd1 vssd1 vccd1 vccd1 HI[183] insts\[183\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[350\] vssd1 vssd1 vccd1 vccd1 HI[350] insts\[350\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[448\] vssd1 vssd1 vccd1 vccd1 HI[448] insts\[448\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_721 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[63\] vssd1 vssd1 vccd1 vccd1 HI[63] insts\[63\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[398\] vssd1 vssd1 vccd1 vccd1 HI[398] insts\[398\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_573 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[146\] vssd1 vssd1 vccd1 vccd1 HI[146] insts\[146\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[313\] vssd1 vssd1 vccd1 vccd1 HI[313] insts\[313\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[26\] vssd1 vssd1 vccd1 vccd1 HI[26] insts\[26\]/LO sky130_fd_sc_hd__conb_1
XFILLER_3_3 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[430\] vssd1 vssd1 vccd1 vccd1 HI[430] insts\[430\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_189 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[263\] vssd1 vssd1 vccd1 vccd1 HI[263] insts\[263\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[380\] vssd1 vssd1 vccd1 vccd1 HI[380] insts\[380\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[109\] vssd1 vssd1 vccd1 vccd1 HI[109] insts\[109\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[93\] vssd1 vssd1 vccd1 vccd1 HI[93] insts\[93\]/LO sky130_fd_sc_hd__conb_1
XFILLER_3_498 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_80 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[226\] vssd1 vssd1 vccd1 vccd1 HI[226] insts\[226\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[343\] vssd1 vssd1 vccd1 vccd1 HI[343] insts\[343\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[176\] vssd1 vssd1 vccd1 vccd1 HI[176] insts\[176\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[56\] vssd1 vssd1 vccd1 vccd1 HI[56] insts\[56\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[460\] vssd1 vssd1 vccd1 vccd1 HI[460] insts\[460\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[293\] vssd1 vssd1 vccd1 vccd1 HI[293] insts\[293\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_541 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_585 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[139\] vssd1 vssd1 vccd1 vccd1 HI[139] insts\[139\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[306\] vssd1 vssd1 vccd1 vccd1 HI[306] insts\[306\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[19\] vssd1 vssd1 vccd1 vccd1 HI[19] insts\[19\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_393 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[423\] vssd1 vssd1 vccd1 vccd1 HI[423] insts\[423\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[256\] vssd1 vssd1 vccd1 vccd1 HI[256] insts\[256\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[373\] vssd1 vssd1 vccd1 vccd1 HI[373] insts\[373\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_617 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[86\] vssd1 vssd1 vccd1 vccd1 HI[86] insts\[86\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[121\] vssd1 vssd1 vccd1 vccd1 HI[121] insts\[121\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[219\] vssd1 vssd1 vccd1 vccd1 HI[219] insts\[219\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[336\] vssd1 vssd1 vccd1 vccd1 HI[336] insts\[336\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[169\] vssd1 vssd1 vccd1 vccd1 HI[169] insts\[169\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[49\] vssd1 vssd1 vccd1 vccd1 HI[49] insts\[49\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[286\] vssd1 vssd1 vccd1 vccd1 HI[286] insts\[286\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[7\] vssd1 vssd1 vccd1 vccd1 HI[7] insts\[7\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[453\] vssd1 vssd1 vccd1 vccd1 HI[453] insts\[453\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_597 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[201\] vssd1 vssd1 vccd1 vccd1 HI[201] insts\[201\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[416\] vssd1 vssd1 vccd1 vccd1 HI[416] insts\[416\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[151\] vssd1 vssd1 vccd1 vccd1 HI[151] insts\[151\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[249\] vssd1 vssd1 vccd1 vccd1 HI[249] insts\[249\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_681 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_8
Xinsts\[31\] vssd1 vssd1 vccd1 vccd1 HI[31] insts\[31\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_629 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[366\] vssd1 vssd1 vccd1 vccd1 HI[366] insts\[366\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[199\] vssd1 vssd1 vccd1 vccd1 HI[199] insts\[199\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[79\] vssd1 vssd1 vccd1 vccd1 HI[79] insts\[79\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[114\] vssd1 vssd1 vccd1 vccd1 HI[114] insts\[114\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[329\] vssd1 vssd1 vccd1 vccd1 HI[329] insts\[329\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[231\] vssd1 vssd1 vccd1 vccd1 HI[231] insts\[231\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[446\] vssd1 vssd1 vccd1 vccd1 HI[446] insts\[446\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[181\] vssd1 vssd1 vccd1 vccd1 HI[181] insts\[181\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[279\] vssd1 vssd1 vccd1 vccd1 HI[279] insts\[279\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[61\] vssd1 vssd1 vccd1 vccd1 HI[61] insts\[61\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[396\] vssd1 vssd1 vccd1 vccd1 HI[396] insts\[396\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[144\] vssd1 vssd1 vccd1 vccd1 HI[144] insts\[144\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[409\] vssd1 vssd1 vccd1 vccd1 HI[409] insts\[409\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[311\] vssd1 vssd1 vccd1 vccd1 HI[311] insts\[311\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[24\] vssd1 vssd1 vccd1 vccd1 HI[24] insts\[24\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[359\] vssd1 vssd1 vccd1 vccd1 HI[359] insts\[359\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_3 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[261\] vssd1 vssd1 vccd1 vccd1 HI[261] insts\[261\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[107\] vssd1 vssd1 vccd1 vccd1 HI[107] insts\[107\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[91\] vssd1 vssd1 vccd1 vccd1 HI[91] insts\[91\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[224\] vssd1 vssd1 vccd1 vccd1 HI[224] insts\[224\]/LO sky130_fd_sc_hd__conb_1
XPHY_0 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[439\] vssd1 vssd1 vccd1 vccd1 HI[439] insts\[439\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[174\] vssd1 vssd1 vccd1 vccd1 HI[174] insts\[174\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[341\] vssd1 vssd1 vccd1 vccd1 HI[341] insts\[341\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[54\] vssd1 vssd1 vccd1 vccd1 HI[54] insts\[54\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[389\] vssd1 vssd1 vccd1 vccd1 HI[389] insts\[389\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[291\] vssd1 vssd1 vccd1 vccd1 HI[291] insts\[291\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[137\] vssd1 vssd1 vccd1 vccd1 HI[137] insts\[137\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[304\] vssd1 vssd1 vccd1 vccd1 HI[304] insts\[304\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[17\] vssd1 vssd1 vccd1 vccd1 HI[17] insts\[17\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[421\] vssd1 vssd1 vccd1 vccd1 HI[421] insts\[421\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[254\] vssd1 vssd1 vccd1 vccd1 HI[254] insts\[254\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[371\] vssd1 vssd1 vccd1 vccd1 HI[371] insts\[371\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[84\] vssd1 vssd1 vccd1 vccd1 HI[84] insts\[84\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[217\] vssd1 vssd1 vccd1 vccd1 HI[217] insts\[217\]/LO sky130_fd_sc_hd__conb_1
XPHY_1 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[334\] vssd1 vssd1 vccd1 vccd1 HI[334] insts\[334\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[167\] vssd1 vssd1 vccd1 vccd1 HI[167] insts\[167\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[47\] vssd1 vssd1 vccd1 vccd1 HI[47] insts\[47\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_309 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[5\] vssd1 vssd1 vccd1 vccd1 HI[5] insts\[5\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[451\] vssd1 vssd1 vccd1 vccd1 HI[451] insts\[451\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[284\] vssd1 vssd1 vccd1 vccd1 HI[284] insts\[284\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_331 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_172 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[247\] vssd1 vssd1 vccd1 vccd1 HI[247] insts\[247\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[414\] vssd1 vssd1 vccd1 vccd1 HI[414] insts\[414\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_470 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_96 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[364\] vssd1 vssd1 vccd1 vccd1 HI[364] insts\[364\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[197\] vssd1 vssd1 vccd1 vccd1 HI[197] insts\[197\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[77\] vssd1 vssd1 vccd1 vccd1 HI[77] insts\[77\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[112\] vssd1 vssd1 vccd1 vccd1 HI[112] insts\[112\]/LO sky130_fd_sc_hd__conb_1
XPHY_2 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[327\] vssd1 vssd1 vccd1 vccd1 HI[327] insts\[327\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_557 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[444\] vssd1 vssd1 vccd1 vccd1 HI[444] insts\[444\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[277\] vssd1 vssd1 vccd1 vccd1 HI[277] insts\[277\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_343 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[394\] vssd1 vssd1 vccd1 vccd1 HI[394] insts\[394\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_118 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_184 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[407\] vssd1 vssd1 vccd1 vccd1 HI[407] insts\[407\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[142\] vssd1 vssd1 vccd1 vccd1 HI[142] insts\[142\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[22\] vssd1 vssd1 vccd1 vccd1 HI[22] insts\[22\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[357\] vssd1 vssd1 vccd1 vccd1 HI[357] insts\[357\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[105\] vssd1 vssd1 vccd1 vccd1 HI[105] insts\[105\]/LO sky130_fd_sc_hd__conb_1
XPHY_3 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[222\] vssd1 vssd1 vccd1 vccd1 HI[222] insts\[222\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[437\] vssd1 vssd1 vccd1 vccd1 HI[437] insts\[437\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[172\] vssd1 vssd1 vccd1 vccd1 HI[172] insts\[172\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_355 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[52\] vssd1 vssd1 vccd1 vccd1 HI[52] insts\[52\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[387\] vssd1 vssd1 vccd1 vccd1 HI[387] insts\[387\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_196 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_8
Xinsts\[135\] vssd1 vssd1 vccd1 vccd1 HI[135] insts\[135\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[302\] vssd1 vssd1 vccd1 vccd1 HI[302] insts\[302\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[15\] vssd1 vssd1 vccd1 vccd1 HI[15] insts\[15\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[252\] vssd1 vssd1 vccd1 vccd1 HI[252] insts\[252\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[82\] vssd1 vssd1 vccd1 vccd1 HI[82] insts\[82\]/LO sky130_fd_sc_hd__conb_1
XPHY_4 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[215\] vssd1 vssd1 vccd1 vccd1 HI[215] insts\[215\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[165\] vssd1 vssd1 vccd1 vccd1 HI[165] insts\[165\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[332\] vssd1 vssd1 vccd1 vccd1 HI[332] insts\[332\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_301 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_367 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[45\] vssd1 vssd1 vccd1 vccd1 HI[45] insts\[45\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_109 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[3\] vssd1 vssd1 vccd1 vccd1 HI[3] insts\[3\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_142 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[282\] vssd1 vssd1 vccd1 vccd1 HI[282] insts\[282\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[128\] vssd1 vssd1 vccd1 vccd1 HI[128] insts\[128\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[412\] vssd1 vssd1 vccd1 vccd1 HI[412] insts\[412\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[245\] vssd1 vssd1 vccd1 vccd1 HI[245] insts\[245\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[362\] vssd1 vssd1 vccd1 vccd1 HI[362] insts\[362\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[195\] vssd1 vssd1 vccd1 vccd1 HI[195] insts\[195\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[75\] vssd1 vssd1 vccd1 vccd1 HI[75] insts\[75\]/LO sky130_fd_sc_hd__conb_1
XPHY_5 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[110\] vssd1 vssd1 vccd1 vccd1 HI[110] insts\[110\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[208\] vssd1 vssd1 vccd1 vccd1 HI[208] insts\[208\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_505 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[158\] vssd1 vssd1 vccd1 vccd1 HI[158] insts\[158\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[325\] vssd1 vssd1 vccd1 vccd1 HI[325] insts\[325\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_379 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[38\] vssd1 vssd1 vccd1 vccd1 HI[38] insts\[38\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[442\] vssd1 vssd1 vccd1 vccd1 HI[442] insts\[442\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[275\] vssd1 vssd1 vccd1 vccd1 HI[275] insts\[275\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_154 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_121 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[392\] vssd1 vssd1 vccd1 vccd1 HI[392] insts\[392\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[405\] vssd1 vssd1 vccd1 vccd1 HI[405] insts\[405\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[140\] vssd1 vssd1 vccd1 vccd1 HI[140] insts\[140\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[238\] vssd1 vssd1 vccd1 vccd1 HI[238] insts\[238\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[20\] vssd1 vssd1 vccd1 vccd1 HI[20] insts\[20\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[355\] vssd1 vssd1 vccd1 vccd1 HI[355] insts\[355\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[188\] vssd1 vssd1 vccd1 vccd1 HI[188] insts\[188\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_709 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[68\] vssd1 vssd1 vccd1 vccd1 HI[68] insts\[68\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_517 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[103\] vssd1 vssd1 vccd1 vccd1 HI[103] insts\[103\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[318\] vssd1 vssd1 vccd1 vccd1 HI[318] insts\[318\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[220\] vssd1 vssd1 vccd1 vccd1 HI[220] insts\[220\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[170\] vssd1 vssd1 vccd1 vccd1 HI[170] insts\[170\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[435\] vssd1 vssd1 vccd1 vccd1 HI[435] insts\[435\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_689 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_645 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_601 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_133 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[268\] vssd1 vssd1 vccd1 vccd1 HI[268] insts\[268\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[50\] vssd1 vssd1 vccd1 vccd1 HI[50] insts\[50\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[385\] vssd1 vssd1 vccd1 vccd1 HI[385] insts\[385\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[98\] vssd1 vssd1 vccd1 vccd1 HI[98] insts\[98\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_442 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_68 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[133\] vssd1 vssd1 vccd1 vccd1 HI[133] insts\[133\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[300\] vssd1 vssd1 vccd1 vccd1 HI[300] insts\[300\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[13\] vssd1 vssd1 vccd1 vccd1 HI[13] insts\[13\]/LO sky130_fd_sc_hd__conb_1
XPHY_7 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[348\] vssd1 vssd1 vccd1 vccd1 HI[348] insts\[348\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[250\] vssd1 vssd1 vccd1 vccd1 HI[250] insts\[250\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[298\] vssd1 vssd1 vccd1 vccd1 HI[298] insts\[298\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_529 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[80\] vssd1 vssd1 vccd1 vccd1 HI[80] insts\[80\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[213\] vssd1 vssd1 vccd1 vccd1 HI[213] insts\[213\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_337 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[428\] vssd1 vssd1 vccd1 vccd1 HI[428] insts\[428\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_657 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_613 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[330\] vssd1 vssd1 vccd1 vccd1 HI[330] insts\[330\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[163\] vssd1 vssd1 vccd1 vccd1 HI[163] insts\[163\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[43\] vssd1 vssd1 vccd1 vccd1 HI[43] insts\[43\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[378\] vssd1 vssd1 vccd1 vccd1 HI[378] insts\[378\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[280\] vssd1 vssd1 vccd1 vccd1 HI[280] insts\[280\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[1\] vssd1 vssd1 vccd1 vccd1 HI[1] insts\[1\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_454 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_421 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_410 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_8
Xinsts\[126\] vssd1 vssd1 vccd1 vccd1 HI[126] insts\[126\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[410\] vssd1 vssd1 vccd1 vccd1 HI[410] insts\[410\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[243\] vssd1 vssd1 vccd1 vccd1 HI[243] insts\[243\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[458\] vssd1 vssd1 vccd1 vccd1 HI[458] insts\[458\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[360\] vssd1 vssd1 vccd1 vccd1 HI[360] insts\[360\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[193\] vssd1 vssd1 vccd1 vccd1 HI[193] insts\[193\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[73\] vssd1 vssd1 vccd1 vccd1 HI[73] insts\[73\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[206\] vssd1 vssd1 vccd1 vccd1 HI[206] insts\[206\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_669 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_625 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_113 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[156\] vssd1 vssd1 vccd1 vccd1 HI[156] insts\[156\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[323\] vssd1 vssd1 vccd1 vccd1 HI[323] insts\[323\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[36\] vssd1 vssd1 vccd1 vccd1 HI[36] insts\[36\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[273\] vssd1 vssd1 vccd1 vccd1 HI[273] insts\[273\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[440\] vssd1 vssd1 vccd1 vccd1 HI[440] insts\[440\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_433 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[390\] vssd1 vssd1 vccd1 vccd1 HI[390] insts\[390\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[119\] vssd1 vssd1 vccd1 vccd1 HI[119] insts\[119\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[403\] vssd1 vssd1 vccd1 vccd1 HI[403] insts\[403\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[236\] vssd1 vssd1 vccd1 vccd1 HI[236] insts\[236\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_701 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[353\] vssd1 vssd1 vccd1 vccd1 HI[353] insts\[353\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[186\] vssd1 vssd1 vccd1 vccd1 HI[186] insts\[186\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[66\] vssd1 vssd1 vccd1 vccd1 HI[66] insts\[66\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[101\] vssd1 vssd1 vccd1 vccd1 HI[101] insts\[101\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[149\] vssd1 vssd1 vccd1 vccd1 HI[149] insts\[149\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_637 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[316\] vssd1 vssd1 vccd1 vccd1 HI[316] insts\[316\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[29\] vssd1 vssd1 vccd1 vccd1 HI[29] insts\[29\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[433\] vssd1 vssd1 vccd1 vccd1 HI[433] insts\[433\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[266\] vssd1 vssd1 vccd1 vccd1 HI[266] insts\[266\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[383\] vssd1 vssd1 vccd1 vccd1 HI[383] insts\[383\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[96\] vssd1 vssd1 vccd1 vccd1 HI[96] insts\[96\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_253 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[131\] vssd1 vssd1 vccd1 vccd1 HI[131] insts\[131\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[229\] vssd1 vssd1 vccd1 vccd1 HI[229] insts\[229\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_713 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[11\] vssd1 vssd1 vccd1 vccd1 HI[11] insts\[11\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[346\] vssd1 vssd1 vccd1 vccd1 HI[346] insts\[346\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[179\] vssd1 vssd1 vccd1 vccd1 HI[179] insts\[179\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[59\] vssd1 vssd1 vccd1 vccd1 HI[59] insts\[59\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_307 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[296\] vssd1 vssd1 vccd1 vccd1 HI[296] insts\[296\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[309\] vssd1 vssd1 vccd1 vccd1 HI[309] insts\[309\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[211\] vssd1 vssd1 vccd1 vccd1 HI[211] insts\[211\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[426\] vssd1 vssd1 vccd1 vccd1 HI[426] insts\[426\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[161\] vssd1 vssd1 vccd1 vccd1 HI[161] insts\[161\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[259\] vssd1 vssd1 vccd1 vccd1 HI[259] insts\[259\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[41\] vssd1 vssd1 vccd1 vccd1 HI[41] insts\[41\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_490 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_722 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[376\] vssd1 vssd1 vccd1 vccd1 HI[376] insts\[376\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_265 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_221 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[89\] vssd1 vssd1 vccd1 vccd1 HI[89] insts\[89\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_60 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[124\] vssd1 vssd1 vccd1 vccd1 HI[124] insts\[124\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_725 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[241\] vssd1 vssd1 vccd1 vccd1 HI[241] insts\[241\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[339\] vssd1 vssd1 vccd1 vccd1 HI[339] insts\[339\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_319 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_8
Xinsts\[456\] vssd1 vssd1 vccd1 vccd1 HI[456] insts\[456\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[289\] vssd1 vssd1 vccd1 vccd1 HI[289] insts\[289\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[191\] vssd1 vssd1 vccd1 vccd1 HI[191] insts\[191\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[71\] vssd1 vssd1 vccd1 vccd1 HI[71] insts\[71\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[204\] vssd1 vssd1 vccd1 vccd1 HI[204] insts\[204\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[419\] vssd1 vssd1 vccd1 vccd1 HI[419] insts\[419\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[154\] vssd1 vssd1 vccd1 vccd1 HI[154] insts\[154\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[321\] vssd1 vssd1 vccd1 vccd1 HI[321] insts\[321\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[34\] vssd1 vssd1 vccd1 vccd1 HI[34] insts\[34\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[369\] vssd1 vssd1 vccd1 vccd1 HI[369] insts\[369\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_277 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_233 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[271\] vssd1 vssd1 vccd1 vccd1 HI[271] insts\[271\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_72 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[117\] vssd1 vssd1 vccd1 vccd1 HI[117] insts\[117\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[234\] vssd1 vssd1 vccd1 vccd1 HI[234] insts\[234\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[401\] vssd1 vssd1 vccd1 vccd1 HI[401] insts\[401\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[351\] vssd1 vssd1 vccd1 vccd1 HI[351] insts\[351\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[449\] vssd1 vssd1 vccd1 vccd1 HI[449] insts\[449\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[184\] vssd1 vssd1 vccd1 vccd1 HI[184] insts\[184\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[64\] vssd1 vssd1 vccd1 vccd1 HI[64] insts\[64\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[399\] vssd1 vssd1 vccd1 vccd1 HI[399] insts\[399\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_673 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[147\] vssd1 vssd1 vccd1 vccd1 HI[147] insts\[147\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[314\] vssd1 vssd1 vccd1 vccd1 HI[314] insts\[314\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[27\] vssd1 vssd1 vccd1 vccd1 HI[27] insts\[27\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[431\] vssd1 vssd1 vccd1 vccd1 HI[431] insts\[431\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_289 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_245 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[264\] vssd1 vssd1 vccd1 vccd1 HI[264] insts\[264\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[381\] vssd1 vssd1 vccd1 vccd1 HI[381] insts\[381\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[94\] vssd1 vssd1 vccd1 vccd1 HI[94] insts\[94\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[227\] vssd1 vssd1 vccd1 vccd1 HI[227] insts\[227\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[344\] vssd1 vssd1 vccd1 vccd1 HI[344] insts\[344\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[177\] vssd1 vssd1 vccd1 vccd1 HI[177] insts\[177\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[57\] vssd1 vssd1 vccd1 vccd1 HI[57] insts\[57\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[461\] vssd1 vssd1 vccd1 vccd1 HI[461] insts\[461\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[294\] vssd1 vssd1 vccd1 vccd1 HI[294] insts\[294\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_641 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_685 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[307\] vssd1 vssd1 vccd1 vccd1 HI[307] insts\[307\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_471 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_8
Xinsts\[424\] vssd1 vssd1 vccd1 vccd1 HI[424] insts\[424\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[257\] vssd1 vssd1 vccd1 vccd1 HI[257] insts\[257\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_85 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_511 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[374\] vssd1 vssd1 vccd1 vccd1 HI[374] insts\[374\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[87\] vssd1 vssd1 vccd1 vccd1 HI[87] insts\[87\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[122\] vssd1 vssd1 vccd1 vccd1 HI[122] insts\[122\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[337\] vssd1 vssd1 vccd1 vccd1 HI[337] insts\[337\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_108 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[8\] vssd1 vssd1 vccd1 vccd1 HI[8] insts\[8\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[454\] vssd1 vssd1 vccd1 vccd1 HI[454] insts\[454\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[287\] vssd1 vssd1 vccd1 vccd1 HI[287] insts\[287\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_653 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_697 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[202\] vssd1 vssd1 vccd1 vccd1 HI[202] insts\[202\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_461 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[417\] vssd1 vssd1 vccd1 vccd1 HI[417] insts\[417\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[152\] vssd1 vssd1 vccd1 vccd1 HI[152] insts\[152\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_97 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[32\] vssd1 vssd1 vccd1 vccd1 HI[32] insts\[32\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[367\] vssd1 vssd1 vccd1 vccd1 HI[367] insts\[367\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[115\] vssd1 vssd1 vccd1 vccd1 HI[115] insts\[115\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[232\] vssd1 vssd1 vccd1 vccd1 HI[232] insts\[232\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[447\] vssd1 vssd1 vccd1 vccd1 HI[447] insts\[447\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[182\] vssd1 vssd1 vccd1 vccd1 HI[182] insts\[182\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[62\] vssd1 vssd1 vccd1 vccd1 HI[62] insts\[62\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_665 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[397\] vssd1 vssd1 vccd1 vccd1 HI[397] insts\[397\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_484 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[145\] vssd1 vssd1 vccd1 vccd1 HI[145] insts\[145\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[312\] vssd1 vssd1 vccd1 vccd1 HI[312] insts\[312\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[25\] vssd1 vssd1 vccd1 vccd1 HI[25] insts\[25\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_281 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[262\] vssd1 vssd1 vccd1 vccd1 HI[262] insts\[262\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_3 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_8
Xinsts\[108\] vssd1 vssd1 vccd1 vccd1 HI[108] insts\[108\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[92\] vssd1 vssd1 vccd1 vccd1 HI[92] insts\[92\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[225\] vssd1 vssd1 vccd1 vccd1 HI[225] insts\[225\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[342\] vssd1 vssd1 vccd1 vccd1 HI[342] insts\[342\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[175\] vssd1 vssd1 vccd1 vccd1 HI[175] insts\[175\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[55\] vssd1 vssd1 vccd1 vccd1 HI[55] insts\[55\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[292\] vssd1 vssd1 vccd1 vccd1 HI[292] insts\[292\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_441 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[138\] vssd1 vssd1 vccd1 vccd1 HI[138] insts\[138\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[305\] vssd1 vssd1 vccd1 vccd1 HI[305] insts\[305\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[18\] vssd1 vssd1 vccd1 vccd1 HI[18] insts\[18\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_293 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_8
Xinsts\[422\] vssd1 vssd1 vccd1 vccd1 HI[422] insts\[422\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[255\] vssd1 vssd1 vccd1 vccd1 HI[255] insts\[255\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[372\] vssd1 vssd1 vccd1 vccd1 HI[372] insts\[372\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[85\] vssd1 vssd1 vccd1 vccd1 HI[85] insts\[85\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[120\] vssd1 vssd1 vccd1 vccd1 HI[120] insts\[120\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[218\] vssd1 vssd1 vccd1 vccd1 HI[218] insts\[218\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[335\] vssd1 vssd1 vccd1 vccd1 HI[335] insts\[335\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[168\] vssd1 vssd1 vccd1 vccd1 HI[168] insts\[168\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[48\] vssd1 vssd1 vccd1 vccd1 HI[48] insts\[48\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[6\] vssd1 vssd1 vccd1 vccd1 HI[6] insts\[6\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[452\] vssd1 vssd1 vccd1 vccd1 HI[452] insts\[452\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[285\] vssd1 vssd1 vccd1 vccd1 HI[285] insts\[285\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[200\] vssd1 vssd1 vccd1 vccd1 HI[200] insts\[200\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_261 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[415\] vssd1 vssd1 vccd1 vccd1 HI[415] insts\[415\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[150\] vssd1 vssd1 vccd1 vccd1 HI[150] insts\[150\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[248\] vssd1 vssd1 vccd1 vccd1 HI[248] insts\[248\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_581 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[30\] vssd1 vssd1 vccd1 vccd1 HI[30] insts\[30\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[365\] vssd1 vssd1 vccd1 vccd1 HI[365] insts\[365\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[198\] vssd1 vssd1 vccd1 vccd1 HI[198] insts\[198\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[78\] vssd1 vssd1 vccd1 vccd1 HI[78] insts\[78\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[113\] vssd1 vssd1 vccd1 vccd1 HI[113] insts\[113\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[230\] vssd1 vssd1 vccd1 vccd1 HI[230] insts\[230\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[328\] vssd1 vssd1 vccd1 vccd1 HI[328] insts\[328\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[445\] vssd1 vssd1 vccd1 vccd1 HI[445] insts\[445\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[278\] vssd1 vssd1 vccd1 vccd1 HI[278] insts\[278\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[180\] vssd1 vssd1 vccd1 vccd1 HI[180] insts\[180\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[60\] vssd1 vssd1 vccd1 vccd1 HI[60] insts\[60\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[395\] vssd1 vssd1 vccd1 vccd1 HI[395] insts\[395\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_273 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[408\] vssd1 vssd1 vccd1 vccd1 HI[408] insts\[408\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[143\] vssd1 vssd1 vccd1 vccd1 HI[143] insts\[143\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[310\] vssd1 vssd1 vccd1 vccd1 HI[310] insts\[310\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[23\] vssd1 vssd1 vccd1 vccd1 HI[23] insts\[23\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[358\] vssd1 vssd1 vccd1 vccd1 HI[358] insts\[358\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[260\] vssd1 vssd1 vccd1 vccd1 HI[260] insts\[260\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[106\] vssd1 vssd1 vccd1 vccd1 HI[106] insts\[106\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[90\] vssd1 vssd1 vccd1 vccd1 HI[90] insts\[90\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[223\] vssd1 vssd1 vccd1 vccd1 HI[223] insts\[223\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[438\] vssd1 vssd1 vccd1 vccd1 HI[438] insts\[438\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[340\] vssd1 vssd1 vccd1 vccd1 HI[340] insts\[340\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[173\] vssd1 vssd1 vccd1 vccd1 HI[173] insts\[173\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[53\] vssd1 vssd1 vccd1 vccd1 HI[53] insts\[53\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[388\] vssd1 vssd1 vccd1 vccd1 HI[388] insts\[388\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[290\] vssd1 vssd1 vccd1 vccd1 HI[290] insts\[290\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_230 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[136\] vssd1 vssd1 vccd1 vccd1 HI[136] insts\[136\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[303\] vssd1 vssd1 vccd1 vccd1 HI[303] insts\[303\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[16\] vssd1 vssd1 vccd1 vccd1 HI[16] insts\[16\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[420\] vssd1 vssd1 vccd1 vccd1 HI[420] insts\[420\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[253\] vssd1 vssd1 vccd1 vccd1 HI[253] insts\[253\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[370\] vssd1 vssd1 vccd1 vccd1 HI[370] insts\[370\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[83\] vssd1 vssd1 vccd1 vccd1 HI[83] insts\[83\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[216\] vssd1 vssd1 vccd1 vccd1 HI[216] insts\[216\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[166\] vssd1 vssd1 vccd1 vccd1 HI[166] insts\[166\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[333\] vssd1 vssd1 vccd1 vccd1 HI[333] insts\[333\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[46\] vssd1 vssd1 vccd1 vccd1 HI[46] insts\[46\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[450\] vssd1 vssd1 vccd1 vccd1 HI[450] insts\[450\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_209 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[283\] vssd1 vssd1 vccd1 vccd1 HI[283] insts\[283\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[4\] vssd1 vssd1 vccd1 vccd1 HI[4] insts\[4\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_710 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_242 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[129\] vssd1 vssd1 vccd1 vccd1 HI[129] insts\[129\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[413\] vssd1 vssd1 vccd1 vccd1 HI[413] insts\[413\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[246\] vssd1 vssd1 vccd1 vccd1 HI[246] insts\[246\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[196\] vssd1 vssd1 vccd1 vccd1 HI[196] insts\[196\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[363\] vssd1 vssd1 vccd1 vccd1 HI[363] insts\[363\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[76\] vssd1 vssd1 vccd1 vccd1 HI[76] insts\[76\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[209\] vssd1 vssd1 vccd1 vccd1 HI[209] insts\[209\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[111\] vssd1 vssd1 vccd1 vccd1 HI[111] insts\[111\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[326\] vssd1 vssd1 vccd1 vccd1 HI[326] insts\[326\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[159\] vssd1 vssd1 vccd1 vccd1 HI[159] insts\[159\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[39\] vssd1 vssd1 vccd1 vccd1 HI[39] insts\[39\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_722 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_8
Xinsts\[443\] vssd1 vssd1 vccd1 vccd1 HI[443] insts\[443\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_221 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_254 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[276\] vssd1 vssd1 vccd1 vccd1 HI[276] insts\[276\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[393\] vssd1 vssd1 vccd1 vccd1 HI[393] insts\[393\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[406\] vssd1 vssd1 vccd1 vccd1 HI[406] insts\[406\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[141\] vssd1 vssd1 vccd1 vccd1 HI[141] insts\[141\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[239\] vssd1 vssd1 vccd1 vccd1 HI[239] insts\[239\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[21\] vssd1 vssd1 vccd1 vccd1 HI[21] insts\[21\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[356\] vssd1 vssd1 vccd1 vccd1 HI[356] insts\[356\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[189\] vssd1 vssd1 vccd1 vccd1 HI[189] insts\[189\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[69\] vssd1 vssd1 vccd1 vccd1 HI[69] insts\[69\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[104\] vssd1 vssd1 vccd1 vccd1 HI[104] insts\[104\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_617 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[221\] vssd1 vssd1 vccd1 vccd1 HI[221] insts\[221\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[319\] vssd1 vssd1 vccd1 vccd1 HI[319] insts\[319\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[436\] vssd1 vssd1 vccd1 vccd1 HI[436] insts\[436\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[171\] vssd1 vssd1 vccd1 vccd1 HI[171] insts\[171\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[269\] vssd1 vssd1 vccd1 vccd1 HI[269] insts\[269\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[51\] vssd1 vssd1 vccd1 vccd1 HI[51] insts\[51\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[386\] vssd1 vssd1 vccd1 vccd1 HI[386] insts\[386\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[99\] vssd1 vssd1 vccd1 vccd1 HI[99] insts\[99\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[134\] vssd1 vssd1 vccd1 vccd1 HI[134] insts\[134\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[301\] vssd1 vssd1 vccd1 vccd1 HI[301] insts\[301\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[14\] vssd1 vssd1 vccd1 vccd1 HI[14] insts\[14\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[349\] vssd1 vssd1 vccd1 vccd1 HI[349] insts\[349\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[251\] vssd1 vssd1 vccd1 vccd1 HI[251] insts\[251\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[299\] vssd1 vssd1 vccd1 vccd1 HI[299] insts\[299\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_629 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_673 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[81\] vssd1 vssd1 vccd1 vccd1 HI[81] insts\[81\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[214\] vssd1 vssd1 vccd1 vccd1 HI[214] insts\[214\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[429\] vssd1 vssd1 vccd1 vccd1 HI[429] insts\[429\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[164\] vssd1 vssd1 vccd1 vccd1 HI[164] insts\[164\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[331\] vssd1 vssd1 vccd1 vccd1 HI[331] insts\[331\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[44\] vssd1 vssd1 vccd1 vccd1 HI[44] insts\[44\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[379\] vssd1 vssd1 vccd1 vccd1 HI[379] insts\[379\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[2\] vssd1 vssd1 vccd1 vccd1 HI[2] insts\[2\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[281\] vssd1 vssd1 vccd1 vccd1 HI[281] insts\[281\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[127\] vssd1 vssd1 vccd1 vccd1 HI[127] insts\[127\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[411\] vssd1 vssd1 vccd1 vccd1 HI[411] insts\[411\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[244\] vssd1 vssd1 vccd1 vccd1 HI[244] insts\[244\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[459\] vssd1 vssd1 vccd1 vccd1 HI[459] insts\[459\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[361\] vssd1 vssd1 vccd1 vccd1 HI[361] insts\[361\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[194\] vssd1 vssd1 vccd1 vccd1 HI[194] insts\[194\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_641 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_685 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[74\] vssd1 vssd1 vccd1 vccd1 HI[74] insts\[74\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_405 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_449 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[207\] vssd1 vssd1 vccd1 vccd1 HI[207] insts\[207\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[157\] vssd1 vssd1 vccd1 vccd1 HI[157] insts\[157\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[324\] vssd1 vssd1 vccd1 vccd1 HI[324] insts\[324\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[37\] vssd1 vssd1 vccd1 vccd1 HI[37] insts\[37\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[441\] vssd1 vssd1 vccd1 vccd1 HI[441] insts\[441\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_533 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[274\] vssd1 vssd1 vccd1 vccd1 HI[274] insts\[274\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[391\] vssd1 vssd1 vccd1 vccd1 HI[391] insts\[391\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[404\] vssd1 vssd1 vccd1 vccd1 HI[404] insts\[404\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[237\] vssd1 vssd1 vccd1 vccd1 HI[237] insts\[237\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_609 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[354\] vssd1 vssd1 vccd1 vccd1 HI[354] insts\[354\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[187\] vssd1 vssd1 vccd1 vccd1 HI[187] insts\[187\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[67\] vssd1 vssd1 vccd1 vccd1 HI[67] insts\[67\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_697 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[102\] vssd1 vssd1 vccd1 vccd1 HI[102] insts\[102\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_417 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[317\] vssd1 vssd1 vccd1 vccd1 HI[317] insts\[317\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[434\] vssd1 vssd1 vccd1 vccd1 HI[434] insts\[434\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_545 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[267\] vssd1 vssd1 vccd1 vccd1 HI[267] insts\[267\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_589 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[384\] vssd1 vssd1 vccd1 vccd1 HI[384] insts\[384\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_386 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[97\] vssd1 vssd1 vccd1 vccd1 HI[97] insts\[97\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[132\] vssd1 vssd1 vccd1 vccd1 HI[132] insts\[132\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[12\] vssd1 vssd1 vccd1 vccd1 HI[12] insts\[12\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[347\] vssd1 vssd1 vccd1 vccd1 HI[347] insts\[347\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_429 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[297\] vssd1 vssd1 vccd1 vccd1 HI[297] insts\[297\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[212\] vssd1 vssd1 vccd1 vccd1 HI[212] insts\[212\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[162\] vssd1 vssd1 vccd1 vccd1 HI[162] insts\[162\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[427\] vssd1 vssd1 vccd1 vccd1 HI[427] insts\[427\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_557 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_502 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[42\] vssd1 vssd1 vccd1 vccd1 HI[42] insts\[42\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[377\] vssd1 vssd1 vccd1 vccd1 HI[377] insts\[377\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_398 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_365 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_321 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[0\] vssd1 vssd1 vccd1 vccd1 HI[0] insts\[0\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[125\] vssd1 vssd1 vccd1 vccd1 HI[125] insts\[125\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[242\] vssd1 vssd1 vccd1 vccd1 HI[242] insts\[242\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[457\] vssd1 vssd1 vccd1 vccd1 HI[457] insts\[457\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[192\] vssd1 vssd1 vccd1 vccd1 HI[192] insts\[192\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[72\] vssd1 vssd1 vccd1 vccd1 HI[72] insts\[72\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[205\] vssd1 vssd1 vccd1 vccd1 HI[205] insts\[205\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_569 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_514 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[155\] vssd1 vssd1 vccd1 vccd1 HI[155] insts\[155\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[322\] vssd1 vssd1 vccd1 vccd1 HI[322] insts\[322\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[35\] vssd1 vssd1 vccd1 vccd1 HI[35] insts\[35\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[272\] vssd1 vssd1 vccd1 vccd1 HI[272] insts\[272\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_377 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_333 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[118\] vssd1 vssd1 vccd1 vccd1 HI[118] insts\[118\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_130 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_141 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[402\] vssd1 vssd1 vccd1 vccd1 HI[402] insts\[402\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[235\] vssd1 vssd1 vccd1 vccd1 HI[235] insts\[235\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_601 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_645 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[352\] vssd1 vssd1 vccd1 vccd1 HI[352] insts\[352\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[185\] vssd1 vssd1 vccd1 vccd1 HI[185] insts\[185\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[65\] vssd1 vssd1 vccd1 vccd1 HI[65] insts\[65\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[100\] vssd1 vssd1 vccd1 vccd1 HI[100] insts\[100\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[148\] vssd1 vssd1 vccd1 vccd1 HI[148] insts\[148\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_526 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[315\] vssd1 vssd1 vccd1 vccd1 HI[315] insts\[315\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[28\] vssd1 vssd1 vccd1 vccd1 HI[28] insts\[28\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[265\] vssd1 vssd1 vccd1 vccd1 HI[265] insts\[265\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[432\] vssd1 vssd1 vccd1 vccd1 HI[432] insts\[432\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_345 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[382\] vssd1 vssd1 vccd1 vccd1 HI[382] insts\[382\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_197 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_153 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[95\] vssd1 vssd1 vccd1 vccd1 HI[95] insts\[95\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[130\] vssd1 vssd1 vccd1 vccd1 HI[130] insts\[130\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[228\] vssd1 vssd1 vccd1 vccd1 HI[228] insts\[228\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_613 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_657 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[10\] vssd1 vssd1 vccd1 vccd1 HI[10] insts\[10\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[178\] vssd1 vssd1 vccd1 vccd1 HI[178] insts\[178\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[345\] vssd1 vssd1 vccd1 vccd1 HI[345] insts\[345\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[58\] vssd1 vssd1 vccd1 vccd1 HI[58] insts\[58\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[462\] vssd1 vssd1 vccd1 vccd1 HI[462] insts\[462\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[295\] vssd1 vssd1 vccd1 vccd1 HI[295] insts\[295\]/LO sky130_fd_sc_hd__conb_1
.ends

.subckt sky130_fd_sc_hd__inv_16 A VGND VPWR Y VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X28 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hvl__conb_1 VGND VNB VPB VPWR HI LO
R0 VGND LO sky130_fd_pr__res_generic_po w=510000u l=45000u
R1 HI VPWR sky130_fd_pr__res_generic_po w=510000u l=45000u
.ends

.subckt sky130_fd_sc_hvl__lsbufhv2lv_1 A VGND VPWR X VNB VPB LVPWR
X0 a_30_1337# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X1 VGND a_30_1337# a_30_207# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X2 VGND a_30_207# a_389_141# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X3 VGND a_30_207# a_389_141# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X4 a_389_1337# a_30_1337# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X5 VGND a_30_207# a_389_141# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X6 VGND A a_30_1337# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X7 VGND a_30_1337# a_389_1337# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X8 a_389_141# a_30_207# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X9 VGND a_30_1337# a_389_1337# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X10 LVPWR a_389_141# X LVPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X11 VGND a_389_141# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X12 a_389_1337# a_30_1337# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X13 LVPWR a_389_1337# a_389_141# LVPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X14 a_30_207# a_30_1337# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X15 a_389_1337# a_389_141# LVPWR LVPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
.ends

.subckt mgmt_protect_hv vccd vssd vdda1 vdda2 mprj2_vdd_logic1 mprj_vdd_logic1 dw_6116_1496#
+ vssa1 dw_13698_1476# vssa2
Xmprj2_logic_high_hvl vssa2 vssa2 vdda2 vdda2 mprj2_logic_high_lv/A mprj2_logic_high_hvl/LO
+ sky130_fd_sc_hvl__conb_1
Xmprj_logic_high_hvl vssa1 vssa1 vdda1 vdda1 mprj_logic_high_lv/A mprj_logic_high_hvl/LO
+ sky130_fd_sc_hvl__conb_1
Xmprj_logic_high_lv mprj_logic_high_lv/A vssd vdda1 mprj_vdd_logic1 vssd vdda1 vccd
+ sky130_fd_sc_hvl__lsbufhv2lv_1
Xmprj2_logic_high_lv mprj2_logic_high_lv/A vssd vdda2 mprj2_vdd_logic1 vssd vdda2
+ vccd sky130_fd_sc_hvl__lsbufhv2lv_1
.ends

.subckt sky130_fd_sc_hd__and2_4 A B VGND VPWR X VNB VPB
X0 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND B a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_110_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VPWR X VNB VPB
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt mgmt_protect caravel_clk caravel_clk2 caravel_rstn la_data_in_core[0] la_data_in_core[100]
+ la_data_in_core[101] la_data_in_core[102] la_data_in_core[103] la_data_in_core[104]
+ la_data_in_core[105] la_data_in_core[106] la_data_in_core[107] la_data_in_core[108]
+ la_data_in_core[109] la_data_in_core[10] la_data_in_core[110] la_data_in_core[111]
+ la_data_in_core[112] la_data_in_core[113] la_data_in_core[114] la_data_in_core[115]
+ la_data_in_core[116] la_data_in_core[117] la_data_in_core[118] la_data_in_core[119]
+ la_data_in_core[11] la_data_in_core[120] la_data_in_core[121] la_data_in_core[122]
+ la_data_in_core[123] la_data_in_core[124] la_data_in_core[125] la_data_in_core[126]
+ la_data_in_core[127] la_data_in_core[12] la_data_in_core[13] la_data_in_core[14]
+ la_data_in_core[15] la_data_in_core[16] la_data_in_core[17] la_data_in_core[18]
+ la_data_in_core[19] la_data_in_core[1] la_data_in_core[20] la_data_in_core[21] la_data_in_core[22]
+ la_data_in_core[23] la_data_in_core[24] la_data_in_core[25] la_data_in_core[26]
+ la_data_in_core[27] la_data_in_core[28] la_data_in_core[29] la_data_in_core[2] la_data_in_core[30]
+ la_data_in_core[31] la_data_in_core[32] la_data_in_core[33] la_data_in_core[34]
+ la_data_in_core[35] la_data_in_core[36] la_data_in_core[37] la_data_in_core[38]
+ la_data_in_core[39] la_data_in_core[3] la_data_in_core[40] la_data_in_core[41] la_data_in_core[42]
+ la_data_in_core[43] la_data_in_core[44] la_data_in_core[45] la_data_in_core[46]
+ la_data_in_core[47] la_data_in_core[48] la_data_in_core[49] la_data_in_core[4] la_data_in_core[50]
+ la_data_in_core[51] la_data_in_core[52] la_data_in_core[53] la_data_in_core[54]
+ la_data_in_core[55] la_data_in_core[56] la_data_in_core[57] la_data_in_core[58]
+ la_data_in_core[59] la_data_in_core[5] la_data_in_core[60] la_data_in_core[61] la_data_in_core[62]
+ la_data_in_core[63] la_data_in_core[64] la_data_in_core[65] la_data_in_core[66]
+ la_data_in_core[67] la_data_in_core[68] la_data_in_core[69] la_data_in_core[6] la_data_in_core[70]
+ la_data_in_core[71] la_data_in_core[72] la_data_in_core[73] la_data_in_core[74]
+ la_data_in_core[75] la_data_in_core[76] la_data_in_core[77] la_data_in_core[78]
+ la_data_in_core[79] la_data_in_core[7] la_data_in_core[80] la_data_in_core[81] la_data_in_core[82]
+ la_data_in_core[83] la_data_in_core[84] la_data_in_core[85] la_data_in_core[86]
+ la_data_in_core[87] la_data_in_core[88] la_data_in_core[89] la_data_in_core[8] la_data_in_core[90]
+ la_data_in_core[91] la_data_in_core[92] la_data_in_core[93] la_data_in_core[94]
+ la_data_in_core[95] la_data_in_core[96] la_data_in_core[97] la_data_in_core[98]
+ la_data_in_core[99] la_data_in_core[9] la_data_in_mprj[0] la_data_in_mprj[100] la_data_in_mprj[101]
+ la_data_in_mprj[102] la_data_in_mprj[103] la_data_in_mprj[104] la_data_in_mprj[105]
+ la_data_in_mprj[106] la_data_in_mprj[107] la_data_in_mprj[108] la_data_in_mprj[109]
+ la_data_in_mprj[10] la_data_in_mprj[110] la_data_in_mprj[111] la_data_in_mprj[112]
+ la_data_in_mprj[113] la_data_in_mprj[114] la_data_in_mprj[115] la_data_in_mprj[116]
+ la_data_in_mprj[117] la_data_in_mprj[118] la_data_in_mprj[119] la_data_in_mprj[11]
+ la_data_in_mprj[120] la_data_in_mprj[121] la_data_in_mprj[122] la_data_in_mprj[123]
+ la_data_in_mprj[124] la_data_in_mprj[125] la_data_in_mprj[126] la_data_in_mprj[127]
+ la_data_in_mprj[12] la_data_in_mprj[13] la_data_in_mprj[14] la_data_in_mprj[15]
+ la_data_in_mprj[16] la_data_in_mprj[17] la_data_in_mprj[18] la_data_in_mprj[19]
+ la_data_in_mprj[1] la_data_in_mprj[20] la_data_in_mprj[21] la_data_in_mprj[22] la_data_in_mprj[23]
+ la_data_in_mprj[24] la_data_in_mprj[25] la_data_in_mprj[26] la_data_in_mprj[27]
+ la_data_in_mprj[28] la_data_in_mprj[29] la_data_in_mprj[2] la_data_in_mprj[30] la_data_in_mprj[31]
+ la_data_in_mprj[32] la_data_in_mprj[33] la_data_in_mprj[34] la_data_in_mprj[35]
+ la_data_in_mprj[36] la_data_in_mprj[37] la_data_in_mprj[38] la_data_in_mprj[39]
+ la_data_in_mprj[3] la_data_in_mprj[40] la_data_in_mprj[41] la_data_in_mprj[42] la_data_in_mprj[43]
+ la_data_in_mprj[44] la_data_in_mprj[45] la_data_in_mprj[46] la_data_in_mprj[47]
+ la_data_in_mprj[48] la_data_in_mprj[49] la_data_in_mprj[4] la_data_in_mprj[50] la_data_in_mprj[51]
+ la_data_in_mprj[52] la_data_in_mprj[53] la_data_in_mprj[54] la_data_in_mprj[55]
+ la_data_in_mprj[56] la_data_in_mprj[57] la_data_in_mprj[58] la_data_in_mprj[59]
+ la_data_in_mprj[5] la_data_in_mprj[60] la_data_in_mprj[61] la_data_in_mprj[62] la_data_in_mprj[63]
+ la_data_in_mprj[64] la_data_in_mprj[65] la_data_in_mprj[66] la_data_in_mprj[67]
+ la_data_in_mprj[68] la_data_in_mprj[69] la_data_in_mprj[6] la_data_in_mprj[70] la_data_in_mprj[71]
+ la_data_in_mprj[72] la_data_in_mprj[73] la_data_in_mprj[74] la_data_in_mprj[75]
+ la_data_in_mprj[76] la_data_in_mprj[77] la_data_in_mprj[78] la_data_in_mprj[79]
+ la_data_in_mprj[7] la_data_in_mprj[80] la_data_in_mprj[81] la_data_in_mprj[82] la_data_in_mprj[83]
+ la_data_in_mprj[84] la_data_in_mprj[85] la_data_in_mprj[86] la_data_in_mprj[87]
+ la_data_in_mprj[88] la_data_in_mprj[89] la_data_in_mprj[8] la_data_in_mprj[90] la_data_in_mprj[91]
+ la_data_in_mprj[92] la_data_in_mprj[93] la_data_in_mprj[94] la_data_in_mprj[95]
+ la_data_in_mprj[96] la_data_in_mprj[97] la_data_in_mprj[98] la_data_in_mprj[99]
+ la_data_in_mprj[9] la_data_out_core[0] la_data_out_core[100] la_data_out_core[101]
+ la_data_out_core[102] la_data_out_core[103] la_data_out_core[104] la_data_out_core[105]
+ la_data_out_core[106] la_data_out_core[107] la_data_out_core[108] la_data_out_core[109]
+ la_data_out_core[10] la_data_out_core[110] la_data_out_core[111] la_data_out_core[112]
+ la_data_out_core[113] la_data_out_core[114] la_data_out_core[115] la_data_out_core[116]
+ la_data_out_core[117] la_data_out_core[118] la_data_out_core[119] la_data_out_core[11]
+ la_data_out_core[120] la_data_out_core[121] la_data_out_core[122] la_data_out_core[123]
+ la_data_out_core[124] la_data_out_core[125] la_data_out_core[126] la_data_out_core[127]
+ la_data_out_core[12] la_data_out_core[13] la_data_out_core[14] la_data_out_core[15]
+ la_data_out_core[16] la_data_out_core[17] la_data_out_core[18] la_data_out_core[19]
+ la_data_out_core[1] la_data_out_core[20] la_data_out_core[21] la_data_out_core[22]
+ la_data_out_core[23] la_data_out_core[24] la_data_out_core[25] la_data_out_core[26]
+ la_data_out_core[27] la_data_out_core[28] la_data_out_core[29] la_data_out_core[2]
+ la_data_out_core[30] la_data_out_core[31] la_data_out_core[32] la_data_out_core[33]
+ la_data_out_core[34] la_data_out_core[35] la_data_out_core[36] la_data_out_core[37]
+ la_data_out_core[38] la_data_out_core[39] la_data_out_core[3] la_data_out_core[40]
+ la_data_out_core[41] la_data_out_core[42] la_data_out_core[43] la_data_out_core[44]
+ la_data_out_core[45] la_data_out_core[46] la_data_out_core[47] la_data_out_core[48]
+ la_data_out_core[49] la_data_out_core[4] la_data_out_core[50] la_data_out_core[51]
+ la_data_out_core[52] la_data_out_core[53] la_data_out_core[54] la_data_out_core[55]
+ la_data_out_core[56] la_data_out_core[57] la_data_out_core[58] la_data_out_core[59]
+ la_data_out_core[5] la_data_out_core[60] la_data_out_core[61] la_data_out_core[62]
+ la_data_out_core[63] la_data_out_core[64] la_data_out_core[65] la_data_out_core[66]
+ la_data_out_core[67] la_data_out_core[68] la_data_out_core[69] la_data_out_core[6]
+ la_data_out_core[70] la_data_out_core[71] la_data_out_core[72] la_data_out_core[73]
+ la_data_out_core[74] la_data_out_core[75] la_data_out_core[76] la_data_out_core[77]
+ la_data_out_core[78] la_data_out_core[79] la_data_out_core[7] la_data_out_core[80]
+ la_data_out_core[81] la_data_out_core[82] la_data_out_core[83] la_data_out_core[84]
+ la_data_out_core[85] la_data_out_core[86] la_data_out_core[87] la_data_out_core[88]
+ la_data_out_core[89] la_data_out_core[8] la_data_out_core[90] la_data_out_core[91]
+ la_data_out_core[92] la_data_out_core[93] la_data_out_core[94] la_data_out_core[95]
+ la_data_out_core[96] la_data_out_core[97] la_data_out_core[98] la_data_out_core[99]
+ la_data_out_core[9] la_data_out_mprj[0] la_data_out_mprj[100] la_data_out_mprj[101]
+ la_data_out_mprj[102] la_data_out_mprj[103] la_data_out_mprj[104] la_data_out_mprj[105]
+ la_data_out_mprj[106] la_data_out_mprj[107] la_data_out_mprj[108] la_data_out_mprj[109]
+ la_data_out_mprj[10] la_data_out_mprj[110] la_data_out_mprj[111] la_data_out_mprj[112]
+ la_data_out_mprj[113] la_data_out_mprj[114] la_data_out_mprj[115] la_data_out_mprj[116]
+ la_data_out_mprj[117] la_data_out_mprj[118] la_data_out_mprj[119] la_data_out_mprj[11]
+ la_data_out_mprj[120] la_data_out_mprj[121] la_data_out_mprj[122] la_data_out_mprj[123]
+ la_data_out_mprj[124] la_data_out_mprj[125] la_data_out_mprj[126] la_data_out_mprj[127]
+ la_data_out_mprj[12] la_data_out_mprj[13] la_data_out_mprj[14] la_data_out_mprj[15]
+ la_data_out_mprj[16] la_data_out_mprj[17] la_data_out_mprj[18] la_data_out_mprj[19]
+ la_data_out_mprj[1] la_data_out_mprj[20] la_data_out_mprj[21] la_data_out_mprj[22]
+ la_data_out_mprj[23] la_data_out_mprj[24] la_data_out_mprj[25] la_data_out_mprj[26]
+ la_data_out_mprj[27] la_data_out_mprj[28] la_data_out_mprj[29] la_data_out_mprj[2]
+ la_data_out_mprj[30] la_data_out_mprj[31] la_data_out_mprj[32] la_data_out_mprj[33]
+ la_data_out_mprj[34] la_data_out_mprj[35] la_data_out_mprj[36] la_data_out_mprj[37]
+ la_data_out_mprj[38] la_data_out_mprj[39] la_data_out_mprj[3] la_data_out_mprj[40]
+ la_data_out_mprj[41] la_data_out_mprj[42] la_data_out_mprj[43] la_data_out_mprj[44]
+ la_data_out_mprj[45] la_data_out_mprj[46] la_data_out_mprj[47] la_data_out_mprj[48]
+ la_data_out_mprj[49] la_data_out_mprj[4] la_data_out_mprj[50] la_data_out_mprj[51]
+ la_data_out_mprj[52] la_data_out_mprj[53] la_data_out_mprj[54] la_data_out_mprj[55]
+ la_data_out_mprj[56] la_data_out_mprj[57] la_data_out_mprj[58] la_data_out_mprj[59]
+ la_data_out_mprj[5] la_data_out_mprj[60] la_data_out_mprj[61] la_data_out_mprj[62]
+ la_data_out_mprj[63] la_data_out_mprj[64] la_data_out_mprj[65] la_data_out_mprj[66]
+ la_data_out_mprj[67] la_data_out_mprj[68] la_data_out_mprj[69] la_data_out_mprj[6]
+ la_data_out_mprj[70] la_data_out_mprj[71] la_data_out_mprj[72] la_data_out_mprj[73]
+ la_data_out_mprj[74] la_data_out_mprj[75] la_data_out_mprj[76] la_data_out_mprj[77]
+ la_data_out_mprj[78] la_data_out_mprj[79] la_data_out_mprj[7] la_data_out_mprj[80]
+ la_data_out_mprj[81] la_data_out_mprj[82] la_data_out_mprj[83] la_data_out_mprj[84]
+ la_data_out_mprj[85] la_data_out_mprj[86] la_data_out_mprj[87] la_data_out_mprj[88]
+ la_data_out_mprj[89] la_data_out_mprj[8] la_data_out_mprj[90] la_data_out_mprj[91]
+ la_data_out_mprj[92] la_data_out_mprj[93] la_data_out_mprj[94] la_data_out_mprj[95]
+ la_data_out_mprj[96] la_data_out_mprj[97] la_data_out_mprj[98] la_data_out_mprj[99]
+ la_data_out_mprj[9] la_iena_mprj[0] la_iena_mprj[100] la_iena_mprj[101] la_iena_mprj[102]
+ la_iena_mprj[103] la_iena_mprj[104] la_iena_mprj[105] la_iena_mprj[106] la_iena_mprj[107]
+ la_iena_mprj[108] la_iena_mprj[109] la_iena_mprj[10] la_iena_mprj[110] la_iena_mprj[111]
+ la_iena_mprj[112] la_iena_mprj[113] la_iena_mprj[114] la_iena_mprj[115] la_iena_mprj[116]
+ la_iena_mprj[117] la_iena_mprj[118] la_iena_mprj[119] la_iena_mprj[11] la_iena_mprj[120]
+ la_iena_mprj[121] la_iena_mprj[122] la_iena_mprj[123] la_iena_mprj[124] la_iena_mprj[125]
+ la_iena_mprj[126] la_iena_mprj[127] la_iena_mprj[12] la_iena_mprj[13] la_iena_mprj[14]
+ la_iena_mprj[15] la_iena_mprj[16] la_iena_mprj[17] la_iena_mprj[18] la_iena_mprj[19]
+ la_iena_mprj[1] la_iena_mprj[20] la_iena_mprj[21] la_iena_mprj[22] la_iena_mprj[23]
+ la_iena_mprj[24] la_iena_mprj[25] la_iena_mprj[26] la_iena_mprj[27] la_iena_mprj[28]
+ la_iena_mprj[29] la_iena_mprj[2] la_iena_mprj[30] la_iena_mprj[31] la_iena_mprj[32]
+ la_iena_mprj[33] la_iena_mprj[34] la_iena_mprj[35] la_iena_mprj[36] la_iena_mprj[37]
+ la_iena_mprj[38] la_iena_mprj[39] la_iena_mprj[3] la_iena_mprj[40] la_iena_mprj[41]
+ la_iena_mprj[42] la_iena_mprj[43] la_iena_mprj[44] la_iena_mprj[45] la_iena_mprj[46]
+ la_iena_mprj[47] la_iena_mprj[48] la_iena_mprj[49] la_iena_mprj[4] la_iena_mprj[50]
+ la_iena_mprj[51] la_iena_mprj[52] la_iena_mprj[53] la_iena_mprj[54] la_iena_mprj[55]
+ la_iena_mprj[56] la_iena_mprj[57] la_iena_mprj[58] la_iena_mprj[59] la_iena_mprj[5]
+ la_iena_mprj[60] la_iena_mprj[61] la_iena_mprj[62] la_iena_mprj[63] la_iena_mprj[64]
+ la_iena_mprj[65] la_iena_mprj[66] la_iena_mprj[67] la_iena_mprj[68] la_iena_mprj[69]
+ la_iena_mprj[6] la_iena_mprj[70] la_iena_mprj[71] la_iena_mprj[72] la_iena_mprj[73]
+ la_iena_mprj[74] la_iena_mprj[75] la_iena_mprj[76] la_iena_mprj[77] la_iena_mprj[78]
+ la_iena_mprj[79] la_iena_mprj[7] la_iena_mprj[80] la_iena_mprj[81] la_iena_mprj[82]
+ la_iena_mprj[83] la_iena_mprj[84] la_iena_mprj[85] la_iena_mprj[86] la_iena_mprj[87]
+ la_iena_mprj[88] la_iena_mprj[89] la_iena_mprj[8] la_iena_mprj[90] la_iena_mprj[91]
+ la_iena_mprj[92] la_iena_mprj[93] la_iena_mprj[94] la_iena_mprj[95] la_iena_mprj[96]
+ la_iena_mprj[97] la_iena_mprj[98] la_iena_mprj[99] la_iena_mprj[9] la_oenb_core[0]
+ la_oenb_core[100] la_oenb_core[101] la_oenb_core[102] la_oenb_core[103] la_oenb_core[104]
+ la_oenb_core[105] la_oenb_core[106] la_oenb_core[107] la_oenb_core[108] la_oenb_core[109]
+ la_oenb_core[10] la_oenb_core[110] la_oenb_core[111] la_oenb_core[112] la_oenb_core[113]
+ la_oenb_core[114] la_oenb_core[115] la_oenb_core[116] la_oenb_core[117] la_oenb_core[118]
+ la_oenb_core[119] la_oenb_core[11] la_oenb_core[120] la_oenb_core[121] la_oenb_core[122]
+ la_oenb_core[123] la_oenb_core[124] la_oenb_core[125] la_oenb_core[126] la_oenb_core[127]
+ la_oenb_core[12] la_oenb_core[13] la_oenb_core[14] la_oenb_core[15] la_oenb_core[16]
+ la_oenb_core[17] la_oenb_core[18] la_oenb_core[19] la_oenb_core[1] la_oenb_core[20]
+ la_oenb_core[21] la_oenb_core[22] la_oenb_core[23] la_oenb_core[24] la_oenb_core[25]
+ la_oenb_core[26] la_oenb_core[27] la_oenb_core[28] la_oenb_core[29] la_oenb_core[2]
+ la_oenb_core[30] la_oenb_core[31] la_oenb_core[32] la_oenb_core[33] la_oenb_core[34]
+ la_oenb_core[35] la_oenb_core[36] la_oenb_core[37] la_oenb_core[38] la_oenb_core[39]
+ la_oenb_core[3] la_oenb_core[40] la_oenb_core[41] la_oenb_core[42] la_oenb_core[43]
+ la_oenb_core[44] la_oenb_core[45] la_oenb_core[46] la_oenb_core[47] la_oenb_core[48]
+ la_oenb_core[49] la_oenb_core[4] la_oenb_core[50] la_oenb_core[51] la_oenb_core[52]
+ la_oenb_core[53] la_oenb_core[54] la_oenb_core[55] la_oenb_core[56] la_oenb_core[57]
+ la_oenb_core[58] la_oenb_core[59] la_oenb_core[5] la_oenb_core[60] la_oenb_core[61]
+ la_oenb_core[62] la_oenb_core[63] la_oenb_core[64] la_oenb_core[65] la_oenb_core[66]
+ la_oenb_core[67] la_oenb_core[68] la_oenb_core[69] la_oenb_core[6] la_oenb_core[70]
+ la_oenb_core[71] la_oenb_core[72] la_oenb_core[73] la_oenb_core[74] la_oenb_core[75]
+ la_oenb_core[76] la_oenb_core[77] la_oenb_core[78] la_oenb_core[79] la_oenb_core[7]
+ la_oenb_core[80] la_oenb_core[81] la_oenb_core[82] la_oenb_core[83] la_oenb_core[84]
+ la_oenb_core[85] la_oenb_core[86] la_oenb_core[87] la_oenb_core[88] la_oenb_core[89]
+ la_oenb_core[8] la_oenb_core[90] la_oenb_core[91] la_oenb_core[92] la_oenb_core[93]
+ la_oenb_core[94] la_oenb_core[95] la_oenb_core[96] la_oenb_core[97] la_oenb_core[98]
+ la_oenb_core[99] la_oenb_core[9] la_oenb_mprj[0] la_oenb_mprj[100] la_oenb_mprj[101]
+ la_oenb_mprj[102] la_oenb_mprj[103] la_oenb_mprj[104] la_oenb_mprj[105] la_oenb_mprj[106]
+ la_oenb_mprj[107] la_oenb_mprj[108] la_oenb_mprj[109] la_oenb_mprj[10] la_oenb_mprj[110]
+ la_oenb_mprj[111] la_oenb_mprj[112] la_oenb_mprj[113] la_oenb_mprj[114] la_oenb_mprj[115]
+ la_oenb_mprj[116] la_oenb_mprj[117] la_oenb_mprj[118] la_oenb_mprj[119] la_oenb_mprj[11]
+ la_oenb_mprj[120] la_oenb_mprj[121] la_oenb_mprj[122] la_oenb_mprj[123] la_oenb_mprj[124]
+ la_oenb_mprj[125] la_oenb_mprj[126] la_oenb_mprj[127] la_oenb_mprj[12] la_oenb_mprj[13]
+ la_oenb_mprj[14] la_oenb_mprj[15] la_oenb_mprj[16] la_oenb_mprj[17] la_oenb_mprj[18]
+ la_oenb_mprj[19] la_oenb_mprj[1] la_oenb_mprj[20] la_oenb_mprj[21] la_oenb_mprj[22]
+ la_oenb_mprj[23] la_oenb_mprj[24] la_oenb_mprj[25] la_oenb_mprj[26] la_oenb_mprj[27]
+ la_oenb_mprj[28] la_oenb_mprj[29] la_oenb_mprj[2] la_oenb_mprj[30] la_oenb_mprj[31]
+ la_oenb_mprj[32] la_oenb_mprj[33] la_oenb_mprj[34] la_oenb_mprj[35] la_oenb_mprj[36]
+ la_oenb_mprj[37] la_oenb_mprj[38] la_oenb_mprj[39] la_oenb_mprj[3] la_oenb_mprj[40]
+ la_oenb_mprj[41] la_oenb_mprj[42] la_oenb_mprj[43] la_oenb_mprj[44] la_oenb_mprj[45]
+ la_oenb_mprj[46] la_oenb_mprj[47] la_oenb_mprj[48] la_oenb_mprj[49] la_oenb_mprj[4]
+ la_oenb_mprj[50] la_oenb_mprj[51] la_oenb_mprj[52] la_oenb_mprj[53] la_oenb_mprj[54]
+ la_oenb_mprj[55] la_oenb_mprj[56] la_oenb_mprj[57] la_oenb_mprj[58] la_oenb_mprj[59]
+ la_oenb_mprj[5] la_oenb_mprj[60] la_oenb_mprj[61] la_oenb_mprj[62] la_oenb_mprj[63]
+ la_oenb_mprj[64] la_oenb_mprj[65] la_oenb_mprj[66] la_oenb_mprj[67] la_oenb_mprj[68]
+ la_oenb_mprj[69] la_oenb_mprj[6] la_oenb_mprj[70] la_oenb_mprj[71] la_oenb_mprj[72]
+ la_oenb_mprj[73] la_oenb_mprj[74] la_oenb_mprj[75] la_oenb_mprj[76] la_oenb_mprj[77]
+ la_oenb_mprj[78] la_oenb_mprj[79] la_oenb_mprj[7] la_oenb_mprj[80] la_oenb_mprj[81]
+ la_oenb_mprj[82] la_oenb_mprj[83] la_oenb_mprj[84] la_oenb_mprj[85] la_oenb_mprj[86]
+ la_oenb_mprj[87] la_oenb_mprj[88] la_oenb_mprj[89] la_oenb_mprj[8] la_oenb_mprj[90]
+ la_oenb_mprj[91] la_oenb_mprj[92] la_oenb_mprj[93] la_oenb_mprj[94] la_oenb_mprj[95]
+ la_oenb_mprj[96] la_oenb_mprj[97] la_oenb_mprj[98] la_oenb_mprj[99] la_oenb_mprj[9]
+ mprj_ack_i_core mprj_ack_i_user mprj_adr_o_core[0] mprj_adr_o_core[10] mprj_adr_o_core[11]
+ mprj_adr_o_core[12] mprj_adr_o_core[13] mprj_adr_o_core[14] mprj_adr_o_core[15]
+ mprj_adr_o_core[16] mprj_adr_o_core[17] mprj_adr_o_core[18] mprj_adr_o_core[19]
+ mprj_adr_o_core[1] mprj_adr_o_core[20] mprj_adr_o_core[21] mprj_adr_o_core[22] mprj_adr_o_core[23]
+ mprj_adr_o_core[24] mprj_adr_o_core[25] mprj_adr_o_core[26] mprj_adr_o_core[27]
+ mprj_adr_o_core[28] mprj_adr_o_core[29] mprj_adr_o_core[2] mprj_adr_o_core[30] mprj_adr_o_core[31]
+ mprj_adr_o_core[3] mprj_adr_o_core[4] mprj_adr_o_core[5] mprj_adr_o_core[6] mprj_adr_o_core[7]
+ mprj_adr_o_core[8] mprj_adr_o_core[9] mprj_adr_o_user[0] mprj_adr_o_user[10] mprj_adr_o_user[11]
+ mprj_adr_o_user[12] mprj_adr_o_user[13] mprj_adr_o_user[14] mprj_adr_o_user[15]
+ mprj_adr_o_user[16] mprj_adr_o_user[17] mprj_adr_o_user[18] mprj_adr_o_user[19]
+ mprj_adr_o_user[1] mprj_adr_o_user[20] mprj_adr_o_user[21] mprj_adr_o_user[22] mprj_adr_o_user[23]
+ mprj_adr_o_user[24] mprj_adr_o_user[25] mprj_adr_o_user[26] mprj_adr_o_user[27]
+ mprj_adr_o_user[28] mprj_adr_o_user[29] mprj_adr_o_user[2] mprj_adr_o_user[30] mprj_adr_o_user[31]
+ mprj_adr_o_user[3] mprj_adr_o_user[4] mprj_adr_o_user[5] mprj_adr_o_user[6] mprj_adr_o_user[7]
+ mprj_adr_o_user[8] mprj_adr_o_user[9] mprj_cyc_o_core mprj_cyc_o_user mprj_dat_i_core[0]
+ mprj_dat_i_core[10] mprj_dat_i_core[11] mprj_dat_i_core[12] mprj_dat_i_core[13]
+ mprj_dat_i_core[14] mprj_dat_i_core[15] mprj_dat_i_core[16] mprj_dat_i_core[17]
+ mprj_dat_i_core[18] mprj_dat_i_core[19] mprj_dat_i_core[1] mprj_dat_i_core[20] mprj_dat_i_core[21]
+ mprj_dat_i_core[22] mprj_dat_i_core[23] mprj_dat_i_core[24] mprj_dat_i_core[25]
+ mprj_dat_i_core[26] mprj_dat_i_core[27] mprj_dat_i_core[28] mprj_dat_i_core[29]
+ mprj_dat_i_core[2] mprj_dat_i_core[30] mprj_dat_i_core[31] mprj_dat_i_core[3] mprj_dat_i_core[4]
+ mprj_dat_i_core[5] mprj_dat_i_core[6] mprj_dat_i_core[7] mprj_dat_i_core[8] mprj_dat_i_core[9]
+ mprj_dat_i_user[0] mprj_dat_i_user[10] mprj_dat_i_user[11] mprj_dat_i_user[12] mprj_dat_i_user[13]
+ mprj_dat_i_user[14] mprj_dat_i_user[15] mprj_dat_i_user[16] mprj_dat_i_user[17]
+ mprj_dat_i_user[18] mprj_dat_i_user[19] mprj_dat_i_user[1] mprj_dat_i_user[20] mprj_dat_i_user[21]
+ mprj_dat_i_user[22] mprj_dat_i_user[23] mprj_dat_i_user[24] mprj_dat_i_user[25]
+ mprj_dat_i_user[26] mprj_dat_i_user[27] mprj_dat_i_user[28] mprj_dat_i_user[29]
+ mprj_dat_i_user[2] mprj_dat_i_user[30] mprj_dat_i_user[31] mprj_dat_i_user[3] mprj_dat_i_user[4]
+ mprj_dat_i_user[5] mprj_dat_i_user[6] mprj_dat_i_user[7] mprj_dat_i_user[8] mprj_dat_i_user[9]
+ mprj_dat_o_core[0] mprj_dat_o_core[10] mprj_dat_o_core[11] mprj_dat_o_core[12] mprj_dat_o_core[13]
+ mprj_dat_o_core[14] mprj_dat_o_core[15] mprj_dat_o_core[16] mprj_dat_o_core[17]
+ mprj_dat_o_core[18] mprj_dat_o_core[19] mprj_dat_o_core[1] mprj_dat_o_core[20] mprj_dat_o_core[21]
+ mprj_dat_o_core[22] mprj_dat_o_core[23] mprj_dat_o_core[24] mprj_dat_o_core[25]
+ mprj_dat_o_core[26] mprj_dat_o_core[27] mprj_dat_o_core[28] mprj_dat_o_core[29]
+ mprj_dat_o_core[2] mprj_dat_o_core[30] mprj_dat_o_core[31] mprj_dat_o_core[3] mprj_dat_o_core[4]
+ mprj_dat_o_core[5] mprj_dat_o_core[6] mprj_dat_o_core[7] mprj_dat_o_core[8] mprj_dat_o_core[9]
+ mprj_dat_o_user[0] mprj_dat_o_user[10] mprj_dat_o_user[11] mprj_dat_o_user[12] mprj_dat_o_user[13]
+ mprj_dat_o_user[14] mprj_dat_o_user[15] mprj_dat_o_user[16] mprj_dat_o_user[17]
+ mprj_dat_o_user[18] mprj_dat_o_user[19] mprj_dat_o_user[1] mprj_dat_o_user[20] mprj_dat_o_user[21]
+ mprj_dat_o_user[22] mprj_dat_o_user[23] mprj_dat_o_user[24] mprj_dat_o_user[25]
+ mprj_dat_o_user[26] mprj_dat_o_user[27] mprj_dat_o_user[28] mprj_dat_o_user[29]
+ mprj_dat_o_user[2] mprj_dat_o_user[30] mprj_dat_o_user[31] mprj_dat_o_user[3] mprj_dat_o_user[4]
+ mprj_dat_o_user[5] mprj_dat_o_user[6] mprj_dat_o_user[7] mprj_dat_o_user[8] mprj_dat_o_user[9]
+ mprj_iena_wb mprj_sel_o_core[0] mprj_sel_o_core[1] mprj_sel_o_core[2] mprj_sel_o_core[3]
+ mprj_sel_o_user[0] mprj_sel_o_user[1] mprj_sel_o_user[2] mprj_sel_o_user[3] mprj_stb_o_core
+ mprj_stb_o_user mprj_we_o_core mprj_we_o_user user1_vcc_powergood user1_vdd_powergood
+ user2_vcc_powergood user2_vdd_powergood user_clock user_clock2 user_irq[0] user_irq[1]
+ user_irq[2] user_irq_core[0] user_irq_core[1] user_irq_core[2] user_irq_ena[0] user_irq_ena[1]
+ user_irq_ena[2] user_reset vccd1 vccd2 vdda1 vdda2 vssd dw_201986_9164# dw_194404_9184#
+ vssa2 vssd2 vssa1 dw_1776_7190# dw_71130_9070# vccd vssd1
XFILLER_45_1385 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_973 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_921 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1145 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_461 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1719 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_965 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_29 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1189 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1009 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2057 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[34\]_A input59/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_527 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1105 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_516 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_ena_buf\[72\] input357/X mprj_logic_high_inst/HI[402] vssd vccd user_to_mprj_in_gates\[72\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_8_1644 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input127_A la_data_out_core[96] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_18_439 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_41 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_501_ _501_/A vssd vccd _501_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
Xla_buf_enable\[50\] _642_/A la_buf_enable\[50\]/B vssd vccd la_buf\[50\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_2_1276 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1808 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_432_ _432_/A vssd vccd _432_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_26_85 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input496_A la_oenb_mprj[82] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_363_ _363_/A vssd vccd _363_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_35_1565 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xla_buf\[36\] _500_/Y la_buf\[36\]/TE vssd vccd la_data_in_core[36] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input92_A la_data_out_core[64] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_2288 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_497 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_851 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[108\] input269/X mprj_logic_high_inst/HI[438] vssd vccd
+ user_to_mprj_in_gates\[108\]/B vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_10_895 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_gates\[8\] input580/X user_wb_ack_gate/B vssd vccd user_wb_dat_gates\[8\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_in_gates\[25\]_A input49/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_1325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1419 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1369 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_593 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_715 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_597 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2008 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_910 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_217 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1329 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[25\] input49/X user_to_mprj_in_gates\[25\]/B vssd vccd user_to_mprj_in_gates\[25\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_53_1665 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_1763 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_1627 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1941 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[100\]_A input5/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[16\]_A input39/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1985 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_1425 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1931 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1469 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1817 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2275 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1563 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1749 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[76\] _339_/Y mprj_logic_high_inst/HI[278] vssd vccd la_oenb_core[76]
+ vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[98\] _361_/A la_buf_enable\[98\]/B vssd vccd la_buf\[98\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
Xmprj_dat_buf\[24\] _456_/Y mprj_dat_buf\[24\]/TE vssd vccd mprj_dat_o_user[24] vssd
+ vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input244_A la_data_out_mprj[86] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_2039 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_501 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_51 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input411_A la_oenb_mprj[120] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[104\]_TE mprj_logic_high_inst/HI[306] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_545 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input509_A la_oenb_mprj[94] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_1062 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_589 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1649 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_415_ _415_/A vssd vccd _415_/Y vssd vccd sky130_fd_sc_hd__inv_12
XFILLER_35_2041 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2085 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_346_ _346_/A vssd vccd _346_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_35_2063 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_173 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1745 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1789 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2001 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output728_A output728/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output630_A output630/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_1177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_2045 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1399 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[122\]_A input285/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_2174 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_1560 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_445 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[4\] _596_/A la_buf_enable\[4\]/B vssd vccd la_buf\[4\]/TE vssd vccd
+ sky130_fd_sc_hd__and2b_1
XFILLER_31_1771 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1793 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1211 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1807 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[127\]_TE mprj_logic_high_inst/HI[329] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_1553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_501 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_2050 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_707 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_589 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[35\] input316/X mprj_logic_high_inst/HI[365] vssd vccd user_to_mprj_in_gates\[35\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_in_ena_buf\[113\]_A input275/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_209 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_405 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xla_buf_enable\[13\] _605_/A la_buf_enable\[13\]/B vssd vccd la_buf\[13\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_23_86 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input194_A la_data_out_mprj[40] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_1833 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input361_A la_iena_mprj[76] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_2007 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input459_A la_oenb_mprj[49] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[41\]_TE la_buf\[41\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_2321 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1929 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input55_A la_data_out_core[30] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[26\]_TE mprj_logic_high_inst/HI[228] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input626_A user_irq_ena[2] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[92\]_A_N _355_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_501 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[104\]_A input265/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_537 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[30\]_A_N _622_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_2325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output678_A output678/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_1891 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_1711 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_798 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_1755 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_329_ _329_/A vssd vccd _329_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_11_1619 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_1799 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[45\]_A_N _637_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[92\] input123/X user_to_mprj_in_gates\[92\]/B vssd vccd user_to_mprj_in_gates\[92\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_48_1597 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1575 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1035 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1901 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1895 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1945 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1759 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1989 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_898 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_356 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1991 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[64\]_TE la_buf\[64\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_2029 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[49\]_TE mprj_logic_high_inst/HI[251] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_1709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput515 la_oenb_mprj[9] vssd vccd _601_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput537 mprj_adr_o_core[28] vssd vccd _428_/A vssd vccd sky130_fd_sc_hd__buf_2
Xinput526 mprj_adr_o_core[18] vssd vccd _418_/A vssd vccd sky130_fd_sc_hd__buf_2
Xinput504 la_oenb_mprj[8] vssd vccd _600_/A vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_29_821 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[109\] _372_/Y mprj_logic_high_inst/HI[311] vssd vccd la_oenb_core[109]
+ vssd vccd sky130_fd_sc_hd__einvp_8
Xinput548 mprj_adr_o_core[9] vssd vccd _409_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput559 mprj_dat_i_user[18] vssd vccd input559/X vssd vccd sky130_fd_sc_hd__buf_12
XANTENNA_user_to_mprj_in_ena_buf\[93\]_A input380/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_515 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[39\] _631_/Y mprj_logic_high_inst/HI[241] vssd vccd la_oenb_core[39]
+ vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_28_353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_397 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1733 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_559 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input207_A la_data_out_mprj[52] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_41 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_85 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1799 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input576_A mprj_dat_i_user[4] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_1939 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_246 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1663 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[13\]_TE mprj_dat_buf\[13\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_441 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__402__A _402_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1895 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_629 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2173 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[84\]_A input370/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2209 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_813 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_662 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[62\] user_to_mprj_in_gates\[62\]/Y vssd vccd output713/A
+ vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_34_345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_805 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[87\]_TE la_buf\[87\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_1421 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_wb_dat_gates\[20\] input562/X user_wb_ack_gate/B vssd vccd user_wb_dat_gates\[20\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_4
XFILLER_50_1465 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1427 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[75\]_A input360/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_621 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_120 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1029 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_304 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_827 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1917 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_540 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1983 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_65 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xinput312 la_iena_mprj[31] vssd vccd input312/X vssd vccd sky130_fd_sc_hd__dlymetal6s2s_1
Xla_buf_enable\[80\] _343_/A la_buf_enable\[80\]/B vssd vccd la_buf\[80\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XANTENNA_input157_A la_data_out_mprj[122] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput301 la_iena_mprj[21] vssd vccd input301/X vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_49_949 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xinput323 la_iena_mprj[41] vssd vccd input323/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput334 la_iena_mprj[51] vssd vccd input334/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput345 la_iena_mprj[61] vssd vccd input345/X vssd vccd sky130_fd_sc_hd__clkbuf_1
XANTENNA_input324_A la_iena_mprj[42] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[66\]_A input350/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput356 la_iena_mprj[71] vssd vccd input356/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput367 la_iena_mprj[81] vssd vccd input367/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput378 la_iena_mprj[91] vssd vccd input378/X vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_29_673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input18_A la_data_out_core[112] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput389 la_oenb_mprj[100] vssd vccd _363_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_40_1645 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1689 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_51 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_594_ _594_/A vssd vccd _594_/Y vssd vccd sky130_fd_sc_hd__clkinv_4
Xla_buf\[66\] _530_/Y la_buf\[66\]/TE vssd vccd la_data_in_core[66] vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_38_1541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_849 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1563 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_893 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1703 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_595 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1747 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1785 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1173 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_599 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[122\] _586_/Y la_buf\[122\]/TE vssd vccd la_data_in_core[122] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_gates\[70\]_B user_to_mprj_in_gates\[70\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1578 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output710_A output710/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[57\]_A input340/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[55\] input82/X user_to_mprj_in_gates\[55\]/B vssd vccd user_to_mprj_in_gates\[55\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_23_1876 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_993 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2017 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1887 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1694 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_613 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_657 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1814 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1273 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[61\]_B user_to_mprj_in_gates\[61\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_28_1721 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1815 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1776 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_1607 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1859 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_908 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[48\]_A input330/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_919 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1447 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1861 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_495 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2150 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_319 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_189 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input274_A la_iena_mprj[112] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[52\]_B user_to_mprj_in_gates\[52\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_11_1791 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_753 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1821 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input441_A la_oenb_mprj[32] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input539_A mprj_adr_o_core[2] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_764 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1303 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput120 la_data_out_core[8] vssd vccd input120/X vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_1_797 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xinput153 la_data_out_mprj[119] vssd vccd _583_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput131 la_data_out_core[9] vssd vccd input131/X vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA_user_to_mprj_in_ena_buf\[39\]_A input320/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput142 la_data_out_mprj[109] vssd vccd _573_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_48_245 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xinput186 la_data_out_mprj[33] vssd vccd _497_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput175 la_data_out_mprj[23] vssd vccd _487_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput164 la_data_out_mprj[13] vssd vccd _477_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_29_481 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1453 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput197 la_data_out_mprj[43] vssd vccd _507_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_17_643 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_646_ _646_/A vssd vccd _646_/Y vssd vccd sky130_fd_sc_hd__inv_2
X_577_ _577_/A vssd vccd _577_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_32_657 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[6\]_A _438_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1257 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_1869 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_1691 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_886 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[25\] user_to_mprj_in_gates\[25\]/Y vssd vccd output672/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_output660_A output660/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output758_A output758/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_1593 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xoutput627 output627/A vssd vccd la_data_in_mprj[0] vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA_user_to_mprj_in_gates\[43\]_B user_to_mprj_in_gates\[43\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xoutput638 output638/A vssd vccd la_data_in_mprj[10] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput649 output649/A vssd vccd la_data_in_mprj[11] vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_45_2065 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[112\]_TE la_buf\[112\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1397 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[27\]_TE mprj_adr_buf\[27\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_933 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_473 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_421 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_19 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_977 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2069 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[34\]_B user_to_mprj_in_gates\[34\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[95\]_A user_to_mprj_in_gates\[95\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_28_2241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1117 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2070 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[65\] input349/X mprj_logic_high_inst/HI[395] vssd vccd user_to_mprj_in_gates\[65\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA__500__A _500_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_749 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_500_ _500_/A vssd vccd _500_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_45_237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_53 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[21\] _613_/Y mprj_logic_high_inst/HI[223] vssd vccd la_oenb_core[21]
+ vssd vccd sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[3\] _595_/Y mprj_logic_high_inst/HI[205] vssd vccd la_oenb_core[3]
+ vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[43\] _635_/A la_buf_enable\[43\]/B vssd vccd la_buf\[43\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
X_431_ _431_/A vssd vccd _431_/Y vssd vccd sky130_fd_sc_hd__inv_8
XFILLER_26_97 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_362_ _362_/A vssd vccd _362_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_42_41 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input489_A la_oenb_mprj[76] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input391_A la_oenb_mprj[102] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_863 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input85_A la_data_out_core[58] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_1820 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_1831 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[29\] _493_/Y la_buf\[29\]/TE vssd vccd la_data_in_core[29] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf\[122\]_A _586_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[86\]_A user_to_mprj_in_gates\[86\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[25\]_B user_to_mprj_in_gates\[25\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_29_1337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_68 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__410__A _410_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_1971 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_204 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1929 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_1261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_922 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_629_ _629_/A vssd vccd _629_/Y vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_user_to_mprj_in_buffers\[10\]_A user_to_mprj_in_gates\[10\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_32_421 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_410 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_605 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[18\] input41/X user_to_mprj_in_gates\[18\]/B vssd vccd user_to_mprj_in_gates\[18\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XANTENNA_user_to_mprj_in_buffers\[124\]_A user_to_mprj_in_gates\[124\]/Y vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[113\]_A _577_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1953 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_buffers\[77\]_A user_to_mprj_in_gates\[77\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[16\]_B user_to_mprj_in_gates\[16\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_buffers\[28\] user_wb_dat_gates\[28\]/Y vssd vccd output776/A vssd vccd
+ sky130_fd_sc_hd__clkinv_8
XANTENNA_user_to_mprj_in_gates\[100\]_B user_to_mprj_in_gates\[100\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[50\]_A _514_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_1437 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[82\]_TE mprj_logic_high_inst/HI[284] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_1943 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1987 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1829 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2287 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_741 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_785 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[115\]_A user_to_mprj_in_gates\[115\]/Y vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[104\]_A _568_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1441 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[68\]_A user_to_mprj_in_gates\[68\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[41\]_A _505_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_314 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_1993 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_oen_buffers\[69\] _332_/Y mprj_logic_high_inst/HI[271] vssd vccd la_oenb_core[69]
+ vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_4_1317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[17\] _449_/Y mprj_dat_buf\[17\]/TE vssd vccd mprj_dat_o_user[17] vssd
+ vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input237_A la_data_out_mprj[7] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_1497 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_557 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input404_A la_oenb_mprj[114] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_1074 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_218 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_414_ _414_/A vssd vccd _414_/Y vssd vccd sky130_fd_sc_hd__clkinv_8
XFILLER_41_273 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_936 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_ena_buf\[120\] input283/X mprj_logic_high_inst/HI[450] vssd vccd
+ user_to_mprj_in_gates\[120\]/B vssd vccd sky130_fd_sc_hd__and2_1
X_345_ _345_/A vssd vccd _345_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_user_to_mprj_in_buffers\[106\]_A user_to_mprj_in_gates\[106\]/Y vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_2097 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__405__A _405_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[59\]_A user_to_mprj_in_gates\[59\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_52_7 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[32\]_A _496_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[12\] _412_/Y mprj_adr_buf\[12\]/TE vssd vccd mprj_adr_o_user[12] vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_42_2013 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1145 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1757 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_buffers\[126\] user_to_mprj_in_gates\[126\]/Y vssd vccd output656/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_la_buf_enable\[50\]_B la_buf_enable\[50\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_1239 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_892 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[92\] user_to_mprj_in_gates\[92\]/Y vssd vccd output746/A
+ vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_42_2057 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1908 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1919 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_557 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[99\]_A _563_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[122\]_B mprj_logic_high_inst/HI[452] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_buffers\[2\] user_wb_dat_gates\[2\]/Y vssd vccd output778/A vssd vccd
+ sky130_fd_sc_hd__clkinv_8
XFILLER_33_741 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_785 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1572 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[23\]_A _487_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1783 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_1223 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[41\]_B la_buf_enable\[41\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_1289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_1565 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2073 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[113\]_B mprj_logic_high_inst/HI[443] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_16_719 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_ena_buf\[28\] input308/X mprj_logic_high_inst/HI[358] vssd vccd user_to_mprj_in_gates\[28\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_23_273 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_907 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_98 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input187_A la_data_out_mprj[34] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[14\]_A _478_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_2019 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input354_A la_iena_mprj[6] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[32\]_B la_buf_enable\[32\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_2333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input48_A la_data_out_core[24] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[1\]_A input299/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input521_A mprj_adr_o_core[13] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input619_A mprj_stb_o_core vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[1\] input299/X mprj_logic_high_inst/HI[331] vssd vccd user_to_mprj_in_gates\[1\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
Xla_buf\[96\] _560_/Y la_buf\[96\]/TE vssd vccd la_data_in_core[96] vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[111\] _374_/A la_buf_enable\[111\]/B vssd vccd la_buf\[111\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_8_1272 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_321 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[104\]_B mprj_logic_high_inst/HI[434] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_34_549 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1425 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[99\]_B la_buf_enable\[99\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_2337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1171 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_991 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1767 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output740_A output740/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1521 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1003 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[85\] input115/X user_to_mprj_in_gates\[85\]/B vssd vccd user_to_mprj_in_gates\[85\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XANTENNA_la_buf_enable\[23\]_B la_buf_enable\[23\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_1047 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_1587 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1913 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1957 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_321 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[92\]_A _355_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_2328 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[14\]_B la_buf_enable\[14\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput516 mprj_ack_i_user vssd vccd input516/X vssd vccd sky130_fd_sc_hd__buf_8
Xinput505 la_oenb_mprj[90] vssd vccd _353_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput527 mprj_adr_o_core[19] vssd vccd _419_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_5_2146 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput538 mprj_adr_o_core[29] vssd vccd _429_/A vssd vccd sky130_fd_sc_hd__buf_2
Xinput549 mprj_cyc_o_core vssd vccd _393_/A vssd vccd sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_user_to_mprj_in_ena_buf\[93\]_B mprj_logic_high_inst/HI[423] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_29_833 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_527 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_869 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input102_A la_data_out_core[73] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_1745 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_53 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1609 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2045 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[83\]_A _346_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_41 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input471_A la_oenb_mprj[5] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_1907 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_85 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[7\] _471_/Y la_buf\[7\]/TE vssd vccd la_data_in_core[7] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input569_A mprj_dat_i_user[27] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf\[11\] _475_/Y la_buf\[11\]/TE vssd vccd la_data_in_core[11] vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_10_1675 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_1705 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_497 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1749 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_107 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_2185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_118 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[4\] _404_/Y mprj_adr_buf\[4\]/TE vssd vccd mprj_adr_o_user[4] vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_19_321 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1091 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[84\]_B mprj_logic_high_inst/HI[414] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_19_365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_825 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1854 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_685 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[55\] user_to_mprj_in_gates\[55\]/Y vssd vccd output705/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_34_357 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output690_A output690/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output788_A output788/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_1233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_2101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1266 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[117\]_TE mprj_logic_high_inst/HI[319] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_1299 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[74\]_A _337_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_gates\[13\] input554/X user_wb_ack_gate/B vssd vccd user_wb_dat_gates\[13\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_4
XFILLER_11_1439 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_781 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_1373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_buffers\[10\] user_wb_dat_gates\[10\]/Y vssd vccd output757/A vssd vccd
+ sky130_fd_sc_hd__clkinv_8
XFILLER_26_2350 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[1\]_A input561/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_1721 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1671 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1765 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[111\] input17/X user_to_mprj_in_gates\[111\]/B vssd vccd user_to_mprj_in_gates\[111\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XANTENNA_user_to_mprj_in_ena_buf\[75\]_B mprj_logic_high_inst/HI[405] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_53_633 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_132 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_677 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[1\]_A input43/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[31\]_TE la_buf\[31\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_1929 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[91\]_A_N _354_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[16\]_TE mprj_logic_high_inst/HI[218] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[65\]_A _657_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_552 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_ena_buf\[95\] input382/X mprj_logic_high_inst/HI[425] vssd vccd user_to_mprj_in_gates\[95\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA__503__A _503_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_77 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2103 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2208 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[121\] _384_/Y mprj_logic_high_inst/HI[323] vssd vccd la_oenb_core[121]
+ vssd vccd sky130_fd_sc_hd__einvp_8
Xmprj_sel_buf\[2\] _398_/Y mprj_sel_buf\[2\]/TE vssd vccd mprj_sel_o_user[2] vssd
+ vccd sky130_fd_sc_hd__einvp_8
Xinput302 la_iena_mprj[22] vssd vccd input302/X vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_40_2325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput313 la_iena_mprj[32] vssd vccd input313/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput324 la_iena_mprj[42] vssd vccd input324/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput335 la_iena_mprj[52] vssd vccd input335/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xuser_to_mprj_oen_buffers\[51\] _643_/Y mprj_logic_high_inst/HI[253] vssd vccd la_oenb_core[51]
+ vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[73\] _336_/A la_buf_enable\[73\]/B vssd vccd la_buf\[73\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XANTENNA_user_to_mprj_in_ena_buf\[66\]_B mprj_logic_high_inst/HI[396] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xinput346 la_iena_mprj[62] vssd vccd input346/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput357 la_iena_mprj[72] vssd vccd input357/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput368 la_iena_mprj[82] vssd vccd input368/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput379 la_iena_mprj[92] vssd vccd input379/X vssd vccd sky130_fd_sc_hd__clkbuf_1
XANTENNA_input317_A la_iena_mprj[36] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_685 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[44\]_A_N _636_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_335 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_593_ _593_/A vssd vccd _593_/Y vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_38_1520 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[59\] _523_/Y la_buf\[59\]/TE vssd vccd la_data_in_core[59] vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_31_305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[59\]_A_N _651_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[56\]_A _648_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_1851 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1715 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1759 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xla_buf\[115\] _579_/Y la_buf\[115\]/TE vssd vccd la_data_in_core[115] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA__413__A _413_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1546 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_405 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1905 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output703_A output703/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[57\]_B mprj_logic_high_inst/HI[387] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_48_961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[54\]_TE la_buf\[54\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_1899 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2029 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1651 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[48\] input74/X user_to_mprj_in_gates\[48\]/B vssd vccd user_to_mprj_in_gates\[48\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XANTENNA_user_to_mprj_oen_buffers\[39\]_TE mprj_logic_high_inst/HI[241] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_669 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[47\]_A _639_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_1241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1203 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1285 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1733 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_1012 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1827 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1619 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2191 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[48\]_B mprj_logic_high_inst/HI[378] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_2_2127 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_1404 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_600 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1873 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[10\] input271/X mprj_logic_high_inst/HI[340] vssd vccd user_to_mprj_in_gates\[10\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_oen_buffers\[38\]_A _630_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_2162 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1461 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[99\] _362_/Y mprj_logic_high_inst/HI[301] vssd vccd la_oenb_core[99]
+ vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_31_87 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input267_A la_iena_mprj[106] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_1833 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj2_vdd_pwrgood mprj2_vdd_pwrgood/A vssd vccd output791/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_46_1877 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput110 la_data_out_core[80] vssd vccd input110/X vssd vccd sky130_fd_sc_hd__buf_4
XANTENNA_input434_A la_oenb_mprj[26] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[77\]_TE la_buf\[77\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput121 la_data_out_core[90] vssd vccd input121/X vssd vccd sky130_fd_sc_hd__buf_4
Xinput154 la_data_out_mprj[11] vssd vccd _475_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput143 la_data_out_mprj[10] vssd vccd _474_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput132 la_data_out_mprj[0] vssd vccd _464_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
XANTENNA_input30_A la_data_out_core[123] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput187 la_data_out_mprj[34] vssd vccd _498_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput176 la_data_out_mprj[24] vssd vccd _488_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput165 la_data_out_mprj[14] vssd vccd _478_/A vssd vccd sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_input601_A mprj_dat_o_core[27] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[39\]_B mprj_logic_high_inst/HI[369] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_40_1465 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_622 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput198 la_data_out_mprj[44] vssd vccd _508_/A vssd vccd sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_45_953 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_655 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_645_ _645_/A vssd vccd _645_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_17_699 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_576_ _576_/A vssd vccd _576_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_31_113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__408__A _408_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_669 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[29\]_A _621_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_1361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_371 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_898 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[18\] user_to_mprj_in_gates\[18\]/Y vssd vccd output664/A
+ vssd vccd sky130_fd_sc_hd__inv_2
XANTENNA_output653_A output653/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput628 output628/A vssd vccd la_data_in_mprj[100] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput639 output639/A vssd vccd la_data_in_mprj[110] vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_45_1321 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_mprj_adr_buf\[25\]_A _425_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_909 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1713 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1663 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1757 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[26\]_TE mprj_dat_buf\[26\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_433 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_945 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_989 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[5\]_TE mprj_logic_high_inst/HI[207] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_50_477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[2\]_A _594_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1781 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1099 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_1129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[16\]_A _416_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_1679 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2082 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[58\] input341/X mprj_logic_high_inst/HI[388] vssd vccd user_to_mprj_in_gates\[58\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_45_205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_65 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_430_ _430_/A vssd vccd _430_/Y vssd vccd sky130_fd_sc_hd__clkinv_8
Xuser_to_mprj_oen_buffers\[14\] _606_/Y mprj_logic_high_inst/HI[216] vssd vccd la_oenb_core[14]
+ vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[36\] _628_/A la_buf_enable\[36\]/B vssd vccd la_buf\[36\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
X_361_ _361_/A vssd vccd _361_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_39_1681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_53 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input384_A la_iena_mprj[97] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_813 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_1843 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_875 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2017 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1887 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input78_A la_data_out_core[51] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input551_A mprj_dat_i_user[10] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_2217 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1145 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1009 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_216 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1803 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_sel_buf\[0\]_TE mprj_sel_buf\[0\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_1251 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_1273 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1295 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_628_ _628_/A vssd vccd _628_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_33_934 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_433 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_2335 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_559_ _559_/A vssd vccd _559_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_32_499 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output770_A output770/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_1911 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__601__A _601_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_1955 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2211 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1999 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_753 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1821 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_797 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_326 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__511__A _511_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_1487 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1329 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_525 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input132_A la_data_out_mprj[0] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_1031 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1593 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
X_413_ _413_/A vssd vccd _413_/Y vssd vccd sky130_fd_sc_hd__inv_6
XFILLER_35_2010 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_41 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input599_A mprj_dat_o_core[25] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf\[41\] _505_/Y la_buf\[41\]/TE vssd vccd la_data_in_core[41] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf\[102\]_TE la_buf\[102\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_344_ _344_/A vssd vccd _344_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_35_2054 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_ena_buf\[113\] input275/X mprj_logic_high_inst/HI[443] vssd vccd
+ user_to_mprj_in_gates\[113\]/B vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_mprj_adr_buf\[17\]_TE mprj_adr_buf\[17\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_1695 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__421__A _421_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[1\]_TE mprj_adr_buf\[1\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_2025 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[119\] user_to_mprj_in_gates\[119\]/Y vssd vccd output648/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_42_2069 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[29\]_A _461_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[85\] user_to_mprj_in_gates\[85\]/Y vssd vccd output738/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_49_385 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[30\] input55/X user_to_mprj_in_gates\[30\]/B vssd vccd user_to_mprj_in_gates\[30\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_33_753 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_775 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_469 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_mprj_adr_buf\[1\]_A _401_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_1257 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__331__A _331_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_dat_buf\[5\]_TE mprj_dat_buf\[5\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_1763 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1577 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2030 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_buffers\[27\]_A user_wb_dat_gates\[27\]/Y vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XFILLER_25_1599 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_517 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[125\]_TE la_buf\[125\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_ack_gate_A input516/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_447 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_919 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__506__A _506_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_1971 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[81\] _344_/Y mprj_logic_high_inst/HI[283] vssd vccd la_oenb_core[81]
+ vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_3_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_2345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input347_A la_iena_mprj[63] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_41 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[1\]_B mprj_logic_high_inst/HI[331] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_4_1104 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_1666 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_85 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input514_A la_oenb_mprj[99] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_buffers\[18\]_A user_wb_dat_gates\[18\]/Y vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XFILLER_46_333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[89\] _553_/Y la_buf\[89\]/TE vssd vccd la_data_in_core[89] vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[104\] _367_/A la_buf_enable\[104\]/B vssd vccd la_buf\[104\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_46_377 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1437 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[72\]_TE mprj_logic_high_inst/HI[274] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_2349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__416__A _416_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_1871 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1533 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output733_A output733/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1015 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[78\] input107/X user_to_mprj_in_gates\[78\]/B vssd vccd user_to_mprj_in_gates\[78\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_42_1121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1925 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1969 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[122\]_B la_buf_enable\[122\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_0_2269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_517 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[91\]_A input122/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj2_pwrgood_A mprj2_pwrgood/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput528 mprj_adr_o_core[1] vssd vccd _401_/A vssd vccd sky130_fd_sc_hd__buf_2
Xinput517 mprj_adr_o_core[0] vssd vccd _400_/A vssd vccd sky130_fd_sc_hd__buf_12
Xinput506 la_oenb_mprj[91] vssd vccd _354_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_40_1806 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2158 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput539 mprj_adr_o_core[2] vssd vccd _402_/A vssd vccd sky130_fd_sc_hd__buf_12
XFILLER_5_1413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_845 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1435 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[40\] input322/X mprj_logic_high_inst/HI[370] vssd vccd user_to_mprj_in_gates\[40\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_la_buf_enable\[113\]_B la_buf_enable\[113\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_539 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[95\]_TE mprj_logic_high_inst/HI[297] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_1757 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_509 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_2193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_65 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2057 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_727 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input297_A la_iena_mprj[18] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_buffers\[4\]_A user_wb_dat_gates\[4\]/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_53 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[82\]_A input112/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_97 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input464_A la_oenb_mprj[53] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input60_A la_data_out_core[35] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1717 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1811 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[7\]_A _471_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[104\]_B la_buf_enable\[104\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_697 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_377 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_572 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[48\] user_to_mprj_in_gates\[48\]/Y vssd vccd output697/A
+ vssd vccd sky130_fd_sc_hd__inv_2
XANTENNA_output683_A output683/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_2113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_2157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[73\]_A input102/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1341 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1385 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1227 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[1\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_1733 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1683 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1777 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2191 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[104\] input9/X user_to_mprj_in_gates\[104\]/B vssd vccd user_to_mprj_in_gates\[104\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_34_881 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[1\]_B user_to_mprj_in_gates\[1\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_40_328 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[64\]_A input92/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_2148 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[88\] input374/X mprj_logic_high_inst/HI[418] vssd vccd user_to_mprj_in_gates\[88\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
Xuser_to_mprj_oen_buffers\[114\] _377_/Y mprj_logic_high_inst/HI[316] vssd vccd la_oenb_core[114]
+ vssd vccd sky130_fd_sc_hd__einvp_8
Xinput303 la_iena_mprj[23] vssd vccd input303/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput325 la_iena_mprj[43] vssd vccd input325/X vssd vccd sky130_fd_sc_hd__dlymetal6s2s_1
Xinput314 la_iena_mprj[33] vssd vccd input314/X vssd vccd sky130_fd_sc_hd__dlymetal6s2s_1
Xinput336 la_iena_mprj[53] vssd vccd input336/X vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_40_2337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput347 la_iena_mprj[63] vssd vccd input347/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput358 la_iena_mprj[73] vssd vccd input358/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput369 la_iena_mprj[83] vssd vccd input369/X vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_1_1107 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_oen_buffers\[44\] _636_/Y mprj_logic_high_inst/HI[246] vssd vccd la_oenb_core[44]
+ vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[66\] _329_/A la_buf_enable\[66\]/B vssd vccd la_buf\[66\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_16_303 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_irq_buffers\[2\] user_irq_gates\[2\]/Y vssd vccd output794/A vssd vccd sky130_fd_sc_hd__clkinv_4
X_592_ _592_/A vssd vccd _592_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_input212_A la_data_out_mprj[57] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_697 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_667 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_347 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1532 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_2119 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_97 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input581_A mprj_dat_i_user[9] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_1727 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[55\]_A input82/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_1142 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1661 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[108\] _572_/Y la_buf\[108\]/TE vssd vccd la_data_in_core[108] vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_45_1569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1558 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[101\] user_to_mprj_in_gates\[101\]/Y vssd vccd output629/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_19_141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1917 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_973 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_461 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1307 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_111 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[5\]_A user_to_mprj_in_gates\[5\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_50_637 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_1253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[46\]_A input72/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__604__A _604_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_1297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1215 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1259 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1024 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2231 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[0\] _432_/Y mprj_dat_buf\[0\]/TE vssd vccd mprj_dat_o_user[0] vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_8_1839 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1057 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_612 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_645 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1841 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1705 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1885 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2174 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1473 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[37\]_A input62/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[121\]_A input28/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__514__A _514_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_99 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_711 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1509 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_1801 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1845 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2017 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input162_A la_data_out_mprj[127] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_1709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput111 la_data_out_core[81] vssd vccd input111/X vssd vccd sky130_fd_sc_hd__buf_4
Xinput100 la_data_out_core[71] vssd vccd input100/X vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_44_2281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput122 la_data_out_core[91] vssd vccd input122/X vssd vccd sky130_fd_sc_hd__buf_4
XANTENNA_input427_A la_oenb_mprj[1] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[107\]_TE mprj_logic_high_inst/HI[309] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
Xinput133 la_data_out_mprj[100] vssd vccd _564_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput144 la_data_out_mprj[110] vssd vccd _574_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput177 la_data_out_mprj[25] vssd vccd _489_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput166 la_data_out_mprj[15] vssd vccd _479_/A vssd vccd sky130_fd_sc_hd__dlymetal6s2s_1
Xinput155 la_data_out_mprj[120] vssd vccd _584_/A vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA_input23_A la_data_out_core[117] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_921 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_461 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput199 la_data_out_mprj[45] vssd vccd _509_/A vssd vccd sky130_fd_sc_hd__dlymetal6s2s_1
Xinput188 la_data_out_mprj[35] vssd vccd _499_/A vssd vccd sky130_fd_sc_hd__dlymetal6s2s_1
X_644_ _644_/A vssd vccd _644_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_45_965 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[71\] _535_/Y la_buf\[71\]/TE vssd vccd la_data_in_core[71] vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_40_1477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_667 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_575_ _575_/A vssd vccd _575_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_31_125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1827 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_811 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_800 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_2241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__424__A _424_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[28\]_A input52/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_383 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[112\]_A input18/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_1579 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xoutput629 output629/A vssd vccd la_data_in_mprj[101] vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA_output646_A output646/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_1281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[21\]_TE la_buf\[21\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_1861 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[60\] input88/X user_to_mprj_in_gates\[60\]/B vssd vccd user_to_mprj_in_gates\[60\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XANTENNA_la_buf_enable\[90\]_A_N _353_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_247 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1725 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_1675 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_781 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1769 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_445 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_489 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[19\]_A input42/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1793 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[103\]_A input8/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__334__A _334_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_1061 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[43\]_A_N _635_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_2265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2107 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1603 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1597 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[58\]_A_N _650_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_2094 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1775 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_217 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_291 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_902 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__509__A _509_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_615 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_360_ _360_/A vssd vccd _360_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_39_1693 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[29\] _621_/A la_buf_enable\[29\]/B vssd vccd la_buf\[29\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_42_65 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1855 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_887 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_869 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input377_A la_iena_mprj[90] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[44\]_TE la_buf\[44\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_2321 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_2029 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1899 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input544_A mprj_adr_o_core[5] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[29\]_TE mprj_logic_high_inst/HI[231] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_1653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2229 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_707 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1815 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_228 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_431 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1859 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_627_ _627_/A vssd vccd _627_/Y vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA__419__A _419_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_1791 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_475 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_558_ _558_/A vssd vccd _558_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_33_946 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_445 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_629 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[30\] user_to_mprj_in_gates\[30\]/Y vssd vccd output678/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
X_489_ _489_/A vssd vccd _489_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_31_1900 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output763_A output763/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_1392 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1381 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[1\]_B la_buf_enable\[1\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_1923 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1967 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2223 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[125\]_A input288/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_209 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__329__A _329_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_721 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_765 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1833 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2280 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1877 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[67\]_TE la_buf\[67\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2073 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[70\] input355/X mprj_logic_high_inst/HI[400] vssd vccd user_to_mprj_in_gates\[70\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_47_1973 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1411 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1455 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[116\]_A input278/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_1561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input125_A la_data_out_core[94] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_1054 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1087 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_412_ _412_/A vssd vccd _412_/Y vssd vccd sky130_fd_sc_hd__inv_12
X_343_ _343_/A vssd vccd _343_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_input494_A la_oenb_mprj[80] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_75 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xla_buf\[34\] _498_/Y la_buf\[34\]/TE vssd vccd la_data_in_core[34] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input90_A la_data_out_core[62] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_1630 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[106\] input267/X mprj_logic_high_inst/HI[436] vssd vccd
+ user_to_mprj_in_gates\[106\]/B vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_13_1663 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_gates\[6\] input578/X user_wb_ack_gate/B vssd vccd user_wb_dat_gates\[6\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_4
XANTENNA_mprj_dat_buf\[16\]_TE mprj_dat_buf\[16\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_861 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[107\]_A input268/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[78\] user_to_mprj_in_gates\[78\]/Y vssd vccd output730/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_40_1093 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_721 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_765 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[23\] input47/X user_to_mprj_in_gates\[23\]/B vssd vccd user_to_mprj_in_gates\[23\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_9_471 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__612__A _612_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_1720 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1775 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2042 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_1589 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1330 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_529 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1385 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_ack_gate_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_573 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_459 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_1803 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_1847 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__522__A _522_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1273 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[74\] _337_/Y mprj_logic_high_inst/HI[276] vssd vccd la_oenb_core[74]
+ vssd vccd sky130_fd_sc_hd__einvp_8
Xoutput790 output790/A vssd vccd user2_vcc_powergood vssd vccd sky130_fd_sc_hd__buf_2
Xla_buf_enable\[96\] _359_/A la_buf_enable\[96\]/B vssd vccd la_buf\[96\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
Xmprj_dat_buf\[22\] _454_/Y mprj_dat_buf\[22\]/TE vssd vccd mprj_dat_o_user[22] vssd
+ vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input242_A la_data_out_mprj[84] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[96\]_A input383/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_53 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_97 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1296 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1932 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1943 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input507_A la_oenb_mprj[92] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_529 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_389 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_724 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[20\]_A input300/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_953 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_2235 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__432__A _432_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output726_A output726/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_1027 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[87\]_A input373/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_1133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_813 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_529 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_573 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__607__A _607_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_1972 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_1273 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[11\]_A input282/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[2\] _594_/A la_buf_enable\[2\]/B vssd vccd la_buf\[2\]/TE vssd vccd
+ sky130_fd_sc_hd__and2b_1
XANTENNA_user_to_mprj_in_gates\[91\]_B user_to_mprj_in_gates\[91\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1593 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__342__A _342_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_1607 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput518 mprj_adr_o_core[10] vssd vccd _410_/A vssd vccd sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_user_to_mprj_in_ena_buf\[78\]_A input363/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput507 la_oenb_mprj[92] vssd vccd _355_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput529 mprj_adr_o_core[20] vssd vccd _420_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_29_857 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1171 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_315 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[33\] input314/X mprj_logic_high_inst/HI[363] vssd vccd user_to_mprj_in_gates\[33\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_44_827 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__517__A _517_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_99 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2069 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_739 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[11\] _603_/A la_buf_enable\[11\]/B vssd vccd la_buf\[11\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XANTENNA_input192_A la_data_out_mprj[39] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_65 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[82\]_B user_to_mprj_in_gates\[82\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1810 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input457_A la_oenb_mprj[47] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input53_A la_data_out_core[29] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[69\]_A input353/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input624_A user_irq_ena[0] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_1442 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1834 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_389 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1845 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__427__A _427_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_595 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1691 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output676_A output676/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_2169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1566 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[73\]_B user_to_mprj_in_gates\[73\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1905 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[90\] input121/X user_to_mprj_in_gates\[90\]/B vssd vccd user_to_mprj_in_gates\[90\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XANTENNA_la_buf\[115\]_TE la_buf\[115\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1397 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1239 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1745 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1609 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1789 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__337__A _337_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_587 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[64\]_B user_to_mprj_in_gates\[64\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_11_1931 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[62\]_TE mprj_logic_high_inst/HI[264] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
Xinput304 la_iena_mprj[24] vssd vccd input304/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput315 la_iena_mprj[34] vssd vccd input315/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput326 la_iena_mprj[44] vssd vccd input326/X vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_40_2349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[107\] _370_/Y mprj_logic_high_inst/HI[309] vssd vccd la_oenb_core[107]
+ vssd vccd sky130_fd_sc_hd__einvp_8
Xinput337 la_iena_mprj[54] vssd vccd input337/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput348 la_iena_mprj[64] vssd vccd input348/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput359 la_iena_mprj[74] vssd vccd input359/X vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_16_315 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[37\] _629_/Y mprj_logic_high_inst/HI[239] vssd vccd la_oenb_core[37]
+ vssd vccd sky130_fd_sc_hd__einvp_8
X_591_ _591_/A vssd vccd _591_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
Xla_buf_enable\[59\] _651_/A la_buf_enable\[59\]/B vssd vccd la_buf\[59\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_44_679 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_359 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input205_A la_data_out_mprj[50] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_503 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1290 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[55\]_B user_to_mprj_in_gates\[55\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_input574_A mprj_dat_i_user[31] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_1739 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1463 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_1673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1929 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1835 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_473 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[40\]_A user_to_mprj_in_gates\[40\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_39_2009 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1319 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_123 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[60\] user_to_mprj_in_gates\[60\]/Y vssd vccd output711/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_mprj_dat_buf\[9\]_A _441_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output793_A output793/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1920 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_863 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1065 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[46\]_B user_to_mprj_in_gates\[46\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[80\]_A _544_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[85\]_TE mprj_logic_high_inst/HI[287] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__620__A _620_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_2243 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1946 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1597 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[31\]_A user_to_mprj_in_gates\[31\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_26_624 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_657 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_307 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1717 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1897 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_buffers\[98\]_A user_to_mprj_in_gates\[98\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[37\]_B user_to_mprj_in_gates\[37\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_33_1485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_517 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[121\]_B user_to_mprj_in_gates\[121\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[71\]_A _535_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_2029 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1813 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__530__A _530_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_1857 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput101 la_data_out_core[72] vssd vccd input101/X vssd vccd sky130_fd_sc_hd__buf_4
XANTENNA_input155_A la_data_out_mprj[120] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_2293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput123 la_data_out_core[92] vssd vccd input123/X vssd vccd sky130_fd_sc_hd__buf_4
Xinput112 la_data_out_core[82] vssd vccd input112/X vssd vccd sky130_fd_sc_hd__buf_4
Xinput145 la_data_out_mprj[111] vssd vccd _575_/A vssd vccd sky130_fd_sc_hd__buf_4
Xinput134 la_data_out_mprj[101] vssd vccd _565_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_40_2157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput156 la_data_out_mprj[121] vssd vccd _585_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput167 la_data_out_mprj[16] vssd vccd _480_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput178 la_data_out_mprj[26] vssd vccd _490_/A vssd vccd sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_input322_A la_iena_mprj[40] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_17_613 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_643_ _643_/A vssd vccd _643_/Y vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_user_to_mprj_in_buffers\[22\]_A user_to_mprj_in_gates\[22\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_input16_A la_data_out_core[110] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput189 la_data_out_mprj[36] vssd vccd _500_/A vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_29_473 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_933 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_421 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1984 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1973 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_977 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_679 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[64\] _528_/Y la_buf\[64\]/TE vssd vccd la_data_in_core[64] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_user_wb_dat_gates\[30\]_A input573/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_574_ _574_/A vssd vccd _574_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_38_1341 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1915 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1904 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1385 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_823 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[125\]_A _589_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_2297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1650 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[89\]_A user_to_mprj_in_gates\[89\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[28\]_B user_to_mprj_in_gates\[28\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[112\]_B user_to_mprj_in_gates\[112\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[62\]_A _526_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf\[120\] _584_/Y la_buf\[120\]/TE vssd vccd la_data_in_core[120] vssd vccd sky130_fd_sc_hd__einvp_8
Xmprj_adr_buf\[28\] _428_/Y mprj_adr_buf\[28\]/TE vssd vccd mprj_adr_o_user[28] vssd
+ vccd sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf_enable\[80\]_B la_buf_enable\[80\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output639_A output639/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__440__A _440_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1481 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1873 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[53\] input80/X user_to_mprj_in_gates\[53\]/B vssd vccd user_to_mprj_in_gates\[53\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XANTENNA_user_to_mprj_in_buffers\[13\]_A user_to_mprj_in_gates\[13\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_3_1737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1687 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[21\]_A input563/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_buffers\[127\]_A user_to_mprj_in_gates\[127\]/Y vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_2028 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[116\]_A _580_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__615__A _615_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_2337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[19\]_B user_to_mprj_in_gates\[19\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[103\]_B user_to_mprj_in_gates\[103\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[53\]_A _517_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[71\]_B la_buf_enable\[71\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_1521 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__350__A _350_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_1615 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1565 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input8_A la_data_out_core[103] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_771 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1787 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_421 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_410 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_wb_dat_gates\[12\]_A input553/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_914 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_925 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_627 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_78 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_buffers\[118\]_A user_to_mprj_in_gates\[118\]/Y vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_1525 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__525__A _525_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[107\]_A _571_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_17_1981 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_77 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[44\]_A _508_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_1867 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2008 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input272_A la_iena_mprj[110] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[62\]_B la_buf_enable\[62\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_1591 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_1621 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_16 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input537_A mprj_adr_o_core[28] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_1665 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[127\] _390_/A la_buf_enable\[127\]/B vssd vccd la_buf\[127\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_29_281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1827 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_741 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_443 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_626_ _626_/A vssd vccd _626_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_45_785 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_487 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_557_ _557_/A vssd vccd _557_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_user_to_mprj_in_buffers\[109\]_A user_to_mprj_in_gates\[109\]/Y vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_1636 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_620 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__435__A _435_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_488_ _488_/A vssd vccd _488_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_13_693 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2050 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[23\] user_to_mprj_in_gates\[23\]/Y vssd vccd output670/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_la_buf\[35\]_A _499_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output756_A output756/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[53\]_B la_buf_enable\[53\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1131 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[120\]_A _383_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_1979 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2235 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1039 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[125\]_B mprj_logic_high_inst/HI[455] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_27_218 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_774 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1812 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1845 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_777 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__345__A _345_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_608 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1889 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[26\]_A _490_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[44\]_B la_buf_enable\[44\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_2041 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_1941 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1805 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2085 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1423 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[111\]_A _374_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_1985 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_1849 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1467 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[63\] input347/X mprj_logic_high_inst/HI[393] vssd vccd user_to_mprj_in_gates\[63\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_4_1309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[116\]_B mprj_logic_high_inst/HI[446] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[1\] _593_/Y mprj_logic_high_inst/HI[203] vssd vccd la_oenb_core[1]
+ vssd vccd sky130_fd_sc_hd__einvp_8
X_411_ _411_/A vssd vccd _411_/Y vssd vccd sky130_fd_sc_hd__inv_4
Xla_buf_enable\[41\] _633_/A la_buf_enable\[41\]/B vssd vccd la_buf\[41\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XANTENNA_input118_A la_data_out_core[88] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_342_ _342_/A vssd vccd _342_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_la_buf\[11\]_TE la_buf\[11\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_601 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input487_A la_oenb_mprj[74] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input83_A la_data_out_core[56] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_1691 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1642 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[27\] _491_/Y la_buf\[27\]/TE vssd vccd la_data_in_core[27] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf\[17\]_A _481_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_1675 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_656 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[35\]_B la_buf_enable\[35\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[4\]_A input332/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[102\]_A _365_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1821 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1771 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[107\]_B mprj_logic_high_inst/HI[437] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_37_549 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_1635 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1061 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_1668 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[42\]_A_N _634_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_609_ _609_/A vssd vccd _609_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_53_2101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_210 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_2145 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_2189 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[16\] input39/X user_to_mprj_in_gates\[16\]/B vssd vccd user_to_mprj_in_gates\[16\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
Xuser_wb_dat_gates\[29\] input571/X user_wb_ack_gate/B vssd vccd user_wb_dat_gates\[29\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_2
XFILLER_53_1477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[57\]_A_N _649_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_buffers\[26\] user_wb_dat_gates\[26\]/Y vssd vccd output774/A vssd vccd
+ sky130_fd_sc_hd__clkinv_8
XANTENNA_la_buf_enable\[26\]_B la_buf_enable\[26\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_2361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_1732 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1787 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1629 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[127\] input34/X user_to_mprj_in_gates\[127\]/B vssd vccd user_to_mprj_in_gates\[127\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_3_2098 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1397 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[34\]_TE la_buf\[34\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[19\]_TE mprj_logic_high_inst/HI[221] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_1631 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[95\]_A _358_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_585 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_57 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_1951 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1859 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[17\]_B la_buf_enable\[17\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput780 output780/A vssd vccd mprj_dat_i_core[31] vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_47_1793 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1231 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[67\] _330_/Y mprj_logic_high_inst/HI[269] vssd vccd la_oenb_core[67]
+ vssd vccd sky130_fd_sc_hd__einvp_8
Xoutput791 output791/A vssd vccd user2_vdd_powergood vssd vccd sky130_fd_sc_hd__buf_2
Xla_buf_enable\[89\] _352_/A la_buf_enable\[89\]/B vssd vccd la_buf\[89\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XANTENNA_user_to_mprj_in_ena_buf\[96\]_B mprj_logic_high_inst/HI[426] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_48_65 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[15\] _447_/Y mprj_dat_buf\[15\]/TE vssd vccd mprj_dat_o_user[15] vssd
+ vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input235_A la_data_out_mprj[78] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_1381 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1955 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_357 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_711 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input402_A la_oenb_mprj[112] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_2129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[86\]_A _349_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_714 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[20\]_B mprj_logic_high_inst/HI[350] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[2\]_TE la_buf\[2\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_921 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_965 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2247 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_2269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[10\] _410_/Y mprj_adr_buf\[10\]/TE vssd vccd mprj_adr_o_user[10] vssd
+ vccd sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_buffers\[124\] user_to_mprj_in_gates\[124\]/Y vssd vccd output654/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_output719_A output719/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[87\]_B mprj_logic_high_inst/HI[417] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[10\]_A _602_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_692 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[57\]_TE la_buf\[57\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[90\] user_to_mprj_in_gates\[90\]/Y vssd vccd output744/A
+ vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_42_1145 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_571 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_wb_dat_buffers\[0\] user_wb_dat_gates\[0\]/Y vssd vccd output756/A vssd vccd
+ sky130_fd_sc_hd__clkinv_8
XANTENNA_user_to_mprj_oen_buffers\[77\]_A _340_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_1940 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_585 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[11\]_B mprj_logic_high_inst/HI[341] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA__623__A _623_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[4\]_A input576/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_1619 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1933 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2055 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput508 la_oenb_mprj[93] vssd vccd _356_/A vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA_user_to_mprj_in_ena_buf\[78\]_B mprj_logic_high_inst/HI[408] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xinput519 mprj_adr_o_core[11] vssd vccd _411_/A vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_9_1551 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_313 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1595 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_869 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[4\]_A input76/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_817 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[26\] input306/X mprj_logic_high_inst/HI[356] vssd vccd user_to_mprj_in_gates\[26\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_43_327 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_861 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[68\]_A _331_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_574 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_279 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1369 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__533__A _533_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_1623 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_77 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input185_A la_data_out_mprj[32] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1822 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1093 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1866 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input352_A la_iena_mprj[68] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[69\]_B mprj_logic_high_inst/HI[399] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_input46_A la_data_out_core[22] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf\[94\] _558_/Y la_buf\[94\]/TE vssd vccd la_data_in_core[94] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input617_A mprj_sel_o_core[2] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[59\]_A _651_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_533 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1578 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output669_A output669/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__443__A _443_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1917 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[83\] input113/X user_to_mprj_in_gates\[83\]/B vssd vccd user_to_mprj_in_gates\[83\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_26_1630 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1757 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_mprj_dat_buf\[29\]_TE mprj_dat_buf\[29\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1492 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__618__A _618_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_809 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[8\]_TE mprj_logic_high_inst/HI[210] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_34_850 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_599 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__353__A _353_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_1943 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_209 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1391 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_905 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1987 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput305 la_iena_mprj[25] vssd vccd input305/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput316 la_iena_mprj[35] vssd vccd input316/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput327 la_iena_mprj[45] vssd vccd input327/X vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_49_909 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_600 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_78 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1201 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput338 la_iena_mprj[55] vssd vccd input338/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput349 la_iena_mprj[65] vssd vccd input349/X vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_5_1245 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_590_ _590_/A vssd vccd _590_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_43_113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__528__A _528_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_327 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input100_A la_data_out_core[71] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_515 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_559 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_49 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xla_buf\[5\] _469_/Y la_buf\[5\]/TE vssd vccd la_data_in_core[5] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_mprj_pwrgood_A mprj_pwrgood/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input567_A mprj_dat_i_user[25] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_2353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_787 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xmprj_adr_buf\[2\] _402_/Y mprj_adr_buf\[2\]/TE vssd vccd mprj_adr_o_user[2] vssd
+ vccd sky130_fd_sc_hd__einvp_8
XANTENNA_mprj_sel_buf\[3\]_TE mprj_sel_buf\[3\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_1273 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_441 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__438__A _438_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_135 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[53\] user_to_mprj_in_gates\[53\]/Y vssd vccd output703/A
+ vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_17_1607 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output786_A output786/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_1509 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[10\]_A _442_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_897 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_341 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_875 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1965 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_wb_dat_gates\[11\] input552/X user_wb_ack_gate/B vssd vccd user_wb_dat_gates\[11\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_4
XANTENNA_mprj_adr_buf\[28\]_A _428_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1173 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2255 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_953 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_931 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1418 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__348__A _348_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_669 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_319 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[5\]_A _597_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_1729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1497 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_529 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[93\] input380/X mprj_logic_high_inst/HI[423] vssd vccd user_to_mprj_in_gates\[93\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_mprj_adr_buf\[19\]_A _419_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_2261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1869 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xinput102 la_data_out_core[73] vssd vccd input102/X vssd vccd sky130_fd_sc_hd__buf_4
Xmprj_sel_buf\[0\] _396_/Y mprj_sel_buf\[0\]/TE vssd vccd mprj_sel_o_user[0] vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_40_2125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1329 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput124 la_data_out_core[93] vssd vccd input124/X vssd vccd sky130_fd_sc_hd__buf_4
Xinput113 la_data_out_core[83] vssd vccd input113/X vssd vccd sky130_fd_sc_hd__buf_4
Xinput135 la_data_out_mprj[102] vssd vccd _566_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
XANTENNA_input148_A la_data_out_mprj[114] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput168 la_data_out_mprj[17] vssd vccd _481_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xla_buf_enable\[71\] _334_/A la_buf_enable\[71\]/B vssd vccd la_buf\[71\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
Xinput146 la_data_out_mprj[112] vssd vccd _576_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput157 la_data_out_mprj[122] vssd vccd _586_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_40_2169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xinput179 la_data_out_mprj[27] vssd vccd _491_/A vssd vccd sky130_fd_sc_hd__dlymetal6s2s_1
X_642_ _642_/A vssd vccd _642_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_29_441 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_945 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input315_A la_iena_mprj[34] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_989 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_433 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[30\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_573_ _573_/A vssd vccd _573_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_44_477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[57\] _521_/Y la_buf\[57\]/TE vssd vccd la_data_in_core[57] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf\[105\]_TE la_buf\[105\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XPHY_130 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1927 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1217 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_835 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1397 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1531 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1662 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_irq_buffers\[2\]_A user_irq_gates\[2\]/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf\[113\] _577_/Y la_buf\[113\]/TE vssd vccd la_data_in_core[113] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_mprj_adr_buf\[4\]_TE mprj_adr_buf\[4\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1493 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1313 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output701_A output701/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_1699 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[21\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[46\] input72/X user_to_mprj_in_gates\[46\]/B vssd vccd user_to_mprj_in_gates\[46\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_2
XFILLER_23_617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_469 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[52\]_TE mprj_logic_high_inst/HI[254] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_1003 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_2349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__631__A _631_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[8\] input120/X user_to_mprj_in_gates\[8\]/B vssd vccd user_to_mprj_in_gates\[8\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_4
XANTENNA_mprj_dat_buf\[8\]_TE mprj_dat_buf\[8\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_1533 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1340 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_433 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[12\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_639 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_937 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1537 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1851 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_981 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1993 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_89 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[97\] _360_/Y mprj_logic_high_inst/HI[299] vssd vccd la_oenb_core[97]
+ vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_13_1879 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__541__A _541_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input265_A la_iena_mprj[104] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_1633 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_28 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1677 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input432_A la_oenb_mprj[24] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_1839 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[90\]_TE la_buf\[90\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_17_411 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_753 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_455 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_625_ _625_/A vssd vccd _625_/Y vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_user_to_mprj_oen_buffers\[75\]_TE mprj_logic_high_inst/HI[277] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
X_556_ _556_/A vssd vccd _556_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_17_499 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_487_ _487_/A vssd vccd _487_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_9_643 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_632 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_2073 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_2062 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[16\] user_to_mprj_in_gates\[16\]/Y vssd vccd output662/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_47_2109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output749_A output749/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output651_A output651/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__451__A _451_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_1853 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1143 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1706 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1728 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1535 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1693 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_786 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__626__A _626_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_1857 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[4\]_A _404_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__361__A _361_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1478 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2097 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1341 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_1953 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1435 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[56\] input339/X mprj_logic_high_inst/HI[386] vssd vccd user_to_mprj_in_gates\[56\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_8_1479 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_2297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[98\]_TE mprj_logic_high_inst/HI[300] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_1067 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_403 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_410_ _410_/A vssd vccd _410_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_14_447 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[12\] _604_/Y mprj_logic_high_inst/HI[214] vssd vccd la_oenb_core[12]
+ vssd vccd sky130_fd_sc_hd__einvp_8
X_341_ _341_/A vssd vccd _341_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
Xla_buf_enable\[34\] _626_/A la_buf_enable\[34\]/B vssd vccd la_buf\[34\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XANTENNA__536__A _536_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_1481 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[8\] user_to_mprj_in_gates\[8\]/Y vssd vccd output743/A vssd
+ vccd sky130_fd_sc_hd__clkinv_4
XFILLER_10_620 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input382_A la_iena_mprj[95] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_613 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1654 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_668 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input76_A la_data_out_core[4] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_1105 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_830 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[4\]_B mprj_logic_high_inst/HI[334] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xmprj_stb_buf _394_/Y mprj_stb_buf/TE vssd vccd mprj_stb_o_user vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_46_1485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1603 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1833 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_517 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_1647 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1877 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2291 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
X_608_ _608_/A vssd vccd _608_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_32_222 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output699_A output699/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__446__A _446_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_539_ _539_/A vssd vccd _539_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_20_417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_buffers\[19\] user_wb_dat_gates\[19\]/Y vssd vccd output766/A vssd vccd
+ sky130_fd_sc_hd__clkinv_8
XFILLER_5_2309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1744 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1799 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[125\]_B la_buf_enable\[125\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_517 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_2055 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__356__A _356_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_597 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1643 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1665 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[94\]_A input125/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_1963 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1761 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xoutput770 output770/A vssd vccd mprj_dat_i_core[22] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput781 output781/A vssd vccd mprj_dat_i_core[3] vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_8_1243 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_1625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xoutput792 output792/A vssd vccd user_irq[0] vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA_la_buf_enable\[116\]_B la_buf_enable\[116\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_517 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1118 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_77 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input130_A la_data_out_core[99] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_1287 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input228_A la_data_out_mprj[71] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_1393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1967 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_594 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_723 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input597_A mprj_dat_o_core[23] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_buffers\[7\]_A user_wb_dat_gates\[7\]/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[111\] input273/X mprj_logic_high_inst/HI[441] vssd vccd
+ user_to_mprj_in_gates\[111\]/B vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_in_gates\[85\]_A input115/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_973 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_977 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_472 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_421 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_clk_buf_A _391_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[30\]_TE mprj_adr_buf\[30\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_2259 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_671 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[117\] user_to_mprj_in_gates\[117\]/Y vssd vccd output646/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_la_buf_enable\[107\]_B la_buf_enable\[107\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_837 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[83\] user_to_mprj_in_gates\[83\]/Y vssd vccd output736/A
+ vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_18_583 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_542 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_597 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1952 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1805 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[76\]_A input105/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_1849 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1013 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[4\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput509 la_oenb_mprj[94] vssd vccd _357_/A vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_25_2045 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_1923 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_1945 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2067 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1989 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[4\]_B user_to_mprj_in_gates\[4\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_24_520 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2005 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[19\] input298/X mprj_logic_high_inst/HI[349] vssd vccd user_to_mprj_in_gates\[19\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_51_1905 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[67\]_A input95/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_1635 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1061 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_936 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_1834 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input178_A la_data_out_mprj[26] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[41\]_A_N _633_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input345_A la_iena_mprj[61] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input39_A la_data_out_core[16] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input512_A la_oenb_mprj[97] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[56\]_A_N _648_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_1961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xla_buf\[87\] _551_/Y la_buf\[87\]/TE vssd vccd la_data_in_core[87] vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[102\] _365_/A la_buf_enable\[102\]/B vssd vccd la_buf\[102\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_46_177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_881 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1775 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_531 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_501 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_545 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[58\]_A input85/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_1860 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_741 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_785 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_2001 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_291 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[24\]_TE la_buf\[24\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_1929 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_2067 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output731_A output731/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[76\] input105/X user_to_mprj_in_gates\[76\]/B vssd vccd user_to_mprj_in_gates\[76\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_38_601 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_645 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[8\]_A user_to_mprj_in_gates\[8\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_4_1471 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1313 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_862 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_391 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[49\]_A input75/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__634__A _634_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_1793 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1955 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1999 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xinput306 la_iena_mprj[26] vssd vccd input306/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput317 la_iena_mprj[36] vssd vccd input317/X vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_9_1371 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput328 la_iena_mprj[46] vssd vccd input328/X vssd vccd sky130_fd_sc_hd__dlymetal6s2s_1
Xinput339 la_iena_mprj[56] vssd vccd input339/X vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_29_57 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1257 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_843 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_865 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_527 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input295_A la_iena_mprj[16] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[124\]_A input31/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__544__A _544_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[47\]_TE la_buf\[47\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_2321 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input462_A la_oenb_mprj[51] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_irq_ena_buf\[2\] input626/X user_irq_ena_buf\[2\]/B vssd vccd user_irq_gates\[2\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_4_799 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1285 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_1995 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1633 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_497 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1001 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1619 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output681_A output681/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[46\] user_to_mprj_in_gates\[46\]/Y vssd vccd output695/A
+ vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_34_1933 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output779_A output779/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[115\]_A input21/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__454__A _454_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_593 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2195 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1049 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_2109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_943 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_965 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__629__A _629_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[102\] input7/X user_to_mprj_in_gates\[102\]/B vssd vccd user_to_mprj_in_gates\[102\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_53_445 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1009 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[106\]_A input11/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__364__A _364_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_386 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1763 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[86\] input372/X mprj_logic_high_inst/HI[416] vssd vccd user_to_mprj_in_gates\[86\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_49_729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput114 la_data_out_core[84] vssd vccd input114/X vssd vccd sky130_fd_sc_hd__buf_4
Xinput103 la_data_out_core[74] vssd vccd input103/X vssd vccd sky130_fd_sc_hd__buf_4
Xuser_to_mprj_oen_buffers\[112\] _375_/Y mprj_logic_high_inst/HI[314] vssd vccd la_oenb_core[112]
+ vssd vccd sky130_fd_sc_hd__einvp_8
Xinput136 la_data_out_mprj[103] vssd vccd _567_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput125 la_data_out_core[94] vssd vccd input125/X vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_5_1021 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput169 la_data_out_mprj[18] vssd vccd _482_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput158 la_data_out_mprj[123] vssd vccd _587_/A vssd vccd sky130_fd_sc_hd__buf_2
Xinput147 la_data_out_mprj[113] vssd vccd _577_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_40_2137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1065 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[42\] _634_/Y mprj_logic_high_inst/HI[244] vssd vccd la_oenb_core[42]
+ vssd vccd sky130_fd_sc_hd__einvp_8
X_641_ _641_/A vssd vccd _641_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
Xla_buf_enable\[64\] _656_/A la_buf_enable\[64\]/B vssd vccd la_buf\[64\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XANTENNA__539__A _539_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_17_637 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2011 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_irq_buffers\[0\] user_irq_gates\[0\]/Y vssd vccd output792/A vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_input210_A la_data_out_mprj[55] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_1942 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
X_572_ _572_/A vssd vccd _572_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_44_445 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input308_A la_iena_mprj[28] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_1997 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_489 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_131 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_120 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1543 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_335 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1674 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[19\]_TE mprj_dat_buf\[19\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf\[106\] _570_/Y la_buf\[106\]/TE vssd vccd la_data_in_core[106] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA__449__A _449_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_2164 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_445 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_0 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_629 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[39\] input64/X user_to_mprj_in_gates\[39\]/B vssd vccd user_to_mprj_in_gates\[39\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_31_673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1605 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_880 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1097 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[4\]_B la_buf_enable\[4\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__359__A _359_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_445 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_489 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_949 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_640 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1549 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_993 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1571 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input160_A la_data_out_mprj[125] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input258_A la_data_out_mprj[99] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_1105 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1645 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1509 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_599 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_1689 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2081 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input425_A la_oenb_mprj[18] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[119\]_A input281/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_1943 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input21_A la_data_out_core[115] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_721 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_624_ _624_/A vssd vccd _624_/Y vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_user_to_mprj_oen_buffers\[120\]_TE mprj_logic_high_inst/HI[322] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_765 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_555_ _555_/A vssd vccd _555_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_17_467 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_1703 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_486_ _486_/A vssd vccd _486_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_38_1173 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_we_buf _395_/Y mprj_we_buf/TE vssd vccd mprj_we_o_user vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_ena_buf\[50\]_A input333/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_611 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2085 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2096 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_655 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_699 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_872 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output644_A output644/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xmprj_pwrgood mprj_pwrgood/A vssd vccd output788/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_29_1865 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1155 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1019 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2290 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1525 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_798 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_245 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[41\]_A input323/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1869 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__642__A _642_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_809 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1397 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_2221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1447 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_2265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_57 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[49\] input331/X mprj_logic_high_inst/HI[379] vssd vccd user_to_mprj_in_gates\[49\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_42_713 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_23 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_415 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_340_ _340_/A vssd vccd _340_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_42_757 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1313 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_908 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_459 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[32\]_A input313/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[27\] _619_/A la_buf_enable\[27\]/B vssd vccd la_buf\[27\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_39_1493 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__552__A _552_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input375_A la_iena_mprj[89] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input69_A la_data_out_core[43] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_1117 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_2132 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[99\]_A input386/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input542_A mprj_adr_o_core[3] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_2187 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1497 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[42\]_TE mprj_logic_high_inst/HI[244] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_1751 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1615 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1845 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_573 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1889 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_607_ _607_/A vssd vccd _607_/Y vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_32_234 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_538_ _538_/A vssd vccd _538_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_user_to_mprj_in_ena_buf\[23\]_A input303/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_1435 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_469_ _469_/A vssd vccd _469_/Y vssd vccd sky130_fd_sc_hd__inv_2
XANTENNA_output761_A output761/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__462__A _462_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[118\]_TE la_buf\[118\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_1756 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_713 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__637__A _637_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[14\]_A input293/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[94\]_B user_to_mprj_in_gates\[94\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_36_1699 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__372__A _372_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[80\]_TE la_buf\[80\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[65\]_TE mprj_logic_high_inst/HI[267] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xoutput771 output771/A vssd vccd mprj_dat_i_core[23] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput760 output760/A vssd vccd mprj_dat_i_core[13] vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_47_1773 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1211 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xoutput793 output793/A vssd vccd user_irq[1] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput782 output782/A vssd vccd mprj_dat_i_core[4] vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_43_1637 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2040 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_529 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_2073 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input123_A la_data_out_core[92] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_1979 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__547__A _547_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_540 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_irq_ena_buf\[1\]_A input625/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_1831 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_1853 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input492_A la_oenb_mprj[79] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_we_buf_A _395_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_901 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[85\]_B user_to_mprj_in_gates\[85\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[104\] input265/X mprj_logic_high_inst/HI[434] vssd vccd
+ user_to_mprj_in_gates\[104\]/B vssd vccd sky130_fd_sc_hd__and2_1
Xla_buf\[32\] _496_/Y la_buf\[32\]/TE vssd vccd la_data_in_core[32] vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_10_484 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_433 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_wb_dat_gates\[4\] input576/X user_wb_ack_gate/B vssd vccd user_wb_dat_gates\[4\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_4
XFILLER_7_989 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_499 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[70\]_A user_to_mprj_in_gates\[70\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_37_337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[76\] user_to_mprj_in_gates\[76\]/Y vssd vccd output728/A
+ vssd vccd sky130_fd_sc_hd__inv_2
XANTENNA__457__A _457_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_18_551 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_882 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_370 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_595 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_554 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[21\] input45/X user_to_mprj_in_gates\[21\]/B vssd vccd user_to_mprj_in_gates\[21\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_33_1817 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[76\]_B user_to_mprj_in_gates\[76\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_31_2253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1552 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[88\]_TE mprj_logic_high_inst/HI[290] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_buffers\[31\] user_wb_dat_gates\[31\]/Y vssd vccd output780/A vssd vccd
+ sky130_fd_sc_hd__inv_6
XFILLER_47_1025 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1069 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[9\] _441_/Y mprj_dat_buf\[9\]/TE vssd vccd mprj_dat_o_user[9] vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_5_2107 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1531 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1957 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2079 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[61\]_A user_to_mprj_in_gates\[61\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA__367__A _367_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_2131 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_727 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1917 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1441 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2017 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[67\]_B user_to_mprj_in_gates\[67\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_36_1485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1603 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1073 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[72\] _335_/Y mprj_logic_high_inst/HI[274] vssd vccd la_oenb_core[72]
+ vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[94\] _357_/A la_buf_enable\[94\]/B vssd vccd la_buf\[94\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_43_1401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[20\] _452_/Y mprj_dat_buf\[20\]/TE vssd vccd mprj_dat_o_user[20] vssd
+ vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input338_A la_iena_mprj[55] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input240_A la_data_out_mprj[82] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[52\]_A user_to_mprj_in_gates\[52\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_19_337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1732 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1973 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input505_A la_oenb_mprj[90] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_893 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_1787 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_510 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_189 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_841 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_543 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_587 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[58\]_B user_to_mprj_in_gates\[58\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[92\]_A _556_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_1872 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_753 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_2013 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2079 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_992 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output724_A output724/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_613 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[43\]_A user_to_mprj_in_gates\[43\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[69\] input97/X user_to_mprj_in_gates\[69\]/B vssd vccd user_to_mprj_in_gates\[69\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_25_307 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_657 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_649 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_370 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_329 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[49\]_B user_to_mprj_in_gates\[49\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[83\]_A _547_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[0\] _592_/A la_buf_enable\[0\]/B vssd vccd la_buf\[0\]/TE vssd vccd
+ sky130_fd_sc_hd__and2b_1
XANTENNA__650__A _650_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_1721 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput307 la_iena_mprj[27] vssd vccd input307/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput318 la_iena_mprj[37] vssd vccd input318/X vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_44_1765 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1383 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[34\]_A user_to_mprj_in_gates\[34\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xinput329 la_iena_mprj[47] vssd vccd input329/X vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_5_1225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_605 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[31\] input312/X mprj_logic_high_inst/HI[361] vssd vccd user_to_mprj_in_gates\[31\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_45_57 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[20\]_TE mprj_adr_buf\[20\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_693 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_855 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[124\]_B user_to_mprj_in_gates\[124\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[74\]_A _538_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_539 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input190_A la_data_out_mprj[37] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_1411 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_29 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input288_A la_iena_mprj[125] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[92\]_B la_buf_enable\[92\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_2333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1591 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__560__A _560_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1621 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input455_A la_oenb_mprj[45] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_1455 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input51_A la_data_out_core[27] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input622_A user_irq_core[1] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[25\]_A user_to_mprj_in_gates\[25\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_23_1827 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_1562 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1945 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[39\] user_to_mprj_in_gates\[39\]/Y vssd vccd output687/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_user_to_mprj_in_gates\[115\]_B user_to_mprj_in_gates\[115\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[65\]_A _529_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output674_A output674/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1989 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[83\]_B la_buf_enable\[83\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__470__A _470_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_1705 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_2213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1749 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_buffers\[16\]_A user_to_mprj_in_gates\[16\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_41_1916 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1409 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_443 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[24\]_A input566/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_671 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__645__A _645_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[40\]_A_N _632_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[119\]_A _583_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[106\]_B user_to_mprj_in_gates\[106\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[56\]_A _520_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[55\]_A_N _647_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[74\]_B la_buf_enable\[74\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_1731 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__380__A _380_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_1775 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[79\] input364/X mprj_logic_high_inst/HI[409] vssd vccd user_to_mprj_in_gates\[79\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
Xinput115 la_data_out_core[85] vssd vccd input115/X vssd vccd sky130_fd_sc_hd__buf_4
Xinput104 la_data_out_core[75] vssd vccd input104/X vssd vccd sky130_fd_sc_hd__buf_4
Xinput126 la_data_out_core[95] vssd vccd input126/X vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_9_1180 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[105\] _368_/Y mprj_logic_high_inst/HI[307] vssd vccd la_oenb_core[105]
+ vssd vccd sky130_fd_sc_hd__einvp_8
Xinput137 la_data_out_mprj[104] vssd vccd _568_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput159 la_data_out_mprj[124] vssd vccd _588_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput148 la_data_out_mprj[114] vssd vccd _578_/A vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_5_1033 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_640_ _640_/A vssd vccd _640_/Y vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_user_wb_dat_gates\[15\]_A input556/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_22_1871 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_oen_buffers\[35\] _627_/Y mprj_logic_high_inst/HI[237] vssd vccd la_oenb_core[35]
+ vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[57\] _649_/A la_buf_enable\[57\]/B vssd vccd la_buf\[57\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_5_1077 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
X_571_ _571_/A vssd vccd _571_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_44_457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2023 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1311 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2045 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input203_A la_data_out_mprj[49] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__555__A _555_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[14\]_TE la_buf\[14\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XPHY_132 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_110 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_303 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_859 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[47\]_A _511_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input99_A la_data_out_core[70] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_1686 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1555 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_347 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[65\]_B la_buf_enable\[65\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input572_A mprj_dat_i_user[2] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_81 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_2185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1821 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1613 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_2121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1061 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_741 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_925 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_273 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1108 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_1 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1464 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output791_A output791/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_671 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__465__A _465_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_641 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_685 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[38\]_A _502_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[56\]_B la_buf_enable\[56\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_2225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[123\]_A _386_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_2269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[37\]_TE la_buf\[37\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_1397 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_785 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_2321 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_405 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_608 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_980 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__375__A _375_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[29\]_A _493_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_818 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[47\]_B la_buf_enable\[47\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_2325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[114\]_A _377_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_1583 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_523 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1117 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input153_A la_data_out_mprj[119] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_2093 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[119\]_B mprj_logic_high_inst/HI[449] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_24_1955 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input320_A la_iena_mprj[39] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_240 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1977 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_623_ _623_/A vssd vccd _623_/Y vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_input418_A la_oenb_mprj[127] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input14_A la_data_out_core[109] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_777 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xla_buf\[62\] _526_/Y la_buf\[62\]/TE vssd vccd la_data_in_core[62] vssd vccd sky130_fd_sc_hd__einvp_8
X_554_ _554_/A vssd vccd _554_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_18_1715 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_485_ _485_/A vssd vccd _485_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_34_1005 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[50\]_B mprj_logic_high_inst/HI[380] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[5\]_TE la_buf\[5\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_1185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1049 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_667 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[38\]_B la_buf_enable\[38\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xmprj_adr_buf\[26\] _426_/Y mprj_adr_buf\[26\]/TE vssd vccd mprj_adr_o_user[26] vssd
+ vccd sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_ena_buf\[7\]_A input365/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_884 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output637_A output637/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[105\]_A _368_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[40\]_A _632_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_1877 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1167 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_1719 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1189 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[51\] input78/X user_to_mprj_in_gates\[51\]/B vssd vccd user_to_mprj_in_gates\[51\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
Xinput490 la_oenb_mprj[77] vssd vccd _340_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_23_405 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_427 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1105 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[41\]_B mprj_logic_high_inst/HI[371] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_31_471 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1425 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[29\]_B la_buf_enable\[29\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[31\]_A _623_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_2233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input6_A la_data_out_core[101] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_2277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[98\]_A _361_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_725 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_427 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[32\]_B mprj_logic_high_inst/HI[362] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_42_769 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_1325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1601 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_637 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input368_A la_iena_mprj[82] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input270_A la_iena_mprj[109] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_2144 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[99\]_B mprj_logic_high_inst/HI[429] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[22\]_A _614_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_1443 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_876 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1421 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input535_A mprj_adr_o_core[26] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_2199 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_397 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1971 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[125\] _388_/A la_buf_enable\[125\]/B vssd vccd la_buf\[125\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_24_1763 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_1857 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_1627 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_606_ _606_/A vssd vccd _606_/Y vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_user_to_mprj_oen_buffers\[89\]_A _352_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_17_265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_537_ _537_/A vssd vccd _537_/Y vssd vccd sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_ena_buf\[23\]_B mprj_logic_high_inst/HI[353] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_32_246 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_468_ _468_/A vssd vccd _468_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_41_780 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_399_ _399_/A vssd vccd _399_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_9_475 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[21\] user_to_mprj_in_gates\[21\]/Y vssd vccd output668/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_output754_A output754/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_2320 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[99\] input130/X user_to_mprj_in_gates\[99\]/B vssd vccd user_to_mprj_in_gates\[99\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XANTENNA_user_to_mprj_oen_buffers\[13\]_A _605_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_2353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1685 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2013 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1481 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_725 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[14\]_B mprj_logic_high_inst/HI[344] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_23_27 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_419 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1509 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_791 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__653__A _653_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[7\]_A input579/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[110\]_TE mprj_logic_high_inst/HI[312] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_629 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xoutput772 output772/A vssd vccd mprj_dat_i_core[24] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput761 output761/A vssd vccd mprj_dat_i_core[14] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput750 output750/A vssd vccd la_data_in_mprj[96] vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_43_1605 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1785 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xoutput794 output794/A vssd vccd user_irq[2] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput783 output783/A vssd vccd mprj_dat_i_core[5] vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_8_1223 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1173 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_ena_buf\[61\] input345/X mprj_logic_high_inst/HI[391] vssd vccd user_to_mprj_in_gates\[61\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_43_1649 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_2085 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2052 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[7\]_A input109/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_511 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_irq_ena_buf\[1\]_B user_irq_ena_buf\[1\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input116_A la_data_out_core[86] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_533 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_279 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_257 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1111 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_1609 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__563__A _563_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_1177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input485_A la_oenb_mprj[72] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input81_A la_data_out_core[54] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_913 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_445 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[25\] _489_/Y la_buf\[25\]/TE vssd vccd la_data_in_core[25] vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_10_496 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1803 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1273 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_809 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1665 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_861 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_buffers\[69\] user_to_mprj_in_gates\[69\]/Y vssd vccd output720/A
+ vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_45_393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_382 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1829 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__473__A _473_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[14\] input37/X user_to_mprj_in_gates\[14\]/B vssd vccd user_to_mprj_in_gates\[14\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_2
Xuser_wb_dat_gates\[27\] input569/X user_wb_ack_gate/B vssd vccd user_wb_dat_gates\[27\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_2
XFILLER_31_2265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1564 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_wb_dat_buffers\[24\] user_wb_dat_gates\[24\]/Y vssd vccd output772/A vssd vccd
+ sky130_fd_sc_hd__clkinv_8
XFILLER_47_1037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1969 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[125\] input32/X user_to_mprj_in_gates\[125\]/B vssd vccd user_to_mprj_in_gates\[125\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XANTENNA__648__A _648_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_809 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_544 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[31\]_A _463_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_1453 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_739 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_2029 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_385 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__383__A _383_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_1929 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1497 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_209 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[32\]_TE mprj_logic_high_inst/HI[234] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_905 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1615 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1085 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_1413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1031 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[65\] _657_/Y mprj_logic_high_inst/HI[267] vssd vccd la_oenb_core[65]
+ vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[87\] _350_/A la_buf_enable\[87\]/B vssd vccd la_buf\[87\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_19_305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_1457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[13\] _445_/Y mprj_dat_buf\[13\]/TE vssd vccd mprj_dat_o_user[13] vssd
+ vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input233_A la_data_out_mprj[76] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__558__A _558_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1985 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input400_A la_oenb_mprj[110] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[108\]_TE la_buf\[108\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_853 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1799 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[22\]_A _454_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_522 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_555 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_525 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_81 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[7\]_TE mprj_adr_buf\[7\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_2025 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_971 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[122\] user_to_mprj_in_gates\[122\]/Y vssd vccd output652/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_output717_A output717/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_2152 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__468__A _468_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_606 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_669 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[70\]_TE la_buf\[70\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_dat_buf\[13\]_A _445_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_18_382 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[55\]_TE mprj_logic_high_inst/HI[257] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_buffers\[20\]_A user_wb_dat_gates\[20\]/Y vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XFILLER_33_385 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1085 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_2073 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1733 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput308 la_iena_mprj[28] vssd vccd input308/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput319 la_iena_mprj[38] vssd vccd input319/X vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_9_1351 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1777 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_647 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1395 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__378__A _378_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[8\]_A _600_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_2205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_105 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_69 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1537 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_ena_buf\[24\] input304/X mprj_logic_high_inst/HI[354] vssd vccd user_to_mprj_in_gates\[24\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_user_wb_dat_buffers\[11\]_A user_wb_dat_gates\[11\]/Y vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XFILLER_12_503 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1423 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_713 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input183_A la_data_out_mprj[30] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_2209 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_757 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_256 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input448_A la_oenb_mprj[39] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input350_A la_iena_mprj[66] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input44_A la_data_out_core[20] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[92\] _556_/Y la_buf\[92\]/TE vssd vccd la_data_in_core[92] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input615_A mprj_sel_o_core[0] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[93\]_TE la_buf\[93\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_1602 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_81 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1793 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_vdd_pwrgood mprj_vdd_pwrgood/A vssd vccd output789/A vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_user_to_mprj_oen_buffers\[78\]_TE mprj_logic_high_inst/HI[280] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_1574 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_363 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_377 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1957 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output667_A output667/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[81\] input111/X user_to_mprj_in_gates\[81\]/B vssd vccd user_to_mprj_in_gates\[81\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_6_1502 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_455 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1568 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[24\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_105 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_683 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_322 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_27 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1754 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1787 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput105 la_data_out_core[76] vssd vccd input105/X vssd vccd sky130_fd_sc_hd__buf_4
Xinput116 la_data_out_core[86] vssd vccd input116/X vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput127 la_data_out_core[96] vssd vccd input127/X vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput149 la_data_out_mprj[115] vssd vccd _579_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput138 la_data_out_mprj[105] vssd vccd _569_/A vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_9_1192 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1045 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[9\]_A_N _601_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_1900 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
X_570_ _570_/A vssd vccd _570_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_user_wb_dat_gates\[15\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_1933 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2035 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XPHY_100 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_650 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2057 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_469 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_oen_buffers\[28\] _620_/Y mprj_logic_high_inst/HI[230] vssd vccd la_oenb_core[28]
+ vssd vccd sky130_fd_sc_hd__einvp_8
XPHY_133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_122 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_111 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[0\]_A _464_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_697 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_315 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input398_A la_oenb_mprj[109] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_359 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__571__A _571_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf\[3\] _467_/Y la_buf\[3\]/TE vssd vccd la_data_in_core[3] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input565_A mprj_dat_i_user[23] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_2164 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1231 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2017 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1833 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_753 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1877 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[0\] _400_/Y mprj_adr_buf\[0\]/TE vssd vccd mprj_adr_o_user[0] vssd
+ vccd sky130_fd_sc_hd__einvp_8
XANTENNA_user_irq_gates\[0\]_A input621/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_1961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_937 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_2 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[51\] user_to_mprj_in_gates\[51\]/Y vssd vccd output701/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_44_981 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_683 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output784_A output784/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_1309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1721 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_697 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1618 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__481__A _481_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_1039 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[10\]_TE mprj_adr_buf\[10\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1861 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__656__A _656_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[7\]_A _407_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_992 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1507 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__391__A _391_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_329 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_ena_buf\[91\] input378/X mprj_logic_high_inst/HI[421] vssd vccd user_to_mprj_in_gates\[91\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_46_2337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1595 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_517 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input146_A la_data_out_mprj[112] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_1967 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_252 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_622_ _622_/A vssd vccd _622_/Y vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_24_1989 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input313_A la_iena_mprj[32] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__566__A _566_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1691 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_553_ _553_/A vssd vccd _553_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_53_2319 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[55\] _519_/Y la_buf\[55\]/TE vssd vccd la_data_in_core[55] vssd vccd sky130_fd_sc_hd__einvp_8
X_484_ _484_/A vssd vccd _484_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_53_1607 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_ena_buf\[127\] input290/X mprj_logic_high_inst/HI[457] vssd vccd
+ user_to_mprj_in_gates\[127\]/B vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_18_1727 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1017 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1905 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_81 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[7\]_B mprj_logic_high_inst/HI[337] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_5_841 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xmprj_adr_buf\[19\] _419_/Y mprj_adr_buf\[19\]/TE vssd vccd mprj_adr_o_user[19] vssd
+ vccd sky130_fd_sc_hd__einvp_8
Xla_buf\[111\] _575_/Y la_buf\[111\]/TE vssd vccd la_data_in_core[111] vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_29_1845 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_2353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_1889 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[99\] user_to_mprj_in_gates\[99\]/Y vssd vccd output753/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_7_1641 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput480 la_oenb_mprj[68] vssd vccd _331_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput491 la_oenb_mprj[78] vssd vccd _341_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XANTENNA__476__A _476_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[54\]_A_N _646_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_buffers\[9\] user_wb_dat_gates\[9\]/Y vssd vccd output787/A vssd vccd
+ sky130_fd_sc_hd__clkinv_8
Xuser_to_mprj_in_gates\[44\] input70/X user_to_mprj_in_gates\[44\]/B vssd vccd user_to_mprj_in_gates\[44\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_35_277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[69\]_A_N _332_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_1117 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_483 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2001 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1871 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2045 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[6\] input98/X user_to_mprj_in_gates\[6\]/B vssd vccd user_to_mprj_in_gates\[6\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_in_gates\[30\]_A input55/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_1377 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_1004 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_550 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__386__A _386_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2049 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[97\]_A input128/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_439 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_601 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_1337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_781 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_634 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1640 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[95\] _358_/Y mprj_logic_high_inst/HI[297] vssd vccd la_oenb_core[95]
+ vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_48_1709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2123 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input263_A la_iena_mprj[102] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[21\]_A input45/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_1455 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input430_A la_oenb_mprj[22] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[119\]_B la_buf_enable\[119\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[8\] input376/X mprj_logic_high_inst/HI[338] vssd vccd user_to_mprj_in_gates\[8\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_input528_A mprj_adr_o_core[1] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_1775 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1983 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[118\] _381_/A la_buf_enable\[118\]/B vssd vccd la_buf\[118\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_40_1076 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_70 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_605_ _605_/A vssd vccd _605_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_17_277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_536_ _536_/A vssd vccd _536_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_user_to_mprj_in_gates\[88\]_A input118/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_467_ _467_/A vssd vccd _467_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_20_409 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_1579 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_398_ _398_/A vssd vccd _398_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_53_1448 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1702 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_487 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[14\] user_to_mprj_in_gates\[14\]/Y vssd vccd output660/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_la_buf\[27\]_TE la_buf\[27\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output747_A output747/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_2332 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_41 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[12\]_A input35/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_85 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2025 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1313 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[79\]_A input108/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_39 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1971 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_wb_dat_gates\[7\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_608 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xoutput762 output762/A vssd vccd mprj_dat_i_core[15] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput740 output740/A vssd vccd la_data_in_mprj[87] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput751 output751/A vssd vccd la_data_in_mprj[97] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput773 output773/A vssd vccd mprj_dat_i_core[25] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput784 output784/A vssd vccd mprj_dat_i_core[6] vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_8_1257 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_ena_buf\[54\] input337/X mprj_logic_high_inst/HI[384] vssd vccd user_to_mprj_in_gates\[54\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_in_gates\[7\]_B user_to_mprj_in_gates\[7\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_41_2064 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_2097 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_545 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[10\] _602_/Y mprj_logic_high_inst/HI[212] vssd vccd la_oenb_core[10]
+ vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input109_A la_data_out_core[7] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_1822 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_523 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_589 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[6\] user_to_mprj_in_gates\[6\]/Y vssd vccd output721/A vssd
+ vccd sky130_fd_sc_hd__clkinv_4
Xla_buf_enable\[32\] _624_/A la_buf_enable\[32\]/B vssd vccd la_buf\[32\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_14_269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_1719 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1189 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1009 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_925 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input380_A la_iena_mprj[93] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input478_A la_oenb_mprj[66] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[18\] _482_/Y la_buf\[18\]/TE vssd vccd la_data_in_core[18] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input74_A la_data_out_core[48] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1790 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1815 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_195 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_173 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_1285 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1859 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2251 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1791 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1633 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1677 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output697_A output697/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_1201 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_519_ _519_/A vssd vccd _519_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_53_1289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_2277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_buffers\[17\] user_wb_dat_gates\[17\]/Y vssd vccd output764/A vssd vccd
+ sky130_fd_sc_hd__clkinv_4
Xuser_to_mprj_in_gates\[118\] input24/X user_to_mprj_in_gates\[118\]/B vssd vccd user_to_mprj_in_gates\[118\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_3_1132 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_501 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_556 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_707 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_589 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1329 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_917 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_405 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1425 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_1043 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[58\] _650_/Y mprj_logic_high_inst/HI[260] vssd vccd la_oenb_core[58]
+ vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_47_637 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_1469 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1817 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_851 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input226_A la_data_out_mprj[6] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_821 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1997 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1229 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[127\]_A input34/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__574__A _574_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_865 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_397 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input595_A mprj_dat_o_core[21] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[100\]_A input261/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_751 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_559 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_1429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_983 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_buffers\[115\] user_to_mprj_in_gates\[115\]/Y vssd vccd output644/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_46_1093 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[81\] user_to_mprj_in_gates\[81\]/Y vssd vccd output734/A
+ vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_38_637 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_2017 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[100\]_TE mprj_logic_high_inst/HI[302] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[118\]_A input24/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__484__A _484_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_2328 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1649 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1974 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2085 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1903 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_29 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput309 la_iena_mprj[29] vssd vccd input309/X vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_44_1745 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_27 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1789 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1609 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_659 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_629 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[109\]_A input14/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__394__A _394_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_1803 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_ena_buf\[17\] input296/X mprj_logic_high_inst/HI[347] vssd vccd user_to_mprj_in_gates\[17\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_40_813 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1705 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_559 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1749 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1435 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_725 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input176_A la_data_out_mprj[24] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_268 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_769 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input343_A la_iena_mprj[5] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_1943 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__569__A _569_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input37_A la_data_out_core[14] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1761 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[85\] _549_/Y la_buf\[85\]/TE vssd vccd la_data_in_core[85] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input510_A la_oenb_mprj[95] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input608_A mprj_dat_o_core[4] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[123\]_TE mprj_logic_high_inst/HI[325] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_629 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[100\] _363_/A la_buf_enable\[100\]/B vssd vccd la_buf\[100\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_35_607 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_1586 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_331 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[80\]_A input366/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_835 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_375 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_389 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2143 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1514 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[74\] input103/X user_to_mprj_in_gates\[74\]/B vssd vccd user_to_mprj_in_gates\[74\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XANTENNA__479__A _479_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[22\]_TE mprj_logic_high_inst/HI[224] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_467 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_489 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_437 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[71\]_A input356/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_695 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1593 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[7\]_B la_buf_enable\[7\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_1782 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput117 la_data_out_core[87] vssd vccd input117/X vssd vccd sky130_fd_sc_hd__buf_4
Xinput106 la_data_out_core[77] vssd vccd input106/X vssd vccd sky130_fd_sc_hd__buf_4
XANTENNA__389__A _389_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_1553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_209 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput128 la_data_out_core[97] vssd vccd input128/X vssd vccd sky130_fd_sc_hd__buf_4
Xinput139 la_data_out_mprj[106] vssd vccd _570_/A vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_44_1597 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1057 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_1851 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[62\]_A input346/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_2069 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XPHY_134 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_123 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_112 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_327 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input293_A la_iena_mprj[14] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_1243 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_533 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input460_A la_oenb_mprj[4] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input558_A mprj_dat_i_user[17] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_2029 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[60\]_TE la_buf\[60\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_2176 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_1287 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_irq_ena_buf\[0\] input624/X user_irq_ena_buf\[0\]/B vssd vccd user_irq_gates\[0\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_oen_buffers\[45\]_TE mprj_logic_high_inst/HI[247] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_1845 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_1637 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1889 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1085 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_905 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_irq_gates\[0\]_B user_irq_gates\[0\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_1433 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_1973 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_949 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_437 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XPHY_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[53\]_A input336/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_993 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_695 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_662 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_654 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[44\] user_to_mprj_in_gates\[44\]/Y vssd vccd output693/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_30_153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output777_A output777/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1733 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_41 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1007 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2001 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1873 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_mprj_sel_buf\[1\]_A _397_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[100\] input5/X user_to_mprj_in_gates\[100\]/B vssd vccd user_to_mprj_in_gates\[100\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_2
XANTENNA_user_to_mprj_in_ena_buf\[44\]_A input326/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_2345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2209 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_816 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1964 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_809 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_1877 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[83\]_TE la_buf\[83\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_1590 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[68\]_TE mprj_logic_high_inst/HI[270] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_2305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1563 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_2349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[84\] input370/X mprj_logic_high_inst/HI[414] vssd vccd user_to_mprj_in_gates\[84\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_49_529 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[110\] _373_/Y mprj_logic_high_inst/HI[312] vssd vccd la_oenb_core[110]
+ vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_29_264 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[40\] _632_/Y mprj_logic_high_inst/HI[242] vssd vccd la_oenb_core[40]
+ vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[62\] _654_/A la_buf_enable\[62\]/B vssd vccd la_buf\[62\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XANTENNA_input139_A la_data_out_mprj[106] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_621_ _621_/A vssd vccd _621_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_44_245 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_552_ _552_/A vssd vccd _552_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_input306_A la_iena_mprj[26] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[35\]_A input316/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_1775 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_483_ _483_/A vssd vccd _483_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_13_643 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[48\] _512_/Y la_buf\[48\]/TE vssd vccd la_data_in_core[48] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA__582__A _582_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1029 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1917 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[2\]_A _434_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_2321 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xla_buf\[104\] _568_/Y la_buf\[104\]/TE vssd vccd la_data_in_core[104] vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_7_1653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput481 la_oenb_mprj[69] vssd vccd _332_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput470 la_oenb_mprj[59] vssd vccd _651_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_36_713 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput492 la_oenb_mprj[79] vssd vccd _342_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XANTENNA_user_to_mprj_in_ena_buf\[26\]_A input306/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_757 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[37\] input62/X user_to_mprj_in_gates\[37\]/B vssd vccd user_to_mprj_in_gates\[37\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_1_1296 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_1129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_985 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__492__A _492_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_462 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[8\]_A_N _600_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_2013 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_1883 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2057 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[91\]_A user_to_mprj_in_gates\[91\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[30\]_B user_to_mprj_in_gates\[30\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_28_1345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1389 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1163 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_27 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1016 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_713 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1049 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[17\]_A input296/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2017 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_749 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[97\]_B user_to_mprj_in_gates\[97\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_22_451 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_793 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_646 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1371 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[88\] _351_/Y mprj_logic_high_inst/HI[290] vssd vccd la_oenb_core[88]
+ vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_46_2113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_2157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input256_A la_data_out_mprj[97] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[21\]_B user_to_mprj_in_gates\[21\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_46_1467 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[82\]_A user_to_mprj_in_gates\[82\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_49_337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1995 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input423_A la_oenb_mprj[16] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__577__A _577_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_1787 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_604_ _604_/A vssd vccd _604_/Y vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_27_82 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_535_ _535_/A vssd vccd _535_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_17_289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[88\]_B user_to_mprj_in_gates\[88\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_53_1405 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_466_ _466_/A vssd vccd _466_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_43_81 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1861 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_397_ _397_/A vssd vccd _397_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_40_292 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1714 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_499 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[31\] _431_/Y mprj_adr_buf\[31\]/TE vssd vccd mprj_adr_o_user[31] vssd
+ vccd sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_buffers\[120\]_A user_to_mprj_in_gates\[120\]/Y vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output642_A output642/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_2344 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_2208 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_53 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[73\]_A user_to_mprj_in_gates\[73\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[12\]_B user_to_mprj_in_gates\[12\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_42_1821 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_97 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__487__A _487_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_521 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_2337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[79\]_B user_to_mprj_in_gates\[79\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_34_2083 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[111\]_A user_to_mprj_in_gates\[111\]/Y vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_1691 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xoutput730 output730/A vssd vccd la_data_in_mprj[78] vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA_la_buf\[100\]_A _564_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput763 output763/A vssd vccd mprj_dat_i_core[16] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput741 output741/A vssd vccd la_data_in_mprj[88] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput752 output752/A vssd vccd la_data_in_mprj[98] vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_48_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xoutput774 output774/A vssd vccd mprj_dat_i_core[26] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput785 output785/A vssd vccd mprj_dat_i_core[7] vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA_user_to_mprj_in_buffers\[64\]_A user_to_mprj_in_gates\[64\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA__397__A _397_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_1916 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_ena_buf\[47\] input329/X mprj_logic_high_inst/HI[377] vssd vccd user_to_mprj_in_gates\[47\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_mprj_adr_buf\[23\]_TE mprj_adr_buf\[23\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_557 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[25\] _617_/A la_buf_enable\[25\]/B vssd vccd la_buf\[25\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_7_937 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input373_A la_iena_mprj[87] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[102\]_A user_to_mprj_in_gates\[102\]/Y vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[53\]_A_N _645_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_469 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input67_A la_data_out_core[41] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input540_A mprj_adr_o_core[30] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[55\]_A user_to_mprj_in_gates\[55\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_26_1827 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[68\]_A_N _331_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_2241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_1297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2263 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1645 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_896 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1689 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_708 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[95\]_A _559_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_518_ _518_/A vssd vccd _518_/Y vssd vccd sky130_fd_sc_hd__inv_2
X_449_ _449_/A vssd vccd _449_/Y vssd vccd sky130_fd_sc_hd__inv_4
XFILLER_31_2289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1599 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_981 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[46\]_A user_to_mprj_in_gates\[46\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_9_1578 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1100 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1144 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_863 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1971 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_2101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[86\]_A _550_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_719 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2105 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[37\]_A user_to_mprj_in_gates\[37\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[10\]_A _474_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_1055 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_863 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1757 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input219_A la_data_out_mprj[63] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[17\]_TE la_buf\[17\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input121_A la_data_out_core[90] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_321 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1631 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[127\]_B user_to_mprj_in_gates\[127\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[77\]_A _541_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input490_A la_oenb_mprj[77] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[100\]_B mprj_logic_high_inst/HI[430] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_input588_A mprj_dat_o_core[15] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[95\]_B la_buf_enable\[95\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[102\] input263/X mprj_logic_high_inst/HI[432] vssd vccd
+ user_to_mprj_in_gates\[102\]/B vssd vccd sky130_fd_sc_hd__and2_1
Xla_buf\[30\] _494_/Y la_buf\[30\]/TE vssd vccd la_data_in_core[30] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA__590__A _590_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_gates\[2\] input572/X user_wb_ack_gate/B vssd vccd user_wb_dat_gates\[2\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_8
XFILLER_6_277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2303 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_buffers\[28\]_A user_to_mprj_in_gates\[28\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_46_1061 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1635 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[108\] user_to_mprj_in_gates\[108\]/Y vssd vccd output636/A
+ vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_24_2071 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_104 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[74\] user_to_mprj_in_gates\[74\]/Y vssd vccd output726/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_45_181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_693 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[118\]_B user_to_mprj_in_gates\[118\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_21_505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[68\]_A _532_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_1043 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[86\]_B la_buf_enable\[86\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_1915 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2097 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1959 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[19\]_A user_to_mprj_in_gates\[19\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xmprj_dat_buf\[7\] _439_/Y mprj_dat_buf\[7\]/TE vssd vccd mprj_dat_o_user[7] vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_44_1757 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_wb_dat_gates\[27\]_A input569/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_39 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[10\]_B la_buf_enable\[10\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_1470 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_27 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[109\]_B user_to_mprj_in_gates\[109\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_24_387 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[59\]_A _523_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_1717 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_869 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1815 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1105 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1859 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[77\]_B la_buf_enable\[77\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_1149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_593 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1613 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_1447 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input169_A la_data_out_mprj[18] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[70\] _333_/Y mprj_logic_high_inst/HI[272] vssd vccd la_oenb_core[70]
+ vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[92\] _355_/A la_buf_enable\[92\]/B vssd vccd la_buf\[92\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_43_1201 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1955 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_925 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1999 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input336_A la_iena_mprj[53] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[18\]_A input559/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_2338 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_1289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1773 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[78\] _542_/Y la_buf\[78\]/TE vssd vccd la_data_in_core[78] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input503_A la_oenb_mprj[89] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__585__A _585_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_1598 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_641 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_343 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[80\]_B mprj_logic_high_inst/HI[410] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[8\]_TE la_buf\[8\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_685 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1038 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_387 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[68\]_B la_buf_enable\[68\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_571 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[70\]_A _333_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output722_A output722/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_2205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2155 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1526 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[67\] input95/X user_to_mprj_in_gates\[67\]/B vssd vccd user_to_mprj_in_gates\[67\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_4_1261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__495__A _495_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[71\]_B mprj_logic_high_inst/HI[401] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_33_1425 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[59\]_B la_buf_enable\[59\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[126\]_A _389_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[61\]_A _653_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_1521 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput118 la_data_out_core[88] vssd vccd input118/X vssd vccd sky130_fd_sc_hd__buf_4
Xinput107 la_data_out_core[78] vssd vccd input107/X vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_44_1565 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput129 la_data_out_core[98] vssd vccd input129/X vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_40_1429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1957 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[62\]_B mprj_logic_high_inst/HI[392] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XPHY_124 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_102 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_685 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_135 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1369 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_335 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1525 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_1623 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_1569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input286_A la_iena_mprj[123] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_51 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[52\]_A _644_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[117\]_A _380_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_545 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input453_A la_oenb_mprj[43] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_589 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1741 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input620_A mprj_we_o_core vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_1649 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1097 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_405 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_917 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1985 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_909 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[53\]_B mprj_logic_high_inst/HI[383] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XPHY_4 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_1701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_buffers\[37\] user_to_mprj_in_gates\[37\]/Y vssd vccd output685/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_31_666 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output672_A output672/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1480 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_895 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[108\]_A _371_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[43\]_A _635_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_2013 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1705 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1841 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1885 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1209 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1378 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_1080 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_29 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[44\]_B mprj_logic_high_inst/HI[374] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_39_1656 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_460 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1943 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_839 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_828 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_2281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1889 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[113\]_TE mprj_logic_high_inst/HI[315] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[34\]_A _626_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[77\] input362/X mprj_logic_high_inst/HI[407] vssd vccd user_to_mprj_in_gates\[77\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_mprj_clk_buf_TE mprj_clk_buf/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_1373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[103\] _366_/Y mprj_logic_high_inst/HI[305] vssd vccd la_oenb_core[103]
+ vssd vccd sky130_fd_sc_hd__einvp_8
X_620_ _620_/A vssd vccd _620_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_29_276 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1671 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[33\] _625_/Y mprj_logic_high_inst/HI[235] vssd vccd la_oenb_core[33]
+ vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_mprj_adr_buf\[30\]_A _430_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_551_ _551_/A vssd vccd _551_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_2_1765 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xla_buf_enable\[55\] _647_/A la_buf_enable\[55\]/B vssd vccd la_buf\[55\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XANTENNA_user_to_mprj_in_ena_buf\[35\]_B mprj_logic_high_inst/HI[365] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
X_482_ _482_/A vssd vccd _482_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_input201_A la_data_out_mprj[47] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_2012 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_780 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_953 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_611 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_699 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input97_A la_data_out_core[69] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1929 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[12\]_TE mprj_logic_high_inst/HI[214] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input570_A mprj_dat_i_user[28] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_821 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[25\]_A _617_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_1665 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput482 la_oenb_mprj[6] vssd vccd _598_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput460 la_oenb_mprj[4] vssd vccd _596_/A vssd vccd sky130_fd_sc_hd__buf_2
Xinput471 la_oenb_mprj[5] vssd vccd _597_/A vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_36_725 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput493 la_oenb_mprj[7] vssd vccd _599_/A vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA_mprj_adr_buf\[21\]_A _421_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[26\]_B mprj_logic_high_inst/HI[356] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_1_1264 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_441 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj2_vdd_pwrgood_A mprj2_vdd_pwrgood/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_997 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1597 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[16\]_A _608_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_1851 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1895 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2069 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1313 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_2361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_1513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1693 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_39 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_725 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_mprj_adr_buf\[12\]_A _412_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[17\]_B mprj_logic_high_inst/HI[347] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_23_1991 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1431 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[50\]_TE la_buf\[50\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_2029 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2321 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[35\]_TE mprj_logic_high_inst/HI[237] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_658 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_117 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1383 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[109\]_A_N _372_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[29\] _461_/Y mprj_dat_buf\[29\]/TE vssd vccd mprj_dat_o_user[29] vssd
+ vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input151_A la_data_out_mprj[117] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_1479 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_389 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input249_A la_data_out_mprj[90] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1799 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input416_A la_oenb_mprj[125] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_603_ _603_/A vssd vccd _603_/Y vssd vccd sky130_fd_sc_hd__inv_2
XANTENNA_input12_A la_data_out_core[107] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_61 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_94 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xla_buf\[60\] _524_/Y la_buf\[60\]/TE vssd vccd la_data_in_core[60] vssd vccd sky130_fd_sc_hd__einvp_8
X_534_ _534_/A vssd vccd _534_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_53_2129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_465_ _465_/A vssd vccd _465_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA__593__A _593_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_761 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_93 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_423 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_396_ _396_/A vssd vccd _396_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_35_1873 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1726 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1759 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[24\] _424_/Y mprj_adr_buf\[24\]/TE vssd vccd mprj_adr_o_user[24] vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_5_673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output635_A output635/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_2141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_65 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2091 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1833 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2196 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1877 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[73\]_TE la_buf\[73\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput290 la_iena_mprj[127] vssd vccd input290/X vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_7_1495 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_555 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[58\]_TE mprj_logic_high_inst/HI[260] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_2305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_2349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_271 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_2095 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[9\] _601_/A la_buf_enable\[9\]/B vssd vccd la_buf\[9\]/TE vssd vccd
+ sky130_fd_sc_hd__and2b_1
Xoutput720 output720/A vssd vccd la_data_in_mprj[69] vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_43_2309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xoutput731 output731/A vssd vccd la_data_in_mprj[79] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput742 output742/A vssd vccd la_data_in_mprj[89] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput753 output753/A vssd vccd la_data_in_mprj[99] vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_28_1121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xoutput775 output775/A vssd vccd mprj_dat_i_core[27] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput764 output764/A vssd vccd mprj_dat_i_core[17] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput786 output786/A vssd vccd mprj_dat_i_core[8] vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA_input4_A la_data_out_core[0] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_1321 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_1332 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[22\]_TE mprj_dat_buf\[22\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[18\] _610_/A la_buf_enable\[18\]/B vssd vccd la_buf\[18\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_7_949 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_1581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input199_A la_data_out_mprj[45] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[1\]_TE mprj_logic_high_inst/HI[203] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_input366_A la_iena_mprj[80] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_irq_gates\[1\] input622/X user_irq_gates\[1\]/B vssd vccd user_irq_gates\[1\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_11_1191 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input533_A mprj_adr_o_core[24] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_1839 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[96\]_TE la_buf\[96\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__588__A _588_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_2325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[123\] _386_/A la_buf_enable\[123\]/B vssd vccd la_buf\[123\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XANTENNA_la_buf_enable\[7\]_A_N _599_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_dat_buf\[25\]_A _457_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_1381 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_517_ _517_/A vssd vccd _517_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
X_448_ _448_/A vssd vccd _448_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
X_379_ _379_/A vssd vccd _379_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_35_1681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output752_A output752/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_2153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[97\] input128/X user_to_mprj_in_gates\[97\]/B vssd vccd user_to_mprj_in_gates\[97\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XANTENNA__498__A _498_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_809 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1112 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_mprj_dat_buf\[16\]_A _448_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_875 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1156 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_buffers\[23\]_A user_wb_dat_gates\[23\]/Y vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XFILLER_37_897 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1983 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1189 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_29 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1467 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_ack_buffer_A user_wb_ack_gate/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_1309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1743 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_1798 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_2253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2117 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_2297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1067 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1769 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_wb_dat_buffers\[14\]_A user_wb_dat_gates\[14\]/Y vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XFILLER_28_897 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input114_A la_data_out_core[84] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_385 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1209 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_377 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1687 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_1409 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_580 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_713 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input483_A la_oenb_mprj[70] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_1810 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_757 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[23\] _487_/Y la_buf\[23\]/TE vssd vccd la_data_in_core[23] vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_6_245 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2326 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_473 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_81 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1073 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1647 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2083 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1421 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_99 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[67\] user_to_mprj_in_gates\[67\]/Y vssd vccd output718/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_45_193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_517 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[12\] input35/X user_to_mprj_in_gates\[12\]/B vssd vccd user_to_mprj_in_gates\[12\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_2
Xuser_wb_dat_gates\[25\] input567/X user_wb_ack_gate/B vssd vccd user_wb_dat_gates\[25\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_2
XFILLER_31_2021 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1927 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_wb_dat_buffers\[22\] user_wb_dat_gates\[22\]/Y vssd vccd output770/A vssd vccd
+ sky130_fd_sc_hd__clkinv_8
XANTENNA_mprj_adr_buf\[13\]_TE mprj_adr_buf\[13\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[123\] input30/X user_to_mprj_in_gates\[123\]/B vssd vccd user_to_mprj_in_gates\[123\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XANTENNA_user_wb_dat_gates\[27\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_39 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[52\]_A_N _644_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_377 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_804 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_1827 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[67\]_A_N _330_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_1117 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_2290 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_buffers\[0\]_A user_wb_dat_gates\[0\]/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_749 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1967 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[63\] _655_/Y mprj_logic_high_inst/HI[265] vssd vccd la_oenb_core[63]
+ vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[85\] _348_/A la_buf_enable\[85\]/B vssd vccd la_buf\[85\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_0_977 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_937 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[11\] _443_/Y mprj_dat_buf\[11\]/TE vssd vccd mprj_dat_o_user[11] vssd
+ vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input231_A la_data_out_mprj[74] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[18\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input329_A la_iena_mprj[47] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_dat_buf\[1\]_TE mprj_dat_buf\[1\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_1785 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[3\]_A _467_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[100\]_B la_buf_enable\[100\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_355 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_697 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_314 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_399 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[121\]_TE la_buf\[121\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_1217 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[127\] _591_/Y la_buf\[127\]/TE vssd vccd la_data_in_core[127] vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_28_1709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1971 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[120\] user_to_mprj_in_gates\[120\]/Y vssd vccd output650/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_26_2167 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output715_A output715/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_1780 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1805 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1273 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1849 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2138 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1437 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1735 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[60\]_A input88/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput108 la_data_out_core[79] vssd vccd input108/X vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_44_1533 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xinput119 la_data_out_core[89] vssd vccd input119/X vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_44_1577 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_981 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_114 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_103 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_601 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_303 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[22\] input302/X mprj_logic_high_inst/HI[352] vssd vccd user_to_mprj_in_gates\[22\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_25_664 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XPHY_136 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_645 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_697 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_483 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_347 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1061 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1083 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input181_A la_data_out_mprj[29] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input279_A la_iena_mprj[117] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_1267 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_557 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[51\]_A input78/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input446_A la_oenb_mprj[37] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input42_A la_data_out_core[19] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_1021 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1775 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput620 mprj_we_o_core vssd vccd _395_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_0_796 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xla_buf\[90\] _554_/Y la_buf\[90\]/TE vssd vccd la_data_in_core[90] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input613_A mprj_dat_o_core[9] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__596__A _596_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_789 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_981 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_5 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_461 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_601 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[91\]_TE mprj_logic_high_inst/HI[293] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[1\]_A user_to_mprj_in_gates\[1\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_7_10 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_188 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1746 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1069 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_2193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output665_A output665/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_391 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[42\]_A input68/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_1313 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_2058 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2025 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1717 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_601 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_472 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1668 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1911 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_645 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_965 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_29 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1201 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_678 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_807 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1245 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1808 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1999 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_2293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput90 la_data_out_core[62] vssd vccd input90/X vssd vccd sky130_fd_sc_hd__buf_4
XANTENNA_user_to_mprj_in_gates\[33\]_A input58/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_1341 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1385 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1227 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_550_ _550_/A vssd vccd _550_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_22_1683 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_461 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[8\] _600_/Y mprj_logic_high_inst/HI[210] vssd vccd la_oenb_core[8]
+ vssd vccd sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[26\] _618_/Y mprj_logic_high_inst/HI[228] vssd vccd la_oenb_core[26]
+ vssd vccd sky130_fd_sc_hd__einvp_8
X_481_ _481_/A vssd vccd _481_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
Xla_buf_enable\[48\] _640_/A la_buf_enable\[48\]/B vssd vccd la_buf\[48\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_13_623 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_965 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input396_A la_oenb_mprj[107] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_1345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[1\] _465_/Y la_buf\[1\]/TE vssd vccd la_data_in_core[1] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input563_A mprj_dat_i_user[21] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_833 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1031 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_321 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[24\]_A input48/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1116 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2251 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1677 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xinput450 la_oenb_mprj[40] vssd vccd _632_/A vssd vccd sky130_fd_sc_hd__buf_4
Xinput461 la_oenb_mprj[50] vssd vccd _642_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput472 la_oenb_mprj[60] vssd vccd _652_/A vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_36_737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput483 la_oenb_mprj[70] vssd vccd _333_/A vssd vccd sky130_fd_sc_hd__buf_2
Xinput494 la_oenb_mprj[80] vssd vccd _343_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_40_1794 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_781 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output782_A output782/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_954 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1565 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_671 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_1429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[15\]_A input38/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1661 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1525 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1443 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_217 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_1752 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2090 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1362 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1395 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_869 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1931 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input144_A la_data_out_mprj[110] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_1193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_602_ _602_/A vssd vccd _602_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_2_1541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input311_A la_iena_mprj[30] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input409_A la_oenb_mprj[119] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_533_ _533_/A vssd vccd _533_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
X_464_ _464_/A vssd vccd _464_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_13_431 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[125\] input288/X mprj_logic_high_inst/HI[455] vssd vccd
+ user_to_mprj_in_gates\[125\]/B vssd vccd sky130_fd_sc_hd__and2_1
Xla_buf\[53\] _517_/Y la_buf\[53\]/TE vssd vccd la_data_in_core[53] vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_13_475 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_435 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_395_ _395_/A vssd vccd _395_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_35_1841 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1885 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_641 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_685 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[17\] _417_/Y mprj_adr_buf\[17\]/TE vssd vccd mprj_adr_o_user[17] vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_4_77 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1801 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1981 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_buffers\[97\] user_to_mprj_in_gates\[97\]/Y vssd vccd output751/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_output628_A output628/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_1845 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1441 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2017 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_1889 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput280 la_iena_mprj[118] vssd vccd input280/X vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_7_1485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[103\]_TE mprj_logic_high_inst/HI[305] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
Xinput291 la_iena_mprj[12] vssd vccd input291/X vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_36_567 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[42\] input68/X user_to_mprj_in_gates\[42\]/B vssd vccd user_to_mprj_in_gates\[42\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_36_589 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_buffers\[7\] user_wb_dat_gates\[7\]/Y vssd vccd output785/A vssd vccd
+ sky130_fd_sc_hd__clkinv_8
XANTENNA_user_to_mprj_in_ena_buf\[121\]_A input284/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_2317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_291 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1985 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_991 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xoutput710 output710/A vssd vccd la_data_in_mprj[5] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput721 output721/A vssd vccd la_data_in_mprj[6] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput732 output732/A vssd vccd la_data_in_mprj[7] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput743 output743/A vssd vccd la_data_in_mprj[8] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput754 output754/A vssd vccd la_data_in_mprj[9] vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_28_1133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[4\] input76/X user_to_mprj_in_gates\[4\]/B vssd vccd user_to_mprj_in_gates\[4\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_4
Xoutput776 output776/A vssd vccd mprj_dat_i_core[28] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput765 output765/A vssd vccd mprj_dat_i_core[18] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput787 output787/A vssd vccd mprj_dat_i_core[9] vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_45_2181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1861 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[112\]_A input274/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_1803 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1284 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_467 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_1593 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_979 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1509 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[93\] _356_/Y mprj_logic_high_inst/HI[295] vssd vccd la_oenb_core[93]
+ vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_2_622 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input261_A la_iena_mprj[100] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input359_A la_iena_mprj[74] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[126\]_TE mprj_logic_high_inst/HI[328] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[6\] input354/X mprj_logic_high_inst/HI[336] vssd vccd user_to_mprj_in_gates\[6\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_input526_A mprj_adr_o_core[18] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1614 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[116\] _379_/A la_buf_enable\[116\]/B vssd vccd la_buf\[116\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XANTENNA_user_to_mprj_in_ena_buf\[103\]_A input264/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_516_ _516_/A vssd vccd _516_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_35_2361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_447_ _447_/A vssd vccd _447_/Y vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_20_209 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_1660 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_378_ _378_/A vssd vccd _378_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_35_1693 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[12\] user_to_mprj_in_gates\[12\]/Y vssd vccd output658/A
+ vssd vccd sky130_fd_sc_hd__clkinv_8
XANTENNA_output745_A output745/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[40\]_TE la_buf\[40\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_2321 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_2198 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1464 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[25\]_TE mprj_logic_high_inst/HI[227] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_1653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1951 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_813 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_887 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1402 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1995 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[108\]_A_N _371_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_2147 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_2169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1479 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1782 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_29 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1923 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1079 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[52\] input335/X mprj_logic_high_inst/HI[382] vssd vccd user_to_mprj_in_gates\[52\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_47_629 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[92\]_A input379/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input107_A la_data_out_core[78] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[4\] user_to_mprj_in_gates\[4\]/Y vssd vccd output699/A vssd
+ vccd sky130_fd_sc_hd__clkinv_4
Xla_buf_enable\[30\] _622_/A la_buf_enable\[30\]/B vssd vccd la_buf\[30\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_24_41 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_389 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_85 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_890 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_592 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_725 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input476_A la_oenb_mprj[64] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_1877 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_769 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[16\] _480_/Y la_buf\[16\]/TE vssd vccd la_data_in_core[16] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf\[63\]_TE la_buf\[63\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input72_A la_data_out_core[46] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_95 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_1317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[48\]_TE mprj_logic_high_inst/HI[250] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__599__A _599_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_2338 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1659 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1085 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_93 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[9\] _409_/Y mprj_adr_buf\[9\]/TE vssd vccd mprj_adr_o_user[9] vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_43_1973 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2095 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1591 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[83\]_A input369/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_813 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1190 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output695_A output695/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_890 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_529 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_2033 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1056 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_1933 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_gates\[18\] input559/X user_wb_ack_gate/B vssd vccd user_wb_dat_gates\[18\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_4
Xuser_wb_dat_buffers\[15\] user_wb_dat_gates\[15\]/Y vssd vccd output762/A vssd vccd
+ sky130_fd_sc_hd__clkinv_4
XFILLER_29_1261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_mprj_dat_buf\[12\]_TE mprj_dat_buf\[12\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[116\] input22/X user_to_mprj_in_gates\[116\]/B vssd vccd user_to_mprj_in_gates\[116\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XANTENNA_user_to_mprj_in_ena_buf\[74\]_A input359/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_695 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1508 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_529 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[86\]_TE la_buf\[86\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_551 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_1839 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[6\]_A_N _598_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1637 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2073 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[126\] _389_/Y mprj_logic_high_inst/HI[328] vssd vccd la_oenb_core[126]
+ vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_47_1361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_905 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[56\] _648_/Y mprj_logic_high_inst/HI[258] vssd vccd la_oenb_core[56]
+ vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[78\] _341_/A la_buf_enable\[78\]/B vssd vccd la_buf\[78\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_48_949 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_85 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input224_A la_data_out_mprj[68] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[65\]_A input349/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_51 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_827 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_665 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input593_A mprj_dat_o_core[1] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_1229 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_61 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_533 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1103 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2102 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_2113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1983 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[113\] user_to_mprj_in_gates\[113\]/Y vssd vccd output642/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_26_2179 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_415 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output708_A output708/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[56\]_A input339/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_1285 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1817 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_860 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1703 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[60\]_B user_to_mprj_in_gates\[60\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_44_2213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput109 la_data_out_core[7] vssd vccd input109/X vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_5_1005 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_1589 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[47\]_A input329/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_1915 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_993 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_985 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_115 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_104 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_462 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_126 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_613 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1603 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_315 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[15\] input294/X mprj_logic_high_inst/HI[345] vssd vccd user_to_mprj_in_gates\[15\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_40_657 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_359 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_503 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input174_A la_data_out_mprj[22] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[51\]_B user_to_mprj_in_gates\[51\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_4_569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input341_A la_iena_mprj[58] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input439_A la_oenb_mprj[30] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput610 mprj_dat_o_core[6] vssd vccd _438_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput621 user_irq_core[0] vssd vccd input621/X vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_43_1033 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_1607 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1787 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input35_A la_data_out_core[12] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_757 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[83\] _547_/Y la_buf\[83\]/TE vssd vccd la_data_in_core[83] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input606_A mprj_dat_o_core[31] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[38\]_A input319/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_993 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_6 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_613 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_473 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1769 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[5\]_A _437_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_1037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_22 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output658_A output658/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[42\]_B user_to_mprj_in_gates\[42\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[51\]_A_N _643_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1990 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1791 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[72\] input101/X user_to_mprj_in_gates\[72\]/B vssd vccd user_to_mprj_in_gates\[72\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_6_2037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[66\]_A_N _329_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[29\]_A input309/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_245 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1060 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_495 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_977 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_1923 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_657 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1382 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1257 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1522 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput91 la_data_out_core[63] vssd vccd input91/X vssd vccd sky130_fd_sc_hd__buf_4
Xinput80 la_data_out_core[53] vssd vccd input80/X vssd vccd sky130_fd_sc_hd__buf_4
XANTENNA_la_buf_enable\[19\]_A_N _611_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_517 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_buffers\[94\]_A user_to_mprj_in_gates\[94\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[33\]_B user_to_mprj_in_gates\[33\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_44_1353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[111\]_TE la_buf\[111\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_1239 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[26\]_TE mprj_adr_buf\[26\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_1756 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1745 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_2181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_480_ _480_/A vssd vccd _480_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_51_2003 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_oen_buffers\[19\] _611_/Y mprj_logic_high_inst/HI[221] vssd vccd la_oenb_core[19]
+ vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_13_635 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_977 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_421 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1313 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1357 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_41 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input291_A la_iena_mprj[12] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input389_A la_oenb_mprj[100] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_63 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_85 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[121\]_A _585_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input556_A mprj_dat_i_user[15] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_1043 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1805 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[85\]_A user_to_mprj_in_gates\[85\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[24\]_B user_to_mprj_in_gates\[24\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_4_377 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2263 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1509 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xinput451 la_oenb_mprj[41] vssd vccd _633_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput440 la_oenb_mprj[31] vssd vccd _623_/A vssd vccd sky130_fd_sc_hd__buf_2
Xinput462 la_oenb_mprj[51] vssd vccd _643_/A vssd vccd sky130_fd_sc_hd__buf_2
Xinput473 la_oenb_mprj[61] vssd vccd _653_/A vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA__400__A _400_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput495 la_oenb_mprj[81] vssd vccd _344_/A vssd vccd sky130_fd_sc_hd__buf_4
Xinput484 la_oenb_mprj[71] vssd vccd _334_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_36_749 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_793 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2201 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[42\] user_to_mprj_in_gates\[42\]/Y vssd vccd output691/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_16_495 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1522 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output775_A output775/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1577 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[123\]_A user_to_mprj_in_gates\[123\]/Y vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[112\]_A _576_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_1905 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[76\]_A user_to_mprj_in_gates\[76\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[15\]_B user_to_mprj_in_gates\[15\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1537 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1155 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1199 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_226 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_421 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1043 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1021 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1775 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[114\]_A user_to_mprj_in_gates\[114\]/Y vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_17_1764 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1065 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[103\]_A _567_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[67\]_A user_to_mprj_in_gates\[67\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_2_837 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[82\] input368/X mprj_logic_high_inst/HI[412] vssd vccd user_to_mprj_in_gates\[82\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_la_buf\[40\]_A _504_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[81\]_TE mprj_logic_high_inst/HI[283] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_1943 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_329 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2232 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_727 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[60\] _652_/A la_buf_enable\[60\]/B vssd vccd la_buf\[60\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XANTENNA_input137_A la_data_out_mprj[104] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_601_ _601_/A vssd vccd _601_/Y vssd vccd sky130_fd_sc_hd__inv_2
X_532_ _532_/A vssd vccd _532_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_input304_A la_iena_mprj[24] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_463_ _463_/A vssd vccd _463_/Y vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_25_281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_443 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1419 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_51 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_785 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[46\] _510_/Y la_buf\[46\]/TE vssd vccd la_data_in_core[46] vssd vccd sky130_fd_sc_hd__einvp_8
X_394_ _394_/A vssd vccd _394_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_51_1121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_487 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_447 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[118\] input280/X mprj_logic_high_inst/HI[448] vssd vccd
+ user_to_mprj_in_gates\[118\]/B vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_in_buffers\[105\]_A user_to_mprj_in_gates\[105\]/Y vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[58\]_A user_to_mprj_in_gates\[58\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_5_697 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[31\]_A _495_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf\[102\] _566_/Y la_buf\[102\]/TE vssd vccd la_data_in_core[102] vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_42_1813 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1453 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_841 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1857 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput270 la_iena_mprj[109] vssd vccd input270/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput281 la_iena_mprj[119] vssd vccd input281/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput292 la_iena_mprj[13] vssd vccd input292/X vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_51_505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[98\]_A _562_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_579 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[35\] input60/X user_to_mprj_in_gates\[35\]/B vssd vccd user_to_mprj_in_gates\[35\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XANTENNA_user_to_mprj_in_ena_buf\[121\]_B mprj_logic_high_inst/HI[451] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_32_730 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1915 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_1341 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_970 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xoutput700 output700/A vssd vccd la_data_in_mprj[50] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput711 output711/A vssd vccd la_data_in_mprj[60] vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA_user_to_mprj_in_buffers\[49\]_A user_to_mprj_in_gates\[49\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xoutput722 output722/A vssd vccd la_data_in_mprj[70] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput733 output733/A vssd vccd la_data_in_mprj[80] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput744 output744/A vssd vccd la_data_in_mprj[90] vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA_la_buf\[22\]_A _486_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput788 output788/A vssd vccd user1_vcc_powergood vssd vccd sky130_fd_sc_hd__buf_2
Xoutput777 output777/A vssd vccd mprj_dat_i_core[29] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput766 output766/A vssd vccd mprj_dat_i_core[19] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput755 output755/A vssd vccd mprj_ack_i_core vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_28_1145 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_29 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[40\]_B la_buf_enable\[40\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1481 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_557 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1873 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[112\]_B mprj_logic_high_inst/HI[442] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[89\]_A _553_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_2175 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1441 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[86\] _349_/Y mprj_logic_high_inst/HI[288] vssd vccd la_oenb_core[86]
+ vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf\[13\]_A _477_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_1201 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_122 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_1223 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input254_A la_data_out_mprj[95] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_645 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_678 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[31\]_B la_buf_enable\[31\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_188 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1565 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1773 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input421_A la_oenb_mprj[14] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[0\]_A input260/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input519_A mprj_adr_o_core[11] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[109\] _372_/A la_buf_enable\[109\]/B vssd vccd la_buf\[109\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_2
XFILLER_46_877 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_515_ _515_/A vssd vccd _515_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_user_to_mprj_in_ena_buf\[103\]_B mprj_logic_high_inst/HI[433] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_2_1394 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_446_ _446_/A vssd vccd _446_/Y vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_la_buf_enable\[98\]_B la_buf_enable\[98\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_593 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_377_ _377_/A vssd vccd _377_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_31_2237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_1525 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1672 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_461 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output640_A output640/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_2177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output738_A output738/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[22\]_B la_buf_enable\[22\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_1621 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_1665 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_321 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_825 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1963 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1414 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[89\]_B la_buf_enable\[89\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_18_1892 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1723 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[91\]_A _354_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_2233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[13\]_B la_buf_enable\[13\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_1935 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_310 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[45\] input327/X mprj_logic_high_inst/HI[375] vssd vccd user_to_mprj_in_gates\[45\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_in_ena_buf\[92\]_B mprj_logic_high_inst/HI[422] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_43_836 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_357 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_1667 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_711 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[23\] _615_/A la_buf_enable\[23\]/B vssd vccd la_buf\[23\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_24_97 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_755 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[82\]_A _345_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_41 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input469_A la_oenb_mprj[58] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input371_A la_iena_mprj[85] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_910 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input65_A la_data_out_core[3] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1307 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_1329 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_497 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_1941 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1445 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_1985 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[83\]_B mprj_logic_high_inst/HI[413] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_34_825 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_869 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1013 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_593 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1609 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output688_A output688/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_429_ _429_/A vssd vccd _429_/Y vssd vccd sky130_fd_sc_hd__inv_8
XFILLER_35_2181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_2045 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1945 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[73\]_A _336_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_1705 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_1367 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_wb_dat_gates\[0\]_A input550/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput1 caravel_clk vssd vccd _391_/A vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_37_641 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[109\] input14/X user_to_mprj_in_gates\[109\]/B vssd vccd user_to_mprj_in_gates\[109\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XANTENNA_user_to_mprj_in_ena_buf\[74\]_B mprj_logic_high_inst/HI[404] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_20_1771 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_313 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[0\]_A input4/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[116\]_TE mprj_logic_high_inst/HI[318] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[64\]_A _656_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_1553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_217 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1649 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2085 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[119\] _382_/Y mprj_logic_high_inst/HI[321] vssd vccd la_oenb_core[119]
+ vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_25_2361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_1237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_917 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2319 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_405 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_97 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[49\] _641_/Y mprj_logic_high_inst/HI[251] vssd vccd la_oenb_core[49]
+ vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_ena_buf\[65\]_B mprj_logic_high_inst/HI[395] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_28_685 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input217_A la_data_out_mprj[61] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[30\]_TE la_buf\[30\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input586_A mprj_dat_o_core[13] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[15\]_TE mprj_logic_high_inst/HI[217] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_51 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_501 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1631 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[55\]_A _647_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_73 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_545 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[100\] input261/X mprj_logic_high_inst/HI[430] vssd vccd
+ user_to_mprj_in_gates\[100\]/B vssd vccd sky130_fd_sc_hd__and2_1
Xuser_wb_dat_gates\[0\] input550/X user_wb_ack_gate/B vssd vccd user_wb_dat_gates\[0\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_4
XFILLER_48_1115 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__403__A _403_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_2125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1995 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[107\]_A_N _370_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[106\] user_to_mprj_in_gates\[106\]/Y vssd vccd output634/A
+ vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_19_641 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_1793 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[72\] user_to_mprj_in_gates\[72\]/Y vssd vccd output724/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_user_to_mprj_in_ena_buf\[56\]_B mprj_logic_high_inst/HI[386] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_47_961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1829 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_wb_dat_gates\[30\] input573/X user_wb_ack_gate/B vssd vccd user_wb_dat_gates\[30\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_2
XFILLER_33_2129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[46\]_A _638_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_2225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[5\] _437_/Y mprj_dat_buf\[5\]/TE vssd vccd mprj_dat_o_user[5] vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_44_2269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_405 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_909 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[47\]_B mprj_logic_high_inst/HI[377] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[53\]_TE la_buf\[53\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_953 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XPHY_116 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_105 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[38\]_TE mprj_logic_high_inst/HI[240] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XPHY_138 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_127 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_327 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_669 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[37\]_A _629_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_1973 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_515 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input167_A la_data_out_mprj[16] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_1711 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xla_buf_enable\[90\] _353_/A la_buf_enable\[90\]/B vssd vccd la_buf\[90\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_7_1805 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput611 mprj_dat_o_core[7] vssd vccd _439_/A vssd vccd sky130_fd_sc_hd__buf_4
Xinput600 mprj_dat_o_core[26] vssd vccd _458_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput622 user_irq_core[1] vssd vccd input622/X vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_7_1849 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input334_A la_iena_mprj[51] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_1799 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_769 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[38\]_B mprj_logic_high_inst/HI[368] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_input28_A la_data_out_core[121] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input501_A la_oenb_mprj[87] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf\[76\] _540_/Y la_buf\[76\]/TE vssd vccd la_data_in_core[76] vssd vccd sky130_fd_sc_hd__einvp_8
XPHY_7 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_441 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_135 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1005 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[28\]_A _620_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_1049 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2209 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output720_A output720/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_725 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[24\]_A _424_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[76\]_TE la_buf\[76\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_1359 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[65\] input93/X user_to_mprj_in_gates\[65\]/B vssd vccd user_to_mprj_in_gates\[65\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XANTENNA_user_to_mprj_in_ena_buf\[29\]_B mprj_logic_high_inst/HI[359] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_4_1072 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_953 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[5\]_A_N _597_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_2073 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2062 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1815 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_1935 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[19\]_A _611_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_1225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1394 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[1\]_A _593_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_1534 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput81 la_data_out_core[54] vssd vccd input81/X vssd vccd sky130_fd_sc_hd__buf_4
Xinput70 la_data_out_core[44] vssd vccd input70/X vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput92 la_data_out_core[64] vssd vccd input92/X vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_24_1939 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_202 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_mprj_adr_buf\[15\]_A _415_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_17_419 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[25\]_TE mprj_dat_buf\[25\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_901 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_934 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2026 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_433 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_989 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_669 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[4\]_TE mprj_logic_high_inst/HI[206] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_32_53 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1369 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_97 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input284_A la_iena_mprj[121] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_1817 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input451_A la_oenb_mprj[41] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_389 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input549_A mprj_cyc_o_core vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[99\]_TE la_buf\[99\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_2325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput430 la_oenb_mprj[22] vssd vccd _614_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_48_533 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput463 la_oenb_mprj[52] vssd vccd _644_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput441 la_oenb_mprj[32] vssd vccd _624_/A vssd vccd sky130_fd_sc_hd__buf_2
Xinput452 la_oenb_mprj[42] vssd vccd _634_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput474 la_oenb_mprj[62] vssd vccd _654_/A vssd vccd sky130_fd_sc_hd__buf_2
Xinput485 la_oenb_mprj[72] vssd vccd _335_/A vssd vccd sky130_fd_sc_hd__buf_2
Xinput496 la_oenb_mprj[82] vssd vccd _345_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_5_1381 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_2213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[35\] user_to_mprj_in_gates\[35\]/Y vssd vccd output683/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_34_1534 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output670_A output670/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output768_A output768/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_1870 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1589 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2017 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1917 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_1549 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_588 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_238 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_761 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_466 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_1743 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1667 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1787 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1618 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1033 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1077 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1055 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_ena_buf\[75\] input360/X mprj_logic_high_inst/HI[405] vssd vccd user_to_mprj_in_gates\[75\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA__501__A _501_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_1861 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1703 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1955 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_1173 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1808 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[101\] _364_/Y mprj_logic_high_inst/HI[303] vssd vccd la_oenb_core[101]
+ vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_40_1037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1015 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_600_ _600_/A vssd vccd _600_/Y vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_18_739 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_oen_buffers\[31\] _623_/Y mprj_logic_high_inst/HI[233] vssd vccd la_oenb_core[31]
+ vssd vccd sky130_fd_sc_hd__einvp_8
X_531_ _531_/A vssd vccd _531_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_33_709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[53\] _645_/A la_buf_enable\[53\]/B vssd vccd la_buf\[53\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_2_1576 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_400 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_462_ _462_/A vssd vccd _462_/Y vssd vccd sky130_fd_sc_hd__inv_6
XANTENNA_la_buf_enable\[50\]_A_N _642_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_393_ _393_/A vssd vccd _393_/Y vssd vccd sky130_fd_sc_hd__inv_6
XFILLER_13_455 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input499_A la_oenb_mprj[85] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_1133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_797 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_499 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_459 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[39\] _503_/Y la_buf\[39\]/TE vssd vccd la_data_in_core[39] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf_enable\[65\]_A_N _657_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input95_A la_data_out_core[67] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_1177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_665 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1647 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__411__A _411_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_893 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_mprj_dat_buf\[28\]_A _460_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_853 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1869 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xinput271 la_iena_mprj[10] vssd vccd input271/X vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput260 la_iena_mprj[0] vssd vccd input260/X vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_40_2261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_897 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput282 la_iena_mprj[11] vssd vccd input282/X vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput293 la_iena_mprj[14] vssd vccd input293/X vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_51_517 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[18\]_A_N _610_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_1607 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1097 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_742 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[28\] input52/X user_to_mprj_in_gates\[28\]/B vssd vccd user_to_mprj_in_gates\[28\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_34_2054 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_1943 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[101\]_TE la_buf\[101\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1927 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[16\]_TE mprj_adr_buf\[16\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[0\]_A _400_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput701 output701/A vssd vccd la_data_in_mprj[51] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput712 output712/A vssd vccd la_data_in_mprj[61] vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_47_1703 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xoutput723 output723/A vssd vccd la_data_in_mprj[71] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput734 output734/A vssd vccd la_data_in_mprj[81] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput745 output745/A vssd vccd la_data_in_mprj[91] vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_12_1684 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xoutput767 output767/A vssd vccd mprj_dat_i_core[1] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput778 output778/A vssd vccd mprj_dat_i_core[2] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput756 output756/A vssd vccd mprj_dat_i_core[0] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput789 output789/A vssd vccd user1_vdd_powergood vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA_mprj_adr_buf\[0\]_TE mprj_adr_buf\[0\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_dat_buf\[19\]_A _451_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1493 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_buffers\[26\]_A user_wb_dat_gates\[26\]/Y vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XFILLER_41_1357 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1841 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_385 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1885 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2187 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_425 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1420 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1453 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_447 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1497 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_602 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[79\] _342_/Y mprj_logic_high_inst/HI[281] vssd vccd la_oenb_core[79]
+ vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_46_1235 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2223 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_105 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xmprj_dat_buf\[27\] _459_/Y mprj_dat_buf\[27\]/TE vssd vccd mprj_dat_o_user[27] vssd
+ vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input247_A la_data_out_mprj[89] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_dat_buf\[4\]_TE mprj_dat_buf\[4\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_2317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1785 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_41 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[0\]_B mprj_logic_high_inst/HI[330] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_18_503 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input414_A la_oenb_mprj[123] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_buffers\[17\]_A user_wb_dat_gates\[17\]/Y vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XANTENNA_input10_A la_data_out_core[105] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_517 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_514_ _514_/A vssd vccd _514_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_2_1373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1905 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1916 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[124\]_TE la_buf\[124\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_445_ _445_/A vssd vccd _445_/Y vssd vccd sky130_fd_sc_hd__clkinv_4
X_376_ _376_/A vssd vccd _376_/Y vssd vccd sky130_fd_sc_hd__inv_2
XANTENNA__406__A _406_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1971 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_941 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[22\] _422_/Y mprj_adr_buf\[22\]/TE vssd vccd mprj_adr_o_user[22] vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_5_473 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output633_A output633/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_1633 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1677 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_837 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[121\]_B la_buf_enable\[121\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_17_580 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_550 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[71\]_TE mprj_logic_high_inst/HI[273] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_18_1871 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_1735 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xla_buf_enable\[7\] _599_/A la_buf_enable\[7\]/B vssd vccd la_buf\[7\]/TE vssd vccd
+ sky130_fd_sc_hd__and2b_1
XANTENNA_user_to_mprj_in_gates\[90\]_A input121/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_1779 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_1500 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1820 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_609 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input2_A caravel_clk2 vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_1831 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1947 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_322 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[38\] input319/X mprj_logic_high_inst/HI[368] vssd vccd user_to_mprj_in_gates\[38\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_la_buf_enable\[112\]_B la_buf_enable\[112\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_1635 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_550 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_723 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1679 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_767 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[16\] _608_/A la_buf_enable\[16\]/B vssd vccd la_buf\[16\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_52_1261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_266 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input197_A la_data_out_mprj[43] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_53 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[81\]_A input111/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_buffers\[3\]_A user_wb_dat_gates\[3\]/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_922 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input364_A la_iena_mprj[79] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_2307 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_421 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input58_A la_data_out_core[33] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_432 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_51 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input531_A mprj_adr_o_core[22] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_2125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1953 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xla_buf_enable\[121\] _384_/A la_buf_enable\[121\]/B vssd vccd la_buf\[121\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_4_2169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1997 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_311 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[6\]_A _470_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[103\]_B la_buf_enable\[103\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[94\]_TE mprj_logic_high_inst/HI[296] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_1779 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_428_ _428_/A vssd vccd _428_/Y vssd vccd sky130_fd_sc_hd__inv_8
XFILLER_31_2057 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_359_ _359_/A vssd vccd _359_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_31_1367 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output750_A output750/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[72\]_A input101/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_1790 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[95\] input126/X user_to_mprj_in_gates\[95\]/B vssd vccd user_to_mprj_in_gates\[95\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_2
XFILLER_9_1324 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_wb_dat_gates\[0\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_1441 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput2 caravel_clk2 vssd vccd _392_/A vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_42_1485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_601 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_645 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1783 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[0\]_B user_to_mprj_in_gates\[0\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_36_1278 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1565 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[63\]_A input91/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_2097 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1385 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_697 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input112_A la_data_out_core[82] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_1490 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1009 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1908 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_531 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input481_A la_oenb_mprj[69] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input579_A mprj_dat_i_user[7] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_557 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_85 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1665 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[21\] _485_/Y la_buf\[21\]/TE vssd vccd la_data_in_core[21] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_gates\[54\]_A input81/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_1643 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_1127 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_785 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_284 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_907 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_973 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_409 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_697 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[65\] user_to_mprj_in_gates\[65\]/Y vssd vccd output716/A
+ vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_user_to_mprj_in_buffers\[4\]_A user_to_mprj_in_gates\[4\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_37_2277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_391 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[10\] input15/X user_to_mprj_in_gates\[10\]/B vssd vccd user_to_mprj_in_gates\[10\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_2
Xuser_wb_dat_gates\[23\] input565/X user_wb_ack_gate/B vssd vccd user_wb_dat_gates\[23\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_2
XFILLER_30_884 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1721 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[45\]_A input71/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_buffers\[20\] user_wb_dat_gates\[20\]/Y vssd vccd output768/A vssd vccd
+ sky130_fd_sc_hd__clkinv_8
XFILLER_44_2237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1093 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[121\] input28/X user_to_mprj_in_gates\[121\]/B vssd vccd user_to_mprj_in_gates\[121\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_53_910 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_461 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_921 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_106 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1329 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1591 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_998 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XPHY_139 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_117 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_128 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_637 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1941 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1985 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[36\]_A input61/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[120\]_A input27/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__504__A _504_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_527 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_1425 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1469 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1817 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_2220 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_oen_buffers\[61\] _653_/Y mprj_logic_high_inst/HI[263] vssd vccd la_oenb_core[61]
+ vssd vccd sky130_fd_sc_hd__einvp_8
Xinput601 mprj_dat_o_core[27] vssd vccd _459_/A vssd vccd sky130_fd_sc_hd__buf_2
Xinput612 mprj_dat_o_core[8] vssd vccd _440_/A vssd vccd sky130_fd_sc_hd__buf_2
Xla_buf_enable\[83\] _346_/A la_buf_enable\[83\]/B vssd vccd la_buf\[83\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_5_2253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput623 user_irq_core[2] vssd vccd input623/X vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_47_225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input327_A la_iena_mprj[45] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_41 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1438 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_85 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1989 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_461 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_8 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_645 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[69\] _533_/Y la_buf\[69\]/TE vssd vccd la_data_in_core[69] vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_43_497 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1017 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_844 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_321 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_57 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__414__A _414_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[111\]_A input17/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[27\]_A input51/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf\[125\] _589_/Y la_buf\[125\]/TE vssd vccd la_data_in_core[125] vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_10_1771 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output713_A output713/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_1305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[106\]_TE mprj_logic_high_inst/HI[308] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[58\] input85/X user_to_mprj_in_gates\[58\]/B vssd vccd user_to_mprj_in_gates\[58\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_39_1605 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_921 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_461 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2041 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2085 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1969 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[102\]_A input7/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[18\]_A input41/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput82 la_data_out_core[55] vssd vccd input82/X vssd vccd sky130_fd_sc_hd__buf_4
Xinput71 la_data_out_core[45] vssd vccd input71/X vssd vccd sky130_fd_sc_hd__buf_4
Xinput60 la_data_out_core[35] vssd vccd input60/X vssd vccd sky130_fd_sc_hd__buf_4
Xinput93 la_data_out_core[65] vssd vccd input93/X vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_48_2181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1609 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2001 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1480 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2045 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[20\]_TE la_buf\[20\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_214 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_781 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_751 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1115 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[20\] input300/X mprj_logic_high_inst/HI[350] vssd vccd user_to_mprj_in_gates\[20\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_53_795 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_659 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_445 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_946 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[106\]_A_N _369_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_2038 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_489 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1793 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input277_A la_iena_mprj[115] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_357 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1829 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input444_A la_oenb_mprj[35] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input40_A la_data_out_core[17] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_501 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput420 la_oenb_mprj[13] vssd vccd _605_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_48_545 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput453 la_oenb_mprj[43] vssd vccd _635_/A vssd vccd sky130_fd_sc_hd__buf_4
Xinput431 la_oenb_mprj[23] vssd vccd _615_/A vssd vccd sky130_fd_sc_hd__buf_2
Xinput442 la_oenb_mprj[33] vssd vccd _625_/A vssd vccd sky130_fd_sc_hd__buf_2
Xinput464 la_oenb_mprj[53] vssd vccd _645_/A vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA_input611_A mprj_dat_o_core[7] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput497 la_oenb_mprj[83] vssd vccd _346_/A vssd vccd sky130_fd_sc_hd__buf_4
Xinput475 la_oenb_mprj[63] vssd vccd _655_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput486 la_oenb_mprj[73] vssd vccd _336_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_5_1393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__409__A _409_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_2361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_209 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[28\] user_to_mprj_in_gates\[28\]/Y vssd vccd output675/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_output663_A output663/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_1882 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2029 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[43\]_TE la_buf\[43\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_2321 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1929 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[0\]_B la_buf_enable\[0\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[28\]_TE mprj_logic_high_inst/HI[230] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_1168 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[124\]_A input287/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_1413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1711 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_489 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1679 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1799 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1089 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1955 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1343 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_817 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1873 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_ena_buf\[68\] input352/X mprj_logic_high_inst/HI[398] vssd vccd user_to_mprj_in_gates\[68\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_2_2201 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_1715 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_1005 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_10 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1027 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_1185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_707 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1049 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2256 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_530_ _530_/A vssd vccd _530_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_user_to_mprj_in_ena_buf\[115\]_A input277/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_1566 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_461_ _461_/A vssd vccd _461_/Y vssd vccd sky130_fd_sc_hd__clkinv_4
Xuser_to_mprj_oen_buffers\[24\] _616_/Y mprj_logic_high_inst/HI[226] vssd vccd la_oenb_core[24]
+ vssd vccd sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[6\] _598_/Y mprj_logic_high_inst/HI[208] vssd vccd la_oenb_core[6]
+ vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[46\] _638_/A la_buf_enable\[46\]/B vssd vccd la_buf\[46\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
X_392_ _392_/A vssd vccd _392_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_13_412 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_721 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_467 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input394_A la_oenb_mprj[105] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[66\]_TE la_buf\[66\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_1145 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input88_A la_data_out_core[60] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_1189 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input561_A mprj_dat_i_user[1] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[4\]_A_N _596_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_2101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_821 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_865 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput250 la_data_out_mprj[91] vssd vccd _555_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput261 la_iena_mprj[100] vssd vccd input261/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput272 la_iena_mprj[110] vssd vccd input272/X vssd vccd sky130_fd_sc_hd__clkbuf_1
XANTENNA_user_to_mprj_in_ena_buf\[106\]_A input267/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput294 la_iena_mprj[15] vssd vccd input294/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput283 la_iena_mprj[120] vssd vccd input283/X vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_51_529 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_209 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1619 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_220 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output780_A output780/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_1999 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_1939 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1229 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_471 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xoutput702 output702/A vssd vccd la_data_in_mprj[52] vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_47_1715 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xoutput713 output713/A vssd vccd la_data_in_mprj[62] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput724 output724/A vssd vccd la_data_in_mprj[72] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput735 output735/A vssd vccd la_data_in_mprj[82] vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA__602__A _602_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_dat_buf\[15\]_TE mprj_dat_buf\[15\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_1737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xoutput779 output779/A vssd vccd mprj_dat_i_core[30] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput768 output768/A vssd vccd mprj_dat_i_core[20] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput757 output757/A vssd vccd mprj_dat_i_core[10] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput746 output746/A vssd vccd la_data_in_mprj[92] vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_41_1314 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1369 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_548 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1897 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[89\]_TE la_buf\[89\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_721 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_1839 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2199 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1465 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_437 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_459 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__512__A _512_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_636 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1247 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2235 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_53 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input142_A la_data_out_mprj[109] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[95\]_A input382/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_2053 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_813 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_515 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_559 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input407_A la_oenb_mprj[117] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_513_ _513_/A vssd vccd _513_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_33_529 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_1928 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_444_ _444_/A vssd vccd _444_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
Xla_buf\[51\] _515_/Y la_buf\[51\]/TE vssd vccd la_data_in_core[51] vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_35_2353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_573 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[123\] input286/X mprj_logic_high_inst/HI[453] vssd vccd
+ user_to_mprj_in_gates\[123\]/B vssd vccd sky130_fd_sc_hd__and2_1
X_375_ _375_/A vssd vccd _375_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_31_1505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_953 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_997 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_1401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1983 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__422__A _422_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_441 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[15\] _415_/Y mprj_adr_buf\[15\]/TE vssd vccd mprj_adr_o_user[15] vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_9_1539 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[95\] user_to_mprj_in_gates\[95\]/Y vssd vccd output749/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_49_651 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1645 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[86\]_A input372/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_813 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_1910 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1689 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_805 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[40\] input66/X user_to_mprj_in_gates\[40\]/B vssd vccd user_to_mprj_in_gates\[40\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_52_849 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_buffers\[5\] user_wb_dat_gates\[5\]/Y vssd vccd output783/A vssd vccd
+ sky130_fd_sc_hd__clkinv_8
XFILLER_32_562 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_713 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[10\]_A input271/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_1747 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[90\]_B user_to_mprj_in_gates\[90\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA__332__A _332_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[2\] input54/X user_to_mprj_in_gates\[2\]/B vssd vccd user_to_mprj_in_gates\[2\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XANTENNA_user_to_mprj_in_ena_buf\[77\]_A input362/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1887 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_813 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[64\]_A_N _656_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1603 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1647 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[79\]_A_N _342_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__507__A _507_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_1273 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1836 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[81\]_B user_to_mprj_in_gates\[81\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_40_65 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[91\] _354_/Y mprj_logic_high_inst/HI[293] vssd vccd la_oenb_core[91]
+ vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_3_934 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[17\]_A_N _609_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input357_A la_iena_mprj[72] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_1618 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[4\] input332/X mprj_logic_high_inst/HI[334] vssd vccd user_to_mprj_in_gates\[4\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
Xla_buf\[99\] _563_/Y la_buf\[99\]/TE vssd vccd la_data_in_core[99] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input524_A mprj_adr_o_core[16] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[68\]_A input352/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_37 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xla_buf_enable\[114\] _377_/A la_buf_enable\[114\]/B vssd vccd la_buf\[114\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_34_805 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1160 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_838 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_551 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_427_ _427_/A vssd vccd _427_/Y vssd vccd sky130_fd_sc_hd__clkinv_8
XANTENNA__417__A _417_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_358_ _358_/A vssd vccd _358_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_31_2069 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_1313 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[10\] user_to_mprj_in_gates\[10\]/Y vssd vccd output638/A
+ vssd vccd sky130_fd_sc_hd__inv_6
XANTENNA_user_to_mprj_in_gates\[72\]_B user_to_mprj_in_gates\[72\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1379 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output743_A output743/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1821 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[88\] input118/X user_to_mprj_in_gates\[88\]/B vssd vccd user_to_mprj_in_gates\[88\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XANTENNA_user_to_mprj_in_ena_buf\[59\]_A input342/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1497 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1093 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput3 caravel_rstn vssd vccd input3/X vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_37_665 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_613 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_657 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1795 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1268 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_510 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1691 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1593 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[63\]_B user_to_mprj_in_gates\[63\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_47_2021 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[114\]_TE la_buf\[114\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_1397 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[50\] input333/X mprj_logic_high_inst/HI[380] vssd vccd user_to_mprj_in_gates\[50\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_mprj_adr_buf\[29\]_TE mprj_adr_buf\[29\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input105_A la_data_out_core[76] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[2\] user_to_mprj_in_gates\[2\]/Y vssd vccd output677/A vssd
+ vccd sky130_fd_sc_hd__clkinv_4
XFILLER_42_189 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_543 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_97 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input474_A la_oenb_mprj[62] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_587 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1677 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[14\] _478_/Y la_buf\[14\]/TE vssd vccd la_data_in_core[14] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_gates\[54\]_B user_to_mprj_in_gates\[54\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_input70_A la_data_out_core[44] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_753 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1139 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_797 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_919 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[61\]_TE mprj_logic_high_inst/HI[263] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
Xmprj_adr_buf\[7\] _407_/Y mprj_adr_buf\[7\]/TE vssd vccd mprj_adr_o_user[7] vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_4_1244 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_985 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[58\] user_to_mprj_in_gates\[58\]/Y vssd vccd output708/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_33_2109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output693_A output693/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_dat_buf\[8\]_A _440_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_2289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1831 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_896 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_gates\[16\] input557/X user_wb_ack_gate/B vssd vccd user_wb_dat_gates\[16\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_8
XFILLER_31_1154 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[45\]_B user_to_mprj_in_gates\[45\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_48_2341 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_wb_dat_buffers\[13\] user_wb_dat_gates\[13\]/Y vssd vccd output760/A vssd vccd
+ sky130_fd_sc_hd__clkinv_8
XFILLER_44_2249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1111 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__610__A _610_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_1971 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[114\] input20/X user_to_mprj_in_gates\[114\]/B vssd vccd user_to_mprj_in_gates\[114\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XANTENNA_user_to_mprj_in_buffers\[30\]_A user_to_mprj_in_gates\[30\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_38_974 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_473 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_602 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_107 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_118 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2209 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1390 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1953 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1997 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[97\]_A user_to_mprj_in_gates\[97\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[36\]_B user_to_mprj_in_gates\[36\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[120\]_B user_to_mprj_in_gates\[120\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_21_89 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_ena_buf\[98\] input385/X mprj_logic_high_inst/HI[428] vssd vccd user_to_mprj_in_gates\[98\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_la_buf\[70\]_A _534_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1437 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[84\]_TE mprj_logic_high_inst/HI[286] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[124\] _387_/Y mprj_logic_high_inst/HI[326] vssd vccd la_oenb_core[124]
+ vssd vccd sky130_fd_sc_hd__einvp_8
Xinput602 mprj_dat_o_core[28] vssd vccd _460_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
XANTENNA__520__A _520_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput613 mprj_dat_o_core[9] vssd vccd _441_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_48_705 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[54\] _646_/Y mprj_logic_high_inst/HI[256] vssd vccd la_oenb_core[54]
+ vssd vccd sky130_fd_sc_hd__einvp_8
Xinput624 user_irq_ena[0] vssd vccd input624/X vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_27_1768 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1069 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xla_buf_enable\[76\] _339_/A la_buf_enable\[76\]/B vssd vccd la_buf\[76\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_1_1417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input222_A la_data_out_mprj[66] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[21\]_A user_to_mprj_in_gates\[21\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_28_473 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_53 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_657 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_9 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_97 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input591_A mprj_dat_o_core[18] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_2142 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_856 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1029 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[124\]_A _588_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_1441 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_buffers\[88\]_A user_to_mprj_in_gates\[88\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[111\]_B user_to_mprj_in_gates\[111\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[27\]_B user_to_mprj_in_gates\[27\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_32_1485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_377 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[61\]_A _525_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf\[118\] _582_/Y la_buf\[118\]/TE vssd vccd la_data_in_core[118] vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_3_561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1783 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_buffers\[111\] user_to_mprj_in_gates\[111\]/Y vssd vccd output640/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA__430__A _430_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_705 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output706_A output706/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_1581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[12\]_A user_to_mprj_in_gates\[12\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_19_473 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_933 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_421 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_925 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[20\]_A input562/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[126\]_A user_to_mprj_in_gates\[126\]/Y vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_2097 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1839 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__605__A _605_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[115\]_A _579_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_1541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[79\]_A user_to_mprj_in_gates\[79\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[102\]_B user_to_mprj_in_gates\[102\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[18\]_B user_to_mprj_in_gates\[18\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_30_693 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xinput50 la_data_out_core[26] vssd vccd input50/X vssd vccd sky130_fd_sc_hd__buf_4
XANTENNA_la_buf\[52\]_A _516_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput61 la_data_out_core[36] vssd vccd input61/X vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput72 la_data_out_core[46] vssd vccd input72/X vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput83 la_data_out_core[56] vssd vccd input83/X vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput94 la_data_out_core[66] vssd vccd input94/X vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_48_2193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2013 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[70\]_B la_buf_enable\[70\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_2057 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__340__A _340_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_1919 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1621 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_793 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1127 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[11\]_A input552/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_2017 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[13\] input292/X mprj_logic_high_inst/HI[343] vssd vccd user_to_mprj_in_gates\[13\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_in_buffers\[117\]_A user_to_mprj_in_gates\[117\]/Y vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[106\]_A _570_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__515__A _515_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_1761 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[43\]_A _507_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1212 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input172_A la_data_out_mprj[20] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1245 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[61\]_B la_buf_enable\[61\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_1565 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput410 la_oenb_mprj[11] vssd vccd _603_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput421 la_oenb_mprj[14] vssd vccd _606_/A vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA_input437_A la_oenb_mprj[29] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput443 la_oenb_mprj[34] vssd vccd _626_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput454 la_oenb_mprj[44] vssd vccd _636_/A vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA_input33_A la_data_out_core[126] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput432 la_oenb_mprj[24] vssd vccd _616_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_48_557 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2073 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[81\] _545_/Y la_buf\[81\]/TE vssd vccd la_data_in_core[81] vssd vccd sky130_fd_sc_hd__einvp_8
Xinput465 la_oenb_mprj[54] vssd vccd _646_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput476 la_oenb_mprj[64] vssd vccd _656_/A vssd vccd sky130_fd_sc_hd__buf_2
Xinput487 la_oenb_mprj[74] vssd vccd _337_/A vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA_input604_A mprj_dat_o_core[2] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_1203 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_1765 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_771 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput498 la_oenb_mprj[84] vssd vccd _347_/A vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_28_281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_925 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[108\]_A user_to_mprj_in_gates\[108\]/Y vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_273 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_671 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__425__A _425_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output656_A output656/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[34\]_A _498_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_1894 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_2333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[52\]_B la_buf_enable\[52\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1621 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1329 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1591 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_881 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[70\] input99/X user_to_mprj_in_gates\[70\]/B vssd vccd user_to_mprj_in_gates\[70\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XANTENNA_user_to_mprj_in_ena_buf\[124\]_B mprj_logic_high_inst/HI[454] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_35_741 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_270 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1469 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_402 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_clk_buf _391_/Y mprj_clk_buf/TE vssd vccd user_clock vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_52_2337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__335__A _335_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1901 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1311 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[25\]_A _489_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1989 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1967 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1399 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[43\]_B la_buf_enable\[43\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_1429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1841 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[110\]_A _373_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_22 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[115\]_B mprj_logic_high_inst/HI[445] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_2_1589 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_460_ _460_/A vssd vccd _460_/Y vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_53_593 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_oen_buffers\[17\] _609_/Y mprj_logic_high_inst/HI[219] vssd vccd la_oenb_core[17]
+ vssd vccd sky130_fd_sc_hd__einvp_8
X_391_ _391_/A vssd vccd _391_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
Xla_buf_enable\[39\] _631_/A la_buf_enable\[39\]/B vssd vccd la_buf\[39\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_40_221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2270 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input387_A la_iena_mprj[9] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[16\]_A _480_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_1591 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_111 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input554_A mprj_dat_i_user[13] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[34\]_B la_buf_enable\[34\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_1605 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[3\]_A input321/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_2157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_833 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[101\]_A _364_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_877 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_321 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput251 la_data_out_mprj[92] vssd vccd _556_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput240 la_data_out_mprj[82] vssd vccd _546_/A vssd vccd sky130_fd_sc_hd__buf_2
Xinput262 la_iena_mprj[101] vssd vccd input262/X vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_48_365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[106\]_B mprj_logic_high_inst/HI[436] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xinput295 la_iena_mprj[16] vssd vccd input295/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput273 la_iena_mprj[111] vssd vccd input273/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput284 la_iena_mprj[121] vssd vccd input284/X vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_1_1044 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_593 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2001 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_589_ _589_/A vssd vccd _589_/Y vssd vccd sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_buffers\[40\] user_to_mprj_in_gates\[40\]/Y vssd vccd output689/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_la_buf\[10\]_TE la_buf\[10\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_1956 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output773_A output773/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_1907 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1377 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_483 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xoutput703 output703/A vssd vccd la_data_in_mprj[53] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput714 output714/A vssd vccd la_data_in_mprj[63] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput725 output725/A vssd vccd la_data_in_mprj[73] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput736 output736/A vssd vccd la_data_in_mprj[83] vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA_la_buf_enable\[25\]_B la_buf_enable\[25\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_1749 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xoutput769 output769/A vssd vccd mprj_dat_i_core[21] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput758 output758/A vssd vccd mprj_dat_i_core[11] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput747 output747/A vssd vccd la_data_in_mprj[93] vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_47_1727 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[105\]_A_N _368_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_2185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_321 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_516 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_571 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[119\]_TE mprj_logic_high_inst/HI[321] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_22_265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[94\]_A _357_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_939 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[16\]_B la_buf_enable\[16\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[80\] input366/X mprj_logic_high_inst/HI[410] vssd vccd user_to_mprj_in_gates\[80\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_28_2361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_659 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[95\]_B mprj_logic_high_inst/HI[425] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_46_825 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1579 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input135_A la_data_out_mprj[102] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_65 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_527 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_869 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
X_512_ _512_/A vssd vccd _512_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_input302_A la_iena_mprj[22] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[33\]_TE la_buf\[33\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_711 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_443_ _443_/A vssd vccd _443_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_41_541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[18\]_TE mprj_logic_high_inst/HI[220] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[44\] _508_/Y la_buf\[44\]/TE vssd vccd la_data_in_core[44] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_oen_buffers\[85\]_A _348_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_585 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
X_374_ _374_/A vssd vccd _374_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_31_2207 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_ena_buf\[116\] input278/X mprj_logic_high_inst/HI[446] vssd vccd
+ user_to_mprj_in_gates\[116\]/B vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_10_983 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1995 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_965 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_497 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1507 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[100\] _564_/Y la_buf\[100\]/TE vssd vccd la_data_in_core[100] vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_42_2325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[86\]_B mprj_logic_high_inst/HI[416] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_49_685 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_825 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[88\] user_to_mprj_in_gates\[88\]/Y vssd vccd output741/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_49_663 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_357 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[33\] input58/X user_to_mprj_in_gates\[33\]/B vssd vccd user_to_mprj_in_gates\[33\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_17_571 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_574 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_725 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[76\]_A _339_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_1753 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1797 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1005 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[10\]_B mprj_logic_high_inst/HI[340] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[1\]_TE la_buf\[1\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_1759 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1049 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_291 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__613__A _613_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_1513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[3\]_A input575/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_1101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[77\]_B mprj_logic_high_inst/HI[407] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_5_1905 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1719 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_825 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[56\]_TE la_buf\[56\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_1877 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_1189 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1899 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_869 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[3\]_A input65/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[3\]_A_N _595_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_1659 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[67\]_A _330_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_1973 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1848 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1285 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_279 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__523__A _523_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_77 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_946 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[84\] _347_/Y mprj_logic_high_inst/HI[286] vssd vccd la_oenb_core[84]
+ vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_2_401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input252_A la_data_out_mprj[93] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_456 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[68\]_B mprj_logic_high_inst/HI[398] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_input517_A mprj_adr_o_core[0] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_1459 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[107\] _370_/A la_buf_enable\[107\]/B vssd vccd la_buf\[107\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_4_1437 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1027 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_426_ _426_/A vssd vccd _426_/Y vssd vccd sky130_fd_sc_hd__inv_12
XANTENNA_user_to_mprj_oen_buffers\[58\]_A _650_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_357_ _357_/A vssd vccd _357_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_35_1483 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__433__A _433_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_773 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1833 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output736_A output736/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_1315 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_1877 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[79\]_TE la_buf\[79\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_990 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[59\]_B mprj_logic_high_inst/HI[389] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_9_1359 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xinput4 la_data_out_core[0] vssd vccd input4/X vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_52_625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__608__A _608_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_669 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[49\]_A _641_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_522 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__343__A _343_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_2033 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1321 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_1229 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_1663 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[28\]_TE mprj_dat_buf\[28\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[43\] input325/X mprj_logic_high_inst/HI[373] vssd vccd user_to_mprj_in_gates\[43\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_27_165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__518__A _518_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[7\]_TE mprj_logic_high_inst/HI[209] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_23_393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[21\] _613_/A la_buf_enable\[21\]/B vssd vccd la_buf\[21\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_11_555 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_1071 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1093 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1689 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input467_A la_oenb_mprj[56] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input63_A la_data_out_core[38] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_765 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_264 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_611 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1256 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_677 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_ack_buffer user_wb_ack_gate/Y vssd vccd output755/A vssd vccd sky130_fd_sc_hd__clkinv_8
XFILLER_33_113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__428__A _428_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_1501 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_371 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output686_A output686/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_409_ _409_/A vssd vccd _409_/Y vssd vccd sky130_fd_sc_hd__inv_8
XFILLER_15_1843 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1707 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1887 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[63\]_A_N _655_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1166 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_mprj_adr_buf\[27\]_A _427_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[78\]_A_N _341_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_1156 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1803 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1009 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_sel_buf\[2\]_TE mprj_sel_buf\[2\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_1983 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1273 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[107\] input12/X user_to_mprj_in_gates\[107\]/B vssd vccd user_to_mprj_in_gates\[107\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_52_433 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__338__A _338_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XPHY_119 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_108 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[16\]_A_N _608_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[4\]_A _596_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_1206 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_385 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_57 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_mprj_adr_buf\[18\]_A _418_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[117\] _380_/Y mprj_logic_high_inst/HI[319] vssd vccd la_oenb_core[117]
+ vssd vccd sky130_fd_sc_hd__einvp_8
Xinput603 mprj_dat_o_core[29] vssd vccd _461_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_25_2161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_717 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput614 mprj_iena_wb vssd vccd input614/X vssd vccd sky130_fd_sc_hd__buf_2
Xinput625 user_irq_ena[1] vssd vccd input625/X vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_47_205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[47\] _639_/Y mprj_logic_high_inst/HI[249] vssd vccd la_oenb_core[47]
+ vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[69\] _332_/A la_buf_enable\[69\]/B vssd vccd la_buf\[69\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_46_65 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input215_A la_data_out_mprj[5] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_1821 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_813 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input584_A mprj_dat_o_core[11] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_363 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_868 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_389 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1497 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_irq_buffers\[1\]_A user_irq_gates\[1\]/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_573 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_717 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[104\] user_to_mprj_in_gates\[104\]/Y vssd vccd output632/A
+ vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_43_1593 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[70\] user_to_mprj_in_gates\[70\]/Y vssd vccd output722/A
+ vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_53_219 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_433 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_945 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_wb_dat_gates\[20\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_937 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_628 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_680 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[104\]_TE la_buf\[104\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_1807 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_1949 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[19\]_TE mprj_adr_buf\[19\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_1553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput40 la_data_out_core[17] vssd vccd input40/X vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_11_1504 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1597 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput73 la_data_out_core[47] vssd vccd input73/X vssd vccd sky130_fd_sc_hd__buf_4
Xinput51 la_data_out_core[27] vssd vccd input51/X vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput62 la_data_out_core[37] vssd vccd input62/X vssd vccd sky130_fd_sc_hd__clkbuf_4
XANTENNA__621__A _621_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput84 la_data_out_core[57] vssd vccd input84/X vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput95 la_data_out_core[67] vssd vccd input95/X vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_44_2025 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[3\]_TE mprj_adr_buf\[3\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_2069 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[3\] _435_/Y mprj_dat_buf\[3\]/TE vssd vccd mprj_dat_o_user[3] vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_45_709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1081 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_wb_dat_gates\[11\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_1139 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_469 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[51\]_TE mprj_logic_high_inst/HI[253] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_1773 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_304 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_1003 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_849 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_1224 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_1257 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input165_A la_data_out_mprj[14] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__531__A _531_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_dat_buf\[7\]_TE mprj_dat_buf\[7\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput411 la_oenb_mprj[120] vssd vccd _383_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput400 la_oenb_mprj[110] vssd vccd _373_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_7_1649 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_2041 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_1577 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_525 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xinput455 la_oenb_mprj[45] vssd vccd _637_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput444 la_oenb_mprj[35] vssd vccd _627_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput422 la_oenb_mprj[15] vssd vccd _607_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput433 la_oenb_mprj[25] vssd vccd _617_/A vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA_input332_A la_iena_mprj[4] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1733 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput477 la_oenb_mprj[65] vssd vccd _657_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput466 la_oenb_mprj[55] vssd vccd _647_/A vssd vccd sky130_fd_sc_hd__buf_2
Xinput488 la_oenb_mprj[75] vssd vccd _338_/A vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA_input26_A la_data_out_core[11] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_2085 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_219 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xinput499 la_oenb_mprj[85] vssd vccd _348_/A vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_40_1777 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_422 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[74\] _538_/Y la_buf\[74\]/TE vssd vccd la_data_in_core[74] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf\[127\]_TE la_buf\[127\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_1640 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_981 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1971 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_683 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_676 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output649_A output649/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__441__A _441_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_893 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_2209 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[63\] input91/X user_to_mprj_in_gates\[63\]/B vssd vccd user_to_mprj_in_gates\[63\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_50_701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[74\]_TE mprj_logic_high_inst/HI[276] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_753 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_285 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_414 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_609 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__616__A _616_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_1003 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_mprj_adr_buf\[3\]_A _403_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1913 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1334 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1979 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__351__A _351_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_1903 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_buffers\[29\]_A user_wb_dat_gates\[29\]/Y vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XFILLER_2_2225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_517 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_34 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_390_ _390_/A vssd vccd _390_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_40_233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__526__A _526_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_480 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_613 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_1169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input282_A la_iena_mprj[11] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_123 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_1021 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1065 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input547_A mprj_adr_o_core[8] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_189 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[3\]_B mprj_logic_high_inst/HI[333] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_1_874 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput252 la_data_out_mprj[93] vssd vccd _557_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput230 la_data_out_mprj[73] vssd vccd _537_/A vssd vccd sky130_fd_sc_hd__buf_2
Xinput241 la_data_out_mprj[83] vssd vccd _547_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput263 la_iena_mprj[102] vssd vccd input263/X vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_48_377 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[97\]_TE mprj_logic_high_inst/HI[299] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
Xinput296 la_iena_mprj[17] vssd vccd input296/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput274 la_iena_mprj[112] vssd vccd input274/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput285 la_iena_mprj[122] vssd vccd input285/X vssd vccd sky130_fd_sc_hd__clkbuf_1
X_657_ _657_/A vssd vccd _657_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_32_701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_588_ _588_/A vssd vccd _588_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_38_2193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2013 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__436__A _436_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[33\] user_to_mprj_in_gates\[33\]/Y vssd vccd output681/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_output766_A output766/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_1681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1389 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_495 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xoutput704 output704/A vssd vccd la_data_in_mprj[54] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput715 output715/A vssd vccd la_data_in_mprj[64] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput726 output726/A vssd vccd la_data_in_mprj[74] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput759 output759/A vssd vccd mprj_dat_i_core[12] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput737 output737/A vssd vccd la_data_in_mprj[84] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput748 output748/A vssd vccd la_data_in_mprj[94] vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_28_1149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2017 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_1305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[124\]_B la_buf_enable\[124\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_528 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_2280 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1201 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1245 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_583 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__346__A _346_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_907 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[93\]_A input124/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1721 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_ena_buf\[73\] input358/X mprj_logic_high_inst/HI[403] vssd vccd user_to_mprj_in_gates\[73\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_4_1608 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[115\]_B la_buf_enable\[115\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_2066 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1861 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_837 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_539 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1490 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input128_A la_data_out_core[97] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_358 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_511_ _511_/A vssd vccd _511_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
Xla_buf_enable\[51\] _643_/A la_buf_enable\[51\]/B vssd vccd la_buf\[51\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_2_1354 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_723 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_442_ _442_/A vssd vccd _442_/Y vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_35_1621 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input497_A la_oenb_mprj[83] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_373_ _373_/A vssd vccd _373_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_41_553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[37\] _501_/Y la_buf\[37\]/TE vssd vccd la_data_in_core[37] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_gates\[84\]_A input114/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_buffers\[6\]_A user_wb_dat_gates\[6\]/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input93_A la_data_out_core[65] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_951 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[109\] input270/X mprj_logic_high_inst/HI[439] vssd vccd
+ user_to_mprj_in_gates\[109\]/B vssd vccd sky130_fd_sc_hd__and2_1
Xuser_wb_dat_gates\[9\] input581/X user_wb_ack_gate/B vssd vccd user_wb_dat_gates\[9\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_4
XFILLER_10_995 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_977 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_1425 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1519 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1761 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_2337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[9\]_A _473_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[106\]_B la_buf_enable\[106\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_697 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1841 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[26\] input50/X user_to_mprj_in_gates\[26\]/B vssd vccd user_to_mprj_in_gates\[26\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_20_737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[75\]_A input104/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1175 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1017 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1525 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_81 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[3\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_1007 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_2353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1641 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_837 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1652 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[3\]_B user_to_mprj_in_gates\[3\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_36_881 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[66\]_A input94/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_1242 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_1985 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_2230 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_218 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[77\] _340_/Y mprj_logic_high_inst/HI[279] vssd vccd la_oenb_core[77]
+ vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[99\] _362_/A la_buf_enable\[99\]/B vssd vccd la_buf\[99\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_28_2181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xmprj_dat_buf\[25\] _457_/Y mprj_dat_buf\[25\]/TE vssd vccd mprj_dat_o_user[25] vssd
+ vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input245_A la_data_out_mprj[87] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_601 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input412_A la_oenb_mprj[121] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_18_303 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_645 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_358 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1705 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_1716 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_425_ _425_/A vssd vccd _425_/Y vssd vccd sky130_fd_sc_hd__inv_12
XFILLER_41_361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[104\]_A_N _367_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_356_ _356_/A vssd vccd _356_/Y vssd vccd sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_gates\[57\]_A input84/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1495 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[20\] _420_/Y mprj_adr_buf\[20\]/TE vssd vccd mprj_adr_o_user[20] vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_48_1801 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_785 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[119\]_A_N _382_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1845 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1889 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1266 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output729_A output729/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output631_A output631/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[109\]_TE mprj_logic_high_inst/HI[311] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_1411 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2189 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1422 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_461 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_100 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput5 la_data_out_core[100] vssd vccd input5/X vssd vccd sky130_fd_sc_hd__clkbuf_4
XANTENNA_user_to_mprj_in_buffers\[7\]_A user_to_mprj_in_gates\[7\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_36_177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_637 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1551 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_1671 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[48\]_A input74/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__624__A _624_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[5\] _597_/A la_buf_enable\[5\]/B vssd vccd la_buf\[5\]/TE vssd vccd
+ sky130_fd_sc_hd__and2b_1
XFILLER_14_1579 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2045 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[23\]_TE la_buf\[23\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_1208 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_1653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_601 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1675 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_645 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[36\] input317/X mprj_logic_high_inst/HI[366] vssd vccd user_to_mprj_in_gates\[36\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_42_125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_2325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[14\] _606_/A la_buf_enable\[14\]/B vssd vccd la_buf\[14\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XANTENNA_user_to_mprj_in_gates\[123\]_A input30/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[39\]_A input64/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__534__A _534_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input195_A la_data_out_mprj[41] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_1083 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input362_A la_iena_mprj[77] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_210 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_243 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input56_A la_data_out_core[31] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_777 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1371 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_645 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_626 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_689 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1535 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_408_ _408_/A vssd vccd _408_/Y vssd vccd sky130_fd_sc_hd__clkinv_16
XFILLER_14_383 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1811 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output679_A output679/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[114\]_A input20/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__444__A _444_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_1855 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_339_ _339_/A vssd vccd _339_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_31_1134 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1899 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1719 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[46\]_TE la_buf\[46\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_1877 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1189 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[93\] input124/X user_to_mprj_in_gates\[93\]/B vssd vccd user_to_mprj_in_gates\[93\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_29_1041 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_1653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[2\]_A_N _594_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_1168 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1995 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1815 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1859 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__619__A _619_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_1285 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_626 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_497 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XPHY_109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[105\]_A input10/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__354__A _354_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_397 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_69 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1218 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput604 mprj_dat_o_core[2] vssd vccd _434_/A vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_5_2212 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xinput615 mprj_sel_o_core[0] vssd vccd _396_/A vssd vccd sky130_fd_sc_hd__dlymetal6s2s_1
Xinput626 user_irq_ena[2] vssd vccd input626/X vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_48_729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_217 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_921 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_1937 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1555 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__529__A _529_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_2289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_77 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_968 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input208_A la_data_out_mprj[53] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input110_A la_data_out_core[80] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_1833 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1811 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1877 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_629 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[69\]_TE la_buf\[69\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_331 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_825 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input577_A mprj_dat_i_user[5] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_1421 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_585 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_2309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__439__A _439_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_1942 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[63\] user_to_mprj_in_gates\[63\]/Y vssd vccd output714/A
+ vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_21_117 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_692 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1521 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_gates\[21\] input563/X user_wb_ack_gate/B vssd vccd user_wb_dat_gates\[21\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_2
XFILLER_15_1663 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput30 la_data_out_core[123] vssd vccd input30/X vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput41 la_data_out_core[18] vssd vccd input41/X vssd vccd sky130_fd_sc_hd__buf_4
XANTENNA_mprj_dat_buf\[18\]_TE mprj_dat_buf\[18\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput52 la_data_out_core[28] vssd vccd input52/X vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput63 la_data_out_core[38] vssd vccd input63/X vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_50_1565 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xinput85 la_data_out_core[58] vssd vccd input85/X vssd vccd sky130_fd_sc_hd__buf_4
Xinput74 la_data_out_core[48] vssd vccd input74/X vssd vccd sky130_fd_sc_hd__buf_4
XANTENNA_la_buf_enable\[3\]_B la_buf_enable\[3\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput96 la_data_out_core[68] vssd vccd input96/X vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_44_2037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[127\]_A input290/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_1781 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_209 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__349__A _349_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_1717 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_286 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_489 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_651 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_684 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1785 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1606 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput401 la_oenb_mprj[111] vssd vccd _374_/A vssd vccd sky130_fd_sc_hd__buf_4
Xla_buf_enable\[81\] _344_/A la_buf_enable\[81\]/B vssd vccd la_buf\[81\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XANTENNA_input158_A la_data_out_mprj[123] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput412 la_oenb_mprj[121] vssd vccd _384_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_27_1589 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput445 la_oenb_mprj[36] vssd vccd _628_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput434 la_oenb_mprj[26] vssd vccd _618_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput423 la_oenb_mprj[16] vssd vccd _608_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
XANTENNA_user_to_mprj_in_ena_buf\[118\]_A input280/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput478 la_oenb_mprj[66] vssd vccd _329_/A vssd vccd sky130_fd_sc_hd__buf_4
Xinput456 la_oenb_mprj[46] vssd vccd _638_/A vssd vccd sky130_fd_sc_hd__buf_4
Xinput467 la_oenb_mprj[56] vssd vccd _648_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
XANTENNA_input325_A la_iena_mprj[43] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_1745 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[62\]_A_N _654_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input19_A la_data_out_core[113] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput489 la_oenb_mprj[76] vssd vccd _339_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_16_434 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[67\] _531_/Y la_buf\[67\]/TE vssd vccd la_data_in_core[67] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf_enable\[77\]_A_N _340_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_611 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_993 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1983 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1803 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_695 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_655 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1273 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_688 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[123\] _587_/Y la_buf\[123\]/TE vssd vccd la_data_in_core[123] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf_enable\[15\]_A_N _607_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1105 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output711_A output711/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[109\]_A input270/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_1149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_1943 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1921 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[56\] input83/X user_to_mprj_in_gates\[56\]/B vssd vccd user_to_mprj_in_gates\[56\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_35_721 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_713 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_757 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[40\]_A input322/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1173 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_2030 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__632__A _632_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_1409 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1821 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1915 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1959 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2248 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_46 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_529 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[31\]_A input312/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_245 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_492 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__542__A _542_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input275_A la_iena_mprj[113] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_135 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_1033 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1077 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_853 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input442_A la_oenb_mprj[33] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[98\]_A input385/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_1425 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xinput220 la_data_out_mprj[64] vssd vccd _528_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_7_1469 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput242 la_data_out_mprj[84] vssd vccd _548_/A vssd vccd sky130_fd_sc_hd__buf_4
Xinput231 la_data_out_mprj[74] vssd vccd _538_/A vssd vccd sky130_fd_sc_hd__buf_2
Xinput253 la_data_out_mprj[94] vssd vccd _558_/A vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_48_345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput297 la_iena_mprj[18] vssd vccd input297/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput264 la_iena_mprj[103] vssd vccd input264/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput275 la_iena_mprj[113] vssd vccd input275/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput286 la_iena_mprj[123] vssd vccd input286/X vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_1_1013 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_389 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2298 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1597 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_656_ _656_/A vssd vccd _656_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_16_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_587_ _587_/A vssd vccd _587_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_34_2025 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_757 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[22\]_A input302/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_1493 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_779 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[26\] user_to_mprj_in_gates\[26\]/Y vssd vccd output673/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_output661_A output661/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_1693 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output759_A output759/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__452__A _452_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput705 output705/A vssd vccd la_data_in_mprj[55] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput716 output716/A vssd vccd la_data_in_mprj[65] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput727 output727/A vssd vccd la_data_in_mprj[75] vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_28_1117 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xoutput738 output738/A vssd vccd la_data_in_mprj[85] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput749 output749/A vssd vccd la_data_in_mprj[95] vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA_user_to_mprj_in_ena_buf\[89\]_A input375/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_2007 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_2029 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[41\]_TE mprj_logic_high_inst/HI[243] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_1213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__627__A _627_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_1257 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_595 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[13\]_A input292/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[93\]_B user_to_mprj_in_gates\[93\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_22_289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1733 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__362__A _362_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_1143 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[117\]_TE la_buf\[117\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[66\] input350/X mprj_logic_high_inst/HI[396] vssd vccd user_to_mprj_in_gates\[66\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_6_2181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1322 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_1873 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_849 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_510_ _510_/A vssd vccd _510_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_45_337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1399 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_441_ _441_/A vssd vccd _441_/Y vssd vccd sky130_fd_sc_hd__clkinv_4
Xuser_to_mprj_oen_buffers\[4\] _596_/Y mprj_logic_high_inst/HI[206] vssd vccd la_oenb_core[4]
+ vssd vccd sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[22\] _614_/Y mprj_logic_high_inst/HI[224] vssd vccd la_oenb_core[22]
+ vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[44\] _636_/A la_buf_enable\[44\]/B vssd vccd la_buf\[44\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XANTENNA__537__A _537_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_irq_ena_buf\[0\]_A input624/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_381 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
X_372_ _372_/A vssd vccd _372_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_13_289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[84\]_B user_to_mprj_in_gates\[84\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_input392_A la_oenb_mprj[103] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input86_A la_data_out_core[59] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_2305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1437 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[64\]_TE mprj_logic_high_inst/HI[266] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_1233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_329 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_639_ _639_/A vssd vccd _639_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA__447__A _447_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_18_1853 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[19\] input42/X user_to_mprj_in_gates\[19\]/B vssd vccd user_to_mprj_in_gates\[19\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_2
XANTENNA_user_to_mprj_in_gates\[75\]_B user_to_mprj_in_gates\[75\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1187 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1029 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_wb_dat_buffers\[29\] user_wb_dat_gates\[29\]/Y vssd vccd output777/A vssd vccd
+ sky130_fd_sc_hd__clkinv_8
XFILLER_47_1537 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1019 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_93 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_buffers\[60\]_A user_to_mprj_in_gates\[60\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_41_1169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1664 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1675 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__357__A _357_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_841 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_893 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1065 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_727 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[66\]_B user_to_mprj_in_gates\[66\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_30_2242 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[87\]_TE mprj_logic_high_inst/HI[289] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_1481 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2079 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xmprj_dat_buf\[18\] _450_/Y mprj_dat_buf\[18\]/TE vssd vccd mprj_dat_o_user[18] vssd
+ vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input238_A la_data_out_mprj[80] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[51\]_A user_to_mprj_in_gates\[51\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_input140_A la_data_out_mprj[107] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_613 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_657 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input405_A la_oenb_mprj[115] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_424_ _424_/A vssd vccd _424_/Y vssd vccd sky130_fd_sc_hd__clkinv_16
XFILLER_33_329 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1728 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[121\] input284/X mprj_logic_high_inst/HI[451] vssd vccd
+ user_to_mprj_in_gates\[121\]/B vssd vccd sky130_fd_sc_hd__and2_1
X_355_ _355_/A vssd vccd _355_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_50_1906 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[57\]_B user_to_mprj_in_gates\[57\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[91\]_A _555_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_797 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1813 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xmprj_adr_buf\[13\] _413_/Y mprj_adr_buf\[13\]/TE vssd vccd mprj_adr_o_user[13] vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_48_1857 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[127\] user_to_mprj_in_gates\[127\]/Y vssd vccd output657/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_46_2293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[93\] user_to_mprj_in_gates\[93\]/Y vssd vccd output747/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_29_1278 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_2157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[42\]_A user_to_mprj_in_gates\[42\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_49_473 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput6 la_data_out_core[101] vssd vccd input6/X vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_36_112 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_841 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_buffers\[3\] user_wb_dat_gates\[3\]/Y vssd vccd output781/A vssd vccd
+ sky130_fd_sc_hd__clkinv_8
XFILLER_36_189 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[48\]_B user_to_mprj_in_gates\[48\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_18_1683 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[82\]_A _546_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1861 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1883 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2057 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__640__A _640_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[0\] input4/X user_to_mprj_in_gates\[0\]/B vssd vccd user_to_mprj_in_gates\[0\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XANTENNA_user_to_mprj_in_buffers\[33\]_A user_to_mprj_in_gates\[33\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_28_613 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_69 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_657 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_635 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_307 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1450 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_ena_buf\[29\] input309/X mprj_logic_high_inst/HI[359] vssd vccd user_to_mprj_in_gates\[29\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_35_57 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_1761 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_2337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[123\]_B user_to_mprj_in_gates\[123\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[39\]_B user_to_mprj_in_gates\[39\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_7_517 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[73\]_A _537_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_2061 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input188_A la_data_out_mprj[35] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[91\]_B la_buf_enable\[91\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__550__A _550_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input355_A la_iena_mprj[70] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input49_A la_data_out_core[25] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input522_A mprj_adr_o_core[14] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[24\]_A user_to_mprj_in_gates\[24\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_8_1383 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[2\] input310/X mprj_logic_high_inst/HI[332] vssd vccd user_to_mprj_in_gates\[2\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
Xla_buf\[97\] _561_/Y la_buf\[97\]/TE vssd vccd la_data_in_core[97] vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[112\] _375_/A la_buf_enable\[112\]/B vssd vccd la_buf\[112\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_46_421 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_638 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_90 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_1569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1547 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[127\]_A _591_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_407_ _407_/A vssd vccd _407_/Y vssd vccd sky130_fd_sc_hd__inv_8
XFILLER_41_181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_338_ _338_/A vssd vccd _338_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_user_to_mprj_in_gates\[114\]_B user_to_mprj_in_gates\[114\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_15_1823 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_693 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1747 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1260 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[64\]_A _528_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_1867 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output741_A output741/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[82\]_B la_buf_enable\[82\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1621 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__460__A _460_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1665 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[86\] input116/X user_to_mprj_in_gates\[86\]/B vssd vccd user_to_mprj_in_gates\[86\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_22_1827 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[15\]_A user_to_mprj_in_gates\[15\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_49_281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_72 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_925 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2357 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_wb_dat_gates\[23\]_A input565/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_638 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_969 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[118\]_A _582_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__635__A _635_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[105\]_B user_to_mprj_in_gates\[105\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_20_321 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[55\]_A _519_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_354 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_376 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[73\]_B la_buf_enable\[73\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__370__A _370_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput616 mprj_sel_o_core[1] vssd vccd _397_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput605 mprj_dat_o_core[30] vssd vccd _462_/A vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_25_2196 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[103\]_A_N _366_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_1949 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_421 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_925 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[14\]_A input555/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[118\]_A_N _381_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input103_A la_data_out_core[74] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_1845 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[0\] user_to_mprj_in_gates\[0\]/Y vssd vccd output627/A vssd
+ vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_la_buf\[109\]_A _573_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__545__A _545_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_490 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1889 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[46\]_A _510_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input472_A la_oenb_mprj[60] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf\[12\] _476_/Y la_buf\[12\]/TE vssd vccd la_data_in_core[12] vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf\[8\] _472_/Y la_buf\[8\]/TE vssd vccd la_data_in_core[8] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf_enable\[64\]_B la_buf_enable\[64\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1941 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1805 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1849 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[5\] _405_/Y mprj_adr_buf\[5\]/TE vssd vccd mprj_adr_o_user[5] vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_47_741 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_421 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_785 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[13\]_TE la_buf\[13\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[56\] user_to_mprj_in_gates\[56\]/Y vssd vccd output706/A
+ vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_37_1311 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output691_A output691/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output789_A output789/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__455__A _455_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[37\]_A _501_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_1675 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1533 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_wb_dat_gates\[14\] input555/X user_wb_ack_gate/B vssd vccd user_wb_dat_gates\[14\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_4
Xinput20 la_data_out_core[114] vssd vccd input20/X vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput31 la_data_out_core[124] vssd vccd input31/X vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_11_1539 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput42 la_data_out_core[19] vssd vccd input42/X vssd vccd sky130_fd_sc_hd__buf_4
XANTENNA_la_buf_enable\[55\]_B la_buf_enable\[55\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput53 la_data_out_core[29] vssd vccd input53/X vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput64 la_data_out_core[39] vssd vccd input64/X vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_48_2141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xinput97 la_data_out_core[69] vssd vccd input97/X vssd vccd sky130_fd_sc_hd__buf_4
Xinput86 la_data_out_core[59] vssd vccd input86/X vssd vccd sky130_fd_sc_hd__buf_4
Xinput75 la_data_out_core[49] vssd vccd input75/X vssd vccd sky130_fd_sc_hd__buf_4
Xuser_wb_dat_buffers\[11\] user_wb_dat_gates\[11\]/Y vssd vccd output758/A vssd vccd
+ sky130_fd_sc_hd__clkinv_8
XANTENNA_user_to_mprj_oen_buffers\[122\]_A _385_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_1832 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[127\]_B mprj_logic_high_inst/HI[457] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_42_1061 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1635 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[112\] input18/X user_to_mprj_in_gates\[112\]/B vssd vccd user_to_mprj_in_gates\[112\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_26_1793 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_722 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__365__A _365_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[28\]_A _492_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_641 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_696 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[46\]_B la_buf_enable\[46\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[96\] input383/X mprj_logic_high_inst/HI[426] vssd vccd user_to_mprj_in_gates\[96\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
Xuser_to_mprj_oen_buffers\[122\] _385_/Y mprj_logic_high_inst/HI[324] vssd vccd la_oenb_core[122]
+ vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_oen_buffers\[113\]_A _376_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xmprj_sel_buf\[3\] _399_/Y mprj_sel_buf\[3\]/TE vssd vccd mprj_sel_o_user[3] vssd
+ vccd sky130_fd_sc_hd__einvp_8
Xinput402 la_oenb_mprj[112] vssd vccd _375_/A vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_7_1629 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[52\] _644_/Y mprj_logic_high_inst/HI[254] vssd vccd la_oenb_core[52]
+ vssd vccd sky130_fd_sc_hd__einvp_8
Xinput446 la_oenb_mprj[37] vssd vccd _629_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput424 la_oenb_mprj[17] vssd vccd _609_/A vssd vccd sky130_fd_sc_hd__buf_2
Xinput435 la_oenb_mprj[27] vssd vccd _619_/A vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA_user_to_mprj_in_ena_buf\[118\]_B mprj_logic_high_inst/HI[448] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xinput413 la_oenb_mprj[122] vssd vccd _385_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput479 la_oenb_mprj[67] vssd vccd _330_/A vssd vccd sky130_fd_sc_hd__buf_4
Xinput457 la_oenb_mprj[47] vssd vccd _639_/A vssd vccd sky130_fd_sc_hd__buf_4
Xinput468 la_oenb_mprj[57] vssd vccd _649_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xla_buf_enable\[74\] _337_/A la_buf_enable\[74\]/B vssd vccd la_buf\[74\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XANTENNA_input318_A la_iena_mprj[37] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input220_A la_data_out_mprj[64] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[36\]_TE la_buf\[36\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_1757 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_785 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_405 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[1\]_A_N _593_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[19\]_A _483_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_1951 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1995 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_667 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_1815 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[37\]_B la_buf_enable\[37\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_1285 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1859 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[116\] _580_/Y la_buf\[116\]/TE vssd vccd la_data_in_core[116] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_ena_buf\[6\]_A input354/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[104\]_A _367_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1602 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_1613 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[109\]_B mprj_logic_high_inst/HI[439] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_clk2_buf_A _392_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_1117 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_538 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output704_A output704/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_1933 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_1381 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1955 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1999 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_2129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[49\] input75/X user_to_mprj_in_gates\[49\]/B vssd vccd user_to_mprj_in_gates\[49\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_50_725 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[40\]_B mprj_logic_high_inst/HI[370] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_50_769 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[4\]_TE la_buf\[4\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_1341 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[28\]_B la_buf_enable\[28\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_1385 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[30\]_A _622_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_1833 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_1719 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1877 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[59\]_TE la_buf\[59\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_2238 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1504 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1548 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_585 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[97\]_A _360_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_1973 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[11\] input282/X mprj_logic_high_inst/HI[341] vssd vccd user_to_mprj_in_gates\[11\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_43_57 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[31\]_B mprj_logic_high_inst/HI[361] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[19\]_B la_buf_enable\[19\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1001 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input170_A la_data_out_mprj[19] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1045 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2011 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_29 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input268_A la_iena_mprj[107] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[21\]_A _613_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1089 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1933 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2055 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[98\]_B mprj_logic_high_inst/HI[428] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xinput210 la_data_out_mprj[55] vssd vccd _519_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
XANTENNA_input435_A la_oenb_mprj[27] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput221 la_data_out_mprj[65] vssd vccd _529_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput232 la_data_out_mprj[75] vssd vccd _539_/A vssd vccd sky130_fd_sc_hd__buf_2
Xinput254 la_data_out_mprj[95] vssd vccd _559_/A vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA_input31_A la_data_out_core[124] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput243 la_data_out_mprj[85] vssd vccd _549_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_48_357 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input602_A mprj_dat_o_core[28] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput265 la_iena_mprj[104] vssd vccd input265/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput276 la_iena_mprj[114] vssd vccd input276/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput287 la_iena_mprj[124] vssd vccd input287/X vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_40_1565 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_711 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput298 la_iena_mprj[19] vssd vccd input298/X vssd vccd sky130_fd_sc_hd__clkbuf_1
X_655_ _655_/A vssd vccd _655_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_16_265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[88\]_A _351_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_586_ _586_/A vssd vccd _586_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_34_2037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_910 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_257 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[22\]_B mprj_logic_high_inst/HI[352] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_40_780 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_471 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1661 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1071 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[19\] user_to_mprj_in_gates\[19\]/Y vssd vccd output665/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_output654_A output654/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_1093 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xoutput706 output706/A vssd vccd la_data_in_mprj[56] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput717 output717/A vssd vccd la_data_in_mprj[66] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput728 output728/A vssd vccd la_data_in_mprj[76] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput739 output739/A vssd vccd la_data_in_mprj[86] vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA_user_to_mprj_oen_buffers\[12\]_A _604_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_2133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[89\]_B mprj_logic_high_inst/HI[419] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_23_1730 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[79\]_A _342_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_1225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_533 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[13\]_B mprj_logic_high_inst/HI[343] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA__643__A _643_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1881 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_1745 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1778 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[61\]_A_N _653_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[6\]_A input578/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_1199 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_1735 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[76\]_A_N _339_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_1685 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_79 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_2193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1841 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_ena_buf\[59\] input342/X mprj_logic_high_inst/HI[389] vssd vccd user_to_mprj_in_gates\[59\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_in_gates\[6\]_A input98/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_1312 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1885 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_irq_ena_buf\[0\]_B user_irq_ena_buf\[0\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_440_ _440_/A vssd vccd _440_/Y vssd vccd sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[15\] _607_/Y mprj_logic_high_inst/HI[217] vssd vccd la_oenb_core[15]
+ vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[37\] _629_/A la_buf_enable\[37\]/B vssd vccd la_buf\[37\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
X_371_ _371_/A vssd vccd _371_/Y vssd vccd sky130_fd_sc_hd__inv_2
XANTENNA_la_buf_enable\[14\]_A_N _606_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__553__A _553_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input385_A la_iena_mprj[98] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_1921 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_1943 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[29\]_A_N _621_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input79_A la_data_out_core[52] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input552_A mprj_dat_i_user[11] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_1449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1201 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1245 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_638_ _638_/A vssd vccd _638_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_32_533 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_511 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_569_ _569_/A vssd vccd _569_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_output771_A output771/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__463__A _463_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1199 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_1549 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_809 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1582 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__638__A _638_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_1022 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1607 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_853 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[30\]_A _462_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_1077 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_897 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_739 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__373__A _373_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1597 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_448 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input133_A la_data_out_mprj[100] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_1693 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__548__A _548_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_669 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input300_A la_iena_mprj[20] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_423_ _423_/A vssd vccd _423_/Y vssd vccd sky130_fd_sc_hd__inv_8
XFILLER_35_2121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_mprj_dat_buf\[21\]_A _453_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf\[42\] _506_/Y la_buf\[42\]/TE vssd vccd la_data_in_core[42] vssd vccd sky130_fd_sc_hd__einvp_8
X_354_ _354_/A vssd vccd _354_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_41_385 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1918 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[114\] input276/X mprj_logic_high_inst/HI[444] vssd vccd
+ user_to_mprj_in_gates\[114\]/B vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_6_721 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[31\]_TE mprj_logic_high_inst/HI[233] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_783 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_242 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1869 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1307 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_441 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[86\] user_to_mprj_in_gates\[86\]/Y vssd vccd output739/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
Xinput7 la_data_out_core[102] vssd vccd input7/X vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_36_124 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__458__A _458_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[31\] input56/X user_to_mprj_in_gates\[31\]/B vssd vccd user_to_mprj_in_gates\[31\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XANTENNA_la_buf\[107\]_TE la_buf\[107\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_831 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1217 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_853 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[12\]_A _444_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_2232 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_897 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1564 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1895 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_mprj_adr_buf\[6\]_TE mprj_adr_buf\[6\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1873 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_1313 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_2069 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1705 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1749 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__368__A _368_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_669 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_319 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[7\]_A _599_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_2305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[54\]_TE mprj_logic_high_inst/HI[256] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_buffers\[10\]_A user_wb_dat_gates\[10\]/Y vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XFILLER_11_503 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1773 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_529 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_2073 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1924 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[82\] _345_/Y mprj_logic_high_inst/HI[284] vssd vccd la_oenb_core[82]
+ vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_2_223 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[30\] _462_/Y mprj_dat_buf\[30\]/TE vssd vccd mprj_dat_o_user[30] vssd
+ vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input250_A la_data_out_mprj[91] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input348_A la_iena_mprj[64] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_1395 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input515_A la_oenb_mprj[9] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_433 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[105\] _368_/A la_buf_enable\[105\]/B vssd vccd la_buf\[105\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_33_149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_91 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_80 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_406_ _406_/A vssd vccd _406_/Y vssd vccd sky130_fd_sc_hd__clkinv_8
XFILLER_37_1559 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1971 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_337_ _337_/A vssd vccd _337_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_35_1272 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1759 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1633 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1021 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output734_A output734/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_1065 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1677 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[79\] input108/X user_to_mprj_in_gates\[79\]/B vssd vccd user_to_mprj_in_gates\[79\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_48_1699 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[92\]_TE la_buf\[92\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1839 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[77\]_TE mprj_logic_high_inst/HI[279] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[23\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_2002 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2073 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_27 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__651__A _651_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput606 mprj_dat_o_core[31] vssd vccd _463_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput617 mprj_sel_o_core[2] vssd vccd _398_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_21_2006 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_433 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[41\] input323/X mprj_logic_high_inst/HI[371] vssd vccd user_to_mprj_in_gates\[41\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_user_wb_dat_gates\[14\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_937 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_mprj_cyc_buf_TE mprj_cyc_buf/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_981 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1857 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input298_A la_iena_mprj[19] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_29 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__561__A _561_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input465_A la_oenb_mprj[54] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input61_A la_data_out_core[36] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1953 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1817 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_433 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1023 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_753 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_403 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1323 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[49\] user_to_mprj_in_gates\[49\]/Y vssd vccd output698/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_50_2213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_631 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output684_A output684/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_1643 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput10 la_data_out_core[105] vssd vccd input10/X vssd vccd sky130_fd_sc_hd__buf_4
Xinput21 la_data_out_core[115] vssd vccd input21/X vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_15_1687 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput54 la_data_out_core[2] vssd vccd input54/X vssd vccd sky130_fd_sc_hd__buf_4
Xinput43 la_data_out_core[1] vssd vccd input43/X vssd vccd sky130_fd_sc_hd__buf_4
XANTENNA__471__A _471_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput32 la_data_out_core[125] vssd vccd input32/X vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput87 la_data_out_core[5] vssd vccd input87/X vssd vccd sky130_fd_sc_hd__buf_2
Xinput65 la_data_out_core[3] vssd vccd input65/X vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput76 la_data_out_core[4] vssd vccd input76/X vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput98 la_data_out_core[6] vssd vccd input98/X vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_48_1485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1844 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1647 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1877 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1073 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_285 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[105\] input10/X user_to_mprj_in_gates\[105\]/B vssd vccd user_to_mprj_in_gates\[105\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_53_767 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__646__A _646_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xmprj2_logic_high_inst mprj2_pwrgood/A vccd2 vssd2 mprj2_logic_high
XFILLER_34_981 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[6\]_A _406_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__381__A _381_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[89\] input375/X mprj_logic_high_inst/HI[419] vssd vccd user_to_mprj_in_gates\[89\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_7_2309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[115\] _378_/Y mprj_logic_high_inst/HI[317] vssd vccd la_oenb_core[115]
+ vssd vccd sky130_fd_sc_hd__einvp_8
Xinput403 la_oenb_mprj[113] vssd vccd _376_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput425 la_oenb_mprj[18] vssd vccd _610_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput436 la_oenb_mprj[28] vssd vccd _620_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput414 la_oenb_mprj[123] vssd vccd _386_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput447 la_oenb_mprj[38] vssd vccd _630_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput458 la_oenb_mprj[48] vssd vccd _640_/A vssd vccd sky130_fd_sc_hd__buf_2
Xinput469 la_oenb_mprj[58] vssd vccd _650_/A vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_29_742 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[45\] _637_/Y mprj_logic_high_inst/HI[247] vssd vccd la_oenb_core[45]
+ vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[67\] _330_/A la_buf_enable\[67\]/B vssd vccd la_buf\[67\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_1_1229 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_797 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input213_A la_data_out_mprj[58] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_907 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_447 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__556__A _556_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1665 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input582_A mprj_dat_o_core[0] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_1963 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1865 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_1827 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_rstn_buf_TE mprj_rstn_buf/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[6\]_B mprj_logic_high_inst/HI[336] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1761 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[109\] _573_/Y la_buf\[109\]/TE vssd vccd la_data_in_core[109] vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_39_517 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2061 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[102\] user_to_mprj_in_gates\[102\]/Y vssd vccd output630/A
+ vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_23_1967 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1741 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1730 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_285 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__466__A _466_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_789 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_439 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1738 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_1153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[102\]_A_N _365_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_1353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1315 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1397 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[117\]_A_N _380_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_1889 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[1\] _433_/Y mprj_dat_buf\[1\]/TE vssd vccd mprj_dat_o_user[1] vssd
+ vccd sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf_enable\[127\]_B la_buf_enable\[127\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xmprj_logic_high_inst mprj_rstn_buf/TE la_buf_enable\[26\]/B la_buf_enable\[27\]/B
+ la_buf_enable\[28\]/B la_buf_enable\[29\]/B la_buf_enable\[30\]/B la_buf_enable\[31\]/B
+ la_buf_enable\[32\]/B la_buf_enable\[33\]/B la_buf_enable\[34\]/B la_buf_enable\[35\]/B
+ mprj_adr_buf\[0\]/TE la_buf_enable\[36\]/B la_buf_enable\[37\]/B la_buf_enable\[38\]/B
+ la_buf_enable\[39\]/B la_buf_enable\[40\]/B la_buf_enable\[41\]/B la_buf_enable\[42\]/B
+ la_buf_enable\[43\]/B la_buf_enable\[44\]/B la_buf_enable\[45\]/B mprj_adr_buf\[1\]/TE
+ la_buf_enable\[46\]/B la_buf_enable\[47\]/B la_buf_enable\[48\]/B la_buf_enable\[49\]/B
+ la_buf_enable\[50\]/B la_buf_enable\[51\]/B la_buf_enable\[52\]/B la_buf_enable\[53\]/B
+ la_buf_enable\[54\]/B la_buf_enable\[55\]/B mprj_adr_buf\[2\]/TE la_buf_enable\[56\]/B
+ la_buf_enable\[57\]/B la_buf_enable\[58\]/B la_buf_enable\[59\]/B la_buf_enable\[60\]/B
+ la_buf_enable\[61\]/B la_buf_enable\[62\]/B la_buf_enable\[63\]/B la_buf_enable\[64\]/B
+ la_buf_enable\[65\]/B mprj_adr_buf\[3\]/TE la_buf_enable\[66\]/B la_buf_enable\[67\]/B
+ la_buf_enable\[68\]/B la_buf_enable\[69\]/B la_buf_enable\[70\]/B la_buf_enable\[71\]/B
+ la_buf_enable\[72\]/B la_buf_enable\[73\]/B la_buf_enable\[74\]/B la_buf_enable\[75\]/B
+ mprj_adr_buf\[4\]/TE la_buf_enable\[76\]/B la_buf_enable\[77\]/B la_buf_enable\[78\]/B
+ la_buf_enable\[79\]/B la_buf_enable\[80\]/B la_buf_enable\[81\]/B la_buf_enable\[82\]/B
+ la_buf_enable\[83\]/B la_buf_enable\[84\]/B la_buf_enable\[85\]/B mprj_adr_buf\[5\]/TE
+ la_buf_enable\[86\]/B la_buf_enable\[87\]/B la_buf_enable\[88\]/B la_buf_enable\[89\]/B
+ la_buf_enable\[90\]/B la_buf_enable\[91\]/B la_buf_enable\[92\]/B la_buf_enable\[93\]/B
+ la_buf_enable\[94\]/B la_buf_enable\[95\]/B mprj_adr_buf\[6\]/TE la_buf_enable\[96\]/B
+ la_buf_enable\[97\]/B la_buf_enable\[98\]/B la_buf_enable\[99\]/B la_buf_enable\[100\]/B
+ la_buf_enable\[101\]/B la_buf_enable\[102\]/B la_buf_enable\[103\]/B la_buf_enable\[104\]/B
+ la_buf_enable\[105\]/B mprj_adr_buf\[7\]/TE la_buf_enable\[106\]/B la_buf_enable\[107\]/B
+ la_buf_enable\[108\]/B la_buf_enable\[109\]/B la_buf_enable\[110\]/B la_buf_enable\[111\]/B
+ la_buf_enable\[112\]/B la_buf_enable\[113\]/B la_buf_enable\[114\]/B la_buf_enable\[115\]/B
+ mprj_adr_buf\[8\]/TE la_buf_enable\[116\]/B la_buf_enable\[117\]/B la_buf_enable\[118\]/B
+ la_buf_enable\[119\]/B la_buf_enable\[120\]/B la_buf_enable\[121\]/B la_buf_enable\[122\]/B
+ la_buf_enable\[123\]/B la_buf_enable\[124\]/B la_buf_enable\[125\]/B mprj_adr_buf\[9\]/TE
+ mprj_clk_buf/TE la_buf_enable\[126\]/B la_buf_enable\[127\]/B mprj_logic_high_inst/HI[202]
+ mprj_logic_high_inst/HI[203] mprj_logic_high_inst/HI[204] mprj_logic_high_inst/HI[205]
+ mprj_logic_high_inst/HI[206] mprj_logic_high_inst/HI[207] mprj_logic_high_inst/HI[208]
+ mprj_logic_high_inst/HI[209] mprj_adr_buf\[10\]/TE mprj_logic_high_inst/HI[210]
+ mprj_logic_high_inst/HI[211] mprj_logic_high_inst/HI[212] mprj_logic_high_inst/HI[213]
+ mprj_logic_high_inst/HI[214] mprj_logic_high_inst/HI[215] mprj_logic_high_inst/HI[216]
+ mprj_logic_high_inst/HI[217] mprj_logic_high_inst/HI[218] mprj_logic_high_inst/HI[219]
+ mprj_adr_buf\[11\]/TE mprj_logic_high_inst/HI[220] mprj_logic_high_inst/HI[221]
+ mprj_logic_high_inst/HI[222] mprj_logic_high_inst/HI[223] mprj_logic_high_inst/HI[224]
+ mprj_logic_high_inst/HI[225] mprj_logic_high_inst/HI[226] mprj_logic_high_inst/HI[227]
+ mprj_logic_high_inst/HI[228] mprj_logic_high_inst/HI[229] mprj_adr_buf\[12\]/TE
+ mprj_logic_high_inst/HI[230] mprj_logic_high_inst/HI[231] mprj_logic_high_inst/HI[232]
+ mprj_logic_high_inst/HI[233] mprj_logic_high_inst/HI[234] mprj_logic_high_inst/HI[235]
+ mprj_logic_high_inst/HI[236] mprj_logic_high_inst/HI[237] mprj_logic_high_inst/HI[238]
+ mprj_logic_high_inst/HI[239] mprj_adr_buf\[13\]/TE mprj_logic_high_inst/HI[240]
+ mprj_logic_high_inst/HI[241] mprj_logic_high_inst/HI[242] mprj_logic_high_inst/HI[243]
+ mprj_logic_high_inst/HI[244] mprj_logic_high_inst/HI[245] mprj_logic_high_inst/HI[246]
+ mprj_logic_high_inst/HI[247] mprj_logic_high_inst/HI[248] mprj_logic_high_inst/HI[249]
+ mprj_adr_buf\[14\]/TE mprj_logic_high_inst/HI[250] mprj_logic_high_inst/HI[251]
+ mprj_logic_high_inst/HI[252] mprj_logic_high_inst/HI[253] mprj_logic_high_inst/HI[254]
+ mprj_logic_high_inst/HI[255] mprj_logic_high_inst/HI[256] mprj_logic_high_inst/HI[257]
+ mprj_logic_high_inst/HI[258] mprj_logic_high_inst/HI[259] mprj_adr_buf\[15\]/TE
+ mprj_logic_high_inst/HI[260] mprj_logic_high_inst/HI[261] mprj_logic_high_inst/HI[262]
+ mprj_logic_high_inst/HI[263] mprj_logic_high_inst/HI[264] mprj_logic_high_inst/HI[265]
+ mprj_logic_high_inst/HI[266] mprj_logic_high_inst/HI[267] mprj_logic_high_inst/HI[268]
+ mprj_logic_high_inst/HI[269] mprj_adr_buf\[16\]/TE mprj_logic_high_inst/HI[270]
+ mprj_logic_high_inst/HI[271] mprj_logic_high_inst/HI[272] mprj_logic_high_inst/HI[273]
+ mprj_logic_high_inst/HI[274] mprj_logic_high_inst/HI[275] mprj_logic_high_inst/HI[276]
+ mprj_logic_high_inst/HI[277] mprj_logic_high_inst/HI[278] mprj_logic_high_inst/HI[279]
+ mprj_adr_buf\[17\]/TE mprj_logic_high_inst/HI[280] mprj_logic_high_inst/HI[281]
+ mprj_logic_high_inst/HI[282] mprj_logic_high_inst/HI[283] mprj_logic_high_inst/HI[284]
+ mprj_logic_high_inst/HI[285] mprj_logic_high_inst/HI[286] mprj_logic_high_inst/HI[288]
+ mprj_logic_high_inst/HI[289] mprj_adr_buf\[18\]/TE mprj_logic_high_inst/HI[290]
+ mprj_logic_high_inst/HI[291] mprj_logic_high_inst/HI[292] mprj_logic_high_inst/HI[293]
+ mprj_logic_high_inst/HI[294] mprj_logic_high_inst/HI[295] mprj_logic_high_inst/HI[296]
+ mprj_logic_high_inst/HI[297] mprj_logic_high_inst/HI[298] mprj_logic_high_inst/HI[299]
+ mprj_adr_buf\[19\]/TE mprj_clk2_buf/TE mprj_logic_high_inst/HI[300] mprj_logic_high_inst/HI[301]
+ mprj_logic_high_inst/HI[302] mprj_logic_high_inst/HI[303] mprj_logic_high_inst/HI[304]
+ mprj_logic_high_inst/HI[305] mprj_logic_high_inst/HI[306] mprj_logic_high_inst/HI[307]
+ mprj_logic_high_inst/HI[308] mprj_logic_high_inst/HI[309] mprj_adr_buf\[20\]/TE
+ mprj_logic_high_inst/HI[310] mprj_logic_high_inst/HI[311] mprj_logic_high_inst/HI[312]
+ mprj_logic_high_inst/HI[313] mprj_logic_high_inst/HI[314] mprj_logic_high_inst/HI[315]
+ mprj_logic_high_inst/HI[316] mprj_logic_high_inst/HI[317] mprj_logic_high_inst/HI[318]
+ mprj_logic_high_inst/HI[319] mprj_adr_buf\[21\]/TE mprj_logic_high_inst/HI[320]
+ mprj_logic_high_inst/HI[321] mprj_logic_high_inst/HI[322] mprj_logic_high_inst/HI[323]
+ mprj_logic_high_inst/HI[324] mprj_logic_high_inst/HI[325] mprj_logic_high_inst/HI[326]
+ mprj_logic_high_inst/HI[327] mprj_logic_high_inst/HI[328] mprj_logic_high_inst/HI[329]
+ mprj_adr_buf\[22\]/TE mprj_logic_high_inst/HI[330] mprj_logic_high_inst/HI[331]
+ mprj_logic_high_inst/HI[332] mprj_logic_high_inst/HI[333] mprj_logic_high_inst/HI[334]
+ mprj_logic_high_inst/HI[335] mprj_logic_high_inst/HI[336] mprj_logic_high_inst/HI[337]
+ mprj_logic_high_inst/HI[338] mprj_logic_high_inst/HI[339] mprj_adr_buf\[23\]/TE
+ mprj_logic_high_inst/HI[340] mprj_logic_high_inst/HI[341] mprj_logic_high_inst/HI[342]
+ mprj_logic_high_inst/HI[343] mprj_logic_high_inst/HI[344] mprj_logic_high_inst/HI[345]
+ mprj_logic_high_inst/HI[346] mprj_logic_high_inst/HI[347] mprj_logic_high_inst/HI[348]
+ mprj_logic_high_inst/HI[349] mprj_adr_buf\[24\]/TE mprj_logic_high_inst/HI[350]
+ mprj_logic_high_inst/HI[351] mprj_logic_high_inst/HI[352] mprj_logic_high_inst/HI[353]
+ mprj_logic_high_inst/HI[354] mprj_logic_high_inst/HI[355] mprj_logic_high_inst/HI[356]
+ mprj_logic_high_inst/HI[357] mprj_logic_high_inst/HI[358] mprj_logic_high_inst/HI[359]
+ mprj_adr_buf\[25\]/TE mprj_logic_high_inst/HI[360] mprj_logic_high_inst/HI[361]
+ mprj_logic_high_inst/HI[362] mprj_logic_high_inst/HI[363] mprj_logic_high_inst/HI[364]
+ mprj_logic_high_inst/HI[365] mprj_logic_high_inst/HI[366] mprj_logic_high_inst/HI[367]
+ mprj_logic_high_inst/HI[368] mprj_logic_high_inst/HI[369] mprj_adr_buf\[26\]/TE
+ mprj_logic_high_inst/HI[370] mprj_logic_high_inst/HI[371] mprj_logic_high_inst/HI[372]
+ mprj_logic_high_inst/HI[373] mprj_logic_high_inst/HI[374] mprj_logic_high_inst/HI[375]
+ mprj_logic_high_inst/HI[376] mprj_logic_high_inst/HI[377] mprj_logic_high_inst/HI[378]
+ mprj_logic_high_inst/HI[379] mprj_adr_buf\[27\]/TE mprj_logic_high_inst/HI[380]
+ mprj_logic_high_inst/HI[381] mprj_logic_high_inst/HI[382] mprj_logic_high_inst/HI[383]
+ mprj_logic_high_inst/HI[384] mprj_logic_high_inst/HI[385] mprj_logic_high_inst/HI[386]
+ mprj_logic_high_inst/HI[387] mprj_logic_high_inst/HI[388] mprj_logic_high_inst/HI[389]
+ mprj_adr_buf\[28\]/TE mprj_logic_high_inst/HI[390] mprj_logic_high_inst/HI[391]
+ mprj_logic_high_inst/HI[392] mprj_logic_high_inst/HI[393] mprj_logic_high_inst/HI[394]
+ mprj_logic_high_inst/HI[395] mprj_logic_high_inst/HI[396] mprj_logic_high_inst/HI[397]
+ mprj_logic_high_inst/HI[398] mprj_logic_high_inst/HI[399] mprj_adr_buf\[29\]/TE
+ mprj_cyc_buf/TE mprj_logic_high_inst/HI[400] mprj_logic_high_inst/HI[401] mprj_logic_high_inst/HI[402]
+ mprj_logic_high_inst/HI[403] mprj_logic_high_inst/HI[404] mprj_logic_high_inst/HI[405]
+ mprj_logic_high_inst/HI[406] mprj_logic_high_inst/HI[407] mprj_logic_high_inst/HI[408]
+ mprj_logic_high_inst/HI[409] mprj_adr_buf\[30\]/TE mprj_logic_high_inst/HI[410]
+ mprj_logic_high_inst/HI[411] mprj_logic_high_inst/HI[412] mprj_logic_high_inst/HI[413]
+ mprj_logic_high_inst/HI[414] mprj_logic_high_inst/HI[415] mprj_logic_high_inst/HI[416]
+ mprj_logic_high_inst/HI[417] mprj_logic_high_inst/HI[418] mprj_logic_high_inst/HI[419]
+ mprj_adr_buf\[31\]/TE mprj_logic_high_inst/HI[420] mprj_logic_high_inst/HI[421]
+ mprj_logic_high_inst/HI[422] mprj_logic_high_inst/HI[423] mprj_logic_high_inst/HI[424]
+ mprj_logic_high_inst/HI[425] mprj_logic_high_inst/HI[426] mprj_logic_high_inst/HI[427]
+ mprj_logic_high_inst/HI[428] mprj_dat_buf\[0\]/TE mprj_logic_high_inst/HI[430] mprj_logic_high_inst/HI[431]
+ mprj_logic_high_inst/HI[432] mprj_logic_high_inst/HI[433] mprj_logic_high_inst/HI[434]
+ mprj_logic_high_inst/HI[435] mprj_logic_high_inst/HI[436] mprj_logic_high_inst/HI[437]
+ mprj_logic_high_inst/HI[438] mprj_logic_high_inst/HI[439] mprj_dat_buf\[1\]/TE mprj_logic_high_inst/HI[440]
+ mprj_logic_high_inst/HI[441] mprj_logic_high_inst/HI[442] mprj_logic_high_inst/HI[443]
+ mprj_logic_high_inst/HI[444] mprj_logic_high_inst/HI[445] mprj_logic_high_inst/HI[446]
+ mprj_logic_high_inst/HI[447] mprj_logic_high_inst/HI[448] mprj_logic_high_inst/HI[449]
+ mprj_dat_buf\[2\]/TE mprj_logic_high_inst/HI[450] mprj_logic_high_inst/HI[451] mprj_logic_high_inst/HI[452]
+ mprj_logic_high_inst/HI[453] mprj_logic_high_inst/HI[454] mprj_logic_high_inst/HI[455]
+ mprj_logic_high_inst/HI[456] mprj_logic_high_inst/HI[457] user_irq_ena_buf\[0\]/B
+ user_irq_ena_buf\[1\]/B mprj_dat_buf\[3\]/TE user_irq_ena_buf\[2\]/B mprj_pwrgood/A
+ user_to_mprj_wb_ena_buf/B mprj_dat_buf\[4\]/TE mprj_dat_buf\[5\]/TE mprj_dat_buf\[6\]/TE
+ mprj_dat_buf\[7\]/TE mprj_stb_buf/TE mprj_dat_buf\[8\]/TE mprj_dat_buf\[9\]/TE mprj_dat_buf\[10\]/TE
+ mprj_dat_buf\[11\]/TE mprj_dat_buf\[12\]/TE mprj_dat_buf\[13\]/TE mprj_dat_buf\[14\]/TE
+ mprj_dat_buf\[15\]/TE mprj_dat_buf\[16\]/TE mprj_dat_buf\[17\]/TE mprj_we_buf/TE
+ mprj_dat_buf\[18\]/TE mprj_dat_buf\[19\]/TE mprj_dat_buf\[20\]/TE mprj_dat_buf\[21\]/TE
+ mprj_dat_buf\[22\]/TE mprj_dat_buf\[23\]/TE mprj_dat_buf\[24\]/TE mprj_dat_buf\[25\]/TE
+ mprj_dat_buf\[26\]/TE mprj_dat_buf\[27\]/TE mprj_sel_buf\[0\]/TE mprj_dat_buf\[28\]/TE
+ mprj_dat_buf\[29\]/TE mprj_dat_buf\[30\]/TE mprj_dat_buf\[31\]/TE la_buf_enable\[0\]/B
+ la_buf_enable\[1\]/B la_buf_enable\[2\]/B la_buf_enable\[3\]/B la_buf_enable\[4\]/B
+ la_buf_enable\[5\]/B mprj_sel_buf\[1\]/TE la_buf_enable\[6\]/B la_buf_enable\[7\]/B
+ la_buf_enable\[8\]/B la_buf_enable\[9\]/B la_buf_enable\[10\]/B la_buf_enable\[11\]/B
+ la_buf_enable\[12\]/B la_buf_enable\[13\]/B la_buf_enable\[14\]/B la_buf_enable\[15\]/B
+ mprj_sel_buf\[2\]/TE la_buf_enable\[16\]/B la_buf_enable\[17\]/B la_buf_enable\[18\]/B
+ la_buf_enable\[19\]/B la_buf_enable\[20\]/B la_buf_enable\[21\]/B la_buf_enable\[22\]/B
+ la_buf_enable\[23\]/B la_buf_enable\[24\]/B la_buf_enable\[25\]/B mprj_sel_buf\[3\]/TE
+ vccd1 mprj_logic_high_inst/HI[287] mprj_logic_high_inst/HI[429] vssd1 mprj_logic_high
XFILLER_26_1591 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_1516 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__376__A _376_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_1985 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1805 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[96\]_A input127/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_69 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1849 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_461 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1551 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_605 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1860 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1057 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1945 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2067 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input163_A la_data_out_mprj[12] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput211 la_data_out_mprj[56] vssd vccd _520_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput200 la_data_out_mprj[46] vssd vccd _510_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
XANTENNA_user_to_mprj_in_gates\[20\]_A input44/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[118\]_B la_buf_enable\[118\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_2201 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_1989 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1500 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput222 la_data_out_mprj[66] vssd vccd _530_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
XANTENNA_input428_A la_oenb_mprj[20] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input330_A la_iena_mprj[48] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput233 la_data_out_mprj[76] vssd vccd _540_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput244 la_data_out_mprj[86] vssd vccd _550_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_36_509 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput255 la_data_out_mprj[96] vssd vccd _560_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
XANTENNA_input24_A la_data_out_core[118] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput266 la_iena_mprj[105] vssd vccd input266/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput277 la_iena_mprj[115] vssd vccd input277/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput288 la_iena_mprj[125] vssd vccd input288/X vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_29_561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1173 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_723 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_654_ _654_/A vssd vccd _654_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
Xinput299 la_iena_mprj[1] vssd vccd input299/X vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_40_1577 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[72\] _536_/Y la_buf\[72\]/TE vssd vccd la_data_in_core[72] vssd vccd sky130_fd_sc_hd__einvp_8
X_585_ _585_/A vssd vccd _585_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_31_225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[87\]_A input117/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_buffers\[9\]_A user_wb_dat_gates\[9\]/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_1927 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_1771 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_792 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_483 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1635 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1083 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xoutput707 output707/A vssd vccd la_data_in_mprj[57] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput718 output718/A vssd vccd la_data_in_mprj[67] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput729 output729/A vssd vccd la_data_in_mprj[77] vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA_output647_A output647/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_2145 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1381 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_693 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[11\]_A input26/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[109\]_B la_buf_enable\[109\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_1742 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[61\] input89/X user_to_mprj_in_gates\[61\]/B vssd vccd user_to_mprj_in_gates\[61\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_48_881 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1775 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_501 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[78\]_A input107/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_545 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_589 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1557 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1123 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[26\]_TE la_buf\[26\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[6\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1757 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2321 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2207 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1703 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[0\]_A_N _592_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_1653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1747 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1697 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_2150 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_807 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[6\]_B user_to_mprj_in_gates\[6\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_2_2058 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1897 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_564 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_370_ _370_/A vssd vccd _370_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_39_1793 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[69\]_A input97/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_903 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1911 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input280_A la_iena_mprj[118] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_2107 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input378_A la_iena_mprj[91] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_1392 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_2129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1999 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input545_A mprj_adr_o_core[6] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_1753 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1257 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_1904 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1341 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1915 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2097 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_1385 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_637_ _637_/A vssd vccd _637_/Y vssd vccd sky130_fd_sc_hd__inv_2
X_568_ _568_/A vssd vccd _568_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_32_589 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[31\] user_to_mprj_in_gates\[31\]/Y vssd vccd output679/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
X_499_ _499_/A vssd vccd _499_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_la_buf\[49\]_TE la_buf\[49\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_2160 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output764_A output764/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_291 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1481 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_51 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1951 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1973 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_807 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_1594 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_821 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1034 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1619 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_865 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__654__A _654_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_1933 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1565 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_427 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2151 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1049 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1016 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[71\] input356/X mprj_logic_high_inst/HI[401] vssd vccd user_to_mprj_in_gates\[71\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_49_57 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1511 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2059 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_637 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input126_A la_data_out_core[95] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_422_ _422_/A vssd vccd _422_/Y vssd vccd sky130_fd_sc_hd__inv_6
XFILLER_39_2291 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[126\]_A input33/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__564__A _564_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_353_ _353_/A vssd vccd _353_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_input495_A la_oenb_mprj[81] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf\[35\] _499_/Y la_buf\[35\]/TE vssd vccd la_data_in_core[35] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input91_A la_data_out_core[63] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_751 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[107\] input268/X mprj_logic_high_inst/HI[437] vssd vccd
+ user_to_mprj_in_gates\[107\]/B vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_5_221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_795 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_gates\[7\] input579/X user_wb_ack_gate/B vssd vccd user_wb_dat_gates\[7\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_8
XFILLER_5_254 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1065 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput8 la_data_out_core[103] vssd vccd input8/X vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_20_1723 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_1870 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_497 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_buffers\[79\] user_to_mprj_in_gates\[79\]/Y vssd vccd output731/A
+ vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_36_136 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[60\]_A_N _652_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_865 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_331 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[117\]_A input23/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__474__A _474_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_1229 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[24\] input48/X user_to_mprj_in_gates\[24\]/B vssd vccd user_to_mprj_in_gates\[24\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XANTENNA_la_buf_enable\[75\]_A_N _338_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_2335 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1831 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[13\]_A_N _605_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_1875 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1717 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__649__A _649_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_1981 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[28\]_A_N _620_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_1474 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_629 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_331 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[108\]_A input13/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__384__A _384_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_515 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1785 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_559 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1936 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2085 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_oen_buffers\[75\] _338_/Y mprj_logic_high_inst/HI[277] vssd vccd la_oenb_core[75]
+ vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_2_235 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_279 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xla_buf_enable\[97\] _360_/A la_buf_enable\[97\]/B vssd vccd la_buf\[97\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_2
XFILLER_47_1892 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xmprj_dat_buf\[23\] _455_/Y mprj_dat_buf\[23\]/TE vssd vccd mprj_dat_o_user[23] vssd
+ vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input243_A la_data_out_mprj[85] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_1756 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__559__A _559_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_946 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input410_A la_oenb_mprj[11] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_445 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input508_A la_oenb_mprj[93] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_489 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_92 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_81 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_70 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_150 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_81 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_405_ _405_/A vssd vccd _405_/Y vssd vccd sky130_fd_sc_hd__inv_16
XFILLER_30_824 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_336_ _336_/A vssd vccd _336_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_19_1983 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_1284 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1705 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_1645 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1033 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_1509 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output727_A output727/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1689 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1138 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__469__A _469_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_63 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[122\]_TE mprj_logic_high_inst/HI[324] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_1761 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1772 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[70\]_A input355/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_183 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xla_buf_enable\[3\] _595_/A la_buf_enable\[3\]/B vssd vccd la_buf\[3\]/TE vssd vccd
+ sky130_fd_sc_hd__and2b_1
XANTENNA_la_buf_enable\[6\]_B la_buf_enable\[6\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_39 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1693 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1199 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2143 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput618 mprj_sel_o_core[3] vssd vccd _399_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput607 mprj_dat_o_core[3] vssd vccd _435_/A vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_5_2237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1525 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__379__A _379_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_957 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[21\]_TE mprj_logic_high_inst/HI[223] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_445 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_489 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[34\] input315/X mprj_logic_high_inst/HI[364] vssd vccd user_to_mprj_in_gates\[34\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_in_ena_buf\[61\]_A input345/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_695 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_993 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_150 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1869 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_839 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_2169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_378 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[12\] _604_/A la_buf_enable\[12\]/B vssd vccd la_buf\[12\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XANTENNA_input193_A la_data_out_mprj[3] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_1468 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input360_A la_iena_mprj[75] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input458_A la_oenb_mprj[48] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1829 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input54_A la_data_out_core[2] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input625_A user_irq_ena[1] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_209 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_721 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_445 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_765 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xpowergood_check vccd vssd vdda1 vdda2 mprj2_vdd_pwrgood/A mprj_vdd_pwrgood/A dw_194404_9184#
+ vssa1 dw_201986_9164# vssa2 mgmt_protect_hv
XFILLER_34_415 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2003 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_489 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1978 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_448 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[52\]_A input335/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_1335 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_2225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output677_A output677/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_2269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput11 la_data_out_core[106] vssd vccd input11/X vssd vccd sky130_fd_sc_hd__buf_4
Xinput22 la_data_out_core[116] vssd vccd input22/X vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_15_1655 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1699 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput55 la_data_out_core[30] vssd vccd input55/X vssd vccd sky130_fd_sc_hd__buf_4
Xinput44 la_data_out_core[20] vssd vccd input44/X vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput33 la_data_out_core[126] vssd vccd input33/X vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput77 la_data_out_core[50] vssd vccd input77/X vssd vccd sky130_fd_sc_hd__buf_4
Xinput66 la_data_out_core[40] vssd vccd input66/X vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput88 la_data_out_core[60] vssd vccd input88/X vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput99 la_data_out_core[70] vssd vccd input99/X vssd vccd sky130_fd_sc_hd__buf_4
Xuser_to_mprj_in_gates\[91\] input122/X user_to_mprj_in_gates\[91\]/B vssd vccd user_to_mprj_in_gates\[91\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_48_1497 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[44\]_TE mprj_logic_high_inst/HI[246] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_1801 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1856 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1659 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1889 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_sel_buf\[0\]_A _396_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[43\]_A input325/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_993 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_278 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1007 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_809 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2227 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput426 la_oenb_mprj[19] vssd vccd _611_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput437 la_oenb_mprj[29] vssd vccd _621_/A vssd vccd sky130_fd_sc_hd__buf_2
Xinput404 la_oenb_mprj[114] vssd vccd _377_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput415 la_oenb_mprj[124] vssd vccd _387_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
Xuser_to_mprj_oen_buffers\[108\] _371_/Y mprj_logic_high_inst/HI[310] vssd vccd la_oenb_core[108]
+ vssd vccd sky130_fd_sc_hd__einvp_8
Xinput448 la_oenb_mprj[39] vssd vccd _631_/A vssd vccd sky130_fd_sc_hd__dlymetal6s2s_1
Xinput459 la_oenb_mprj[49] vssd vccd _641_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_29_754 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1208 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_713 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[38\] _630_/Y mprj_logic_high_inst/HI[240] vssd vccd la_oenb_core[38]
+ vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_44_757 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_919 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_2209 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_459 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input206_A la_data_out_mprj[51] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[34\]_A input315/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_1677 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_1833 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1390 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__572__A _572_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_1839 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[82\]_TE la_buf\[82\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input575_A mprj_dat_i_user[3] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_dat_buf\[1\]_A _433_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[67\]_TE mprj_logic_high_inst/HI[269] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1773 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1637 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_529 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_573 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1979 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1419 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_201 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[61\] user_to_mprj_in_gates\[61\]/Y vssd vccd output712/A
+ vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_19_297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[25\]_A input305/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output794_A output794/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_749 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1619 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_2066 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__482__A _482_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_1327 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_mprj_dat_buf\[31\]_TE mprj_dat_buf\[31\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1283 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[90\]_A user_to_mprj_in_gates\[90\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_2_2207 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_1653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_713 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_573 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__657__A _657_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_576 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[16\]_A input295/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_749 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[96\]_B user_to_mprj_in_gates\[96\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_39_1997 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1817 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_473 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__392__A _392_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_1563 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_105 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1913 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1957 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2079 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput201 la_data_out_mprj[47] vssd vccd _511_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
XANTENNA_user_to_mprj_in_buffers\[81\]_A user_to_mprj_in_gates\[81\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_input156_A la_data_out_mprj[121] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[20\]_B user_to_mprj_in_gates\[20\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_40_2213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput245 la_data_out_mprj[87] vssd vccd _551_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput234 la_data_out_mprj[77] vssd vccd _541_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput223 la_data_out_mprj[67] vssd vccd _531_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput212 la_data_out_mprj[57] vssd vccd _521_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_44_1681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1512 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput256 la_data_out_mprj[97] vssd vccd _561_/A vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA_input323_A la_iena_mprj[41] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput267 la_iena_mprj[106] vssd vccd input267/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput278 la_iena_mprj[116] vssd vccd input278/X vssd vccd sky130_fd_sc_hd__clkbuf_1
XANTENNA__567__A _567_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input17_A la_data_out_core[111] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput289 la_iena_mprj[126] vssd vccd input289/X vssd vccd sky130_fd_sc_hd__clkbuf_1
X_653_ _653_/A vssd vccd _653_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_17_735 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1589 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_565 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xla_buf\[65\] _529_/Y la_buf\[65\]/TE vssd vccd la_data_in_core[65] vssd vccd sky130_fd_sc_hd__einvp_8
X_584_ _584_/A vssd vccd _584_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_38_1441 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[87\]_B user_to_mprj_in_gates\[87\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_51_2353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_934 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_440 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1603 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_956 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_495 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1647 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[121\] _585_/Y la_buf\[121\]/TE vssd vccd la_data_in_core[121] vssd vccd sky130_fd_sc_hd__einvp_8
Xmprj_adr_buf\[29\] _429_/Y mprj_adr_buf\[29\]/TE vssd vccd mprj_adr_o_user[29] vssd
+ vccd sky130_fd_sc_hd__einvp_8
Xoutput708 output708/A vssd vccd la_data_in_mprj[58] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput719 output719/A vssd vccd la_data_in_mprj[68] vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_10_1393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_2157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[72\]_A user_to_mprj_in_gates\[72\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[11\]_B user_to_mprj_in_gates\[11\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_39_337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1973 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1754 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[54\] input81/X user_to_mprj_in_gates\[54\]/B vssd vccd user_to_mprj_in_gates\[54\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XANTENNA__477__A _477_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_893 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_521 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1787 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1583 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_557 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_226 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[78\]_B user_to_mprj_in_gates\[78\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_17_1569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1173 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1135 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1179 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[110\]_A user_to_mprj_in_gates\[110\]/Y vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_609 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1621 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2219 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1715 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[63\]_A user_to_mprj_in_gates\[63\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_38_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2090 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input9_A la_data_out_core[104] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__387__A _387_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_329 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_576 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_727 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[69\]_B user_to_mprj_in_gates\[69\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_35_1636 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input273_A la_iena_mprj[111] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[101\]_A user_to_mprj_in_gates\[101\]/Y vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_2119 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1691 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input440_A la_oenb_mprj[31] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[54\]_A user_to_mprj_in_gates\[54\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_input538_A mprj_adr_o_core[29] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_1721 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_1765 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[101\]_A_N _364_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_1353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1927 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_189 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_841 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1397 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_636_ _636_/A vssd vccd _636_/Y vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_17_587 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_567_ _567_/A vssd vccd _567_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_mprj_adr_buf\[22\]_TE mprj_adr_buf\[22\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[116\]_A_N _379_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_498_ _498_/A vssd vccd _498_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_la_buf\[94\]_A _558_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_1769 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_1591 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[24\] user_to_mprj_in_gates\[24\]/Y vssd vccd output671/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_51_1493 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output757_A output757/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_981 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1190 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_491 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[45\]_A user_to_mprj_in_gates\[45\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_29_1985 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1689 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1046 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_833 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_321 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1901 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1945 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_877 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[85\]_A _549_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_1956 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1989 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1577 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1028 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_69 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1905 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1523 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[36\]_A user_to_mprj_in_gates\[36\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_8_1567 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1409 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[64\] input348/X mprj_logic_high_inst/HI[394] vssd vccd user_to_mprj_in_gates\[64\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_45_137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[2\] _594_/Y mprj_logic_high_inst/HI[204] vssd vccd la_oenb_core[2]
+ vssd vccd sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[20\] _612_/Y mprj_logic_high_inst/HI[222] vssd vccd la_oenb_core[20]
+ vssd vccd sky130_fd_sc_hd__einvp_8
X_421_ _421_/A vssd vccd _421_/Y vssd vccd sky130_fd_sc_hd__inv_12
Xla_buf_enable\[42\] _634_/A la_buf_enable\[42\]/B vssd vccd la_buf\[42\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XANTENNA_input119_A la_data_out_core[89] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_844 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_352_ _352_/A vssd vccd _352_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_user_to_mprj_in_gates\[126\]_B user_to_mprj_in_gates\[126\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_35_2167 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[76\]_A _540_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input390_A la_oenb_mprj[101] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_763 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input488_A la_oenb_mprj[75] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[94\]_B la_buf_enable\[94\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input84_A la_data_out_core[57] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_1731 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[28\] _492_/Y la_buf\[28\]/TE vssd vccd la_data_in_core[28] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA__580__A _580_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_1775 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_60 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_266 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_93 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_1237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[27\]_A user_to_mprj_in_gates\[27\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_7_1022 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1077 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput9 la_data_out_core[104] vssd vccd input9/X vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_40_1161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[16\]_TE la_buf\[16\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_619_ _619_/A vssd vccd _619_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_17_351 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[117\]_B user_to_mprj_in_gates\[117\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[67\]_A _531_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_387 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[17\] input40/X user_to_mprj_in_gates\[17\]/B vssd vccd user_to_mprj_in_gates\[17\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_9_550 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[85\]_B la_buf_enable\[85\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__490__A _490_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_buffers\[27\] user_wb_dat_gates\[27\]/Y vssd vccd output775/A vssd vccd
+ sky130_fd_sc_hd__clkinv_8
XFILLER_25_2347 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1843 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[18\]_A user_to_mprj_in_gates\[18\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_29_1793 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2110 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1887 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[26\]_A input568/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_1729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_27 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_641 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[108\]_B user_to_mprj_in_gates\[108\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[58\]_A _522_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_685 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1797 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[76\]_B la_buf_enable\[76\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1341 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_1959 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1320 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[68\] _331_/Y mprj_logic_high_inst/HI[270] vssd vccd la_oenb_core[68]
+ vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_43_1768 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[16\] _448_/Y mprj_dat_buf\[16\]/TE vssd vccd mprj_dat_o_user[16] vssd
+ vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input236_A la_data_out_mprj[79] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[39\]_TE la_buf\[39\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[17\]_A input558/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input403_A la_oenb_mprj[113] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_2218 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__575__A _575_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_2229 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XPHY_82 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_71 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_60 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[49\]_A _513_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_404_ _404_/A vssd vccd _404_/Y vssd vccd sky130_fd_sc_hd__inv_2
XPHY_93 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_836 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_93 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_335_ _335_/A vssd vccd _335_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_41_162 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_869 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[67\]_B la_buf_enable\[67\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_571 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xmprj_adr_buf\[11\] _411_/Y mprj_adr_buf\[11\]/TE vssd vccd mprj_adr_o_user[11] vssd
+ vccd sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_buffers\[125\] user_to_mprj_in_gates\[125\]/Y vssd vccd output655/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_38_903 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[91\] user_to_mprj_in_gates\[91\]/Y vssd vccd output745/A
+ vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_38_925 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_424 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_273 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_939 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_671 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1784 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__485__A _485_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_buffers\[1\] user_wb_dat_gates\[1\]/Y vssd vccd output767/A vssd vccd
+ sky130_fd_sc_hd__clkinv_8
XANTENNA_user_to_mprj_in_ena_buf\[70\]_B mprj_logic_high_inst/HI[400] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_36_1005 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[7\]_TE la_buf\[7\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_663 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1049 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_685 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_2097 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[58\]_B la_buf_enable\[58\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1661 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[125\]_A _388_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[60\]_A _652_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_1145 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2111 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2155 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1009 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1651 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput608 mprj_dat_o_core[4] vssd vccd _436_/A vssd vccd sky130_fd_sc_hd__buf_4
Xinput619 mprj_stb_o_core vssd vccd _394_/A vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_5_1504 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1537 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_969 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_405 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_917 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__395__A _395_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[27\] input307/X mprj_logic_high_inst/HI[357] vssd vccd user_to_mprj_in_gates\[27\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_in_ena_buf\[61\]_B mprj_logic_high_inst/HI[391] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_52_961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_162 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_335 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[49\]_B la_buf_enable\[49\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input186_A la_data_out_mprj[33] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[116\]_A _379_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[51\]_A _643_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input353_A la_iena_mprj[69] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input47_A la_data_out_core[23] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_2277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input520_A mprj_adr_o_core[12] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[0\] input260/X mprj_logic_high_inst/HI[330] vssd vccd user_to_mprj_in_gates\[0\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
Xla_buf\[95\] _559_/Y la_buf\[95\]/TE vssd vccd la_data_in_core[95] vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[110\] _373_/A la_buf_enable\[110\]/B vssd vccd la_buf\[110\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XANTENNA_input618_A mprj_sel_o_core[3] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[74\]_A_N _337_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_777 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1957 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[89\]_A_N _352_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[52\]_B mprj_logic_high_inst/HI[382] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_43_983 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[12\]_A_N _604_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput12 la_data_out_core[107] vssd vccd input12/X vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_11_891 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[9\]_A input387/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput45 la_data_out_core[21] vssd vccd input45/X vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput23 la_data_out_core[117] vssd vccd input23/X vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput34 la_data_out_core[127] vssd vccd input34/X vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput89 la_data_out_core[61] vssd vccd input89/X vssd vccd sky130_fd_sc_hd__buf_4
Xinput78 la_data_out_core[51] vssd vccd input78/X vssd vccd sky130_fd_sc_hd__buf_4
Xinput67 la_data_out_core[41] vssd vccd input67/X vssd vccd sky130_fd_sc_hd__buf_4
XANTENNA_user_to_mprj_oen_buffers\[42\]_A _634_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[107\]_A _370_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput56 la_data_out_core[31] vssd vccd input56/X vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_48_1421 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[27\]_A_N _619_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1329 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[84\] input114/X user_to_mprj_in_gates\[84\]/B vssd vccd user_to_mprj_in_gates\[84\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_6_1813 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_232 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1868 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_1097 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_799 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_405 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_257 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[43\]_B mprj_logic_high_inst/HI[373] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_21_611 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1019 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[33\]_A _625_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_2239 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput427 la_oenb_mprj[1] vssd vccd _593_/A vssd vccd sky130_fd_sc_hd__buf_2
Xinput405 la_oenb_mprj[115] vssd vccd _378_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput416 la_oenb_mprj[125] vssd vccd _388_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_5_1301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput449 la_oenb_mprj[3] vssd vccd _595_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput438 la_oenb_mprj[2] vssd vccd _594_/A vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_5_1345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_725 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_769 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1601 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[34\]_B mprj_logic_high_inst/HI[364] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_input101_A la_data_out_core[72] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_1689 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_942 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1845 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_615 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input470_A la_oenb_mprj[59] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[6\] _470_/Y la_buf\[6\]/TE vssd vccd la_data_in_core[6] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_oen_buffers\[24\]_A _616_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[112\]_TE mprj_logic_high_inst/HI[314] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input568_A mprj_dat_i_user[26] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf\[10\] _474_/Y la_buf\[10\]/TE vssd vccd la_data_in_core[10] vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_49_1785 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1649 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[3\] _403_/Y mprj_adr_buf\[3\]/TE vssd vccd mprj_adr_o_user[3] vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_47_541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_we_buf_TE mprj_we_buf/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[20\]_A _420_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_585 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_235 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[54\] user_to_mprj_in_gates\[54\]/Y vssd vccd output704/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_user_to_mprj_in_ena_buf\[25\]_B mprj_logic_high_inst/HI[355] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_output787_A output787/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_430 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_953 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_2045 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2078 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_gates\[12\] input553/X user_wb_ack_gate/B vssd vccd user_wb_dat_gates\[12\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_oen_buffers\[11\]_TE mprj_logic_high_inst/HI[213] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[15\]_A _607_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1295 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1665 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[110\] input16/X user_to_mprj_in_gates\[110\]/B vssd vccd user_to_mprj_in_gates\[110\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XANTENNA_mprj_adr_buf\[11\]_A _411_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_533 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_585 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1932 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[16\]_B mprj_logic_high_inst/HI[346] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_43_27 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_268 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_419 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1829 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[9\]_A input581/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_629 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[94\] input381/X mprj_logic_high_inst/HI[424] vssd vccd user_to_mprj_in_gates\[94\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_46_1925 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_oen_buffers\[120\] _383_/Y mprj_logic_high_inst/HI[322] vssd vccd la_oenb_core[120]
+ vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_44_2361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_1969 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_sel_buf\[1\] _397_/Y mprj_sel_buf\[1\]/TE vssd vccd mprj_sel_o_user[1] vssd
+ vccd sky130_fd_sc_hd__einvp_8
Xinput202 la_data_out_mprj[48] vssd vccd _512_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_40_2225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput224 la_data_out_mprj[68] vssd vccd _532_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput213 la_data_out_mprj[58] vssd vccd _522_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput235 la_data_out_mprj[78] vssd vccd _542_/A vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA_user_to_mprj_in_gates\[9\]_A input131/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input149_A la_data_out_mprj[115] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_2269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_530 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_1693 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1524 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[50\] _642_/Y mprj_logic_high_inst/HI[252] vssd vccd la_oenb_core[50]
+ vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[72\] _335_/A la_buf_enable\[72\]/B vssd vccd la_buf\[72\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
Xinput246 la_data_out_mprj[88] vssd vccd _552_/A vssd vccd sky130_fd_sc_hd__buf_2
Xinput257 la_data_out_mprj[98] vssd vccd _562_/A vssd vccd sky130_fd_sc_hd__buf_2
Xinput268 la_iena_mprj[107] vssd vccd input268/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput279 la_iena_mprj[117] vssd vccd input279/X vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_5_1153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input316_A la_iena_mprj[35] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_652_ _652_/A vssd vccd _652_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_44_533 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_583_ _583_/A vssd vccd _583_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_16_279 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[58\] _522_/Y la_buf\[58\]/TE vssd vccd la_data_in_core[58] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA__583__A _583_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_1453 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1620 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[34\]_TE mprj_logic_high_inst/HI[236] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_979 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_946 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_1615 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1659 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xoutput709 output709/A vssd vccd la_data_in_mprj[59] vssd vccd sky130_fd_sc_hd__buf_2
Xla_buf\[114\] _578_/Y la_buf\[114\]/TE vssd vccd la_data_in_core[114] vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_45_2169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1805 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output702_A output702/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_1711 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1985 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_1766 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1849 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1799 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_533 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[47\] input73/X user_to_mprj_in_gates\[47\]/B vssd vccd user_to_mprj_in_gates\[47\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_50_525 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_238 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__493__A _493_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[9\]_TE mprj_adr_buf\[9\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_1141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1147 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[9\] input131/X user_to_mprj_in_gates\[9\]/B vssd vccd user_to_mprj_in_gates\[9\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_4
XFILLER_8_1727 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_511 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[72\]_TE la_buf\[72\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_533 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_739 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[57\]_TE mprj_logic_high_inst/HI[259] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_2327 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1648 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2073 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[98\] _361_/Y mprj_logic_high_inst/HI[300] vssd vccd la_oenb_core[98]
+ vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input266_A la_iena_mprj[105] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_632 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_1777 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input433_A la_oenb_mprj[25] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__578__A _578_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input600_A mprj_dat_o_core[26] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_1939 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_831 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_1365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_853 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_635_ _635_/A vssd vccd _635_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_mprj_dat_buf\[24\]_A _456_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_897 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_buffers\[31\]_A user_wb_dat_gates\[31\]/Y vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
X_566_ _566_/A vssd vccd _566_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_17_599 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_mprj_dat_buf\[21\]_TE mprj_dat_buf\[21\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_1261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_1737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_497_ _497_/A vssd vccd _497_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_8_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[0\]_TE mprj_logic_high_inst/HI[202] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[17\] user_to_mprj_in_gates\[17\]/Y vssd vccd output663/A
+ vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_47_2209 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output652_A output652/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_993 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[95\]_TE la_buf\[95\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_1997 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2314 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__488__A _488_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_dat_buf\[15\]_A _447_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_buffers\[22\]_A user_wb_dat_gates\[22\]/Y vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XFILLER_50_333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1913 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_29 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_385 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1058 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_377 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1589 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1441 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1535 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1917 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_1485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__398__A _398_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_1641 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1579 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[57\] input340/X mprj_logic_high_inst/HI[387] vssd vccd user_to_mprj_in_gates\[57\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_41_2353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_503 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_420_ _420_/A vssd vccd _420_/Y vssd vccd sky130_fd_sc_hd__clkinv_8
XANTENNA_user_wb_dat_buffers\[13\]_A user_wb_dat_gates\[13\]/Y vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XFILLER_2_1178 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_856 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[13\] _605_/Y mprj_logic_high_inst/HI[215] vssd vccd la_oenb_core[13]
+ vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[35\] _627_/A la_buf_enable\[35\]/B vssd vccd la_buf\[35\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
X_351_ _351_/A vssd vccd _351_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_39_1581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[9\] user_to_mprj_in_gates\[9\]/Y vssd vccd output754/A vssd
+ vccd sky130_fd_sc_hd__inv_6
XANTENNA_input383_A la_iena_mprj[96] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_1743 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_735 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_713 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_775 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_757 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input77_A la_data_out_core[50] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input550_A mprj_dat_i_user[0] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_72 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_985 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_1541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1089 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1703 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1933 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1173 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_190 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_363 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_618_ _618_/A vssd vccd _618_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_32_300 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_549_ _549_/A vssd vccd _549_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_9_562 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1761 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2326 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1811 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1855 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_29 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1899 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[26\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_39 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_609 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_683 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1721 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_697 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_27 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[100\]_A_N _363_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[12\]_TE mprj_adr_buf\[12\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_215 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_248 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_1861 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[115\]_A_N _378_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[17\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_1229 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_926 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input131_A la_data_out_core[9] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input229_A la_data_out_mprj[72] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_108 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_469 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_403_ _403_/A vssd vccd _403_/Y vssd vccd sky130_fd_sc_hd__inv_12
XPHY_83 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_50 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_72 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_61 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input598_A mprj_dat_o_core[24] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[2\]_A _466_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_804 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XPHY_94 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_848 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[40\] _504_/Y la_buf\[40\]/TE vssd vccd la_data_in_core[40] vssd vccd sky130_fd_sc_hd__einvp_8
X_334_ _334_/A vssd vccd _334_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
Xuser_to_mprj_in_ena_buf\[112\] input274/X mprj_logic_high_inst/HI[442] vssd vccd
+ user_to_mprj_in_gates\[112\]/B vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA__591__A _591_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1117 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[118\] user_to_mprj_in_gates\[118\]/Y vssd vccd output647/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_1_281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_irq_gates\[2\]_A input623/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_915 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_1257 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_937 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[84\] user_to_mprj_in_gates\[84\]/Y vssd vccd output737/A
+ vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_37_436 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1691 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[0\]_TE mprj_dat_buf\[0\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_1796 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_981 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_683 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1017 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_152 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1905 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_697 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[120\]_TE la_buf\[120\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1102 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2123 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1630 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput609 mprj_dat_o_core[5] vssd vccd _437_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_25_2167 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1663 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1549 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1251 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[9\]_A _409_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_973 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_303 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_347 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1871 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1735 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[80\] _343_/Y mprj_logic_high_inst/HI[282] vssd vccd la_oenb_core[80]
+ vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input179_A la_data_out_mprj[27] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1978 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[50\]_A input77/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input346_A la_iena_mprj[62] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_2289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input513_A la_oenb_mprj[98] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1831 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1048 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[88\] _552_/Y la_buf\[88\]/TE vssd vccd la_data_in_core[88] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA__586__A _586_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[103\] _366_/A la_buf_enable\[103\]/B vssd vccd la_buf\[103\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_46_277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_981 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_995 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_461 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1602 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_1771 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_645 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[0\]_A user_to_mprj_in_gates\[0\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xinput13 la_data_out_core[108] vssd vccd input13/X vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_50_2249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_841 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput46 la_data_out_core[22] vssd vccd input46/X vssd vccd sky130_fd_sc_hd__buf_4
Xinput35 la_data_out_core[12] vssd vccd input35/X vssd vccd sky130_fd_sc_hd__clkbuf_2
XANTENNA_user_to_mprj_in_ena_buf\[9\]_B mprj_logic_high_inst/HI[339] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xinput24 la_data_out_core[118] vssd vccd input24/X vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_48_2101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1993 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput79 la_data_out_core[52] vssd vccd input79/X vssd vccd sky130_fd_sc_hd__buf_4
Xinput57 la_data_out_core[32] vssd vccd input57/X vssd vccd sky130_fd_sc_hd__buf_4
Xinput68 la_data_out_core[42] vssd vccd input68/X vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_10_391 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output732_A output732/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[41\]_A input67/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1308 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[77\] input106/X user_to_mprj_in_gates\[77\]/B vssd vccd user_to_mprj_in_gates\[77\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_22_1606 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__496__A _496_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_2261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_266 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_244 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_491 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_461 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[90\]_TE mprj_logic_high_inst/HI[292] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_973 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_29 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_111 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1172 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[29\]_TE la_buf\[29\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1481 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[32\]_A input57/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput428 la_oenb_mprj[20] vssd vccd _612_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput406 la_oenb_mprj[116] vssd vccd _379_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput417 la_oenb_mprj[126] vssd vccd _389_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_5_1313 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput439 la_oenb_mprj[30] vssd vccd _622_/A vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_5_1357 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[99\]_A input130/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_2314 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1613 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_781 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_954 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_623 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_667 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input296_A la_iena_mprj[17] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_627 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_844 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input463_A la_oenb_mprj[52] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[23\]_A input47/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_81 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_597 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_247 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_781 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_921 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_932 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output682_A output682/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_17_1719 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[47\] user_to_mprj_in_gates\[47\]/Y vssd vccd output696/A
+ vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_33_1009 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_987 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_442 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[14\]_A input37/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_1127 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1105 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2251 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1677 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[103\] input8/X user_to_mprj_in_gates\[103\]/B vssd vccd user_to_mprj_in_gates\[103\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_39_1922 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1944 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_39 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_781 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[73\]_A_N _336_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[9\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[87\] input373/X mprj_logic_high_inst/HI[417] vssd vccd user_to_mprj_in_gates\[87\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_la_buf_enable\[88\]_A_N _351_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[113\] _376_/Y mprj_logic_high_inst/HI[315] vssd vccd la_oenb_core[113]
+ vssd vccd sky130_fd_sc_hd__einvp_8
Xmprj_clk2_buf _392_/Y mprj_clk2_buf/TE vssd vccd user_clock2 vssd vccd sky130_fd_sc_hd__einvp_8
Xinput225 la_data_out_mprj[69] vssd vccd _533_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput214 la_data_out_mprj[59] vssd vccd _523_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput203 la_data_out_mprj[49] vssd vccd _513_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
XANTENNA_user_to_mprj_in_gates\[9\]_B user_to_mprj_in_gates\[9\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xinput236 la_data_out_mprj[79] vssd vccd _543_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_5_1121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput258 la_data_out_mprj[99] vssd vccd _563_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput247 la_data_out_mprj[89] vssd vccd _553_/A vssd vccd sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_la_buf_enable\[11\]_A_N _603_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput269 la_iena_mprj[108] vssd vccd input269/X vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_40_1536 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[43\] _635_/Y mprj_logic_high_inst/HI[245] vssd vccd la_oenb_core[43]
+ vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[65\] _657_/A la_buf_enable\[65\]/B vssd vccd la_buf\[65\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_5_1165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
X_651_ _651_/A vssd vccd _651_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_44_501 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_irq_buffers\[1\] user_irq_gates\[1\]/Y vssd vccd output793/A vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_input211_A la_data_out_mprj[56] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_582_ _582_/A vssd vccd _582_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_44_545 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input309_A la_iena_mprj[29] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[26\]_A_N _618_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_2322 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1465 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1329 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input580_A mprj_dat_i_user[8] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_1627 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_2273 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_1561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1425 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[107\] _571_/Y la_buf\[107\]/TE vssd vccd la_data_in_core[107] vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_45_1469 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[100\] user_to_mprj_in_gates\[100\]/Y vssd vccd output628/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_3_1817 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_545 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[120\]_A input283/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_1429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_991 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_1981 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_1441 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2028 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[102\]_TE mprj_logic_high_inst/HI[304] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_523 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_545 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[111\]_A input273/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_2339 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1785 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_924 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2085 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_405 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input259_A la_data_out_mprj[9] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input161_A la_data_out_mprj[126] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_1609 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2001 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1789 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input426_A la_oenb_mprj[19] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_2045 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input22_A la_data_out_core[116] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_2089 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
X_634_ _634_/A vssd vccd _634_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_45_865 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[70\] _534_/Y la_buf\[70\]/TE vssd vccd la_data_in_core[70] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA__594__A _594_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_565_ _565_/A vssd vccd _565_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_53_1705 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_1803 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_496_ _496_/A vssd vccd _496_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_user_to_mprj_in_ena_buf\[102\]_A input263/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_711 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_755 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_788 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output645_A output645/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[125\]_TE mprj_logic_high_inst/HI[327] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_1761 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_2326 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1004 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1925 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_389 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_29 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_27 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1453 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_2321 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1929 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1547 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[24\]_TE mprj_logic_high_inst/HI[226] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_1653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[91\]_A input378/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_813 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_802 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_515 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_350_ _350_/A vssd vccd _350_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_35_1413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1593 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[28\] _620_/A la_buf_enable\[28\]/B vssd vccd la_buf\[28\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_13_1755 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input376_A la_iena_mprj[8] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_747 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1206 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input543_A mprj_adr_o_core[4] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_975 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__589__A _589_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_1597 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1901 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_629 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1945 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1715 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_1989 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[82\]_A input368/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_1737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_617_ _617_/A vssd vccd _617_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_17_375 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_2203 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_548_ _548_/A vssd vccd _548_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_53_1535 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_479_ _479_/A vssd vccd _479_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_53_1579 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output762_A output762/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_574 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[62\]_TE la_buf\[62\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[47\]_TE mprj_logic_high_inst/HI[249] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__499__A _499_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_1773 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1867 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_117 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[73\]_A input358/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_695 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_665 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_378 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1733 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_39 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1619 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[9\]_B la_buf_enable\[9\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_1261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_mprj_dat_buf\[11\]_TE mprj_dat_buf\[11\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_1737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_629 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1399 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_938 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[64\]_A input348/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input124_A la_data_out_core[93] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XPHY_40 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_402_ _402_/A vssd vccd _402_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_25_51 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XPHY_62 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_51 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_73 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_95 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_84 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_333_ _333_/A vssd vccd _333_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_input493_A la_oenb_mprj[7] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[85\]_TE la_buf\[85\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_511 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[105\] input266/X mprj_logic_high_inst/HI[435] vssd vccd
+ user_to_mprj_in_gates\[105\]/B vssd vccd sky130_fd_sc_hd__and2_1
Xla_buf\[33\] _497_/Y la_buf\[33\]/TE vssd vccd la_data_in_core[33] vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_10_551 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_533 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_gates\[5\] input577/X user_wb_ack_gate/B vssd vccd user_wb_dat_gates\[5\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_4
XFILLER_2_783 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_33 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1946 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_irq_gates\[2\]_B user_irq_gates\[2\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[77\] user_to_mprj_in_gates\[77\]/Y vssd vccd output729/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_user_to_mprj_in_ena_buf\[55\]_A input338/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_971 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_695 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[22\] input46/X user_to_mprj_in_gates\[22\]/B vssd vccd user_to_mprj_in_gates\[22\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_36_1029 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1917 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_2353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_1114 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1642 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1675 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2179 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_mprj_sel_buf\[3\]_A _399_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_949 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[46\]_A input328/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_440 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_359 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_1883 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1173 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1747 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[50\]_B user_to_mprj_in_gates\[50\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[73\] _336_/Y mprj_logic_high_inst/HI[275] vssd vccd la_oenb_core[73]
+ vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[95\] _358_/A la_buf_enable\[95\]/B vssd vccd la_buf\[95\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
Xoutput690 output690/A vssd vccd la_data_in_mprj[41] vssd vccd sky130_fd_sc_hd__buf_2
Xmprj_dat_buf\[21\] _453_/Y mprj_dat_buf\[21\]/TE vssd vccd mprj_dat_o_user[21] vssd
+ vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input339_A la_iena_mprj[56] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input241_A la_data_out_mprj[83] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_1005 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_1843 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_245 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input506_A la_oenb_mprj[91] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[37\]_A input318/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_61 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2017 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_993 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_643 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_657 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[4\]_A _436_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput36 la_data_out_core[13] vssd vccd input36/X vssd vccd sky130_fd_sc_hd__buf_4
Xinput14 la_data_out_core[109] vssd vccd input14/X vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput25 la_data_out_core[119] vssd vccd input25/X vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_7_853 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput47 la_data_out_core[23] vssd vccd input47/X vssd vccd sky130_fd_sc_hd__buf_4
Xinput58 la_data_out_core[33] vssd vccd input58/X vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput69 la_data_out_core[43] vssd vccd input69/X vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_48_2113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_2157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2146 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[41\]_B user_to_mprj_in_gates\[41\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1456 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output725_A output725/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_1033 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_713 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_757 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[28\]_A input308/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_256 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_473 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[114\]_A_N _377_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_1861 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_123 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[1\] _593_/A la_buf_enable\[1\]/B vssd vccd la_buf\[1\]/TE vssd vccd
+ sky130_fd_sc_hd__and2b_1
XFILLER_31_1493 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[93\]_A user_to_mprj_in_gates\[93\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[32\]_B user_to_mprj_in_gates\[32\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_44_1821 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput407 la_oenb_mprj[117] vssd vccd _380_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput418 la_oenb_mprj[127] vssd vccd _390_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_9_1483 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2059 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput429 la_oenb_mprj[21] vssd vccd _613_/A vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_5_1325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1369 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[19\]_A input298/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_749 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_ena_buf\[32\] input313/X mprj_logic_high_inst/HI[362] vssd vccd user_to_mprj_in_gates\[32\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_43_237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[99\]_B user_to_mprj_in_gates\[99\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_52_793 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_635 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_966 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_105 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_41 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[10\] _602_/A la_buf_enable\[10\]/B vssd vccd la_buf\[10\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XANTENNA_input191_A la_data_out_mprj[38] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_22_85 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1511 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input289_A la_iena_mprj[126] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[120\]_A _584_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input456_A la_oenb_mprj[46] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[84\]_A user_to_mprj_in_gates\[84\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[23\]_B user_to_mprj_in_gates\[23\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_input52_A la_data_out_core[28] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input623_A user_irq_core[2] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__597__A _597_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[110\]_TE la_buf\[110\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_1712 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_93 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[25\]_TE mprj_adr_buf\[25\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_1113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_944 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_1591 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output675_A output675/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_999 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_buffers\[122\]_A user_to_mprj_in_gates\[122\]/Y vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[111\]_A _575_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[75\]_A user_to_mprj_in_gates\[75\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[14\]_B user_to_mprj_in_gates\[14\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_28_1805 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2263 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1849 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1117 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1623 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1139 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1689 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2081 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_215 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1956 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_793 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2245 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_buffers\[113\]_A user_to_mprj_in_gates\[113\]/Y vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_1599 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1831 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[102\]_A _566_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_1875 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[66\]_A user_to_mprj_in_gates\[66\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_27_2049 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_837 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xinput226 la_data_out_mprj[6] vssd vccd _470_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput215 la_data_out_mprj[5] vssd vccd _469_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput204 la_data_out_mprj[4] vssd vccd _468_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_40_2249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[106\] _369_/Y mprj_logic_high_inst/HI[308] vssd vccd la_oenb_core[106]
+ vssd vccd sky130_fd_sc_hd__einvp_8
Xinput259 la_data_out_mprj[9] vssd vccd _473_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput237 la_data_out_mprj[7] vssd vccd _471_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput248 la_data_out_mprj[8] vssd vccd _472_/A vssd vccd sky130_fd_sc_hd__dlymetal6s2s_1
X_650_ _650_/A vssd vccd _650_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_22_1971 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_576 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[36\] _628_/Y mprj_logic_high_inst/HI[238] vssd vccd la_oenb_core[36]
+ vssd vccd sky130_fd_sc_hd__einvp_8
X_581_ _581_/A vssd vccd _581_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
Xla_buf_enable\[58\] _650_/A la_buf_enable\[58\]/B vssd vccd la_buf\[58\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_44_557 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input204_A la_data_out_mprj[4] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_403 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2334 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_447 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[104\]_A user_to_mprj_in_gates\[104\]/Y vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input573_A mprj_dat_i_user[30] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_2105 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_2241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[57\]_A user_to_mprj_in_gates\[57\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[30\]_A _494_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1437 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[80\]_TE mprj_logic_high_inst/HI[282] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_1871 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_841 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1829 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[19\]_TE la_buf\[19\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output792_A output792/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[97\]_A _561_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_2109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[120\]_B mprj_logic_high_inst/HI[450] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_31_741 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1853 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_785 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[48\]_A user_to_mprj_in_gates\[48\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[21\]_A _485_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1061 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_29 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_841 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1453 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[88\]_A _552_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[111\]_B mprj_logic_high_inst/HI[441] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_10_947 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_2097 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1959 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_929 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[39\]_A user_to_mprj_in_gates\[39\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[12\]_A _476_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_1217 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input154_A la_data_out_mprj[11] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_2193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2013 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[30\]_B la_buf_enable\[30\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input321_A la_iena_mprj[3] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_2057 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input419_A la_oenb_mprj[12] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input15_A la_data_out_core[10] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_633_ _633_/A vssd vccd _633_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_17_535 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[63\] _527_/Y la_buf\[63\]/TE vssd vccd la_data_in_core[63] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf\[79\]_A _543_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_877 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_888 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
X_564_ _564_/A vssd vccd _564_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_2_1884 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_538 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_495_ _495_/A vssd vccd _495_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_user_to_mprj_in_ena_buf\[102\]_B mprj_logic_high_inst/HI[432] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1105 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_590 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[97\]_B la_buf_enable\[97\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_2120 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_1859 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_723 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_767 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[27\] _427_/Y mprj_adr_buf\[27\]/TE vssd vccd mprj_adr_o_user[27] vssd
+ vccd sky130_fd_sc_hd__einvp_8
XANTENNA_output638_A output638/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1381 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1245 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1808 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_ack_gate input516/X user_wb_ack_gate/B vssd vccd user_wb_ack_gate/Y vssd
+ vccd sky130_fd_sc_hd__nand2_4
XANTENNA_la_buf_enable\[21\]_B la_buf_enable\[21\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2338 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[52\] input79/X user_to_mprj_in_gates\[52\]/B vssd vccd user_to_mprj_in_gates\[52\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
Xinput590 mprj_dat_o_core[17] vssd vccd _449_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
XANTENNA_la_buf_enable\[72\]_A_N _335_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_1565 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_332 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_2004 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[87\]_A_N _350_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_357 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[88\]_B la_buf_enable\[88\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_1205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_2204 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1503 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[10\]_A_N _602_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[90\]_A _353_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[25\]_A_N _617_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_2019 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_39 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[29\]_A input571/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_2333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[12\]_B la_buf_enable\[12\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input7_A la_data_out_core[102] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_1559 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1621 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_1665 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1272 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_693 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1136 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[91\]_B mprj_logic_high_inst/HI[421] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_26_365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_313 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_398 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_527 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_825 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_869 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[79\]_B la_buf_enable\[79\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_1425 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_571 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_700 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1881 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[81\]_A _344_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_41 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_1767 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input271_A la_iena_mprj[10] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input369_A la_iena_mprj[83] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_85 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_1521 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input536_A mprj_adr_o_core[27] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_486 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[126\] _389_/A la_buf_enable\[126\]/B vssd vccd la_buf\[126\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_4_1913 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_1957 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[82\]_B mprj_logic_high_inst/HI[412] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_4_1979 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_1197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_641 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_616_ _616_/A vssd vccd _616_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_45_685 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_387 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_547_ _547_/A vssd vccd _547_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
X_478_ _478_/A vssd vccd _478_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_9_531 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[22\] user_to_mprj_in_gates\[22\]/Y vssd vccd output669/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_user_to_mprj_oen_buffers\[72\]_A _335_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_1271 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output755_A output755/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_781 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_1785 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1445 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[73\]_B mprj_logic_high_inst/HI[403] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_50_121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2001 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2045 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[63\]_A _655_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1377 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_1841 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_2141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[62\] input346/X mprj_logic_high_inst/HI[392] vssd vccd user_to_mprj_in_gates\[62\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_43_1727 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_2185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_641 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[64\]_B mprj_logic_high_inst/HI[394] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XPHY_30 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_685 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[0\] _592_/Y mprj_logic_high_inst/HI[202] vssd vccd la_oenb_core[0]
+ vssd vccd sky130_fd_sc_hd__einvp_8
X_401_ _401_/A vssd vccd _401_/Y vssd vccd sky130_fd_sc_hd__inv_12
Xla_buf_enable\[40\] _632_/A la_buf_enable\[40\]/B vssd vccd la_buf\[40\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XANTENNA_input117_A la_data_out_core[87] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XPHY_74 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_63 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_52 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_41 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_335 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_96 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_85 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1943 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_332_ _332_/A vssd vccd _332_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_35_1233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_2281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_390 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input486_A la_oenb_mprj[73] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[54\]_A _646_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[119\]_A _382_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[115\]_TE mprj_logic_high_inst/HI[317] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input82_A la_data_out_core[55] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_51 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_1553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_545 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[26\] _490_/Y la_buf\[26\]/TE vssd vccd la_data_in_core[26] vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_6_523 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_589 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2052 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1958 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_795 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_1237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_405 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1721 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_89 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_1557 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[55\]_B mprj_logic_high_inst/HI[385] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_20_1579 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_2045 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1929 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[15\] input38/X user_to_mprj_in_gates\[15\]/B vssd vccd user_to_mprj_in_gates\[15\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_2
Xuser_wb_dat_gates\[28\] input570/X user_wb_ack_gate/B vssd vccd user_wb_dat_gates\[28\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_2
XFILLER_53_1377 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[14\]_TE mprj_logic_high_inst/HI[216] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[45\]_A _637_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_383 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_372 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_wb_dat_buffers\[25\] user_wb_dat_gates\[25\]/Y vssd vccd output773/A vssd vccd
+ sky130_fd_sc_hd__inv_6
XFILLER_29_2250 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1593 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1687 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[126\] input33/X user_to_mprj_in_gates\[126\]/B vssd vccd user_to_mprj_in_gates\[126\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_46_29 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[46\]_B mprj_logic_high_inst/HI[376] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_36_1553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[36\]_A _628_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_1851 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1895 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1704 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1759 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_2225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xoutput680 output680/A vssd vccd la_data_in_mprj[32] vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_43_1513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[66\] _329_/Y mprj_logic_high_inst/HI[268] vssd vccd la_oenb_core[66]
+ vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[88\] _351_/A la_buf_enable\[88\]/B vssd vccd la_buf\[88\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
Xoutput691 output691/A vssd vccd la_data_in_mprj[42] vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_19_405 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1175 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[14\] _446_/Y mprj_dat_buf\[14\]/TE vssd vccd mprj_dat_o_user[14] vssd
+ vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input234_A la_data_out_mprj[77] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_1164 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_1811 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1916 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_909 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1855 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[37\]_B mprj_logic_high_inst/HI[367] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_15_600 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input401_A la_oenb_mprj[111] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[52\]_TE la_buf\[52\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_953 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2029 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_633 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[37\]_TE mprj_logic_high_inst/HI[239] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_1751 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_699 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_61 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_1637 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_669 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput37 la_data_out_core[14] vssd vccd input37/X vssd vccd sky130_fd_sc_hd__buf_4
Xinput26 la_data_out_core[11] vssd vccd input26/X vssd vccd sky130_fd_sc_hd__clkbuf_2
XANTENNA_user_to_mprj_oen_buffers\[27\]_A _619_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput15 la_data_out_core[10] vssd vccd input15/X vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput48 la_data_out_core[24] vssd vccd input48/X vssd vccd sky130_fd_sc_hd__buf_4
Xinput59 la_data_out_core[34] vssd vccd input59/X vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_48_2169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1468 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[123\] user_to_mprj_in_gates\[123\]/Y vssd vccd output653/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_46_1181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output718_A output718/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[23\]_A _423_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_2191 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_725 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_769 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[28\]_B mprj_logic_high_inst/HI[358] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_34_920 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1704 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_1873 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_135 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2151 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[0\]_A _592_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[18\]_A _610_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_2195 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2209 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1833 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput419 la_oenb_mprj[12] vssd vccd _604_/A vssd vccd sky130_fd_sc_hd__buf_2
Xinput408 la_oenb_mprj[118] vssd vccd _381_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_9_1451 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1495 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[14\]_A _414_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[75\]_TE la_buf\[75\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_1877 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[19\]_B mprj_logic_high_inst/HI[349] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_43_205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[25\] input305/X mprj_logic_high_inst/HI[355] vssd vccd user_to_mprj_in_gates\[25\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_24_441 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_1902 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_647 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_53 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_97 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1523 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_813 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input184_A la_data_out_mprj[31] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_2309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1567 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input449_A la_oenb_mprj[3] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input351_A la_iena_mprj[67] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input45_A la_data_out_core[21] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf\[93\] _557_/Y la_buf\[93\]/TE vssd vccd la_data_in_core[93] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input616_A mprj_sel_o_core[1] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_1685 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[24\]_TE mprj_dat_buf\[24\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[3\]_TE mprj_logic_high_inst/HI[205] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_30_477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_466 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output668_A output668/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1817 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[98\]_TE la_buf\[98\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_2325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[82\] input112/X user_to_mprj_in_gates\[82\]/B vssd vccd user_to_mprj_in_gates\[82\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_26_2242 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_890 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2275 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1635 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_2093 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_547 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_411 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2257 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1843 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1887 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_809 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput216 la_data_out_mprj[60] vssd vccd _524_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput205 la_data_out_mprj[50] vssd vccd _514_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput227 la_data_out_mprj[70] vssd vccd _534_/A vssd vccd sky130_fd_sc_hd__buf_2
Xinput238 la_data_out_mprj[80] vssd vccd _544_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput249 la_data_out_mprj[90] vssd vccd _554_/A vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_29_588 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1189 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_580_ _580_/A vssd vccd _580_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_38_2113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_525 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_208 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[29\] _621_/Y mprj_logic_high_inst/HI[231] vssd vccd la_oenb_core[29]
+ vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_9_927 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2346 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_63 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_426 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input399_A la_oenb_mprj[10] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_96 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_459 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[4\] _468_/Y la_buf\[4\]/TE vssd vccd la_data_in_core[4] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input566_A mprj_dat_i_user[24] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_2253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__401__A _401_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[113\]_A_N _376_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_1883 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1933 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[1\] _401_/Y mprj_adr_buf\[1\]/TE vssd vccd mprj_adr_o_user[1] vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_48_853 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[27\]_A _459_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_1521 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_385 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[52\] user_to_mprj_in_gates\[52\]/Y vssd vccd output702/A
+ vssd vccd sky130_fd_sc_hd__inv_2
XANTENNA_output785_A output785/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_753 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1821 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_gates\[10\] input551/X user_wb_ack_gate/B vssd vccd user_wb_dat_gates\[10\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_4
XFILLER_28_2304 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_853 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1465 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[18\]_A _450_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_buffers\[25\]_A user_wb_dat_gates\[25\]/Y vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XFILLER_41_517 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[100\]_TE la_buf\[100\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1651 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[92\] input379/X mprj_logic_high_inst/HI[422] vssd vccd user_to_mprj_in_gates\[92\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_mprj_adr_buf\[15\]_TE mprj_adr_buf\[15\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_0_145 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1229 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_639 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input147_A la_data_out_mprj[113] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_2025 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xla_buf_enable\[70\] _333_/A la_buf_enable\[70\]/B vssd vccd la_buf\[70\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_28_41 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_341 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_632_ _632_/A vssd vccd _632_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_user_wb_dat_buffers\[16\]_A user_wb_dat_gates\[16\]/Y vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XFILLER_28_85 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_547 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input314_A la_iena_mprj[33] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_563_ _563_/A vssd vccd _563_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_44_377 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[56\] _520_/Y la_buf\[56\]/TE vssd vccd la_data_in_core[56] vssd vccd sky130_fd_sc_hd__einvp_8
X_494_ _494_/A vssd vccd _494_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_38_1253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2154 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1117 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_735 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_wb_ena_buf input614/X user_to_mprj_wb_ena_buf/B vssd vccd user_wb_ack_gate/B
+ vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_51_1453 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_779 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1901 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xla_buf\[112\] _576_/Y la_buf\[112\]/TE vssd vccd la_data_in_core[112] vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_49_1393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1257 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output700_A output700/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_dat_buf\[3\]_TE mprj_dat_buf\[3\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput591 mprj_dat_o_core[18] vssd vccd _450_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput580 mprj_dat_i_user[8] vssd vccd input580/X vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_47_193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_856 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[120\]_B la_buf_enable\[120\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[45\] input71/X user_to_mprj_in_gates\[45\]/B vssd vccd user_to_mprj_in_gates\[45\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_2
XFILLER_23_517 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[123\]_TE la_buf\[123\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1515 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1971 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[7\] input109/X user_to_mprj_in_gates\[7\]/B vssd vccd user_to_mprj_in_gates\[7\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_4
XANTENNA_user_wb_dat_gates\[29\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_2345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1677 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_2241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_303 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_539 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[111\]_B la_buf_enable\[111\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_1437 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[70\]_TE mprj_logic_high_inst/HI[272] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_22_583 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_881 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_712 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1795 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[96\] _359_/Y mprj_logic_high_inst/HI[298] vssd vccd la_oenb_core[96]
+ vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_user_wb_dat_buffers\[2\]_A user_wb_dat_gates\[2\]/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[80\]_A input110/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input264_A la_iena_mprj[103] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_443 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_1533 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_51 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input431_A la_oenb_mprj[23] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_1831 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[9\] input387/X mprj_logic_high_inst/HI[339] vssd vccd user_to_mprj_in_gates\[9\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_input529_A mprj_adr_o_core[20] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_1588 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_1132 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_95 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[119\] _382_/A la_buf_enable\[119\]/B vssd vccd la_buf\[119\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_2
XFILLER_37_609 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1969 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_1728 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[5\]_A _469_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_615_ _615_/A vssd vccd _615_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_45_697 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_546_ _546_/A vssd vccd _546_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_la_buf_enable\[102\]_B la_buf_enable\[102\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_17_399 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_358 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1061 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1635 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_477_ _477_/A vssd vccd _477_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_41_881 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_587 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1283 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[15\] user_to_mprj_in_gates\[15\]/Y vssd vccd output661/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_output748_A output748/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output650_A output650/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[71\]_A input100/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1021 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1065 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[93\]_TE mprj_logic_high_inst/HI[295] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2013 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_881 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[62\]_A input90/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1389 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj2_pwrgood mprj2_pwrgood/A vssd vccd output790/A vssd vccd sky130_fd_sc_hd__buf_12
XFILLER_8_1335 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[55\] input338/X mprj_logic_high_inst/HI[385] vssd vccd user_to_mprj_in_gates\[55\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_41_2197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1441 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_31 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_20 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_601 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_303 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_400_ _400_/A vssd vccd _400_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_27_697 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XPHY_64 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_53 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_42 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_645 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_347 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[11\] _603_/Y mprj_logic_high_inst/HI[213] vssd vccd la_oenb_core[11]
+ vssd vccd sky130_fd_sc_hd__einvp_8
X_331_ _331_/A vssd vccd _331_/Y vssd vccd sky130_fd_sc_hd__inv_2
XPHY_97 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_86 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_75 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1381 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1201 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1955 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[7\] user_to_mprj_in_gates\[7\]/Y vssd vccd output732/A vssd
+ vccd sky130_fd_sc_hd__clkinv_4
Xla_buf_enable\[33\] _625_/A la_buf_enable\[33\]/B vssd vccd la_buf\[33\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_19_1999 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input381_A la_iena_mprj[94] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input479_A la_oenb_mprj[67] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[71\]_A_N _334_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_2329 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1565 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_557 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[19\] _483_/Y la_buf\[19\]/TE vssd vccd la_data_in_core[19] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_gates\[53\]_A input80/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input75_A la_data_out_core[49] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_1005 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_2064 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1341 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[86\]_A_N _349_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_1915 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1385 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1733 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_461 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_409 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_buffers\[3\]_A user_to_mprj_in_gates\[3\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_output698_A output698/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[24\]_A_N _616_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_529_ _529_/A vssd vccd _529_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_32_133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1621 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[39\]_A_N _631_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_395 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[44\]_A input70/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_2262 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_buffers\[18\] user_wb_dat_gates\[18\]/Y vssd vccd output765/A vssd vccd
+ sky130_fd_sc_hd__inv_6
XFILLER_25_2104 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_mprj_vdd_pwrgood_A mprj_vdd_pwrgood/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_1561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1699 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[119\] input25/X user_to_mprj_in_gates\[119\]/B vssd vccd user_to_mprj_in_gates\[119\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_52_921 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_601 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_645 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_634 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1521 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1565 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1716 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[35\]_A input60/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xoutput670 output670/A vssd vccd la_data_in_mprj[23] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput681 output681/A vssd vccd la_data_in_mprj[33] vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_43_2237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_1661 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1525 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xoutput692 output692/A vssd vccd la_data_in_mprj[43] vssd vccd sky130_fd_sc_hd__buf_2
Xuser_to_mprj_oen_buffers\[59\] _651_/Y mprj_logic_high_inst/HI[261] vssd vccd la_oenb_core[59]
+ vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_19_417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_1569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1187 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input227_A la_data_out_mprj[70] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_1293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_41 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_461 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1867 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_965 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input596_A mprj_dat_o_core[22] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_1763 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_851 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[110\] input272/X mprj_logic_high_inst/HI[440] vssd vccd
+ user_to_mprj_in_gates\[110\]/B vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_35_1053 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_895 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput16 la_data_out_core[110] vssd vccd input16/X vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput27 la_data_out_core[120] vssd vccd input27/X vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_7_833 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_321 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput49 la_data_out_core[25] vssd vccd input49/X vssd vccd sky130_fd_sc_hd__buf_4
Xinput38 la_data_out_core[15] vssd vccd input38/X vssd vccd sky130_fd_sc_hd__buf_4
XANTENNA_user_to_mprj_in_gates\[26\]_A input50/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__404__A _404_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[110\]_A input16/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[116\] user_to_mprj_in_gates\[116\]/Y vssd vccd output645/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_46_1193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[82\] user_to_mprj_in_gates\[82\]/Y vssd vccd output735/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_4_1541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_rstn_buf_A input3/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_497 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1885 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1749 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2163 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[17\]_A input40/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[101\]_A input6/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_1801 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2017 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1981 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xinput409 la_oenb_mprj[119] vssd vccd _382_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_44_1845 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1463 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[105\]_TE mprj_logic_high_inst/HI[307] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_759 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_217 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2063 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_464 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[18\] input297/X mprj_logic_high_inst/HI[348] vssd vccd user_to_mprj_in_gates\[18\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_36_1373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_1805 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_659 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1849 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1248 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_65 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1535 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1723 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_869 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input177_A la_data_out_mprj[25] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_1579 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_379 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input344_A la_iena_mprj[60] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input38_A la_data_out_core[15] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input511_A la_oenb_mprj[96] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_247 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1631 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1861 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[86\] _550_/Y la_buf\[86\]/TE vssd vccd la_data_in_core[86] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input609_A mprj_dat_o_core[5] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_258 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[101\] _364_/A la_buf_enable\[101\]/B vssd vccd la_buf\[101\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_21_1697 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_431 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_486 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_489 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_641 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_685 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output730_A output730/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[75\] input104/X user_to_mprj_in_gates\[75\]/B vssd vccd user_to_mprj_in_gates\[75\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_6_1647 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2061 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_589 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[123\]_A input286/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_1914 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_291 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_209 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_423 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1693 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1579 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1991 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[42\]_TE la_buf\[42\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1899 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_2321 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_828 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[27\]_TE mprj_logic_high_inst/HI[229] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
Xinput217 la_data_out_mprj[61] vssd vccd _525_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput206 la_data_out_mprj[51] vssd vccd _515_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_48_309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1271 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput228 la_data_out_mprj[71] vssd vccd _535_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput239 la_data_out_mprj[81] vssd vccd _545_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_38_2125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1984 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[114\]_A input276/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_2169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input294_A la_iena_mprj[15] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_438 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_2221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1343 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input461_A la_oenb_mprj[50] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input559_A mprj_dat_i_user[18] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_2265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_irq_ena_buf\[1\] input625/X user_irq_ena_buf\[1\]/B vssd vccd user_irq_gates\[1\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_49_2287 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1901 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1945 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1989 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_865 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_2223 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1544 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[105\]_A input266/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_22_209 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_721 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_buffers\[45\] user_to_mprj_in_gates\[45\]/Y vssd vccd output694/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_output680_A output680/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1833 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_765 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output778_A output778/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_798 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[65\]_TE la_buf\[65\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_1107 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1637 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2051 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1973 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_865 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[101\] input6/X user_to_mprj_in_gates\[101\]/B vssd vccd user_to_mprj_in_gates\[101\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_39_1733 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_529 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1933 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1939 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1663 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[85\] input371/X mprj_logic_high_inst/HI[415] vssd vccd user_to_mprj_in_gates\[85\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA__502__A _502_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_dat_buf\[14\]_TE mprj_dat_buf\[14\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_2151 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[111\] _374_/Y mprj_logic_high_inst/HI[313] vssd vccd la_oenb_core[111]
+ vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_ena_buf\[94\]_A input381/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[41\] _633_/Y mprj_logic_high_inst/HI[243] vssd vccd la_oenb_core[41]
+ vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[63\] _655_/A la_buf_enable\[63\]/B vssd vccd la_buf\[63\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
X_631_ _631_/A vssd vccd _631_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_28_97 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_562_ _562_/A vssd vccd _562_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_44_334 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_559 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input307_A la_iena_mprj[27] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_389 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_41 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_493_ _493_/A vssd vccd _493_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_44_85 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1817 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[88\]_TE la_buf\[88\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_2133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[49\] _513_/Y la_buf\[49\]/TE vssd vccd la_data_in_core[49] vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_51_1421 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_747 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_279 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_920 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2073 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_57 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__412__A _412_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf\[105\] _569_/Y la_buf\[105\]/TE vssd vccd la_data_in_core[105] vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_45_1269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[85\]_A input371/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_813 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput581 mprj_dat_i_user[9] vssd vccd input581/X vssd vccd sky130_fd_sc_hd__buf_8
Xinput570 mprj_dat_i_user[28] vssd vccd input570/X vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_47_161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xinput592 mprj_dat_o_core[19] vssd vccd _451_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_1_1341 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[38\] input63/X user_to_mprj_in_gates\[38\]/B vssd vccd user_to_mprj_in_gates\[38\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_23_529 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1527 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1983 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[76\]_A input361/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_1241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_1116 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_2253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_893 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[112\]_A_N _375_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_1741 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[80\]_B user_to_mprj_in_gates\[80\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[127\]_A_N _390_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_2213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[89\] _352_/Y mprj_logic_high_inst/HI[291] vssd vccd la_oenb_core[89]
+ vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_1_411 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input257_A la_data_out_mprj[98] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_1005 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1049 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_1854 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input424_A la_oenb_mprj[17] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[67\]_A input351/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input20_A la_data_out_core[114] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_1144 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_614_ _614_/A vssd vccd _614_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_2_1672 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_665 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_545_ _545_/A vssd vccd _545_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_44_197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1647 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_476_ _476_/A vssd vccd _476_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA__407__A _407_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_1073 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_893 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_511 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_599 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[71\]_B user_to_mprj_in_gates\[71\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_5_761 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output643_A output643/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1033 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1607 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1077 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[58\]_A input341/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_189 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1059 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2025 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1313 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[62\]_B user_to_mprj_in_gates\[62\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_8_1347 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_2165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[49\]_A input331/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_1453 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_ena_buf\[48\] input330/X mprj_logic_high_inst/HI[378] vssd vccd user_to_mprj_in_gates\[48\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_6_1093 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_21 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_10 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_613 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_665 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XPHY_54 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_65 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_43 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_32 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_315 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_330_ _330_/A vssd vccd _330_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XPHY_98 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_87 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_76 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_657 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_359 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1967 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_2261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xla_buf_enable\[26\] _618_/A la_buf_enable\[26\]/B vssd vccd la_buf\[26\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_39_1393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input374_A la_iena_mprj[88] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[53\]_B user_to_mprj_in_gates\[53\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_6_569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input68_A la_data_out_core[42] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input541_A mprj_adr_o_core[31] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_2076 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[113\]_TE la_buf\[113\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_764 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_775 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1397 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[28\]_TE mprj_adr_buf\[28\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_1701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1745 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_473 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1302 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_1313 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_528_ _528_/A vssd vccd _528_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_mprj_dat_buf\[7\]_A _439_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_2058 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_459_ _459_/A vssd vccd _459_/Y vssd vccd sky130_fd_sc_hd__inv_6
XANTENNA_output760_A output760/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_363 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[44\]_B user_to_mprj_in_gates\[44\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_29_2274 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__600__A _600_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[60\]_TE mprj_logic_high_inst/HI[262] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_1233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_613 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_454 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_657 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_307 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1533 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1577 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[96\]_A user_to_mprj_in_gates\[96\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[35\]_B user_to_mprj_in_gates\[35\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1905 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_517 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1728 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xoutput660 output660/A vssd vccd la_data_in_mprj[14] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput671 output671/A vssd vccd la_data_in_mprj[24] vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_47_1673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xoutput682 output682/A vssd vccd la_data_in_mprj[34] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput693 output693/A vssd vccd la_data_in_mprj[44] vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA__510__A _510_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_1537 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1982 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1199 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input122_A la_data_out_core[91] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_1824 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1879 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_buffers\[20\]_A user_to_mprj_in_gates\[20\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_36_53 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_473 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_624 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_605 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1731 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_668 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1021 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input491_A la_oenb_mprj[78] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_85 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1775 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input589_A mprj_dat_o_core[16] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_863 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1087 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1920 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[103\] input264/X mprj_logic_high_inst/HI[433] vssd vccd
+ user_to_mprj_in_gates\[103\]/B vssd vccd sky130_fd_sc_hd__and2_1
Xla_buf\[31\] _495_/Y la_buf\[31\]/TE vssd vccd la_data_in_core[31] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf\[123\]_A _587_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput17 la_data_out_core[111] vssd vccd input17/X vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput28 la_data_out_core[121] vssd vccd input28/X vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_6_333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_gates\[3\] input575/X user_wb_ack_gate/B vssd vccd user_wb_dat_gates\[3\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_in_buffers\[87\]_A user_to_mprj_in_gates\[87\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[26\]_B user_to_mprj_in_gates\[26\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xinput39 la_data_out_core[16] vssd vccd input39/X vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_7_878 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_377 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[110\]_B user_to_mprj_in_gates\[110\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[60\]_A _524_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[83\]_TE mprj_logic_high_inst/HI[285] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__420__A _420_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[109\] user_to_mprj_in_gates\[109\]/Y vssd vccd output637/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_4_1553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[75\] user_to_mprj_in_gates\[75\]/Y vssd vccd output727/A
+ vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_38_749 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_buffers\[11\]_A user_to_mprj_in_gates\[11\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_4_1597 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1820 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[20\] input44/X user_to_mprj_in_gates\[20\]/B vssd vccd user_to_mprj_in_gates\[20\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_53_1143 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1717 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[125\]_A user_to_mprj_in_gates\[125\]/Y vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_1897 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1187 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[114\]_A _578_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[17\]_B user_to_mprj_in_gates\[17\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_31_2175 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_wb_dat_buffers\[30\] user_wb_dat_gates\[30\]/Y vssd vccd output779/A vssd vccd
+ sky130_fd_sc_hd__clkinv_8
XANTENNA_user_to_mprj_in_buffers\[78\]_A user_to_mprj_in_gates\[78\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[101\]_B user_to_mprj_in_gates\[101\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[51\]_A _515_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_1813 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xmprj_dat_buf\[8\] _440_/Y mprj_dat_buf\[8\]/TE vssd vccd mprj_dat_o_user[8] vssd
+ vccd sky130_fd_sc_hd__einvp_8
XANTENNA__330__A _330_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_1475 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_1857 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1381 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2029 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[70\]_A_N _333_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_2020 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_273 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[85\]_A_N _348_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[10\]_A input551/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_925 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1341 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_1915 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[116\]_A user_to_mprj_in_gates\[116\]/Y vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_1817 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1828 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[105\]_A _569_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__505__A _505_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_693 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_buffers\[69\]_A user_to_mprj_in_gates\[69\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_10_1503 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_77 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1547 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[42\]_A _506_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_859 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[71\] _334_/Y mprj_logic_high_inst/HI[273] vssd vccd la_oenb_core[71]
+ vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[93\] _356_/A la_buf_enable\[93\]/B vssd vccd la_buf\[93\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XANTENNA_la_buf_enable\[23\]_A_N _615_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[60\]_B la_buf_enable\[60\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_1301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input337_A la_iena_mprj[54] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[38\]_A_N _630_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_1643 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1873 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[79\] _543_/Y la_buf\[79\]/TE vssd vccd la_data_in_core[79] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input504_A la_oenb_mprj[8] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_741 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_443 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_785 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_2006 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_498 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[107\]_A user_to_mprj_in_gates\[107\]/Y vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_671 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__415__A _415_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_697 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[33\]_A _497_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_2305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output723_A output723/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[51\]_B la_buf_enable\[51\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_391 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_380 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_2349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_1565 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1615 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[68\] input96/X user_to_mprj_in_gates\[68\]/B vssd vccd user_to_mprj_in_gates\[68\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_4_2073 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_229 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[123\]_B mprj_logic_high_inst/HI[453] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_37_1661 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_435 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_273 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1009 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[24\]_A _488_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[42\]_B la_buf_enable\[42\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput218 la_data_out_mprj[62] vssd vccd _526_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput207 la_data_out_mprj[52] vssd vccd _516_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_9_1283 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput229 la_data_out_mprj[72] vssd vccd _536_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_29_535 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1996 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[30\] input311/X mprj_logic_high_inst/HI[360] vssd vccd user_to_mprj_in_gates\[30\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_in_ena_buf\[114\]_B mprj_logic_high_inst/HI[444] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_38_2137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_601 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input287_A la_iena_mprj[124] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[15\]_A _479_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_645 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input454_A la_oenb_mprj[44] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_1399 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[33\]_B la_buf_enable\[33\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input50_A la_data_out_core[26] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1587 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[2\]_A input310/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input621_A user_irq_core[0] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_1957 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[100\]_A _363_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_2257 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[105\]_B mprj_logic_high_inst/HI[435] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_30_221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[38\] user_to_mprj_in_gates\[38\]/Y vssd vccd output686/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_34_1845 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_777 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output673_A output673/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_2281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_461 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[24\]_B la_buf_enable\[24\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_1649 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_1941 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1805 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2063 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1412 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_321 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_833 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1849 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_877 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_357 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1901 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[93\]_A _356_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_2067 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1945 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1989 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1675 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[15\]_B la_buf_enable\[15\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[78\] input363/X mprj_logic_high_inst/HI[408] vssd vccd user_to_mprj_in_gates\[78\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
Xuser_to_mprj_oen_buffers\[104\] _367_/Y mprj_logic_high_inst/HI[306] vssd vccd la_oenb_core[104]
+ vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_ena_buf\[94\]_B mprj_logic_high_inst/HI[424] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
X_630_ _630_/A vssd vccd _630_/Y vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_29_365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1771 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_561_ _561_/A vssd vccd _561_/Y vssd vccd sky130_fd_sc_hd__clkinv_4
Xuser_to_mprj_oen_buffers\[34\] _626_/Y mprj_logic_high_inst/HI[236] vssd vccd la_oenb_core[34]
+ vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[56\] _648_/A la_buf_enable\[56\]/B vssd vccd la_buf\[56\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_2_1821 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_346 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_53 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_711 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input202_A la_data_out_mprj[48] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_492_ _492_/A vssd vccd _492_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_53_1709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_1829 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_97 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2145 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[118\]_TE mprj_logic_high_inst/HI[320] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[84\]_A _347_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_1433 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input98_A la_data_out_core[6] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input571_A mprj_dat_i_user[29] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_932 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2041 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1130 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2085 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_69 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1936 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1204 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_107 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1721 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1765 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput582 mprj_dat_o_core[0] vssd vccd _432_/A vssd vccd sky130_fd_sc_hd__clkbuf_8
Xinput560 mprj_dat_i_user[19] vssd vccd input560/X vssd vccd sky130_fd_sc_hd__buf_8
Xinput571 mprj_dat_i_user[29] vssd vccd input571/X vssd vccd sky130_fd_sc_hd__clkbuf_16
XANTENNA_user_to_mprj_in_ena_buf\[85\]_B mprj_logic_high_inst/HI[415] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_36_825 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput593 mprj_dat_o_core[1] vssd vccd _433_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_1_1353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_869 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_2098 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output790_A output790/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[32\]_TE la_buf\[32\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_571 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[17\]_TE mprj_logic_high_inst/HI[219] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[75\]_A _338_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1951 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__603__A _603_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_1995 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1507 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[2\]_A input572/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_1457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1793 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[76\]_B mprj_logic_high_inst/HI[406] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_39_641 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_2221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[2\]_A input54/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_850 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[66\]_A _329_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_1704 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[0\]_TE la_buf\[0\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_55 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__513__A _513_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_2225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1483 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_2269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_946 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_456 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_405 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input152_A la_data_out_mprj[118] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[67\]_B mprj_logic_high_inst/HI[397] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_2_2341 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_613_ _613_/A vssd vccd _613_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_input417_A la_oenb_mprj[126] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[55\]_TE la_buf\[55\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input13_A la_data_out_core[108] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[61\] _525_/Y la_buf\[61\]/TE vssd vccd la_data_in_core[61] vssd vccd sky130_fd_sc_hd__einvp_8
X_544_ _544_/A vssd vccd _544_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_2_1695 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_475_ _475_/A vssd vccd _475_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_53_1506 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_1659 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[57\]_A _649_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_523 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1837 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xmprj_adr_buf\[25\] _425_/Y mprj_adr_buf\[25\]/TE vssd vccd mprj_adr_o_user[25] vssd
+ vccd sky130_fd_sc_hd__einvp_8
XANTENNA__423__A _423_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_773 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_1001 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output636_A output636/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1045 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2252 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1619 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_1089 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1933 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[58\]_B mprj_logic_high_inst/HI[388] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[50\] input77/X user_to_mprj_in_gates\[50\]/B vssd vccd user_to_mprj_in_gates\[50\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
Xinput390 la_oenb_mprj[101] vssd vccd _364_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_3_1437 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1005 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_861 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[48\]_A _640_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__333__A _333_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[78\]_TE la_buf\[78\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_1359 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input5_A la_data_out_core[100] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1590 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[49\]_B mprj_logic_high_inst/HI[379] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_41_2177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XPHY_22 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_11 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_2084 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XPHY_55 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_44 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_33 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__508__A _508_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_102 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_327 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XPHY_88 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_77 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_66 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_669 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_99 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[39\]_A _631_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_1225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xla_buf_enable\[19\] _611_/A la_buf_enable\[19\]/B vssd vccd la_buf\[19\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_13_1589 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input367_A la_iena_mprj[81] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_irq_gates\[2\] input623/X user_irq_gates\[2\]/B vssd vccd user_irq_gates\[2\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_46_2088 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input534_A mprj_adr_o_core[25] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2331 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_1365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1871 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[124\] _387_/A la_buf_enable\[124\]/B vssd vccd la_buf\[124\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_24_1663 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[27\]_TE mprj_dat_buf\[27\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_2182 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_655 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_441 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1481 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_527_ _527_/A vssd vccd _527_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA__418__A _418_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[6\]_TE mprj_logic_high_inst/HI[208] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
X_458_ _458_/A vssd vccd _458_/Y vssd vccd sky130_fd_sc_hd__inv_4
XFILLER_31_2324 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_331 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_389_ _389_/A vssd vccd _389_/Y vssd vccd sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_buffers\[20\] user_to_mprj_in_gates\[20\]/Y vssd vccd output667/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_output753_A output753/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[98\] input129/X user_to_mprj_in_gates\[98\]/B vssd vccd user_to_mprj_in_gates\[98\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_29_2286 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_mprj_adr_buf\[26\]_A _426_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_909 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[111\]_A_N _374_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_1201 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_953 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1267 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[126\]_A_N _389_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_669 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2235 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_466 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_319 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[3\]_A _595_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_1409 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1589 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1917 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_529 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xoutput661 output661/A vssd vccd la_data_in_mprj[15] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput672 output672/A vssd vccd la_data_in_mprj[25] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput650 output650/A vssd vccd la_data_in_mprj[120] vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_8_1123 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xoutput683 output683/A vssd vccd la_data_in_mprj[35] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput694 output694/A vssd vccd la_data_in_mprj[45] vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA_mprj_adr_buf\[17\]_A _417_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[60\] input344/X mprj_logic_high_inst/HI[390] vssd vccd user_to_mprj_in_gates\[60\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_43_1549 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_mprj_sel_buf\[1\]_TE mprj_sel_buf\[1\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_1994 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_953 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_901 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input115_A la_data_out_core[85] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1509 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_499 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1033 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1787 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1607 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_802 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_97 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1099 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input484_A la_oenb_mprj[71] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input80_A la_data_out_core[53] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput18 la_data_out_core[112] vssd vccd input18/X vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_6_301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_190 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1965 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xla_buf\[24\] _488_/Y la_buf\[24\]/TE vssd vccd la_data_in_core[24] vssd vccd sky130_fd_sc_hd__einvp_8
Xinput29 la_data_out_core[122] vssd vccd input29/X vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_6_345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_389 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_irq_buffers\[0\]_A user_irq_gates\[0\]/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_584 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1703 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1769 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1565 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[68\] user_to_mprj_in_gates\[68\]/Y vssd vccd output719/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_45_293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1832 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_gates\[26\] input568/X user_wb_ack_gate/B vssd vccd user_wb_dat_gates\[26\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_4
Xuser_to_mprj_in_gates\[13\] input36/X user_to_mprj_in_gates\[13\]/B vssd vccd user_to_mprj_in_gates\[13\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_33_1729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_wb_dat_buffers\[23\] user_wb_dat_gates\[23\]/Y vssd vccd output771/A vssd vccd
+ sky130_fd_sc_hd__inv_6
XANTENNA__611__A _611_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_1393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_80 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1869 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[124\] input31/X user_to_mprj_in_gates\[124\]/B vssd vccd user_to_mprj_in_gates\[124\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_37_761 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1031 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2032 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[10\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_2076 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1927 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[103\]_TE la_buf\[103\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[18\]_TE mprj_adr_buf\[18\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_1559 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[2\]_TE mprj_adr_buf\[2\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__521__A _521_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_2025 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1313 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[64\] _656_/Y mprj_logic_high_inst/HI[266] vssd vccd la_oenb_core[64]
+ vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[86\] _349_/A la_buf_enable\[86\]/B vssd vccd la_buf\[86\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_43_1357 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[12\] _444_/Y mprj_dat_buf\[12\]/TE vssd vccd mprj_dat_o_user[12] vssd
+ vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input232_A la_data_out_mprj[75] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_cyc_buf_A _393_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_1841 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1655 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1885 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_411 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_455 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2018 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_797 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[50\]_TE mprj_logic_high_inst/HI[252] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_694 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__431__A _431_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[121\] user_to_mprj_in_gates\[121\]/Y vssd vccd output651/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_mprj_dat_buf\[6\]_TE mprj_dat_buf\[6\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_2317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output716_A output716/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[126\]_TE la_buf\[126\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_1905 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__606__A _606_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_1673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_981 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[2\]_A _402_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__341__A _341_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_819 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2209 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xinput208 la_data_out_mprj[53] vssd vccd _517_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput219 la_data_out_mprj[63] vssd vccd _527_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
XANTENNA_user_wb_dat_buffers\[28\]_A user_wb_dat_gates\[28\]/Y vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XFILLER_9_1251 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1295 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_547 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1931 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[23\] input303/X mprj_logic_high_inst/HI[353] vssd vccd user_to_mprj_in_gates\[23\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_oen_buffers\[73\]_TE mprj_logic_high_inst/HI[275] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__516__A _516_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_1161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_447 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1637 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1047 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_613 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input182_A la_data_out_mprj[2] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_657 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_145 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input447_A la_oenb_mprj[38] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input43_A la_data_out_core[1] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_1831 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_1121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[2\]_B mprj_logic_high_inst/HI[332] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_buffers\[19\]_A user_wb_dat_gates\[19\]/Y vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
Xla_buf\[91\] _555_/Y la_buf\[91\]/TE vssd vccd la_data_in_core[91] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input614_A mprj_iena_wb vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_1693 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__426__A _426_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output666_A output666/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_473 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_2125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[80\] input110/X user_to_mprj_in_gates\[80\]/B vssd vccd user_to_mprj_in_gates\[80\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_45_1953 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[84\]_A_N _347_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_2075 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1424 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1817 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_377 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[96\]_TE mprj_logic_high_inst/HI[298] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[123\]_B la_buf_enable\[123\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_889 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1713 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[99\]_A_N _362_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[22\]_A_N _614_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_2057 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1913 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_244 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__336__A _336_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_907 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[92\]_A input123/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_1979 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[37\]_A_N _629_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_609 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_1441 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_377 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_560_ _560_/A vssd vccd _560_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_la_buf_enable\[114\]_B la_buf_enable\[114\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_1833 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1877 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1783 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_358 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_oen_buffers\[27\] _619_/Y mprj_logic_high_inst/HI[229] vssd vccd la_oenb_core[27]
+ vssd vccd sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[9\] _601_/Y mprj_logic_high_inst/HI[211] vssd vccd la_oenb_core[9]
+ vssd vccd sky130_fd_sc_hd__einvp_8
X_491_ _491_/A vssd vccd _491_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
Xla_buf_enable\[49\] _641_/A la_buf_enable\[49\]/B vssd vccd la_buf\[49\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_53_881 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_65 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_723 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input397_A la_oenb_mprj[108] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_buffers\[5\]_A user_wb_dat_gates\[5\]/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_1565 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[83\]_A input113/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_1445 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xla_buf\[2\] _466_/Y la_buf\[2\]/TE vssd vccd la_data_in_core[2] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input564_A mprj_dat_i_user[22] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_2053 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1142 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_421 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_944 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_1175 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1733 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1788 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1619 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput550 mprj_dat_i_user[0] vssd vccd input550/X vssd vccd sky130_fd_sc_hd__buf_8
Xinput561 mprj_dat_i_user[1] vssd vccd input561/X vssd vccd sky130_fd_sc_hd__buf_8
Xinput572 mprj_dat_i_user[2] vssd vccd input572/X vssd vccd sky130_fd_sc_hd__buf_8
XANTENNA_la_buf\[8\]_A _472_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_837 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput594 mprj_dat_o_core[20] vssd vccd _452_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
XANTENNA_la_buf_enable\[105\]_B la_buf_enable\[105\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput583 mprj_dat_o_core[10] vssd vccd _442_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_39_1009 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_buffers\[50\] user_to_mprj_in_gates\[50\]/Y vssd vccd output700/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_output783_A output783/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1632 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1621 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1665 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[74\]_A input103/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1963 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1425 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1469 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[2\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1761 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_130 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1287 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[2\]_B user_to_mprj_in_gates\[2\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_39_1565 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_862 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[65\]_A input93/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[90\] input377/X mprj_logic_high_inst/HI[420] vssd vccd user_to_mprj_in_gates\[90\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_46_2237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_925 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input145_A la_data_out_mprj[111] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_163 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_601 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_612_ _612_/A vssd vccd _612_/Y vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_input312_A la_iena_mprj[31] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_543_ _543_/A vssd vccd _543_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_53_2219 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_474_ _474_/A vssd vccd _474_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_13_531 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[126\] input289/X mprj_logic_high_inst/HI[456] vssd vccd
+ user_to_mprj_in_gates\[126\]/B vssd vccd sky130_fd_sc_hd__and2_1
Xla_buf\[54\] _518_/Y la_buf\[54\]/TE vssd vccd la_data_in_core[54] vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_35_1941 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1974 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1805 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[56\]_A input83/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1849 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_785 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[110\] _574_/Y la_buf\[110\]/TE vssd vccd la_data_in_core[110] vssd vccd sky130_fd_sc_hd__einvp_8
Xmprj_adr_buf\[18\] _418_/Y mprj_adr_buf\[18\]/TE vssd vccd mprj_adr_o_user[18] vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_7_2264 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1901 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1057 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_buffers\[98\] user_to_mprj_in_gates\[98\]/Y vssd vccd output752/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_output629_A output629/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_1945 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1989 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_601 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1416 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput380 la_iena_mprj[93] vssd vccd input380/X vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_36_645 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[6\]_A user_to_mprj_in_gates\[6\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xinput391 la_oenb_mprj[102] vssd vccd _365_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
Xuser_to_mprj_in_gates\[43\] input69/X user_to_mprj_in_gates\[43\]/B vssd vccd user_to_mprj_in_gates\[43\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_2
Xuser_wb_dat_buffers\[8\] user_wb_dat_gates\[8\]/Y vssd vccd output786/A vssd vccd
+ sky130_fd_sc_hd__clkinv_8
XFILLER_16_391 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1017 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_895 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[47\]_A input73/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_2185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__614__A _614_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_1771 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[5\] input87/X user_to_mprj_in_gates\[5\]/B vssd vccd user_to_mprj_in_gates\[5\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_4
XFILLER_45_2281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[108\]_TE mprj_logic_high_inst/HI[310] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_461 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1051 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1972 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_12 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_56 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_45 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_23 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_34 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_637 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XPHY_89 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_78 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_67 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1248 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_383 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[38\]_A input63/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[122\]_A input29/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__524__A _524_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1609 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[94\] _357_/Y mprj_logic_high_inst/HI[296] vssd vccd la_oenb_core[94]
+ vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input262_A la_iena_mprj[101] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_733 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[22\]_TE la_buf\[22\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_1907 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_1631 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[7\] input365/X mprj_logic_high_inst/HI[337] vssd vccd user_to_mprj_in_gates\[7\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_input527_A mprj_adr_o_core[19] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_1883 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[117\] _380_/A la_buf_enable\[117\]/B vssd vccd la_buf\[117\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_24_1675 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_667 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_497 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_526_ _526_/A vssd vccd _526_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_20_309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_457_ _457_/A vssd vccd _457_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_31_2336 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_343 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_388_ _388_/A vssd vccd _388_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_user_to_mprj_in_gates\[29\]_A input53/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_1793 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__434__A _434_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[113\]_A input19/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1613 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[13\] user_to_mprj_in_gates\[13\]/Y vssd vccd output659/A
+ vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_29_2210 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output746_A output746/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_593 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_409 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_943 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_965 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__609__A _609_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_497 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2247 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_478 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[104\]_A input9/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__344__A _344_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1134 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[45\]_TE la_buf\[45\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1929 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xoutput662 output662/A vssd vccd la_data_in_mprj[16] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput640 output640/A vssd vccd la_data_in_mprj[111] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput651 output651/A vssd vccd la_data_in_mprj[121] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput673 output673/A vssd vccd la_data_in_mprj[26] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput684 output684/A vssd vccd la_data_in_mprj[36] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput695 output695/A vssd vccd la_data_in_mprj[46] vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_8_1135 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[53\] input336/X mprj_logic_high_inst/HI[383] vssd vccd user_to_mprj_in_gates\[53\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_28_921 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1909 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_965 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__519__A _519_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_913 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_497 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input108_A la_data_out_core[79] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[5\] user_to_mprj_in_gates\[5\]/Y vssd vccd output710/A vssd
+ vccd sky130_fd_sc_hd__clkinv_4
Xla_buf_enable\[31\] _623_/A la_buf_enable\[31\]/B vssd vccd la_buf\[31\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_19_1799 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_1619 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1933 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput19 la_data_out_core[113] vssd vccd input19/X vssd vccd sky130_fd_sc_hd__clkbuf_4
XANTENNA_input477_A la_oenb_mprj[65] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf\[17\] _481_/Y la_buf\[17\]/TE vssd vccd la_data_in_core[17] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input73_A la_data_out_core[47] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_357 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_1715 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1005 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1049 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2195 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1691 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1577 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__429__A _429_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_209 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1844 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_629 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output696_A output696/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_509_ _509_/A vssd vccd _509_/Y vssd vccd sky130_fd_sc_hd__inv_2
XANTENNA_la_buf\[68\]_TE la_buf\[68\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_gates\[19\] input560/X user_wb_ack_gate/B vssd vccd user_wb_dat_gates\[19\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_4
XFILLER_6_891 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_buffers\[16\] user_wb_dat_gates\[16\]/Y vssd vccd output763/A vssd vccd
+ sky130_fd_sc_hd__clkinv_4
XANTENNA_la_buf_enable\[2\]_B la_buf_enable\[2\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_2095 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2009 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_92 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[117\] input23/X user_to_mprj_in_gates\[117\]/B vssd vccd user_to_mprj_in_gates\[117\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XANTENNA_user_to_mprj_in_ena_buf\[126\]_A input289/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_1583 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1043 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__339__A _339_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_1065 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_905 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_607 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2088 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_489 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1939 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[17\]_TE mprj_dat_buf\[17\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_oen_buffers\[127\] _390_/Y mprj_logic_high_inst/HI[329] vssd vccd la_oenb_core[127]
+ vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_43_2037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[57\] _649_/Y mprj_logic_high_inst/HI[259] vssd vccd la_oenb_core[57]
+ vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[79\] _342_/A la_buf_enable\[79\]/B vssd vccd la_buf\[79\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_43_1369 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[117\]_A input279/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input225_A la_data_out_mprj[69] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_795 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1897 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_721 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_467 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input594_A mprj_dat_o_core[20] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_1329 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[110\]_A_N _373_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[125\]_A_N _388_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[114\] user_to_mprj_in_gates\[114\]/Y vssd vccd output643/A
+ vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_38_537 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output709_A output709/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[108\]_A input269/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[80\] user_to_mprj_in_gates\[80\]/Y vssd vccd output733/A
+ vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_4_1341 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_529 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_518 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1385 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2217 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_993 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1803 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__622__A _622_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput209 la_data_out_mprj[54] vssd vccd _518_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_42_2081 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1943 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_713 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1703 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_404 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[16\] input295/X mprj_logic_high_inst/HI[346] vssd vccd user_to_mprj_in_gates\[16\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_40_768 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_459 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[30\]_A input311/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_757 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1649 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1173 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1747 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1059 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__532__A _532_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input175_A la_data_out_mprj[23] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_669 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input342_A la_iena_mprj[59] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[97\]_A input384/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_1133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1887 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input36_A la_data_out_core[13] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_2237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_1177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[84\] _548_/Y la_buf\[84\]/TE vssd vccd la_data_in_core[84] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input607_A mprj_dat_o_core[3] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_573 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_275 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[21\]_A input301/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_245 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_931 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_492 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1593 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output659_A output659/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__442__A _442_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[73\] input102/X user_to_mprj_in_gates\[73\]/B vssd vccd user_to_mprj_in_gates\[73\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XANTENNA_user_to_mprj_in_ena_buf\[88\]_A input374/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_1829 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_389 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1013 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__617__A _617_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_1725 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_713 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1925 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[12\]_A input291/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_1313 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_256 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[92\]_B user_to_mprj_in_gates\[92\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA__352__A _352_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[79\]_A input364/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_1453 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1497 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[40\]_TE mprj_logic_high_inst/HI[242] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_1812 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1981 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_389 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_1856 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_1795 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__527__A _527_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_490_ _490_/A vssd vccd _490_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_25_573 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_77 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_735 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input292_A la_iena_mprj[13] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[83\]_B user_to_mprj_in_gates\[83\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_5_27 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_433 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input557_A mprj_dat_i_user[16] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_1905 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1154 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2065 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[116\]_TE la_buf\[116\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_2170 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput540 mprj_adr_o_core[30] vssd vccd _430_/A vssd vccd sky130_fd_sc_hd__buf_2
Xinput551 mprj_dat_i_user[10] vssd vccd input551/X vssd vccd sky130_fd_sc_hd__buf_8
Xinput562 mprj_dat_i_user[20] vssd vccd input562/X vssd vccd sky130_fd_sc_hd__clkbuf_16
Xinput573 mprj_dat_i_user[30] vssd vccd input573/X vssd vccd sky130_fd_sc_hd__buf_12
Xinput595 mprj_dat_o_core[21] vssd vccd _453_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput584 mprj_dat_o_core[11] vssd vccd _443_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_35_337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__437__A _437_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_551 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_521 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[43\] user_to_mprj_in_gates\[43\]/Y vssd vccd output692/A
+ vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_31_565 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output776_A output776/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1644 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1677 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[74\]_B user_to_mprj_in_gates\[74\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_8_783 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[63\]_TE mprj_logic_high_inst/HI[265] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1773 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__347__A _347_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_17_1831 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_727 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1154 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1777 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[65\]_B user_to_mprj_in_gates\[65\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_46_2249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[83\] input369/X mprj_logic_high_inst/HI[413] vssd vccd user_to_mprj_in_gates\[83\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_49_429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_613 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_611_ _611_/A vssd vccd _611_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
Xla_buf_enable\[61\] _653_/A la_buf_enable\[61\]/B vssd vccd la_buf\[61\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XANTENNA_user_to_mprj_in_buffers\[50\]_A user_to_mprj_in_gates\[50\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_input138_A la_data_out_mprj[105] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_17_359 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_819 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_542_ _542_/A vssd vccd _542_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_input305_A la_iena_mprj[25] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_1686 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_189 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_473_ _473_/A vssd vccd _473_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_13_543 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_340 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[47\] _511_/Y la_buf\[47\]/TE vssd vccd la_data_in_core[47] vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_35_1986 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1817 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_587 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[119\] input281/X mprj_logic_high_inst/HI[449] vssd vccd
+ user_to_mprj_in_gates\[119\]/B vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_in_gates\[56\]_B user_to_mprj_in_gates\[56\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[83\]_A_N _346_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_1953 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[90\]_A _554_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[98\]_A_N _361_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[86\]_TE mprj_logic_high_inst/HI[288] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_797 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[103\] _567_/Y la_buf\[103\]/TE vssd vccd la_data_in_core[103] vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_27_2160 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[21\]_A_N _613_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_1913 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_992 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1957 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[41\]_A user_to_mprj_in_gates\[41\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xinput370 la_iena_mprj[84] vssd vccd input370/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput381 la_iena_mprj[94] vssd vccd input381/X vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_3_1428 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_613 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput392 la_oenb_mprj[103] vssd vccd _366_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_1_1152 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[36\]_A_N _628_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[36\] input61/X user_to_mprj_in_gates\[36\]/B vssd vccd user_to_mprj_in_gates\[36\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_52_1029 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1441 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[47\]_B user_to_mprj_in_gates\[47\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1463 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[81\]_A _545_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__630__A _630_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_1245 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1063 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[32\]_A user_to_mprj_in_gates\[32\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_39_440 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_473 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_13 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_189 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XPHY_46 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_35 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_24 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1937 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XPHY_79 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_68 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_57 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_57 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_693 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_buffers\[99\]_A user_to_mprj_in_gates\[99\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[38\]_B user_to_mprj_in_gates\[38\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_52_1574 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[122\]_B user_to_mprj_in_gates\[122\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[72\]_A _536_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[90\]_B la_buf_enable\[90\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_200 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1009 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1271 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[87\] _350_/Y mprj_logic_high_inst/HI[289] vssd vccd la_oenb_core[87]
+ vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA__540__A _540_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_211 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input255_A la_data_out_mprj[96] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_39 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input422_A la_oenb_mprj[15] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[23\]_A user_to_mprj_in_gates\[23\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_8_1895 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_1687 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_wb_dat_gates\[31\]_A input574/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_525_ _525_/A vssd vccd _525_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_53_2028 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_456_ _456_/A vssd vccd _456_/Y vssd vccd sky130_fd_sc_hd__inv_4
XANTENNA_la_buf\[126\]_A _590_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_387_ _387_/A vssd vccd _387_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_31_2348 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[113\]_B user_to_mprj_in_gates\[113\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[29\]_B user_to_mprj_in_gates\[29\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_9_355 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xmprj_adr_buf\[30\] _430_/Y mprj_adr_buf\[30\]/TE vssd vccd mprj_adr_o_user[30] vssd
+ vccd sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf\[63\]_A _527_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_2222 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output641_A output641/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__450__A _450_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[81\]_B la_buf_enable\[81\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output739_A output739/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_1721 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2073 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2062 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_buffers\[14\]_A user_to_mprj_in_gates\[14\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_42_1765 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_977 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_432 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_925 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[22\]_A input564/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[117\]_A _581_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_2259 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__625__A _625_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[104\]_B user_to_mprj_in_gates\[104\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[54\]_A _518_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_1591 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[72\]_B la_buf_enable\[72\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput652 output652/A vssd vccd la_data_in_mprj[122] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput663 output663/A vssd vccd la_data_in_mprj[17] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput630 output630/A vssd vccd la_data_in_mprj[102] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput641 output641/A vssd vccd la_data_in_mprj[112] vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA__360__A _360_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_wb_ena_buf_A input614/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_1031 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1103 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xoutput674 output674/A vssd vccd la_data_in_mprj[27] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput685 output685/A vssd vccd la_data_in_mprj[37] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput696 output696/A vssd vccd la_data_in_mprj[47] vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA_mprj_stb_buf_A _394_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_1147 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1097 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[46\] input328/X mprj_logic_high_inst/HI[376] vssd vccd user_to_mprj_in_gates\[46\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_28_977 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1781 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_925 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[13\]_A input554/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[119\]_A user_to_mprj_in_gates\[119\]/Y vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[108\]_A _572_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_833 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xla_buf_enable\[24\] _616_/A la_buf_enable\[24\]/B vssd vccd la_buf\[24\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XANTENNA__535__A _535_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_1945 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[45\]_A _509_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_387 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input372_A la_iena_mprj[86] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[63\]_B la_buf_enable\[63\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input66_A la_data_out_core[40] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_597 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_1727 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_925 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_402 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1589 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_273 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_508_ _508_/A vssd vccd _508_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
X_439_ _439_/A vssd vccd _439_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_output689_A output689/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__445__A _445_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[36\]_A _500_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1444 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_881 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[54\]_B la_buf_enable\[54\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_2041 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[121\]_A _384_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[126\]_B mprj_logic_high_inst/HI[456] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_37_741 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_785 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_240 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1088 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1055 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1077 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[12\]_TE la_buf\[12\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_917 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_991 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__355__A _355_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_641 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[27\]_A _491_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[45\]_B la_buf_enable\[45\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1749 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2152 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_328 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_2185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2049 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[112\]_A _375_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_11 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[117\]_B mprj_logic_high_inst/HI[447] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_28_741 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input218_A la_data_out_mprj[62] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input120_A la_data_out_core[8] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_273 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input587_A mprj_dat_o_core[14] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[18\]_A _482_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_645 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[101\] input262/X mprj_logic_high_inst/HI[431] vssd vccd
+ user_to_mprj_in_gates\[101\]/B vssd vccd sky130_fd_sc_hd__and2_1
Xuser_wb_dat_gates\[1\] input561/X user_wb_ack_gate/B vssd vccd user_wb_dat_gates\[1\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_8
XFILLER_6_177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[36\]_B la_buf_enable\[36\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[5\]_A input343/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[103\]_A _366_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[107\] user_to_mprj_in_gates\[107\]/Y vssd vccd output635/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_38_505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1579 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[108\]_B mprj_logic_high_inst/HI[438] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_4_1353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_549 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[73\] user_to_mprj_in_gates\[73\]/Y vssd vccd output725/A
+ vssd vccd sky130_fd_sc_hd__inv_2
XANTENNA_la_buf\[35\]_TE la_buf\[35\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_1397 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_gates\[31\] input574/X user_wb_ack_gate/B vssd vccd user_wb_dat_gates\[31\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_2
XFILLER_21_449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1815 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[27\]_B la_buf_enable\[27\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_2325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[6\] _438_/Y mprj_dat_buf\[6\]/TE vssd vccd mprj_dat_o_user[6] vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_44_1657 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1128 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2093 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_1955 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_210 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_733 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[96\]_A _359_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_725 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_416 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1715 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[30\]_B mprj_logic_high_inst/HI[360] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_36_1185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1759 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[3\]_TE la_buf\[3\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_482 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[18\]_B la_buf_enable\[18\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_637 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1369 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input168_A la_data_out_mprj[17] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[91\] _354_/A la_buf_enable\[91\]/B vssd vccd la_buf\[91\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XANTENNA_user_to_mprj_oen_buffers\[20\]_A _612_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_1905 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[97\]_B mprj_logic_high_inst/HI[427] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_43_1145 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1899 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input335_A la_iena_mprj[52] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[58\]_TE la_buf\[58\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_1719 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_869 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1189 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input29_A la_data_out_core[122] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf\[77\] _541_/Y la_buf\[77\]/TE vssd vccd la_data_in_core[77] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input502_A la_oenb_mprj[88] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[87\]_A _350_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_585 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_287 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[21\]_B mprj_logic_high_inst/HI[351] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_8_943 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1900 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output721_A output721/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[11\]_A _603_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_803 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[88\]_B mprj_logic_high_inst/HI[418] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_24_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[66\] input94/X user_to_mprj_in_gates\[66\]/B vssd vccd user_to_mprj_in_gates\[66\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_4_1161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_357 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_725 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[78\]_A _341_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[12\]_B mprj_logic_high_inst/HI[342] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_33_1325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_268 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__633__A _633_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_1623 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[5\]_A input577/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[79\]_B mprj_logic_high_inst/HI[409] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_44_1465 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1072 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1329 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1307 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_79 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[5\]_A input87/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_1868 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_585 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[124\]_A_N _387_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[69\]_A _332_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_279 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1469 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__543__A _543_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input285_A la_iena_mprj[122] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_957 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1917 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_39 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_445 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input452_A la_oenb_mprj[42] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_1166 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_611 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1663 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput530 mprj_adr_o_core[21] vssd vccd _421_/A vssd vccd sky130_fd_sc_hd__buf_2
Xinput541 mprj_adr_o_core[31] vssd vccd _431_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput552 mprj_dat_i_user[11] vssd vccd input552/X vssd vccd sky130_fd_sc_hd__buf_12
Xinput563 mprj_dat_i_user[21] vssd vccd input563/X vssd vccd sky130_fd_sc_hd__buf_12
XFILLER_48_677 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xinput596 mprj_dat_o_core[22] vssd vccd _454_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput574 mprj_dat_i_user[31] vssd vccd input574/X vssd vccd sky130_fd_sc_hd__buf_12
Xinput585 mprj_dat_o_core[12] vssd vccd _444_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_51_809 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[9\]_TE mprj_logic_high_inst/HI[211] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_1_1389 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_533 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_577 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[36\] user_to_mprj_in_gates\[36\]/Y vssd vccd output684/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_output671_A output671/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output769_A output769/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__453__A _453_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1689 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2081 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_751 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_600 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1785 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__628__A _628_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_872 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_533 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1843 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_1887 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_739 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__363__A _363_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_2181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_209 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[76\] input361/X mprj_logic_high_inst/HI[406] vssd vccd user_to_mprj_in_gates\[76\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_28_1961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1273 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[102\] _365_/Y mprj_logic_high_inst/HI[304] vssd vccd la_oenb_core[102]
+ vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_44_1251 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
X_610_ _610_/A vssd vccd _610_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
Xuser_to_mprj_oen_buffers\[32\] _624_/Y mprj_logic_high_inst/HI[234] vssd vccd la_oenb_core[32]
+ vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA__538__A _538_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_1632 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
X_541_ _541_/A vssd vccd _541_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_2_1643 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xla_buf_enable\[54\] _646_/A la_buf_enable\[54\]/B vssd vccd la_buf\[54\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XANTENNA_input200_A la_data_out_mprj[46] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_472_ _472_/A vssd vccd _472_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_18_1629 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_511 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_853 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_mprj_dat_buf\[20\]_A _452_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_691 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_352 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_555 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_190 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_599 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input96_A la_data_out_core[68] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_1998 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1829 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_721 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1819 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_953 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1565 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1969 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput360 la_iena_mprj[75] vssd vccd input360/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput371 la_iena_mprj[85] vssd vccd input371/X vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_36_625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput393 la_oenb_mprj[104] vssd vccd _367_/A vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA__448__A _448_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput382 la_iena_mprj[95] vssd vccd input382/X vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_51_617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_371 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[29\] input53/X user_to_mprj_in_gates\[29\]/B vssd vccd user_to_mprj_in_gates\[29\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XANTENNA_mprj_dat_buf\[11\]_A _443_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_691 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_2132 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1453 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_385 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1475 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[30\]_TE mprj_logic_high_inst/HI[232] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[29\]_A _429_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_1257 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_1457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_102 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1941 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1075 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__358__A _358_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XPHY_47 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_36 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_25 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_14 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1331 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[6\]_A _598_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XPHY_58 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_69 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_69 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[106\]_TE la_buf\[106\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_503 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_57 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1586 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_mprj_adr_buf\[5\]_TE mprj_adr_buf\[5\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_1283 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_757 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[28\] _460_/Y mprj_dat_buf\[28\]/TE vssd vccd mprj_dat_o_user[28] vssd
+ vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input150_A la_data_out_mprj[116] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input248_A la_data_out_mprj[8] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input415_A la_oenb_mprj[124] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_2163 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input11_A la_data_out_core[106] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_989 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[31\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_524_ _524_/A vssd vccd _524_/Y vssd vccd sky130_fd_sc_hd__inv_2
X_455_ _455_/A vssd vccd _455_/Y vssd vccd sky130_fd_sc_hd__inv_6
XFILLER_53_1317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[53\]_TE mprj_logic_high_inst/HI[255] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_363 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_386_ _386_/A vssd vccd _386_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_31_2305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_1773 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1637 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[23\] _423_/Y mprj_adr_buf\[23\]/TE vssd vccd mprj_adr_o_user[23] vssd
+ vccd sky130_fd_sc_hd__einvp_8
XANTENNA_mprj_dat_buf\[9\]_TE mprj_dat_buf\[9\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_573 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_2234 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output634_A output634/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_2041 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1733 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2085 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1777 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput190 la_data_out_mprj[37] vssd vccd _501_/A vssd vccd sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_444 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_937 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_989 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[22\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_691 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1840 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[8\] _600_/A la_buf_enable\[8\]/B vssd vccd la_buf\[8\]/TE vssd vccd
+ sky130_fd_sc_hd__and2b_1
XANTENNA__641__A _641_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_1600 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xoutput653 output653/A vssd vccd la_data_in_mprj[123] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput631 output631/A vssd vccd la_data_in_mprj[103] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput642 output642/A vssd vccd la_data_in_mprj[113] vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA_user_to_mprj_wb_ena_buf_B user_to_mprj_wb_ena_buf/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_2209 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_1115 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xoutput664 output664/A vssd vccd la_data_in_mprj[18] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput675 output675/A vssd vccd la_data_in_mprj[28] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput686 output686/A vssd vccd la_data_in_mprj[38] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput697 output697/A vssd vccd la_data_in_mprj[48] vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA_input3_A caravel_rstn vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_1065 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[82\]_A_N _345_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[91\]_TE la_buf\[91\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_1793 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[39\] input320/X mprj_logic_high_inst/HI[369] vssd vccd user_to_mprj_in_gates\[39\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_oen_buffers\[76\]_TE mprj_logic_high_inst/HI[278] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[13\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_937 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_425 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[97\]_A_N _360_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_2040 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_67 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_867 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[17\] _609_/A la_buf_enable\[17\]/B vssd vccd la_buf\[17\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XANTENNA_la_buf_enable\[20\]_A_N _612_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input198_A la_data_out_mprj[44] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_1957 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_399 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__551__A _551_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input365_A la_iena_mprj[7] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[35\]_A_N _627_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_irq_gates\[0\] input621/X user_irq_gates\[0\]/B vssd vccd user_irq_gates\[0\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XANTENNA_input59_A la_data_out_core[34] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_1739 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input532_A mprj_adr_o_core[23] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_2203 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_2225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[122\] _385_/A la_buf_enable\[122\]/B vssd vccd la_buf\[122\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_4_2269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_499 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_937 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_414 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_507_ _507_/A vssd vccd _507_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_42_981 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1114 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_438_ _438_/A vssd vccd _438_/Y vssd vccd sky130_fd_sc_hd__inv_2
X_369_ _369_/A vssd vccd _369_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_31_1401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output751_A output751/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__461__A _461_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_2053 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[96\] input127/X user_to_mprj_in_gates\[96\]/B vssd vccd user_to_mprj_in_gates\[96\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_42_2253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_219 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[99\]_TE mprj_logic_high_inst/HI[301] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_1181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_753 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_1883 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_797 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__636__A _636_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[5\]_A _405_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_1378 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1209 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__371__A _371_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_1698 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_2164 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_517 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_23 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1051 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_753 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input113_A la_data_out_core[83] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__546__A _546_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_613 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input482_A la_oenb_mprj[6] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_657 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[22\] _486_/Y la_buf\[22\]/TE vssd vccd la_data_in_core[22] vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_32_1787 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_189 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[5\]_B mprj_logic_high_inst/HI[335] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_3_841 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1861 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_517 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[66\] user_to_mprj_in_gates\[66\]/Y vssd vccd output717/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_mprj_stb_buf_TE mprj_stb_buf/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__456__A _456_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[11\] input26/X user_to_mprj_in_gates\[11\]/B vssd vccd user_to_mprj_in_gates\[11\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_2
Xuser_wb_dat_gates\[24\] input566/X user_wb_ack_gate/B vssd vccd user_wb_dat_gates\[24\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_2
XFILLER_50_1821 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_wb_dat_buffers\[21\] user_wb_dat_gates\[21\]/Y vssd vccd output769/A vssd vccd
+ sky130_fd_sc_hd__clkinv_8
XFILLER_44_2337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1182 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1669 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[122\] input29/X user_to_mprj_in_gates\[122\]/B vssd vccd user_to_mprj_in_gates\[122\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XANTENNA_la_buf_enable\[126\]_B la_buf_enable\[126\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_22_1967 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1691 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__366__A _366_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_428 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_47 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_1727 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[95\]_A input126/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_1197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1525 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_104 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_mprj_adr_buf\[31\]_TE mprj_adr_buf\[31\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_1917 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[62\] _654_/Y mprj_logic_high_inst/HI[264] vssd vccd la_oenb_core[62]
+ vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[84\] _347_/A la_buf_enable\[84\]/B vssd vccd la_buf\[84\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_43_1157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[10\] _442_/Y mprj_dat_buf\[10\]/TE vssd vccd mprj_dat_o_user[10] vssd
+ vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input230_A la_data_out_mprj[73] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[117\]_B la_buf_enable\[117\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_2353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1641 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input328_A la_iena_mprj[46] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_509 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_wb_dat_buffers\[8\]_A user_wb_dat_gates\[8\]/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_597 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1805 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[86\]_A input116/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_299 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_421 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_999 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xla_buf\[126\] _590_/Y la_buf\[126\]/TE vssd vccd la_data_in_core[126] vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_28_1609 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1871 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1079 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_682 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_303 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_815 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[10\]_A input15/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output714_A output714/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[108\]_B la_buf_enable\[108\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[59\] input86/X user_to_mprj_in_gates\[59\]/B vssd vccd user_to_mprj_in_gates\[59\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_19_572 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1173 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1705 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1749 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[77\]_A input106/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_2185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1635 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1679 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[5\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_2281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[5\]_B user_to_mprj_in_gates\[5\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_2_1847 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_501 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[21\] input301/X mprj_logic_high_inst/HI[351] vssd vccd user_to_mprj_in_gates\[21\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_25_553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[68\]_A input96/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_589 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1579 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input180_A la_data_out_mprj[28] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input278_A la_iena_mprj[116] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[25\]_TE la_buf\[25\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_969 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1929 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1631 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input445_A la_oenb_mprj[36] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input41_A la_data_out_core[18] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_1090 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1675 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput520 mprj_adr_o_core[12] vssd vccd _412_/A vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_48_645 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_623 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput531 mprj_adr_o_core[22] vssd vccd _422_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput542 mprj_adr_o_core[3] vssd vccd _403_/A vssd vccd sky130_fd_sc_hd__buf_2
Xinput553 mprj_dat_i_user[12] vssd vccd input553/X vssd vccd sky130_fd_sc_hd__buf_8
Xinput564 mprj_dat_i_user[22] vssd vccd input564/X vssd vccd sky130_fd_sc_hd__buf_12
XANTENNA_input612_A mprj_dat_o_core[8] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_2036 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xinput597 mprj_dat_o_core[23] vssd vccd _455_/A vssd vccd sky130_fd_sc_hd__buf_2
Xinput575 mprj_dat_i_user[3] vssd vccd input575/X vssd vccd sky130_fd_sc_hd__buf_6
Xinput586 mprj_dat_o_core[13] vssd vccd _445_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_1_2069 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_881 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_501 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[59\]_A input86/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_589 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[29\] user_to_mprj_in_gates\[29\]/Y vssd vccd output676/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_11_291 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_763 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output664_A output664/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_2093 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_612 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_buffers\[9\]_A user_to_mprj_in_gates\[9\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_38_177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_884 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_501 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1811 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_545 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__644__A _644_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_17_1855 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_589 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1719 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[48\]_TE la_buf\[48\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_1281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_2193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1899 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1167 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1189 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1590 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_57 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1973 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[69\] input353/X mprj_logic_high_inst/HI[399] vssd vccd user_to_mprj_in_gates\[69\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_40_1105 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_1285 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1859 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_1149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_540_ _540_/A vssd vccd _540_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_22_1594 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_339 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_2091 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[25\] _617_/Y mprj_logic_high_inst/HI[227] vssd vccd la_oenb_core[25]
+ vssd vccd sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[7\] _599_/Y mprj_logic_high_inst/HI[209] vssd vccd la_oenb_core[7]
+ vssd vccd sky130_fd_sc_hd__einvp_8
X_471_ _471_/A vssd vccd _471_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
Xla_buf_enable\[47\] _639_/A la_buf_enable\[47\]/B vssd vccd la_buf\[47\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_13_523 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1201 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_567 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__554__A _554_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[125\]_A input32/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input395_A la_oenb_mprj[106] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input89_A la_data_out_core[61] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_1289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[0\] _464_/Y la_buf\[0\]/TE vssd vccd la_data_in_core[0] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input562_A mprj_dat_i_user[20] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_1737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_2004 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_965 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput350 la_iena_mprj[66] vssd vccd input350/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput361 la_iena_mprj[76] vssd vccd input361/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput372 la_iena_mprj[86] vssd vccd input372/X vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_29_90 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput394 la_oenb_mprj[105] vssd vccd _368_/A vssd vccd sky130_fd_sc_hd__buf_4
Xinput383 la_iena_mprj[96] vssd vccd input383/X vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_36_637 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_629 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_383 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2144 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output781_A output781/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[116\]_A input22/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__464__A _464_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1329 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[123\]_A_N _386_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_1308 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1010 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__639__A _639_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_1087 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1469 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_114 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1953 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_497 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XPHY_26 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_37 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_59 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_48 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[107\]_A input12/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__374__A _374_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_515 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1554 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1663 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_559 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_69 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_2026 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_268 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2335 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_217 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input143_A la_data_out_mprj[10] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_2120 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__549__A _549_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_2153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_1093 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_615 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input310_A la_iena_mprj[2] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input408_A la_oenb_mprj[118] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_523_ _523_/A vssd vccd _523_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_26_681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_454_ _454_/A vssd vccd _454_/Y vssd vccd sky130_fd_sc_hd__inv_4
XFILLER_33_629 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_331 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[124\] input287/X mprj_logic_high_inst/HI[454] vssd vccd
+ user_to_mprj_in_gates\[124\]/B vssd vccd sky130_fd_sc_hd__and2_1
Xla_buf\[52\] _516_/Y la_buf\[52\]/TE vssd vccd la_data_in_core[52] vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_41_673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_385_ _385_/A vssd vccd _385_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_41_662 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_1763 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1785 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1649 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1501 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xmprj_adr_buf\[16\] _416_/Y mprj_adr_buf\[16\]/TE vssd vccd mprj_adr_o_user[16] vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_42_1701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_buffers\[96\] user_to_mprj_in_gates\[96\]/Y vssd vccd output750/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_output627_A output627/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_2097 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1341 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1745 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__459__A _459_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xmprj_rstn_buf input3/X mprj_rstn_buf/TE vssd vccd user_reset vssd vccd sky130_fd_sc_hd__einvp_8
Xinput180 la_data_out_mprj[28] vssd vccd _492_/A vssd vccd sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_42_1789 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput191 la_data_out_mprj[38] vssd vccd _502_/A vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_36_456 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[41\] input67/X user_to_mprj_in_gates\[41\]/B vssd vccd user_to_mprj_in_gates\[41\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_52_949 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_buffers\[6\] user_wb_dat_gates\[6\]/Y vssd vccd output784/A vssd vccd
+ sky130_fd_sc_hd__clkinv_8
XFILLER_31_161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_1803 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1273 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[5\]_B la_buf_enable\[5\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_2324 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1612 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xoutput654 output654/A vssd vccd la_data_in_mprj[124] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput632 output632/A vssd vccd la_data_in_mprj[104] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput643 output643/A vssd vccd la_data_in_mprj[114] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput665 output665/A vssd vccd la_data_in_mprj[19] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput676 output676/A vssd vccd la_data_in_mprj[29] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput687 output687/A vssd vccd la_data_in_mprj[39] vssd vccd sky130_fd_sc_hd__buf_2
Xuser_to_mprj_in_gates\[3\] input65/X user_to_mprj_in_gates\[3\]/B vssd vccd user_to_mprj_in_gates\[3\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_2
Xoutput698 output698/A vssd vccd la_data_in_mprj[49] vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_25_1943 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__369__A _369_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_1233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_209 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[121\]_TE mprj_logic_high_inst/HI[323] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_445 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_949 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_437 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1703 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1004 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[60\]_A input344/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_79 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_879 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1409 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1682 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[92\] _355_/Y mprj_logic_high_inst/HI[294] vssd vccd la_oenb_core[92]
+ vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input260_A la_iena_mprj[0] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input358_A la_iena_mprj[73] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_2237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[5\] input343/X mprj_logic_high_inst/HI[335] vssd vccd user_to_mprj_in_gates\[5\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_input525_A mprj_adr_o_core[17] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[115\] _378_/A la_buf_enable\[115\]/B vssd vccd la_buf\[115\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XANTENNA_user_to_mprj_oen_buffers\[20\]_TE mprj_logic_high_inst/HI[222] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_949 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_426 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_506_ _506_/A vssd vccd _506_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_user_to_mprj_in_ena_buf\[51\]_A input334/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_651 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_993 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_437_ _437_/A vssd vccd _437_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_53_1159 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_368_ _368_/A vssd vccd _368_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_31_1413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[11\] user_to_mprj_in_gates\[11\]/Y vssd vccd output649/A
+ vssd vccd sky130_fd_sc_hd__inv_6
XANTENNA_output744_A output744/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_2065 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[89\] input119/X user_to_mprj_in_gates\[89\]/B vssd vccd user_to_mprj_in_gates\[89\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_3_40 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1597 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1851 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_713 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_757 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1302 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[42\]_A input324/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_1895 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__652__A _652_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_2176 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[43\]_TE mprj_logic_high_inst/HI[245] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_529 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_35 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1740 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_209 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[51\] input334/X mprj_logic_high_inst/HI[381] vssd vccd user_to_mprj_in_gates\[51\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_25_1795 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_57 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_cyc_buf _393_/Y mprj_cyc_buf/TE vssd vccd mprj_cyc_o_user vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_ena_buf\[33\]_A input314/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input106_A la_data_out_core[77] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_245 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_buffers\[3\] user_to_mprj_in_gates\[3\]/Y vssd vccd output688/A vssd
+ vccd sky130_fd_sc_hd__clkinv_4
XFILLER_42_289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1566 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_470 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_632 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_643 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__562__A _562_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input475_A la_oenb_mprj[63] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_669 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xla_buf\[15\] _479_/Y la_buf\[15\]/TE vssd vccd la_data_in_core[15] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf\[119\]_TE la_buf\[119\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input71_A la_data_out_core[45] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1217 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[0\]_A _432_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_831 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_897 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1609 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_396 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2001 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xmprj_adr_buf\[8\] _408_/Y mprj_adr_buf\[8\]/TE vssd vccd mprj_adr_o_user[8] vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_43_1873 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_713 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_757 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[24\]_A input304/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[59\] user_to_mprj_in_gates\[59\]/Y vssd vccd output709/A
+ vssd vccd sky130_fd_sc_hd__inv_2
XANTENNA_output694_A output694/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__472__A _472_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_1811 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_wb_dat_gates\[17\] input558/X user_wb_ack_gate/B vssd vccd user_wb_dat_gates\[17\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_4
XANTENNA_la_buf_enable\[81\]_A_N _344_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_1877 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[81\]_TE la_buf\[81\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_680 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_wb_dat_buffers\[14\] user_wb_dat_gates\[14\]/Y vssd vccd output761/A vssd vccd
+ sky130_fd_sc_hd__clkinv_8
XANTENNA_la_buf_enable\[96\]_A_N _359_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[66\]_TE mprj_logic_high_inst/HI[268] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_2349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1194 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1108 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[115\] input21/X user_to_mprj_in_gates\[115\]/B vssd vccd user_to_mprj_in_gates\[115\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XANTENNA__647__A _647_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_510 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_573 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[15\]_A input294/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[34\]_A_N _626_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_1419 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1608 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[95\]_B user_to_mprj_in_gates\[95\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_40_749 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[49\]_A_N _641_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__382__A _382_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_1739 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_ena_buf\[99\] input386/X mprj_logic_high_inst/HI[429] vssd vccd user_to_mprj_in_gates\[99\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_mprj_clk2_buf_TE mprj_clk2_buf/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1537 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[125\] _388_/Y mprj_logic_high_inst/HI[327] vssd vccd la_oenb_core[125]
+ vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_mprj_dat_buf\[30\]_TE mprj_dat_buf\[30\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_1929 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_2321 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_889 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_oen_buffers\[55\] _647_/Y mprj_logic_high_inst/HI[257] vssd vccd la_oenb_core[55]
+ vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_buffers\[80\]_A user_to_mprj_in_gates\[80\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_47_337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xla_buf_enable\[77\] _340_/A la_buf_enable\[77\]/B vssd vccd la_buf\[77\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_5_1653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input223_A la_data_out_mprj[67] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_573 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__557__A _557_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_irq_ena_buf\[2\]_A input626/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1817 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input592_A mprj_dat_o_core[19] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[86\]_B user_to_mprj_in_gates\[86\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_32_1541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_433 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[89\]_TE mprj_logic_high_inst/HI[291] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_411 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_967 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[119\] _583_/Y la_buf\[119\]/TE vssd vccd la_data_in_core[119] vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_10_1883 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_694 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[112\] user_to_mprj_in_gates\[112\]/Y vssd vccd output641/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_39_827 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[10\]_B user_to_mprj_in_gates\[10\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[71\]_A user_to_mprj_in_gates\[71\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_output707_A output707/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_1681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1130 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__467__A _467_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_2017 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[77\]_B user_to_mprj_in_gates\[77\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_30_793 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1647 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_1073 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_2293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[62\]_A user_to_mprj_in_gates\[62\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_28_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__377__A _377_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_852 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[14\] input293/X mprj_logic_high_inst/HI[344] vssd vccd user_to_mprj_in_gates\[14\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_in_gates\[68\]_B user_to_mprj_in_gates\[68\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_40_557 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2002 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1861 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input173_A la_data_out_mprj[21] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[100\]_A user_to_mprj_in_gates\[100\]/Y vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_469 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input340_A la_iena_mprj[57] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_1643 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput521 mprj_adr_o_core[13] vssd vccd _413_/A vssd vccd sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_input438_A la_oenb_mprj[2] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[53\]_A user_to_mprj_in_gates\[53\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xinput510 la_oenb_mprj[95] vssd vccd _358_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_27_1687 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput532 mprj_adr_o_core[23] vssd vccd _423_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput554 mprj_dat_i_user[13] vssd vccd input554/X vssd vccd sky130_fd_sc_hd__buf_8
Xinput543 mprj_adr_o_core[4] vssd vccd _404_/A vssd vccd sky130_fd_sc_hd__buf_12
XANTENNA_input34_A la_data_out_core[127] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_635 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_657 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1821 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1461 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput587 mprj_dat_o_core[14] vssd vccd _446_/A vssd vccd sky130_fd_sc_hd__buf_4
Xla_buf\[82\] _546_/Y la_buf\[82\]/TE vssd vccd la_data_in_core[82] vssd vccd sky130_fd_sc_hd__einvp_8
Xinput598 mprj_dat_o_core[24] vssd vccd _456_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput576 mprj_dat_i_user[4] vssd vccd input576/X vssd vccd sky130_fd_sc_hd__buf_6
Xinput565 mprj_dat_i_user[23] vssd vccd input565/X vssd vccd sky130_fd_sc_hd__buf_12
XANTENNA_input605_A mprj_dat_o_core[30] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_1314 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_893 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[59\]_B user_to_mprj_in_gates\[59\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[93\]_A _557_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_1961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output657_A output657/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_775 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_981 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[71\] input100/X user_to_mprj_in_gates\[71\]/B vssd vccd user_to_mprj_in_gates\[71\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XANTENNA_user_to_mprj_in_buffers\[44\]_A user_to_mprj_in_gates\[44\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_41_1629 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_841 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_189 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_mprj_adr_buf\[21\]_TE mprj_adr_buf\[21\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_1525 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1703 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_557 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1823 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_1867 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[84\]_A _548_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_1113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1769 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1411 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_907 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_428 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_buffers\[35\]_A user_to_mprj_in_gates\[35\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_28_1985 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_1827 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_1297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_178 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_307 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1573 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_690 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
X_470_ _470_/A vssd vccd _470_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_25_373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[18\] _610_/Y mprj_logic_high_inst/HI[220] vssd vccd la_oenb_core[18]
+ vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_40_321 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[125\]_B user_to_mprj_in_gates\[125\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_40_365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[75\]_A _539_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_579 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input388_A la_oenb_mprj[0] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input290_A la_iena_mprj[127] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[93\]_B la_buf_enable\[93\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__570__A _570_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input555_A mprj_dat_i_user[14] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_1716 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1749 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2235 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_buffers\[26\]_A user_to_mprj_in_gates\[26\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_49_977 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_421 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput340 la_iena_mprj[57] vssd vccd input340/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput351 la_iena_mprj[67] vssd vccd input351/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput362 la_iena_mprj[77] vssd vccd input362/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput395 la_oenb_mprj[106] vssd vccd _369_/A vssd vccd sky130_fd_sc_hd__buf_2
Xinput373 la_iena_mprj[87] vssd vccd input373/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput384 la_iena_mprj[97] vssd vccd input384/X vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_35_137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_599_ _599_/A vssd vccd _599_/Y vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_38_2281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[41\] user_to_mprj_in_gates\[41\]/Y vssd vccd output690/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_user_to_mprj_in_gates\[116\]_B user_to_mprj_in_gates\[116\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_output774_A output774/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[66\]_A _530_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[84\]_B la_buf_enable\[84\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__480__A _480_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_1805 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1849 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[17\]_A user_to_mprj_in_gates\[17\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_6_1022 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[25\]_A input567/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_126 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_27 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_38 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_16 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_27 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[15\]_TE la_buf\[15\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XPHY_49 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__655__A _655_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_22_321 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[107\]_B user_to_mprj_in_gates\[107\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_52_1533 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1631 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[57\]_A _521_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_1090 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1675 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_527 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[75\]_B la_buf_enable\[75\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__390__A _390_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_2038 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_ena_buf\[81\] input367/X mprj_logic_high_inst/HI[411] vssd vccd user_to_mprj_in_gates\[81\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_24_2303 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2347 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1793 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1635 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2143 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2132 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_925 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_627 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input136_A la_data_out_mprj[103] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[16\]_A input557/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input303_A la_iena_mprj[23] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_522_ _522_/A vssd vccd _522_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_26_693 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_453_ _453_/A vssd vccd _453_/Y vssd vccd sky130_fd_sc_hd__inv_4
XANTENNA__565__A _565_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_343 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_685 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[45\] _509_/Y la_buf\[45\]/TE vssd vccd la_data_in_core[45] vssd vccd sky130_fd_sc_hd__einvp_8
X_384_ _384_/A vssd vccd _384_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_la_buf\[48\]_A _512_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_1021 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[117\] input279/X mprj_logic_high_inst/HI[447] vssd vccd
+ user_to_mprj_in_gates\[117\]/B vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_51_1065 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[66\]_B la_buf_enable\[66\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_70 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1607 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[101\] _565_/Y la_buf\[101\]/TE vssd vccd la_data_in_core[101] vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_49_741 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1397 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_785 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1757 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_buffers\[89\] user_to_mprj_in_gates\[89\]/Y vssd vccd output742/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
Xinput181 la_data_out_mprj[29] vssd vccd _493_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput170 la_data_out_mprj[19] vssd vccd _483_/A vssd vccd sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_la_buf\[38\]_TE la_buf\[38\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput192 la_data_out_mprj[39] vssd vccd _503_/A vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_36_468 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_405 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[34\] input59/X user_to_mprj_in_gates\[34\]/B vssd vccd user_to_mprj_in_gates\[34\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XANTENNA__475__A _475_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[39\]_A _503_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_1815 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1285 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1859 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[57\]_B la_buf_enable\[57\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_391 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2336 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xoutput633 output633/A vssd vccd la_data_in_mprj[105] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput644 output644/A vssd vccd la_data_in_mprj[115] vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA_user_to_mprj_oen_buffers\[124\]_A _387_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput655 output655/A vssd vccd la_data_in_mprj[125] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput666 output666/A vssd vccd la_data_in_mprj[1] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput677 output677/A vssd vccd la_data_in_mprj[2] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput688 output688/A vssd vccd la_data_in_mprj[3] vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_25_1911 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xoutput699 output699/A vssd vccd la_data_in_mprj[4] vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_41_1201 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1955 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1245 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_925 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1999 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__385__A _385_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_1715 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_641 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[60\]_B mprj_logic_high_inst/HI[390] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_23_685 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[6\]_TE la_buf\[6\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_807 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1330 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_335 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2097 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[48\]_B la_buf_enable\[48\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[85\] _348_/Y mprj_logic_high_inst/HI[287] vssd vccd la_oenb_core[85]
+ vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_oen_buffers\[50\]_A _642_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[115\]_A _378_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input253_A la_data_out_mprj[94] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_2111 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1504 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input420_A la_oenb_mprj[13] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input518_A mprj_adr_o_core[10] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[108\] _371_/A la_buf_enable\[108\]/B vssd vccd la_buf\[108\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_2_1261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1283 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_479 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_505_ _505_/A vssd vccd _505_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_33_449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[51\]_B mprj_logic_high_inst/HI[381] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_33_438 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_436_ _436_/A vssd vccd _436_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_la_buf_enable\[122\]_A_N _385_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_367_ _367_/A vssd vccd _367_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_la_buf_enable\[39\]_B la_buf_enable\[39\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1469 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[8\]_A input376/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[106\]_A _369_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[41\]_A _633_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1933 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output737_A output737/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_766 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_725 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_405 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_769 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[42\]_B mprj_logic_high_inst/HI[372] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_32_471 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_1093 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[32\]_A _624_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_1752 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_69 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_47 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_ena_buf\[44\] input326/X mprj_logic_high_inst/HI[374] vssd vccd user_to_mprj_in_gates\[44\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_oen_buffers\[99\]_A _362_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_1581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_769 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_909 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[33\]_B mprj_logic_high_inst/HI[363] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_23_482 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[22\] _614_/A la_buf_enable\[22\]/B vssd vccd la_buf\[22\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_11_655 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_699 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input468_A la_oenb_mprj[57] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input370_A la_iena_mprj[84] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[23\]_A _615_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input64_A la_data_out_core[39] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_821 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_1229 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1491 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_854 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1885 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1367 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_725 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_769 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[24\]_B mprj_logic_high_inst/HI[354] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_30_920 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1509 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_471 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output687_A output687/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_419_ _419_/A vssd vccd _419_/Y vssd vccd sky130_fd_sc_hd__inv_16
XFILLER_30_964 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1943 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[111\]_TE mprj_logic_high_inst/HI[313] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[14\]_A _606_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_692 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1212 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[108\] input13/X user_to_mprj_in_gates\[108\]/B vssd vccd user_to_mprj_in_gates\[108\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_37_585 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[10\]_A _410_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_235 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_533 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[15\]_B mprj_logic_high_inst/HI[345] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_20_1682 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_522 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_27 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[8\]_A input580/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[10\]_TE mprj_logic_high_inst/HI[212] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1549 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1847 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[118\] _381_/Y mprj_logic_high_inst/HI[320] vssd vccd la_oenb_core[118]
+ vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_48_817 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[8\]_A input120/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1665 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[48\] _640_/Y mprj_logic_high_inst/HI[250] vssd vccd la_oenb_core[48]
+ vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_28_585 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input216_A la_data_out_mprj[60] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_irq_ena_buf\[2\]_B user_irq_ena_buf\[2\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__573__A _573_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input585_A mprj_dat_o_core[12] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_445 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1575 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_979 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_489 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1895 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_1429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[105\] user_to_mprj_in_gates\[105\]/Y vssd vccd output633/A
+ vssd vccd sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_buffers\[71\] user_to_mprj_in_gates\[71\]/Y vssd vccd output723/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_43_1693 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_1142 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1991 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2143 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2029 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__483__A _483_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_2321 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[33\]_TE mprj_logic_high_inst/HI[235] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_761 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1030 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1697 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1085 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[4\] _436_/Y mprj_dat_buf\[4\]/TE vssd vccd mprj_dat_o_user[4] vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_29_305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1170 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1722 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[109\]_TE la_buf\[109\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1217 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_897 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__393__A _393_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_525 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1873 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[8\]_TE mprj_adr_buf\[8\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_1103 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1313 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1357 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input166_A la_data_out_mprj[15] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_1705 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xinput500 la_oenb_mprj[86] vssd vccd _349_/A vssd vccd sky130_fd_sc_hd__buf_4
Xinput511 la_oenb_mprj[96] vssd vccd _359_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_27_1655 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_1699 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1749 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput533 mprj_adr_o_core[24] vssd vccd _424_/A vssd vccd sky130_fd_sc_hd__buf_4
Xinput522 mprj_adr_o_core[14] vssd vccd _414_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput555 mprj_dat_i_user[14] vssd vccd input555/X vssd vccd sky130_fd_sc_hd__buf_12
XANTENNA_input333_A la_iena_mprj[50] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__568__A _568_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput544 mprj_adr_o_core[5] vssd vccd _405_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_25_2091 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1833 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput588 mprj_dat_o_core[15] vssd vccd _447_/A vssd vccd sky130_fd_sc_hd__buf_4
Xinput577 mprj_dat_i_user[5] vssd vccd input577/X vssd vccd sky130_fd_sc_hd__buf_8
Xinput566 mprj_dat_i_user[24] vssd vccd input566/X vssd vccd sky130_fd_sc_hd__buf_12
XANTENNA_la_buf_enable\[80\]_A_N _343_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input27_A la_data_out_core[120] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_2185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_669 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1484 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_1877 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput599 mprj_dat_o_core[25] vssd vccd _457_/A vssd vccd sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_input500_A la_oenb_mprj[86] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[71\]_TE la_buf\[71\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf\[75\] _539_/Y la_buf\[75\]/TE vssd vccd la_data_in_core[75] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_mprj_dat_buf\[23\]_A _455_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[56\]_TE mprj_logic_high_inst/HI[258] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[95\]_A_N _358_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_buffers\[30\]_A user_wb_dat_gates\[30\]/Y vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XFILLER_16_588 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_385 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1973 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[33\]_A_N _625_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_1692 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_993 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_669 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[64\] input92/X user_to_mprj_in_gates\[64\]/B vssd vccd user_to_mprj_in_gates\[64\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XANTENNA__478__A _478_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[48\]_A_N _640_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_dat_buf\[14\]_A _446_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_897 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_buffers\[21\]_A user_wb_dat_gates\[21\]/Y vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XFILLER_22_525 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_mprj_dat_buf\[20\]_TE mprj_dat_buf\[20\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_2140 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1423 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2091 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[94\]_TE la_buf\[94\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_102 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_124 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__388__A _388_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_319 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[79\]_TE mprj_logic_high_inst/HI[281] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_1624 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[9\]_A _601_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_buffers\[12\]_A user_wb_dat_gates\[12\]/Y vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XFILLER_25_385 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_377 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1247 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input283_A la_iena_mprj[120] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input450_A la_oenb_mprj[40] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_245 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input548_A mprj_adr_o_core[9] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1728 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_2197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput330 la_iena_mprj[48] vssd vccd input330/X vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_48_433 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput341 la_iena_mprj[58] vssd vccd input341/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput352 la_iena_mprj[68] vssd vccd input352/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput363 la_iena_mprj[78] vssd vccd input363/X vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_49_989 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput396 la_oenb_mprj[107] vssd vccd _370_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput374 la_iena_mprj[88] vssd vccd input374/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput385 la_iena_mprj[98] vssd vccd input385/X vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_1_1112 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_105 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_609 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_598_ _598_/A vssd vccd _598_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_43_193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_322 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[34\] user_to_mprj_in_gates\[34\]/Y vssd vccd output682/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_output767_A output767/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_551 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_41 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_74 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_63 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_1817 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_96 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_2253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_2297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[25\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_606 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XPHY_28 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_17 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_2057 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1977 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_39 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_39 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_377 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_27 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1687 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_539 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1654 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_248 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_ena_buf\[74\] input359/X mprj_logic_high_inst/HI[404] vssd vccd user_to_mprj_in_gates\[74\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_28_1761 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_1603 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_1647 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[100\] _363_/Y mprj_logic_high_inst/HI[302] vssd vccd la_oenb_core[100]
+ vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_user_wb_dat_gates\[16\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_1084 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_1983 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_959 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_937 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[30\] _622_/Y mprj_logic_high_inst/HI[232] vssd vccd la_oenb_core[30]
+ vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input129_A la_data_out_core[98] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_18_639 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xla_buf_enable\[52\] _644_/A la_buf_enable\[52\]/B vssd vccd la_buf\[52\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
X_521_ _521_/A vssd vccd _521_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_2_1465 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2188 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_609 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_452_ _452_/A vssd vccd _452_/Y vssd vccd sky130_fd_sc_hd__inv_4
XFILLER_25_193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[1\]_A _465_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_383_ _383_/A vssd vccd _383_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_40_141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input498_A la_oenb_mprj[84] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_355 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1033 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_697 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[38\] _502_/Y la_buf\[38\]/TE vssd vccd la_data_in_core[38] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA__581__A _581_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input94_A la_data_out_core[66] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_1077 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1525 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[11\]_TE mprj_adr_buf\[11\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_1619 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_753 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput160 la_data_out_mprj[125] vssd vccd _589_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput171 la_data_out_mprj[1] vssd vccd _465_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
XANTENNA_user_irq_gates\[1\]_A input622/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_797 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput193 la_data_out_mprj[3] vssd vccd _467_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput182 la_data_out_mprj[2] vssd vccd _466_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_51_417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[27\] input51/X user_to_mprj_in_gates\[27\]/B vssd vccd user_to_mprj_in_gates\[27\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_32_697 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__491__A _491_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_196 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1827 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1898 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2348 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xoutput634 output634/A vssd vccd la_data_in_mprj[106] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput645 output645/A vssd vccd la_data_in_mprj[116] vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_47_1625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xoutput656 output656/A vssd vccd la_data_in_mprj[126] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput667 output667/A vssd vccd la_data_in_mprj[20] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput678 output678/A vssd vccd la_data_in_mprj[30] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput689 output689/A vssd vccd la_data_in_mprj[40] vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_41_1213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1923 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1967 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1257 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_285 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_263 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_937 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_981 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[8\]_A _408_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1342 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_697 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_303 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_347 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[78\] _341_/Y mprj_logic_high_inst/HI[280] vssd vccd la_oenb_core[78]
+ vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_46_1157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2123 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_568 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[26\] _458_/Y mprj_dat_buf\[26\]/TE vssd vccd mprj_dat_o_user[26] vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_8_1630 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2167 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input246_A la_data_out_mprj[88] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1516 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_403 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input413_A la_oenb_mprj[122] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__576__A _576_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_18_447 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
X_504_ _504_/A vssd vccd _504_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_37_1849 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_675 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_973 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_435_ _435_/A vssd vccd _435_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_41_461 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_366_ _366_/A vssd vccd _366_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_35_1573 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_830 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[21\] _421_/Y mprj_adr_buf\[21\]/TE vssd vccd mprj_adr_o_user[21] vssd
+ vccd sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_ena_buf\[8\]_B mprj_logic_high_inst/HI[338] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1901 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1945 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output632_A output632/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1989 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1427 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[40\]_A input66/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1004 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1173 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__486__A _486_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_778 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_29 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_645 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1635 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[6\] _598_/A la_buf_enable\[6\]/B vssd vccd la_buf\[6\]/TE vssd vccd
+ sky130_fd_sc_hd__and2b_1
XFILLER_31_1993 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_2009 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[31\]_A input56/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input1_A caravel_clk vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_1764 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_1775 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1065 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_767 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__396__A _396_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[37\] input318/X mprj_logic_high_inst/HI[367] vssd vccd user_to_mprj_in_gates\[37\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_3_1593 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[98\]_A input129/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_1579 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_667 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1713 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[15\] _607_/A la_buf_enable\[15\]/B vssd vccd la_buf\[15\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_7_605 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_494 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_678 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_1161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input196_A la_data_out_mprj[42] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[28\]_TE la_buf\[28\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input363_A la_iena_mprj[78] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_2207 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_866 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[22\]_A input46/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input57_A la_data_out_core[32] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input530_A mprj_adr_o_core[21] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[120\] _383_/A la_buf_enable\[120\]/B vssd vccd la_buf\[120\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_19_701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1897 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[89\]_A input119/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_748 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_483 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_418_ _418_/A vssd vccd _418_/Y vssd vccd sky130_fd_sc_hd__inv_12
XFILLER_15_1911 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_976 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1201 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1955 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_349_ _349_/A vssd vccd _349_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_31_1245 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1819 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1999 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_1690 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_1289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[94\] input125/X user_to_mprj_in_gates\[94\]/B vssd vccd user_to_mprj_in_gates\[94\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XANTENNA_user_to_mprj_in_gates\[13\]_A input36/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_1224 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_509 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1341 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1385 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_545 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_597 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1145 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_589 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_39 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_wb_dat_gates\[8\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_1263 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1859 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[8\]_B user_to_mprj_in_gates\[8\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[121\]_A_N _384_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_2345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_829 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1677 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input209_A la_data_out_mprj[54] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input111_A la_data_out_core[81] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_1933 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_431 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1521 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input480_A la_oenb_mprj[68] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input578_A mprj_dat_i_user[6] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf\[20\] _484_/Y la_buf\[20\]/TE vssd vccd la_data_in_core[20] vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_32_1565 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_1005 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1049 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_641 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_542 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_862 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[64\] user_to_mprj_in_gates\[64\]/Y vssd vccd output715/A
+ vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_37_2155 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_567 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_217 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_589 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_291 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_gates\[22\] input564/X user_wb_ack_gate/B vssd vccd user_wb_dat_gates\[22\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_2
XFILLER_50_1621 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_773 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1665 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1042 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1097 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1425 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_1087 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[120\] input27/X user_to_mprj_in_gates\[120\]/B vssd vccd user_to_mprj_in_gates\[120\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_22_1734 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_873 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_501 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1182 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_2253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1229 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2108 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[110\]_A input272/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_397 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_272 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1841 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1115 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1885 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1601 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_1369 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2335 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[60\] _652_/Y mprj_logic_high_inst/HI[262] vssd vccd la_oenb_core[60]
+ vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[82\] _345_/A la_buf_enable\[82\]/B vssd vccd la_buf\[82\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XANTENNA_input159_A la_data_out_mprj[124] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput501 la_oenb_mprj[87] vssd vccd _350_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput512 la_oenb_mprj[97] vssd vccd _360_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput545 mprj_adr_o_core[6] vssd vccd _406_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput523 mprj_adr_o_core[15] vssd vccd _415_/A vssd vccd sky130_fd_sc_hd__buf_2
Xinput534 mprj_adr_o_core[25] vssd vccd _425_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_47_125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1981 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xinput578 mprj_dat_i_user[6] vssd vccd input578/X vssd vccd sky130_fd_sc_hd__buf_8
Xinput556 mprj_dat_i_user[15] vssd vccd input556/X vssd vccd sky130_fd_sc_hd__buf_12
Xinput567 mprj_dat_i_user[25] vssd vccd input567/X vssd vccd sky130_fd_sc_hd__buf_12
XANTENNA_input326_A la_iena_mprj[44] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1845 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput589 mprj_dat_o_core[16] vssd vccd _448_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_28_361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_1889 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[101\]_TE mprj_logic_high_inst/HI[303] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
Xla_buf\[68\] _532_/Y la_buf\[68\]/TE vssd vccd la_data_in_core[68] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA__584__A _584_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[101\]_A input262/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_2041 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_700 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1941 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1985 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[124\] _588_/Y la_buf\[124\]/TE vssd vccd la_data_in_core[124] vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_43_2181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_1205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output712_A output712/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[57\] input84/X user_to_mprj_in_gates\[57\]/B vssd vccd user_to_mprj_in_gates\[57\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_19_361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[119\]_A input25/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__494__A _494_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_813 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1251 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2152 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_29 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_419 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_1509 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_27 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1807 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[124\]_TE mprj_logic_high_inst/HI[326] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_136 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_1553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_629 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[90\]_A input377/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_1037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_1259 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_389 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1693 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input276_A la_iena_mprj[114] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input443_A la_oenb_mprj[34] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__579__A _579_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2310 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1525 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput320 la_iena_mprj[39] vssd vccd input320/X vssd vccd sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_42_1929 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_445 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input610_A mprj_dat_o_core[6] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[23\]_TE mprj_logic_high_inst/HI[225] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
Xinput331 la_iena_mprj[49] vssd vccd input331/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput342 la_iena_mprj[59] vssd vccd input342/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput353 la_iena_mprj[69] vssd vccd input353/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput397 la_oenb_mprj[108] vssd vccd _371_/A vssd vccd sky130_fd_sc_hd__buf_4
Xinput364 la_iena_mprj[79] vssd vccd input364/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput375 la_iena_mprj[89] vssd vccd input375/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput386 la_iena_mprj[99] vssd vccd input386/X vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_48_489 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[81\]_A input367/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_81 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_813 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_597_ _597_/A vssd vccd _597_/Y vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_38_2261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_buffers\[27\] user_to_mprj_in_gates\[27\]/Y vssd vccd output674/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_output662_A output662/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_1181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_1793 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1788 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1829 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1217 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__489__A _489_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_2129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_629 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_29 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_18 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[72\]_A input357/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_1989 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_2069 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1357 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_39 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[8\]_B la_buf_enable\[8\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_17_1699 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1877 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[61\]_TE la_buf\[61\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1866 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1287 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[94\]_A_N _357_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__399__A _399_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[46\]_TE mprj_logic_high_inst/HI[248] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_1709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[67\] input351/X mprj_logic_high_inst/HI[397] vssd vccd user_to_mprj_in_gates\[67\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_24_1659 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_2281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_607 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1580 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_520_ _520_/A vssd vccd _520_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_41_1995 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[63\]_A input347/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_150 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[5\] _597_/Y mprj_logic_high_inst/HI[207] vssd vccd la_oenb_core[5]
+ vssd vccd sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[23\] _615_/Y mprj_logic_high_inst/HI[225] vssd vccd la_oenb_core[23]
+ vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[45\] _637_/A la_buf_enable\[45\]/B vssd vccd la_buf\[45\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
X_451_ _451_/A vssd vccd _451_/Y vssd vccd sky130_fd_sc_hd__inv_4
XFILLER_13_301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_621 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_382_ _382_/A vssd vccd _382_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_la_buf_enable\[32\]_A_N _624_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1001 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input393_A la_oenb_mprj[104] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_1045 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[47\]_A_N _639_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input87_A la_data_out_core[5] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_1089 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input560_A mprj_dat_i_user[19] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_1537 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2001 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2045 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_mprj_dat_buf\[10\]_TE mprj_dat_buf\[10\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_721 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_916 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_765 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput161 la_data_out_mprj[126] vssd vccd _590_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput150 la_data_out_mprj[116] vssd vccd _580_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput172 la_data_out_mprj[20] vssd vccd _484_/A vssd vccd sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_user_irq_gates\[1\]_B user_irq_gates\[1\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput194 la_data_out_mprj[40] vssd vccd _504_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput183 la_data_out_mprj[30] vssd vccd _494_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
XANTENNA_user_to_mprj_in_ena_buf\[54\]_A input337/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
X_649_ _649_/A vssd vccd _649_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_38_2080 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_632 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1811 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_1975 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1839 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[84\]_TE la_buf\[84\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_371 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[69\]_TE mprj_logic_high_inst/HI[271] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
Xoutput635 output635/A vssd vccd la_data_in_mprj[107] vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_47_1637 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xoutput657 output657/A vssd vccd la_data_in_mprj[127] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput668 output668/A vssd vccd la_data_in_mprj[21] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput679 output679/A vssd vccd la_data_in_mprj[31] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput646 output646/A vssd vccd la_data_in_mprj[117] vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_45_2073 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1935 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_275 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_949 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_1269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_sel_buf\[2\]_A _398_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[45\]_A input327/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_437 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_481 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_993 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_805 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_665 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2077 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_315 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1354 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_359 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1630 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2135 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_1169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1675 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2179 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[19\] _451_/Y mprj_dat_buf\[19\]/TE vssd vccd mprj_dat_o_user[19] vssd
+ vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input239_A la_data_out_mprj[81] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input141_A la_data_out_mprj[108] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_713 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_415 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1528 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1230 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_757 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_908 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input406_A la_oenb_mprj[116] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[36\]_A input317/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_503_ _503_/A vssd vccd _503_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_2_1296 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_434_ _434_/A vssd vccd _434_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_26_470 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_2253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[50\] _514_/Y la_buf\[50\]/TE vssd vccd la_data_in_core[50] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA__592__A _592_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_473 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2106 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_687 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[122\] input285/X mprj_logic_high_inst/HI[452] vssd vccd
+ user_to_mprj_in_gates\[122\]/B vssd vccd sky130_fd_sc_hd__and2_1
X_365_ _365_/A vssd vccd _365_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_35_1585 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_mprj_dat_buf\[3\]_A _435_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_842 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_886 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_1913 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1957 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[14\] _414_/Y mprj_adr_buf\[14\]/TE vssd vccd mprj_adr_o_user[14] vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_29_1345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1439 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[40\]_B user_to_mprj_in_gates\[40\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[94\] user_to_mprj_in_gates\[94\]/Y vssd vccd output748/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_49_573 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[27\]_A input307/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_749 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_wb_dat_buffers\[4\] user_wb_dat_gates\[4\]/Y vssd vccd output782/A vssd vccd
+ sky130_fd_sc_hd__clkinv_8
XFILLER_20_657 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1603 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1794 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1073 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1647 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[1\] input43/X user_to_mprj_in_gates\[1\]/B vssd vccd user_to_mprj_in_gates\[1\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XANTENNA_user_to_mprj_in_buffers\[92\]_A user_to_mprj_in_gates\[92\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[31\]_B user_to_mprj_in_gates\[31\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_28_713 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1607 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1787 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_1077 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[18\]_A input297/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_779 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[98\]_B user_to_mprj_in_gates\[98\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_52_1173 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input189_A la_data_out_mprj[36] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[90\] _353_/Y mprj_logic_high_inst/HI[292] vssd vccd la_oenb_core[90]
+ vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_3_878 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input356_A la_iena_mprj[71] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[83\]_A user_to_mprj_in_gates\[83\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[22\]_B user_to_mprj_in_gates\[22\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_43_1832 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[3\] input321/X mprj_logic_high_inst/HI[333] vssd vccd user_to_mprj_in_gates\[3\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
Xla_buf\[98\] _562_/Y la_buf\[98\]/TE vssd vccd la_data_in_core[98] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_input523_A mprj_adr_o_core[15] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_713 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[113\] _376_/A la_buf_enable\[113\]/B vssd vccd la_buf\[113\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XANTENNA__587__A _587_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_2326 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[89\]_B user_to_mprj_in_gates\[89\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_37_1625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1603 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1093 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_417_ _417_/A vssd vccd _417_/Y vssd vccd sky130_fd_sc_hd__inv_6
XFILLER_15_1923 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_348_ _348_/A vssd vccd _348_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_14_495 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1847 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1967 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1257 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[121\]_A user_to_mprj_in_gates\[121\]/Y vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output742_A output742/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1721 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[110\]_A _574_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1765 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[74\]_A user_to_mprj_in_gates\[74\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[13\]_B user_to_mprj_in_gates\[13\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_44_1629 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[87\] input117/X user_to_mprj_in_gates\[87\]/B vssd vccd user_to_mprj_in_gates\[87\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_42_1353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__497__A _497_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_705 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_mprj_adr_buf\[24\]_TE mprj_adr_buf\[24\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_1870 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_557 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_2161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_421 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1591 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_498 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[112\]_A user_to_mprj_in_gates\[112\]/Y vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[101\]_A _565_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[65\]_A user_to_mprj_in_gates\[65\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_47_1275 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1117 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_2252 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_329 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_543 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_727 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1901 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input104_A la_data_out_core[75] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_1967 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[1\] user_to_mprj_in_gates\[1\]/Y vssd vccd output666/A vssd
+ vccd sky130_fd_sc_hd__clkinv_4
XFILLER_23_281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_410 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_51 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_443 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_62 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input473_A la_oenb_mprj[61] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[103\]_A user_to_mprj_in_gates\[103\]/Y vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_1533 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xla_buf\[13\] _477_/Y la_buf\[13\]/TE vssd vccd la_data_in_core[13] vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf\[9\] _473_/Y la_buf\[9\]/TE vssd vccd la_data_in_core[9] vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_48_1017 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[56\]_A user_to_mprj_in_gates\[56\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1905 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2027 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_163 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[6\] _406_/Y mprj_adr_buf\[6\]/TE vssd vccd mprj_adr_o_user[6] vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_8_1280 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_841 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_830 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_554 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2112 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[57\] user_to_mprj_in_gates\[57\]/Y vssd vccd output707/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_37_2167 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output692_A output692/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[96\]_A _560_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_579 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2009 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1731 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1633 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1775 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_gates\[15\] input556/X user_wb_ack_gate/B vssd vccd user_wb_dat_gates\[15\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_4
XFILLER_30_785 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1021 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1677 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_1054 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_981 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_buffers\[47\]_A user_to_mprj_in_gates\[47\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_44_2127 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_wb_dat_buffers\[12\] user_wb_dat_gates\[12\]/Y vssd vccd output759/A vssd vccd
+ sky130_fd_sc_hd__clkinv_8
XANTENNA_la_buf\[20\]_A _484_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_1871 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_29 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1099 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[113\] input19/X user_to_mprj_in_gates\[113\]/B vssd vccd user_to_mprj_in_gates\[113\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XANTENNA_la_buf\[18\]_TE la_buf\[18\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_1194 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_332 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[110\]_B mprj_logic_high_inst/HI[440] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[87\]_A _551_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[97\] input384/X mprj_logic_high_inst/HI[427] vssd vccd user_to_mprj_in_gates\[97\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_49_1337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_buffers\[38\]_A user_to_mprj_in_gates\[38\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_27_2347 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[123\] _386_/Y mprj_logic_high_inst/HI[325] vssd vccd la_oenb_core[123]
+ vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf\[11\]_A _475_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput502 la_oenb_mprj[88] vssd vccd _351_/A vssd vccd sky130_fd_sc_hd__buf_4
Xuser_to_mprj_oen_buffers\[53\] _645_/Y mprj_logic_high_inst/HI[255] vssd vccd la_oenb_core[53]
+ vssd vccd sky130_fd_sc_hd__einvp_8
Xinput546 mprj_adr_o_core[7] vssd vccd _407_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput524 mprj_adr_o_core[16] vssd vccd _416_/A vssd vccd sky130_fd_sc_hd__buf_2
Xinput513 la_oenb_mprj[98] vssd vccd _361_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput535 mprj_adr_o_core[26] vssd vccd _426_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_47_137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[75\] _338_/A la_buf_enable\[75\]/B vssd vccd la_buf\[75\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
Xinput568 mprj_dat_i_user[26] vssd vccd input568/X vssd vccd sky130_fd_sc_hd__buf_8
Xinput579 mprj_dat_i_user[7] vssd vccd input579/X vssd vccd sky130_fd_sc_hd__buf_8
Xinput557 mprj_dat_i_user[16] vssd vccd input557/X vssd vccd sky130_fd_sc_hd__clkbuf_16
XFILLER_5_1453 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_1857 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input319_A la_iena_mprj[38] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input221_A la_data_out_mprj[65] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_844 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[101\]_B mprj_logic_high_inst/HI[431] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[78\]_A _542_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input590_A mprj_dat_o_core[17] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_712 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[96\]_B la_buf_enable\[96\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_1953 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_1915 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1997 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1385 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_962 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[117\] _581_/Y la_buf\[117\]/TE vssd vccd la_data_in_core[117] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_buffers\[29\]_A user_to_mprj_in_gates\[29\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1871 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_461 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[110\] user_to_mprj_in_gates\[110\]/Y vssd vccd output639/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_6_1217 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[20\]_B la_buf_enable\[20\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output705_A output705/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_1481 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_321 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[119\]_B user_to_mprj_in_gates\[119\]/B vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[69\]_A _533_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_869 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[87\]_B la_buf_enable\[87\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[120\]_A_N _383_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_1138 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_1441 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_593 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1933 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_39 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[11\]_B la_buf_enable\[11\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[28\]_A input570/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_1819 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_148 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1565 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1005 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[90\]_B mprj_logic_high_inst/HI[420] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[9\]_TE la_buf\[9\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_1049 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[12\] input291/X mprj_logic_high_inst/HI[342] vssd vccd user_to_mprj_in_gates\[12\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_41_869 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2340 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[78\]_B la_buf_enable\[78\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_1661 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[80\]_A _343_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_41 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input171_A la_data_out_mprj[1] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_2133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_1145 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_85 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input269_A la_iena_mprj[108] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1009 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1537 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_925 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput321 la_iena_mprj[3] vssd vccd input321/X vssd vccd sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_input436_A la_oenb_mprj[28] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[19\]_A input560/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput310 la_iena_mprj[2] vssd vccd input310/X vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_7_1504 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xinput354 la_iena_mprj[6] vssd vccd input354/X vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput332 la_iena_mprj[4] vssd vccd input332/X vssd vccd sky130_fd_sc_hd__buf_2
Xinput343 la_iena_mprj[5] vssd vccd input343/X vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA_input32_A la_data_out_core[125] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1621 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[80\] _544_/Y la_buf\[80\]/TE vssd vccd la_data_in_core[80] vssd vccd sky130_fd_sc_hd__einvp_8
Xinput387 la_iena_mprj[9] vssd vccd input387/X vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA_input603_A mprj_dat_o_core[29] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput365 la_iena_mprj[7] vssd vccd input365/X vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput376 la_iena_mprj[8] vssd vccd input376/X vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_40_1665 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA__595__A _595_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput398 la_oenb_mprj[109] vssd vccd _372_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_1_1136 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1147 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[81\]_B mprj_logic_high_inst/HI[411] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_32_825 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_596_ _596_/A vssd vccd _596_/Y vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_32_803 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1425 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_869 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[69\]_B la_buf_enable\[69\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_571 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1761 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_575 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output655_A output655/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[71\]_A _334_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_1229 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_1491 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_1429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1852 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_641 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XPHY_19 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[72\]_B mprj_logic_high_inst/HI[402] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_39_1369 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_685 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_357 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1970 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[127\]_A _390_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[62\]_A _654_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1889 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1299 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1329 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1592 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_405 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[63\]_B mprj_logic_high_inst/HI[393] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
X_450_ _450_/A vssd vccd _450_/Y vssd vccd sky130_fd_sc_hd__inv_4
Xuser_to_mprj_oen_buffers\[16\] _608_/Y mprj_logic_high_inst/HI[218] vssd vccd la_oenb_core[16]
+ vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[38\] _630_/A la_buf_enable\[38\]/B vssd vccd la_buf\[38\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
X_381_ _381_/A vssd vccd _381_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_25_162 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1057 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input386_A la_iena_mprj[99] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[118\]_A _381_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[53\]_A _645_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input553_A mprj_dat_i_user[12] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_2013 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_1549 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_740 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_777 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xinput162 la_data_out_mprj[127] vssd vccd _591_/A vssd vccd sky130_fd_sc_hd__buf_2
Xinput140 la_data_out_mprj[107] vssd vccd _571_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput151 la_data_out_mprj[117] vssd vccd _581_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_48_265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_405 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput195 la_data_out_mprj[41] vssd vccd _505_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput184 la_data_out_mprj[31] vssd vccd _495_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput173 la_data_out_mprj[21] vssd vccd _485_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_7_1389 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_909 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[54\]_B mprj_logic_high_inst/HI[384] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
X_648_ _648_/A vssd vccd _648_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_36_1509 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_579_ _579_/A vssd vccd _579_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_38_2092 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output772_A output772/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[114\]_TE mprj_logic_high_inst/HI[316] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_18_1987 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[44\]_A _636_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[109\]_A _372_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_1553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_383 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xoutput636 output636/A vssd vccd la_data_in_mprj[108] vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_47_1649 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2041 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xoutput658 output658/A vssd vccd la_data_in_mprj[12] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput669 output669/A vssd vccd la_data_in_mprj[22] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput647 output647/A vssd vccd la_data_in_mprj[118] vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_28_1037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2085 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_405 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_29 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[45\]_B mprj_logic_high_inst/HI[375] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_36_961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_600 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_953 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2045 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_839 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1366 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_327 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[35\]_A _627_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[13\]_TE mprj_logic_high_inst/HI[215] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1642 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_537 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1593 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_725 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input134_A la_data_out_mprj[101] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[31\]_A _431_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_1220 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1793 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_769 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_427 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[36\]_B mprj_logic_high_inst/HI[366] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_input301_A la_iena_mprj[21] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_502_ _502_/A vssd vccd _502_/Y vssd vccd sky130_fd_sc_hd__inv_2
X_433_ _433_/A vssd vccd _433_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_35_2221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_441 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2276 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_699 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[43\] _507_/Y la_buf\[43\]/TE vssd vccd la_data_in_core[43] vssd vccd sky130_fd_sc_hd__einvp_8
X_364_ _364_/A vssd vccd _364_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_31_2118 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_2265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_ena_buf\[115\] input277/X mprj_logic_high_inst/HI[445] vssd vccd
+ user_to_mprj_in_gates\[115\]/B vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_oen_buffers\[26\]_A _618_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_854 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1313 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1925 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_11 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_1969 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1357 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1407 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_585 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1568 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_buffers\[87\] user_to_mprj_in_gates\[87\]/Y vssd vccd output740/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_mprj_adr_buf\[22\]_A _422_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[27\]_B mprj_logic_high_inst/HI[357] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[51\]_TE la_buf\[51\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[32\] input57/X user_to_mprj_in_gates\[32\]/B vssd vccd user_to_mprj_in_gates\[32\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_51_249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_953 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[36\]_TE mprj_logic_high_inst/HI[238] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[93\]_A_N _356_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_1615 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_669 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[17\]_A _609_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_1659 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1085 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1973 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[31\]_A_N _623_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_1805 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1001 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1619 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1849 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[13\]_A _413_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_2241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_2263 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[46\]_A_N _638_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_1089 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1551 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[18\]_B mprj_logic_high_inst/HI[348] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_15_419 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_629 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_117 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[83\] _346_/Y mprj_logic_high_inst/HI[285] vssd vccd la_oenb_core[83]
+ vssd vccd sky130_fd_sc_hd__einvp_8
XFILLER_5_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[31\] _463_/Y mprj_dat_buf\[31\]/TE vssd vccd mprj_dat_o_user[31] vssd
+ vccd sky130_fd_sc_hd__einvp_8
XFILLER_2_334 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input349_A la_iena_mprj[65] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input251_A la_data_out_mprj[92] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_1844 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2027 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[74\]_TE la_buf\[74\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input516_A mprj_ack_i_user vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_725 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_533 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[106\] _369_/A la_buf_enable\[106\]/B vssd vccd la_buf\[106\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XANTENNA_user_to_mprj_oen_buffers\[59\]_TE mprj_logic_high_inst/HI[261] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_2338 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_279 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1615 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1637 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_416_ _416_/A vssd vccd _416_/Y vssd vccd sky130_fd_sc_hd__inv_12
XFILLER_35_2073 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_347_ _347_/A vssd vccd _347_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_15_1935 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1859 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_1979 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1733 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_output735_A output735/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1777 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1259 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[23\]_TE mprj_dat_buf\[23\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_1125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_433 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[2\]_TE mprj_logic_high_inst/HI[204] vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
XFILLER_49_2209 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1817 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[97\]_TE la_buf\[97\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_2264 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_555 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_ena_buf\[42\] input324/X mprj_logic_high_inst/HI[372] vssd vccd user_to_mprj_in_gates\[42\]/B
+ vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_31_709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1924 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_2213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[20\] _612_/A la_buf_enable\[20\]/B vssd vccd la_buf\[20\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_23_293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input299_A la_iena_mprj[1] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_74 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1990 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input466_A la_oenb_mprj[55] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input62_A la_data_out_core[37] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1029 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_120 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_1917 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2039 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_665 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__598__A _598_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_2353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_533 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_mprj_dat_buf\[26\]_A _458_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_897 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_599 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2124 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2179 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output685_A output685/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_1489 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1743 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1607 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1645 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1787 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1563 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2139 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1933 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1850 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_1883 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1703 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_2222 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_1747 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[17\]_A _449_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_823 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_886 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[106\] input11/X user_to_mprj_in_gates\[106\]/B vssd vccd user_to_mprj_in_gates\[106\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XANTENNA_user_wb_dat_buffers\[24\]_A user_wb_dat_gates\[24\]/Y vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XFILLER_37_385 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_344 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_29 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_720 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1409 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2017 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_908 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2359 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput503 la_oenb_mprj[89] vssd vccd _352_/A vssd vccd sky130_fd_sc_hd__buf_4
Xuser_to_mprj_oen_buffers\[116\] _379_/Y mprj_logic_high_inst/HI[318] vssd vccd la_oenb_core[116]
+ vssd vccd sky130_fd_sc_hd__einvp_8
Xinput525 mprj_adr_o_core[17] vssd vccd _417_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput536 mprj_adr_o_core[27] vssd vccd _427_/A vssd vccd sky130_fd_sc_hd__buf_2
Xinput514 la_oenb_mprj[99] vssd vccd _362_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_9_1590 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1421 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_105 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xinput569 mprj_dat_i_user[27] vssd vccd input569/X vssd vccd sky130_fd_sc_hd__buf_8
Xinput558 mprj_dat_i_user[17] vssd vccd input558/X vssd vccd sky130_fd_sc_hd__buf_12
Xinput547 mprj_adr_o_core[8] vssd vccd _408_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_47_149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_341 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[46\] _638_/Y mprj_logic_high_inst/HI[248] vssd vccd la_oenb_core[46]
+ vssd vccd sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[68\] _331_/A la_buf_enable\[68\]/B vssd vccd la_buf\[68\]/TE vssd
+ vccd sky130_fd_sc_hd__and2b_1
XFILLER_29_897 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_503 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input214_A la_data_out_mprj[59] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_buffers\[15\]_A user_wb_dat_gates\[15\]/Y vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XFILLER_40_1869 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_856 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1721 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1787 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input583_A mprj_dat_o_core[10] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_1927 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_234 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1397 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1651 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[14\]_TE mprj_adr_buf\[14\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_974 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1883 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_473 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1229 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[103\] user_to_mprj_in_gates\[103\]/Y vssd vccd output631/A
+ vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_43_1493 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_650 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_801 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1885 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_1729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1453 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_790 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1901 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1989 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[2\] _434_/Y mprj_dat_buf\[2\]/TE vssd vccd mprj_dat_o_user[2] vssd
+ vccd sky130_fd_sc_hd__einvp_8
XANTENNA_user_wb_dat_gates\[28\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_2306 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_mprj_dat_buf\[2\]_TE mprj_dat_buf\[2\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_1691 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_664 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1017 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[110\]_B la_buf_enable\[110\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_1905 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[122\]_TE la_buf\[122\]/TE vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1971 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_749 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_wb_dat_buffers\[1\]_A user_wb_dat_gates\[1\]/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_53 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input164_A la_data_out_mprj[13] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_97 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2167 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_wb_dat_gates\[19\]_B user_wb_ack_gate/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput300 la_iena_mprj[20] vssd vccd input300/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput311 la_iena_mprj[30] vssd vccd input311/X vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_29_51 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_999 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_937 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input429_A la_oenb_mprj[21] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input331_A la_iena_mprj[49] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput322 la_iena_mprj[40] vssd vccd input322/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput333 la_iena_mprj[50] vssd vccd input333/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput344 la_iena_mprj[60] vssd vccd input344/X vssd vccd sky130_fd_sc_hd__clkbuf_1
XFILLER_40_1633 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_469 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xinput388 la_oenb_mprj[0] vssd vccd _592_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
XANTENNA_input25_A la_data_out_core[119] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput355 la_iena_mprj[70] vssd vccd input355/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput366 la_iena_mprj[80] vssd vccd input366/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput377 la_iena_mprj[90] vssd vccd input377/X vssd vccd sky130_fd_sc_hd__clkbuf_1
Xinput399 la_oenb_mprj[10] vssd vccd _602_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_40_1677 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[73\] _537_/Y la_buf\[73\]/TE vssd vccd la_data_in_core[73] vssd vccd sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf\[4\]_A _468_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[101\]_B la_buf_enable\[101\]/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_595_ _595_/A vssd vccd _595_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_32_837 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_881 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_583 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1773 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_587 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[70\]_A input99/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output648_A output648/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[62\] input90/X user_to_mprj_in_gates\[62\]/B vssd vccd user_to_mprj_in_gates\[62\]/Y
+ vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_48_981 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1864 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_601 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_697 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_645 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1050 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_892 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1802 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1982 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[61\]_A input89/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_2307 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1803 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1847 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_992 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[92\]_TE mprj_logic_high_inst/HI[294] vssd vccd
+ vccd vssd sky130_fd_sc_hd__diode_2
X_380_ _380_/A vssd vccd _380_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_9_307 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_input281_A la_iena_mprj[119] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input379_A la_iena_mprj[92] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[52\]_A input79/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input546_A mprj_adr_o_core[7] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1357 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput130 la_data_out_core[99] vssd vccd input130/X vssd vccd sky130_fd_sc_hd__buf_4
Xinput152 la_data_out_mprj[118] vssd vccd _582_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput163 la_data_out_mprj[12] vssd vccd _476_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput141 la_data_out_mprj[108] vssd vccd _572_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_36_417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1441 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xinput196 la_data_out_mprj[42] vssd vccd _506_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput185 la_data_out_mprj[32] vssd vccd _496_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
Xinput174 la_data_out_mprj[22] vssd vccd _486_/A vssd vccd sky130_fd_sc_hd__clkbuf_2
XFILLER_40_1485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
X_647_ _647_/A vssd vccd _647_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
X_578_ _578_/A vssd vccd _578_/Y vssd vccd sky130_fd_sc_hd__inv_4
XFILLER_32_601 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_645 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[2\]_A user_to_mprj_in_gates\[2\]/Y vssd vccd vccd
+ vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[32\] user_to_mprj_in_gates\[32\]/Y vssd vccd output680/A
+ vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_output765_A output765/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_874 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1565 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[43\]_A input69/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput659 output659/A vssd vccd la_data_in_mprj[13] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput637 output637/A vssd vccd la_data_in_mprj[109] vssd vccd sky130_fd_sc_hd__buf_2
Xoutput648 output648/A vssd vccd la_data_in_mprj[119] vssd vccd sky130_fd_sc_hd__buf_2
XFILLER_45_2053 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1049 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2097 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
.ends

.subckt sky130_fd_sc_hvl__decap_4 VGND VPWR VNB VPB
X0 VGND VPWR VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=1e+06u
X1 VPWR VGND VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
.ends

.subckt sky130_fd_sc_hvl__decap_8 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=1e+06u
X2 VPWR VGND VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3 VGND VPWR VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=1e+06u
.ends

.subckt sky130_fd_sc_hvl__diode_2 DIODE VGND VPB VPWR VNB
D0 VNB DIODE sky130_fd_pr__diode_pw2nd_11v0 pj=5.88e+06u area=6.072e+11p
.ends

.subckt xres_buf A X VPWR LVPWR LVGND VGND
XFILLER_0_24 VGND VPWR VGND VPWR sky130_fd_sc_hvl__decap_4
XFILLER_1_0 VGND VPWR VGND VPWR sky130_fd_sc_hvl__decap_8
XFILLER_0_16 VGND VPWR VGND VPWR sky130_fd_sc_hvl__decap_8
XFILLER_1_8 VGND VPWR VGND VPWR sky130_fd_sc_hvl__decap_4
XANTENNA_lvlshiftdown_A A VGND VPWR VPWR VGND sky130_fd_sc_hvl__diode_2
XFILLER_2_0 VGND VPWR VGND VPWR sky130_fd_sc_hvl__decap_8
XFILLER_0_0 VGND VPWR VGND VPWR sky130_fd_sc_hvl__decap_8
Xlvlshiftdown A VGND VPWR X VGND VPWR LVPWR sky130_fd_sc_hvl__lsbufhv2lv_1
XFILLER_0_8 VGND VPWR VGND VPWR sky130_fd_sc_hvl__decap_8
.ends

* Black-box entry subcircuit for user_project_wrapper abstract view
.subckt user_project_wrapper analog_io[0] analog_io[10] analog_io[11] analog_io[12]
+ analog_io[13] analog_io[14] analog_io[15] analog_io[16] analog_io[17] analog_io[18]
+ analog_io[19] analog_io[1] analog_io[20] analog_io[21] analog_io[22] analog_io[23]
+ analog_io[24] analog_io[25] analog_io[26] analog_io[27] analog_io[28] analog_io[2]
+ analog_io[3] analog_io[4] analog_io[5] analog_io[6] analog_io[7] analog_io[8] analog_io[9]
+ io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17]
+ io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23] io_in[24] io_in[25]
+ io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31] io_in[32] io_in[33]
+ io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14]
+ io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21]
+ io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29]
+ io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36]
+ io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9]
+ io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15] io_out[16]
+ io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22] io_out[23]
+ io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29] io_out[2] io_out[30]
+ io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36] io_out[37] io_out[3]
+ io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100]
+ la_data_in[101] la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105]
+ la_data_in[106] la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110]
+ la_data_in[111] la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115]
+ la_data_in[116] la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120]
+ la_data_in[121] la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125]
+ la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15]
+ la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20]
+ la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26]
+ la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31]
+ la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37]
+ la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42]
+ la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48]
+ la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53]
+ la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59]
+ la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64]
+ la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6]
+ la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75]
+ la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80]
+ la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86]
+ la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91]
+ la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97]
+ la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101]
+ la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106]
+ la_data_out[107] la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110]
+ la_data_out[111] la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115]
+ la_data_out[116] la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11]
+ la_data_out[120] la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124]
+ la_data_out[125] la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13]
+ la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18]
+ la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23]
+ la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28]
+ la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33]
+ la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38]
+ la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43]
+ la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48]
+ la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53]
+ la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58]
+ la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63]
+ la_data_out[64] la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68]
+ la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73]
+ la_data_out[74] la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78]
+ la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83]
+ la_data_out[84] la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88]
+ la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93]
+ la_data_out[94] la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98]
+ la_data_out[99] la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102]
+ la_oenb[103] la_oenb[104] la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109]
+ la_oenb[10] la_oenb[110] la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115]
+ la_oenb[116] la_oenb[117] la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121]
+ la_oenb[122] la_oenb[123] la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12]
+ la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19]
+ la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25]
+ la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31]
+ la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38]
+ la_oenb[39] la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44]
+ la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50]
+ la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57]
+ la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63]
+ la_oenb[64] la_oenb[65] la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6]
+ la_oenb[70] la_oenb[71] la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76]
+ la_oenb[77] la_oenb[78] la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82]
+ la_oenb[83] la_oenb[84] la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89]
+ la_oenb[8] la_oenb[90] la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95]
+ la_oenb[96] la_oenb[97] la_oenb[98] la_oenb[99] la_oenb[9] user_clock2 user_irq[0]
+ user_irq[1] user_irq[2] vccd1 vccd2 vdda1 vdda2 vssa1 vssa2 vssd1 vssd2 wb_clk_i
+ wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13]
+ wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19]
+ wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24]
+ wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2]
+ wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6]
+ wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11]
+ wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17]
+ wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22]
+ wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28]
+ wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4]
+ wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10]
+ wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16]
+ wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21]
+ wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27]
+ wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3]
+ wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0]
+ wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
.ends

.subckt sky130_fd_sc_hd__or2_4 A B VGND VPWR X VNB VPB
X0 a_121_297# B a_35_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR a_35_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 X a_35_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_35_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 X a_35_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR a_35_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 X a_35_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR A a_121_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND A a_35_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_35_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VPWR X VNB VPB
X0 a_27_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_27_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_277_297# B a_205_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR A a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_205_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND C a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_109_297# D a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VGND A a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VPWR X VNB VPB
X0 a_78_199# B1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VPWR A1 a_493_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_493_297# A2 a_78_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR a_78_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A2 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_78_199# B2 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_215_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_215_47# B2 a_78_199# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_292_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND a_78_199# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__or3_1 A B C VGND VPWR X VNB VPB
X0 X a_29_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_111_297# C a_29_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 X a_29_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_183_297# B a_111_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VPWR A a_183_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_29_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VGND C a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VGND A a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VPWR X VNB VPB
X0 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_27_297# B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VGND A2 a_373_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_27_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_373_47# A1 a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_109_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_109_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VPWR X VNB VPB
X0 a_240_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 X a_51_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VGND A1 a_240_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_51_297# B2 a_245_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_149_47# C1 a_51_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_240_47# B1 a_149_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR A1 a_512_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X a_51_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_149_47# B2 a_240_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_245_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR C1 a_51_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_512_297# A2 a_51_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VPWR X VNB VPB
X0 a_103_199# B1 a_253_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VPWR a_103_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_337_297# A2 a_253_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_103_199# A3 a_337_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_253_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR B1 a_103_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND a_103_199# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_253_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_253_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VGND A2 a_253_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and3_1 A B C VGND VPWR X VNB VPB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VPWR C a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_181_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VGND C a_181_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_27_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__or3_4 A B C VGND VPWR X VNB VPB
X0 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR A a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_193_297# B a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_109_297# C a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VGND C a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VPWR Y VNB VPB
X0 a_27_47# C a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_27_47# C a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_445_47# B a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_445_47# B a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_27_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_27_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 Y A a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 Y A a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_803_47# B a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_803_47# B a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VGND D a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_445_47# C a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_803_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 a_445_47# C a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 a_803_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 VGND D a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VPWR Y VNB VPB
X0 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_471_47# B a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_27_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_27_47# C a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_277_47# B a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 Y A a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_277_47# C a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_471_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND D a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VPWR X VNB VPB
X0 a_206_369# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_206_369# A2_N a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND B2 a_489_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_585_369# B2 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_489_47# a_206_369# a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_489_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR A2_N a_206_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_76_199# a_206_369# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_205_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR B1 a_585_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VPWR Y VNB VPB
X0 a_199_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_113_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A1 a_113_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_113_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND A2 a_199_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VPWR Y VNB VPB
X0 a_110_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y A2 a_110_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_326_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y C1 a_326_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VPWR X VNB VPB
X0 a_27_47# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_197_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_303_47# C a_197_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR D a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VGND D a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VPWR X VNB VPB
X0 VPWR A a_304_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_304_297# B a_220_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND C a_32_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_220_297# C a_114_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_32_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_32_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR a_32_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X a_32_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND A a_32_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR a_32_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 X a_32_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 X a_32_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 X a_32_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_114_297# D a_32_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VGND a_32_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VGND a_32_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VPWR X VNB VPB
X0 a_93_21# A1 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_93_21# B1 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_584_47# B1 a_93_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR a_93_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND B2 a_584_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_256_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_250_297# B2 a_93_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND a_93_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_250_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR A2 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_250_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_346_47# A2 a_256_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VPWR X VNB VPB
X0 a_75_199# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_208_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_315_47# A2 a_208_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND B1 a_75_199# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_75_199# A1 a_315_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_75_199# C1 a_544_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_544_297# B1 a_201_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR a_75_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_201_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR A2 a_201_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_201_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND a_75_199# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VPWR Y VNB VPB
X0 Y A1 a_181_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_181_47# A2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Y B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_109_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_109_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VPWR X VNB VPB
X0 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_109_53# D_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_215_297# a_109_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_392_297# C a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_465_297# B a_392_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_215_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR A a_465_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_297_297# a_109_53# a_215_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_109_53# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VGND C a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VGND A a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VPWR X VNB VPB
X0 VPWR B1 a_566_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_484_47# B1 a_96_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X a_96_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR a_96_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_96_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_566_297# B2 a_96_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR a_96_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X a_96_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VGND a_96_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_96_21# B2 a_566_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR A1 a_918_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_484_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_566_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_484_47# B2 a_96_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_96_21# A2 a_918_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_918_297# A2 a_96_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_484_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_918_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_96_21# B1 a_484_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 VGND A2 a_484_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_96_21# B2 a_484_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 VGND A1 a_484_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 X a_96_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VGND a_96_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VPWR X VNB VPB
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_209_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_303_47# A2 a_209_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_209_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_80_21# A1 a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR A2 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_80_21# B1 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_209_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VPWR X VNB VPB
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_80_21# C1 a_472_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A2 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_300_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_217_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_80_21# A1 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_472_297# B1 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_80_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VPWR Y VNB VPB
X0 a_27_47# B a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_27_47# B a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Y A a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y A a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_27_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_27_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_445_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_445_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND C a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_445_47# B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_445_47# B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VGND C a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VPWR X VNB VPB
X0 a_676_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_512_47# B1 a_409_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_306_47# D1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND A2 a_512_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR C1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR A1 a_676_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_512_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_409_47# C1 a_306_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_79_21# D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VPWR Y VNB VPB
X0 a_471_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_471_47# B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_471_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR A1 a_1241_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_471_47# B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_471_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_1241_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_27_47# B2 a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR B1 a_553_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND A2 a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_553_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_27_47# B2 a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VGND A2 a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_27_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VGND A1 a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 Y C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_27_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_1241_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 VPWR B1 a_553_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 VPWR A1 a_1241_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 Y B2 a_553_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 a_1241_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 a_553_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_471_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X28 Y A2 a_1241_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 a_553_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 a_27_47# B1 a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 VGND A1 a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X32 Y B2 a_553_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 a_1241_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 a_27_47# B1 a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X35 a_553_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 Y A2 a_1241_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X37 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 a_471_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X39 a_471_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VPWR X VNB VPB
X0 a_176_21# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VGND D_N a_27_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND a_176_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 X a_176_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR a_176_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_555_297# C a_483_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_176_21# a_27_53# a_555_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 X a_176_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_387_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_483_297# B a_387_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VGND B a_176_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VGND a_27_53# a_176_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 VPWR D_N a_27_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 a_176_21# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VPWR X VNB VPB
X0 VPWR a_315_380# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X a_315_380# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_315_380# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND C_N a_27_410# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VPWR C_N a_27_410# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR A a_583_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND a_27_410# a_315_380# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_583_297# B a_499_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND A a_315_380# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_397_297# a_205_93# a_315_380# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 X a_315_380# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 X a_315_380# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_499_297# a_27_410# a_397_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VPWR a_315_380# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_205_93# D_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_205_93# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 VGND a_315_380# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VGND a_315_380# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_315_380# a_205_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 X a_315_380# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__ebufn_2 A TE_B VGND VPWR Z VNB VPB
X0 a_320_309# a_27_47# Z VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Z a_27_47# a_320_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 VGND a_214_47# a_392_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_214_47# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5 a_320_309# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X6 a_392_47# a_214_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR TE_B a_320_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X8 Z a_27_47# a_392_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_214_47# TE_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_392_47# a_27_47# Z VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VPWR Y VNB VPB
X0 a_286_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_286_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y A2 a_487_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A1 a_286_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND A2 a_286_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_487_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_27_47# B1 a_286_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR A1 a_487_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_27_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_487_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_286_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VPWR Y VNB VPB
X0 a_27_47# C1 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_803_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_27_47# C1 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND A2 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_1163_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND A2 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Y A2 a_1163_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_1163_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_445_47# B1 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR D1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_445_47# B1 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 Y D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VPWR A1 a_1163_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_27_47# D1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_27_47# D1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VGND A1 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_1163_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_803_47# B1 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 VPWR A1 a_1163_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 a_803_47# B1 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 Y D1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_445_47# C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 a_803_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 a_1163_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 Y A2 a_1163_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 a_445_47# C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X34 a_803_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X35 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 a_803_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X37 VPWR D1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 Y D1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X39 VGND A1 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VPWR Y VNB VPB
X0 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_27_47# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR A1 a_307_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_307_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_109_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VPWR X VNB VPB
X0 a_465_47# A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_109_297# B1 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_205_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR A2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_193_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_27_47# B1 a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_109_297# C1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VGND C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND A2 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VPWR Y VNB VPB
X0 a_109_47# B1 a_213_123# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Y B2 a_295_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A1 a_493_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_213_123# B2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_295_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_493_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND A2 a_213_123# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_213_123# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_109_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VPWR Y VNB VPB
X0 Y B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Y B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_381_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_109_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_109_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND A2 a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VPWR X VNB VPB
X0 VGND A2 a_660_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VGND C1 a_85_193# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_414_297# C1 a_334_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND a_85_193# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_334_297# D1 a_85_193# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_516_297# B1 a_414_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_516_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_660_47# A1 a_85_193# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_85_193# D1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR A1 a_516_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_85_193# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR a_85_193# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor2_4 A B VGND VPWR Y VNB VPB
X0 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VPWR X VNB VPB
X0 a_381_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR A2 a_381_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_465_47# A4 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_549_47# A3 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_665_47# A2 a_549_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_381_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR A4 a_381_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_381_297# B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_79_21# A1 a_665_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VPWR X VNB VPB
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X a_80_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_80_21# D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR C1 a_80_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 X a_80_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_80_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_674_297# A2 a_80_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_386_47# D1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR A1 a_674_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_566_47# B1 a_458_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND A2 a_566_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_566_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_458_47# C1 a_386_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VPWR X VNB VPB
X0 a_77_199# B2 a_227_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_323_297# A2 a_227_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_227_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_227_47# B1 a_77_199# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND a_77_199# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR B1 a_539_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_227_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR a_77_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_77_199# A3 a_323_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND A2 a_227_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_227_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_539_297# B2 a_77_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VPWR X VNB VPB
X0 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_79_21# A0 a_792_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_1259_199# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_1302_47# A0 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X8 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_792_297# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_1259_199# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND a_1259_199# a_1302_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X14 a_79_21# A1 a_792_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X15 a_79_21# A0 a_1302_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X16 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VPWR S a_792_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_792_297# A0 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_1302_47# a_1259_199# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X23 VPWR a_1259_199# a_1302_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 a_1302_297# a_1259_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 a_792_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X27 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_1302_297# A1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VGND S a_792_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X30 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 a_79_21# A1 a_1302_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X33 a_792_47# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VPWR Y VNB VPB
X0 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_115_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_115_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR A1 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A2 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y B1 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND A1 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_32_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 Y B1 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y A2 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_32_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_32_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_32_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_115_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_32_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_32_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VGND A2 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VPWR A1 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 Y A2 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 VGND A1 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_115_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VPWR X VNB VPB
X0 a_226_47# A2_N a_226_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_489_413# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_226_297# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR B2 a_489_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_489_413# a_226_47# a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_76_199# a_226_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VGND B1 a_556_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_556_47# B2 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VGND A2_N a_226_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_226_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VPWR X VNB VPB
X0 a_109_93# C_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_215_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND a_109_93# a_215_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VGND A a_215_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VPWR A a_369_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_369_297# B a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 X a_215_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_297_297# a_109_93# a_215_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_109_93# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 X a_215_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkinvlp_2 A VGND VPWR Y VNB VPB
X0 Y A a_150_67# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=250000u
X2 a_150_67# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X3 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=250000u
.ends

.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VPWR Y VNB VPB
X0 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_193_47# C a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y A a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_277_47# B a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_109_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VPWR X VNB VPB
X0 a_585_47# B1 a_266_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VGND A2 a_266_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_81_21# C1 a_585_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_266_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_368_297# A2 a_266_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_266_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_266_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_81_21# A3 a_368_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_81_21# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VPWR B1 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VPWR Y VNB VPB
X0 a_281_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_475_297# D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y D a_475_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND D Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_475_297# C a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_281_297# C a_475_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_27_297# B a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VPWR Y VNB VPB
X0 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_449_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_27_297# B a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y C a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_449_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y C a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_449_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_27_297# B a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 a_449_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VPWR X VNB VPB
X0 VPWR D a_343_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_223_47# B_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_515_93# a_223_47# a_429_93# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_223_47# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 X a_343_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_429_93# a_27_47# a_343_93# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VGND D a_615_93# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_343_93# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_343_93# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_615_93# C a_515_93# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 X a_343_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VPWR a_223_47# a_343_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VPWR X VNB VPB
X0 a_204_297# A1 a_396_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR a_396_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 X a_396_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR S a_314_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_204_297# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_396_47# A0 a_314_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_206_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 X a_396_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 X a_396_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR a_396_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_490_47# A1 a_396_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND S a_490_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND a_396_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_396_47# A0 a_206_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VGND a_396_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VPWR S a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 X a_396_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VGND S a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VPWR X VNB VPB
X0 a_27_47# B1 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_109_47# A2 a_717_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_717_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND A2 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_277_297# B2 a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_109_47# B2 a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_277_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_277_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_277_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VPWR C1 a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_27_47# C1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_27_47# B2 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VGND A1 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_277_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_277_47# B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 VPWR B1 a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 VPWR A1 a_717_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 a_109_47# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 a_717_297# A2 a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_109_47# C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VPWR X VNB VPB
X0 X a_79_204# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR A1 a_473_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_473_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_79_204# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND C1 a_79_204# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_79_204# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR a_79_204# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_473_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_473_297# B1 a_727_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X a_79_204# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND B1 a_79_204# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_79_204# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND a_79_204# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_1123_47# A1 a_79_204# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_555_297# B1 a_473_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VPWR A2 a_473_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VGND A2 a_1123_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_951_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VPWR a_79_204# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND a_79_204# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_79_204# A1 a_951_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 a_79_204# C1 a_555_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_727_297# C1 a_79_204# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 X a_79_204# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VPWR X VNB VPB
X0 VGND A a_311_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VPWR A a_561_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_393_413# a_205_93# a_311_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VGND C_N a_27_410# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VPWR C_N a_27_410# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 X a_311_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND a_27_410# a_311_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_561_297# B a_489_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_205_93# D_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_205_93# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_489_297# a_27_410# a_393_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_311_413# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_311_413# a_205_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 X a_311_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VPWR Y VNB VPB
X0 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_191_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_297_297# B a_191_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_109_297# D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VPWR Y VNB VPB
X0 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_235_47# C1 a_163_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_343_47# B1 a_235_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_454_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR A1 a_454_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_163_47# D1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VGND A2 a_343_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_343_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VPWR X VNB VPB
X0 VPWR a_86_235# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND C1 a_86_235# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X a_86_235# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_86_235# D1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 X a_86_235# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_715_47# A1 a_86_235# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND A2 a_715_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_499_297# C1 a_427_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND a_86_235# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_86_235# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_607_297# B1 a_499_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_427_297# D1 a_86_235# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VPWR A1 a_607_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_607_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VPWR Y VNB VPB
X0 Y A1 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_641_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_109_297# B1 a_641_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_277_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_109_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR A3 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_27_47# A2 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_641_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_277_47# A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_109_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 Y C1 a_641_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VPWR X VNB VPB
X0 VPWR A a_300_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_218_297# a_27_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND B_N a_27_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_300_297# a_27_53# a_218_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 X a_218_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR a_218_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 X a_218_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND a_218_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_27_53# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VGND A a_218_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VPWR X VNB VPB
X0 a_176_21# a_27_47# a_626_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_626_297# B a_542_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR C_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VGND a_176_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_542_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR a_176_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 X a_176_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X a_176_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 X a_176_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_176_21# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VPWR a_176_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 X a_176_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_176_21# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND a_176_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VGND B a_176_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VGND C_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VPWR X VNB VPB
X0 a_222_93# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VPWR A1 a_544_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND a_79_199# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_222_93# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VGND A2 a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_448_47# a_222_93# a_79_199# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_79_199# a_222_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_544_297# A2 a_79_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_448_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR a_79_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VPWR Y VNB VPB
X0 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y A1 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 Y A1 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND A2 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_27_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_27_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_803_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_803_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_803_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_803_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 VGND B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 VGND A2 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 VGND B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VPWR X VNB VPB
X0 a_465_47# A2 a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VGND A4 a_561_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR A3 a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_297_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_297_297# A4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR A1 a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_381_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_297_297# B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_79_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_561_47# A3 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VPWR Y VNB VPB
X0 Y A1 a_194_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_194_47# A2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y C1 a_376_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_376_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_109_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_109_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VPWR Y VNB VPB
X0 Y C a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_281_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_281_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_27_297# B a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VPWR X VNB VPB
X0 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND a_215_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR a_215_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_109_93# D_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_215_297# a_109_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND C a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND A a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_215_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_109_93# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VPWR A a_487_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND a_215_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_487_297# B a_403_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_403_297# C a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VPWR a_215_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_297_297# a_109_93# a_215_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VPWR X VNB VPB
X0 a_109_93# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 X a_209_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_109_93# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_296_53# a_109_93# a_209_311# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VPWR C a_209_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_368_53# B a_296_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 X a_209_311# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_209_311# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VPWR a_109_93# a_209_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VGND C a_368_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor2_8 A B VGND VPWR Y VNB VPB
X0 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VPWR Y VNB VPB
X0 a_991_47# C a_633_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_991_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_991_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_633_47# B a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_633_47# B a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND D a_991_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND D a_991_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_215_47# a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_215_47# B a_633_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_215_47# B a_633_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 a_633_47# C a_991_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 a_633_47# C a_991_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_215_47# a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 a_991_47# C a_633_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X32 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand4bb_1 A_N B_N C D VGND VPWR Y VNB VPB
X0 VGND B_N a_27_93# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_496_21# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 Y a_496_21# a_426_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR a_496_21# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_426_47# a_27_93# a_326_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR B_N a_27_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_496_21# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 Y a_27_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_218_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_326_47# C a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VPWR X VNB VPB
X0 a_388_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VPWR C_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND a_176_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 X a_176_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR a_176_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND B a_176_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 X a_176_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_176_21# a_27_47# a_472_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_472_297# B a_388_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_176_21# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_176_21# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VGND C_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VPWR X VNB VPB
X0 a_297_47# a_27_47# a_193_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_369_47# B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VPWR D a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 X a_193_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND D a_469_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 X a_193_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR B a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_193_413# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_193_413# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_469_47# C a_369_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VPWR Y VNB VPB
X0 Y A3 a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_449_297# A3 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y A3 a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A1 a_31_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y B1 a_31_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_449_297# A3 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Y B1 a_31_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_31_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_27_297# A2 a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND A1 a_31_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_31_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_31_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_31_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_449_297# A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VGND A2 a_31_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 VGND A2 a_31_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 VGND A3 a_31_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 a_31_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 a_27_297# A2 a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 VGND A3 a_31_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 a_31_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X28 a_449_297# A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 a_31_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 a_31_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and3_4 A B C VGND VPWR X VNB VPB
X0 VPWR A a_94_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_294_47# B a_185_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_185_47# A a_94_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR a_94_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND C a_294_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_94_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 X a_94_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X a_94_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR C a_94_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X a_94_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND a_94_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR a_94_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND a_94_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 X a_94_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VPWR Y VNB VPB
X0 a_33_47# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VGND A1 a_33_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VGND A2 a_33_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_33_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_797_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y A2 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_797_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y B2 a_797_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_115_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR B1 a_797_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_33_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND A1 a_33_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_33_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_33_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 Y A2 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_33_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_797_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_115_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 VPWR A1 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VPWR B1 a_797_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VGND A2 a_33_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 a_33_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 a_797_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR A1 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 Y B2 a_33_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 Y B2 a_797_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 Y B1 a_33_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 Y B2 a_33_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X28 a_115_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 Y B1 a_33_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 a_33_47# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 a_115_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt housekeeping debug_in debug_mode debug_oeb debug_out irq[0] irq[1] irq[2]
+ mask_rev_in[0] mask_rev_in[10] mask_rev_in[11] mask_rev_in[12] mask_rev_in[13] mask_rev_in[14]
+ mask_rev_in[15] mask_rev_in[16] mask_rev_in[17] mask_rev_in[18] mask_rev_in[19]
+ mask_rev_in[1] mask_rev_in[20] mask_rev_in[21] mask_rev_in[22] mask_rev_in[23] mask_rev_in[24]
+ mask_rev_in[25] mask_rev_in[26] mask_rev_in[27] mask_rev_in[28] mask_rev_in[29]
+ mask_rev_in[2] mask_rev_in[30] mask_rev_in[31] mask_rev_in[3] mask_rev_in[4] mask_rev_in[5]
+ mask_rev_in[6] mask_rev_in[7] mask_rev_in[8] mask_rev_in[9] mgmt_gpio_in[0] mgmt_gpio_in[10]
+ mgmt_gpio_in[11] mgmt_gpio_in[12] mgmt_gpio_in[13] mgmt_gpio_in[14] mgmt_gpio_in[15]
+ mgmt_gpio_in[16] mgmt_gpio_in[17] mgmt_gpio_in[18] mgmt_gpio_in[19] mgmt_gpio_in[1]
+ mgmt_gpio_in[20] mgmt_gpio_in[21] mgmt_gpio_in[22] mgmt_gpio_in[23] mgmt_gpio_in[24]
+ mgmt_gpio_in[25] mgmt_gpio_in[26] mgmt_gpio_in[27] mgmt_gpio_in[28] mgmt_gpio_in[29]
+ mgmt_gpio_in[2] mgmt_gpio_in[30] mgmt_gpio_in[31] mgmt_gpio_in[32] mgmt_gpio_in[33]
+ mgmt_gpio_in[34] mgmt_gpio_in[35] mgmt_gpio_in[36] mgmt_gpio_in[37] mgmt_gpio_in[3]
+ mgmt_gpio_in[4] mgmt_gpio_in[5] mgmt_gpio_in[6] mgmt_gpio_in[7] mgmt_gpio_in[8]
+ mgmt_gpio_in[9] mgmt_gpio_oeb[0] mgmt_gpio_oeb[10] mgmt_gpio_oeb[11] mgmt_gpio_oeb[12]
+ mgmt_gpio_oeb[13] mgmt_gpio_oeb[14] mgmt_gpio_oeb[15] mgmt_gpio_oeb[16] mgmt_gpio_oeb[17]
+ mgmt_gpio_oeb[18] mgmt_gpio_oeb[19] mgmt_gpio_oeb[1] mgmt_gpio_oeb[20] mgmt_gpio_oeb[21]
+ mgmt_gpio_oeb[22] mgmt_gpio_oeb[23] mgmt_gpio_oeb[24] mgmt_gpio_oeb[25] mgmt_gpio_oeb[26]
+ mgmt_gpio_oeb[27] mgmt_gpio_oeb[28] mgmt_gpio_oeb[29] mgmt_gpio_oeb[2] mgmt_gpio_oeb[30]
+ mgmt_gpio_oeb[31] mgmt_gpio_oeb[32] mgmt_gpio_oeb[33] mgmt_gpio_oeb[34] mgmt_gpio_oeb[35]
+ mgmt_gpio_oeb[36] mgmt_gpio_oeb[37] mgmt_gpio_oeb[3] mgmt_gpio_oeb[4] mgmt_gpio_oeb[5]
+ mgmt_gpio_oeb[6] mgmt_gpio_oeb[7] mgmt_gpio_oeb[8] mgmt_gpio_oeb[9] mgmt_gpio_out[0]
+ mgmt_gpio_out[10] mgmt_gpio_out[11] mgmt_gpio_out[12] mgmt_gpio_out[13] mgmt_gpio_out[14]
+ mgmt_gpio_out[15] mgmt_gpio_out[16] mgmt_gpio_out[17] mgmt_gpio_out[18] mgmt_gpio_out[19]
+ mgmt_gpio_out[1] mgmt_gpio_out[20] mgmt_gpio_out[21] mgmt_gpio_out[22] mgmt_gpio_out[23]
+ mgmt_gpio_out[24] mgmt_gpio_out[25] mgmt_gpio_out[26] mgmt_gpio_out[27] mgmt_gpio_out[28]
+ mgmt_gpio_out[29] mgmt_gpio_out[2] mgmt_gpio_out[30] mgmt_gpio_out[31] mgmt_gpio_out[32]
+ mgmt_gpio_out[33] mgmt_gpio_out[34] mgmt_gpio_out[35] mgmt_gpio_out[36] mgmt_gpio_out[37]
+ mgmt_gpio_out[3] mgmt_gpio_out[4] mgmt_gpio_out[5] mgmt_gpio_out[6] mgmt_gpio_out[7]
+ mgmt_gpio_out[8] mgmt_gpio_out[9] pad_flash_clk pad_flash_clk_oeb pad_flash_csb
+ pad_flash_csb_oeb pad_flash_io0_di pad_flash_io0_do pad_flash_io0_ieb pad_flash_io0_oeb
+ pad_flash_io1_di pad_flash_io1_do pad_flash_io1_ieb pad_flash_io1_oeb pll90_sel[0]
+ pll90_sel[1] pll90_sel[2] pll_bypass pll_dco_ena pll_div[0] pll_div[1] pll_div[2]
+ pll_div[3] pll_div[4] pll_ena pll_sel[0] pll_sel[1] pll_sel[2] pll_trim[0] pll_trim[10]
+ pll_trim[11] pll_trim[12] pll_trim[13] pll_trim[14] pll_trim[15] pll_trim[16] pll_trim[17]
+ pll_trim[18] pll_trim[19] pll_trim[1] pll_trim[20] pll_trim[21] pll_trim[22] pll_trim[23]
+ pll_trim[24] pll_trim[25] pll_trim[2] pll_trim[3] pll_trim[4] pll_trim[5] pll_trim[6]
+ pll_trim[7] pll_trim[8] pll_trim[9] porb pwr_ctrl_out[0] pwr_ctrl_out[1] pwr_ctrl_out[2]
+ pwr_ctrl_out[3] qspi_enabled reset ser_rx ser_tx serial_clock serial_data_1 serial_data_2
+ serial_load serial_resetn spi_csb spi_enabled spi_sck spi_sdi spi_sdo spi_sdoenb
+ spimemio_flash_clk spimemio_flash_csb spimemio_flash_io0_di spimemio_flash_io0_do
+ spimemio_flash_io0_oeb spimemio_flash_io1_di spimemio_flash_io1_do spimemio_flash_io1_oeb
+ spimemio_flash_io2_di spimemio_flash_io2_do spimemio_flash_io2_oeb spimemio_flash_io3_di
+ spimemio_flash_io3_do spimemio_flash_io3_oeb sram_ro_addr[0] sram_ro_addr[1] sram_ro_addr[2]
+ sram_ro_addr[3] sram_ro_addr[4] sram_ro_addr[5] sram_ro_addr[6] sram_ro_addr[7]
+ sram_ro_clk sram_ro_csb sram_ro_data[0] sram_ro_data[10] sram_ro_data[11] sram_ro_data[12]
+ sram_ro_data[13] sram_ro_data[14] sram_ro_data[15] sram_ro_data[16] sram_ro_data[17]
+ sram_ro_data[18] sram_ro_data[19] sram_ro_data[1] sram_ro_data[20] sram_ro_data[21]
+ sram_ro_data[22] sram_ro_data[23] sram_ro_data[24] sram_ro_data[25] sram_ro_data[26]
+ sram_ro_data[27] sram_ro_data[28] sram_ro_data[29] sram_ro_data[2] sram_ro_data[30]
+ sram_ro_data[31] sram_ro_data[3] sram_ro_data[4] sram_ro_data[5] sram_ro_data[6]
+ sram_ro_data[7] sram_ro_data[8] sram_ro_data[9] trap uart_enabled user_clock usr1_vcc_pwrgood
+ usr1_vdd_pwrgood usr2_vcc_pwrgood usr2_vdd_pwrgood wb_ack_o wb_adr_i[0] wb_adr_i[10]
+ wb_adr_i[11] wb_adr_i[12] wb_adr_i[13] wb_adr_i[14] wb_adr_i[15] wb_adr_i[16] wb_adr_i[17]
+ wb_adr_i[18] wb_adr_i[19] wb_adr_i[1] wb_adr_i[20] wb_adr_i[21] wb_adr_i[22] wb_adr_i[23]
+ wb_adr_i[24] wb_adr_i[25] wb_adr_i[26] wb_adr_i[27] wb_adr_i[28] wb_adr_i[29] wb_adr_i[2]
+ wb_adr_i[30] wb_adr_i[31] wb_adr_i[3] wb_adr_i[4] wb_adr_i[5] wb_adr_i[6] wb_adr_i[7]
+ wb_adr_i[8] wb_adr_i[9] wb_clk_i wb_cyc_i wb_dat_i[0] wb_dat_i[10] wb_dat_i[11]
+ wb_dat_i[12] wb_dat_i[13] wb_dat_i[14] wb_dat_i[15] wb_dat_i[16] wb_dat_i[17] wb_dat_i[18]
+ wb_dat_i[19] wb_dat_i[1] wb_dat_i[20] wb_dat_i[21] wb_dat_i[22] wb_dat_i[23] wb_dat_i[24]
+ wb_dat_i[25] wb_dat_i[26] wb_dat_i[27] wb_dat_i[28] wb_dat_i[29] wb_dat_i[2] wb_dat_i[30]
+ wb_dat_i[31] wb_dat_i[3] wb_dat_i[4] wb_dat_i[5] wb_dat_i[6] wb_dat_i[7] wb_dat_i[8]
+ wb_dat_i[9] wb_dat_o[0] wb_dat_o[10] wb_dat_o[11] wb_dat_o[12] wb_dat_o[13] wb_dat_o[14]
+ wb_dat_o[15] wb_dat_o[16] wb_dat_o[17] wb_dat_o[18] wb_dat_o[19] wb_dat_o[1] wb_dat_o[20]
+ wb_dat_o[21] wb_dat_o[22] wb_dat_o[23] wb_dat_o[24] wb_dat_o[25] wb_dat_o[26] wb_dat_o[27]
+ wb_dat_o[28] wb_dat_o[29] wb_dat_o[2] wb_dat_o[30] wb_dat_o[31] wb_dat_o[3] wb_dat_o[4]
+ wb_dat_o[5] wb_dat_o[6] wb_dat_o[7] wb_dat_o[8] wb_dat_o[9] wb_rstn_i wb_sel_i[0]
+ wb_sel_i[1] wb_sel_i[2] wb_sel_i[3] wb_stb_i wb_we_i VGND VPWR
XFILLER_67_553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_288 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7963_ _7979_/A _7994_/B VGND VPWR _8096_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_9702_ _4446_/A1 _9702_/D _4981_/X VGND VPWR _9702_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6914_ _9287_/Q VGND VPWR _6914_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_82_556 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7894_ _8583_/A _7894_/B _7903_/C _8193_/A VGND VPWR _7895_/A VGND VPWR sky130_fd_sc_hd__or4_1
XFILLER_52_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_111 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6845_ _9537_/Q VGND VPWR _6845_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9633_ _9639_/CLK _9633_/D _9633_/SET_B VGND VPWR _9633_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_50_453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_144 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6776_ _6774_/Y _5121_/B _6775_/Y _5949_/B VGND VPWR _6776_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_9564_ _9617_/CLK _9564_/D _9295_/SET_B VGND VPWR _9564_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_9495_ _9534_/CLK _9495_/D _9647_/SET_B VGND VPWR _9495_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_8515_ _8515_/A _8515_/B VGND VPWR _8703_/B VGND VPWR sky130_fd_sc_hd__nor2_1
X_5727_ _7041_/A _7127_/C VGND VPWR _5728_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_108_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_8446_ _7864_/X _8341_/B _8009_/X _8445_/X _8013_/X VGND VPWR _8448_/C VGND VPWR
+ sky130_fd_sc_hd__o2111ai_2
XFILLER_175_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8377_ _8583_/C _8377_/B _8377_/C VGND VPWR _8565_/A VGND VPWR sky130_fd_sc_hd__or3_1
X_5589_ _9316_/Q _5585_/A _8925_/A1 _5585_/Y VGND VPWR _9316_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_4609_ _9727_/Q _4604_/A _5966_/B1 _4604_/Y VGND VPWR _9727_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_104_400 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7328_ _6812_/Y _7126_/X _6868_/Y _7128_/X VGND VPWR _7328_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_7259_ _6218_/Y _7059_/D _6152_/Y _7116_/X _7258_/X VGND VPWR _7264_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_131_263 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_488 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_48 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA_202 input83/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_213 _6073_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_26_472 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_108 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_396 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_219 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_61 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_571 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_92 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_331 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_556 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4960_ _6022_/A _6022_/B _6022_/C _9708_/Q VGND VPWR _4960_/X VGND VPWR sky130_fd_sc_hd__o31a_1
X_4891_ _4891_/A _4911_/A VGND VPWR _5450_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_6630_ _6149_/A _6629_/Y _9039_/Q _6149_/Y VGND VPWR _9039_/D VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_165_609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6561_ _6561_/A VGND VPWR _6561_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_164_108 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5512_ _9369_/Q _5509_/A _8844_/X _5509_/Y VGND VPWR _9369_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8300_ _8496_/A _8300_/B VGND VPWR _8301_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_145_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_9280_ _9280_/CLK _9280_/D _9757_/SET_B VGND VPWR _9280_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6492_ _9207_/Q VGND VPWR _8751_/A VGND VPWR sky130_fd_sc_hd__inv_6
XFILLER_172_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8231_ _8231_/A _8676_/B _8658_/B _8573_/B VGND VPWR _8237_/A VGND VPWR sky130_fd_sc_hd__or4_1
X_5443_ _5443_/A VGND VPWR _5444_/A VGND VPWR sky130_fd_sc_hd__clkbuf_2
X_8162_ _8162_/A _8370_/A VGND VPWR _8163_/B VGND VPWR sky130_fd_sc_hd__or2_1
X_5374_ _5671_/A _5374_/B VGND VPWR _5375_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_7113_ _4742_/Y _7112_/X _4668_/Y _7077_/B VGND VPWR _7113_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_141_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_252 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8093_ _8093_/A _8093_/B VGND VPWR _8431_/A VGND VPWR sky130_fd_sc_hd__nor2_1
X_7044_ _7075_/A _7115_/B VGND VPWR _7045_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_82_320 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_534 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8995_ _9563_/Q _8767_/A VGND VPWR mgmt_gpio_out[18] VGND VPWR sky130_fd_sc_hd__ebufn_8
XFILLER_82_386 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7946_ _8379_/C _8195_/A VGND VPWR _8079_/C VGND VPWR sky130_fd_sc_hd__or2_1
X_7877_ _8515_/B _8232_/B VGND VPWR _7877_/X VGND VPWR sky130_fd_sc_hd__or2_2
X_6828_ _6823_/Y _6027_/B _6824_/Y _5336_/B _6827_/X VGND VPWR _6829_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_2
X_9616_ _9788_/CLK _9616_/D _9646_/SET_B VGND VPWR _9616_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_156_609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_514 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_9547_ _9639_/CLK _9547_/D _9757_/SET_B VGND VPWR _9547_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6759_ _6759_/A _6759_/B _6759_/C VGND VPWR _6784_/C VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_148_182 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_118 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9478_ _9483_/CLK _9478_/D _9685_/SET_B VGND VPWR _9478_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_163_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_152 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_8429_ _8703_/A _8585_/B VGND VPWR _8560_/B VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_163_174 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_302 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_320 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_247 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_73 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_62 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_191 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_386 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_439 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_491 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_550 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5090_ _5090_/A VGND VPWR _5091_/A VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_96_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7800_ _8379_/C _7839_/A _8379_/D VGND VPWR _8093_/A VGND VPWR sky130_fd_sc_hd__or3_4
X_5992_ _9698_/Q _5992_/B VGND VPWR _7008_/B VGND VPWR sky130_fd_sc_hd__nand2_1
X_8780_ _8780_/A VGND VPWR _8780_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_24_239 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4943_ _6022_/A _6022_/D _6022_/C VGND VPWR _4944_/A VGND VPWR sky130_fd_sc_hd__or3_1
X_5848__6 _8924_/X VGND VPWR _5893_/A1 VGND VPWR sky130_fd_sc_hd__inv_4
X_7731_ _7731_/A _8975_/S VGND VPWR _7732_/A VGND VPWR sky130_fd_sc_hd__and2_1
X_7662_ _7662_/A _7662_/B _7662_/C _7662_/D VGND VPWR _7662_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
X_4874_ _9726_/Q VGND VPWR _4874_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_6613_ _8771_/A _5420_/B _6612_/Y _5442_/B VGND VPWR _6613_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_9401_ _9758_/CLK _9401_/D _7011_/B VGND VPWR _9401_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_7593_ _6129_/Y _7419_/X _6116_/Y _7421_/X VGND VPWR _7593_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_20_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9332_ _9545_/CLK _9332_/D _4628_/A VGND VPWR _9332_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6544_ _9635_/Q VGND VPWR _6544_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_145_152 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_19 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6475_ _6475_/A _6475_/B _6475_/C _6475_/D VGND VPWR _6475_/Y VGND VPWR sky130_fd_sc_hd__nand4_2
X_9263_ _9601_/CLK _9263_/D _9295_/SET_B VGND VPWR _9263_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_8214_ _8311_/B VGND VPWR _8214_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_5426_ _9428_/Q _5422_/A _8925_/A1 _5422_/Y VGND VPWR _9428_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_145_196 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_9194_ _9378_/CLK _9194_/D _9646_/SET_B VGND VPWR _9194_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
Xoutput253 _7010_/Y VGND VPWR pad_flash_csb_oeb VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput242 _7700_/X VGND VPWR mgmt_gpio_oeb[7] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput220 _8774_/X VGND VPWR mgmt_gpio_oeb[21] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput231 _8794_/X VGND VPWR mgmt_gpio_oeb[31] VGND VPWR sky130_fd_sc_hd__buf_2
X_8145_ _7987_/Y _8390_/B _8144_/X VGND VPWR _8145_/X VGND VPWR sky130_fd_sc_hd__a21o_1
Xoutput264 _9720_/Q VGND VPWR pll_dco_ena VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput275 _9742_/Q VGND VPWR pll_trim[10] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput286 _9752_/Q VGND VPWR pll_trim[20] VGND VPWR sky130_fd_sc_hd__buf_2
X_5357_ _5357_/A VGND VPWR _5357_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_5288_ _9520_/Q _5280_/A _8916_/A1 _5280_/Y VGND VPWR _9520_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8076_ _8515_/B _8437_/B _8075_/Y VGND VPWR _8078_/A VGND VPWR sky130_fd_sc_hd__o21ai_1
Xoutput297 _9739_/Q VGND VPWR pll_trim[7] VGND VPWR sky130_fd_sc_hd__buf_2
X_7027_ _7027_/A VGND VPWR _7073_/C VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_15_206 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8978_ _7482_/X _4875_/Y _8978_/S VGND VPWR _8978_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_7929_ _7929_/A _7929_/B VGND VPWR _7929_/Y VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_11_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_119 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_214 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_344 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_388 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_483 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_24 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xnet299_3 _8837_/A1 VGND VPWR _6359_/A1 VGND VPWR sky130_fd_sc_hd__inv_4
XFILLER_159_244 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_294 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4590_ _5960_/A _4590_/B VGND VPWR _4591_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_143_612 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6260_ _6258_/Y _4590_/B _6259_/Y _6086_/X VGND VPWR _6260_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_5211_ _9570_/Q _5203_/Y _8916_/X _5203_/A VGND VPWR _9570_/D VGND VPWR sky130_fd_sc_hd__o22a_1
X_6191_ input41/X _8930_/S _6190_/Y _5431_/B VGND VPWR _6191_/X VGND VPWR sky130_fd_sc_hd__o2bb2a_1
XFILLER_111_531 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_423 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5142_ _9620_/Q _5136_/A _8955_/A1 _5136_/Y VGND VPWR _9620_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_96_231 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5073_ _5073_/A VGND VPWR _9662_/D VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_8901_ _7728_/X _9698_/Q _9048_/Q VGND VPWR _8901_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_84_448 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_8832_ _6544_/Y _9058_/Q _8977_/S VGND VPWR _8832_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_12_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5975_ _9096_/Q _5970_/A _8929_/A1 _5970_/Y VGND VPWR _9096_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8763_ _8763_/A VGND VPWR _8764_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_7714_ _9084_/Q _7713_/B _9085_/Q VGND VPWR _7715_/B VGND VPWR sky130_fd_sc_hd__a21oi_1
X_8694_ _8496_/A _8216_/X _8312_/D _7905_/X VGND VPWR _8695_/B VGND VPWR sky130_fd_sc_hd__o211ai_1
X_4926_ _9502_/Q VGND VPWR _4926_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
X_4857_ _9778_/Q VGND VPWR _4857_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7645_ _6729_/Y _7408_/X _6685_/Y _7410_/X VGND VPWR _7645_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_176_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7576_ _6182_/Y _7415_/X _6215_/Y _7417_/X _7575_/X VGND VPWR _7590_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_193_578 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4788_ _4784_/Y _5941_/B _4786_/Y _5488_/B VGND VPWR _4788_/X VGND VPWR sky130_fd_sc_hd__o22a_2
X_9315_ _9535_/CLK _9315_/D _9647_/SET_B VGND VPWR _9315_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6527_ _9367_/Q VGND VPWR _8799_/A VGND VPWR sky130_fd_sc_hd__inv_6
XFILLER_106_303 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_9246_ _9278_/CLK _9246_/D _9779_/SET_B VGND VPWR _9246_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
X_6458_ _9105_/Q VGND VPWR _6458_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
XFILLER_121_306 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5409_ _9439_/Q _5406_/A _5965_/B1 _5406_/Y VGND VPWR _9439_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_9177_ _9613_/CLK _9177_/D _9646_/SET_B VGND VPWR _9177_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6389_ _6384_/Y _4564_/B _6385_/Y _4907_/X _6388_/X VGND VPWR _6408_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_2
XFILLER_161_497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8128_ _8130_/B _8640_/B VGND VPWR _8676_/A VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_125_77 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_275 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_8059_ _8085_/A VGND VPWR _8064_/B VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_18_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_98 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_96 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_247 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_246 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_567 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_100 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_62 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_61 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_320 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5760_ _9238_/Q _5759_/A _8846_/X _5759_/Y VGND VPWR _9238_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_187_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_91 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4711_ _4931_/A _4780_/B VGND VPWR _5632_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_5691_ _5691_/A _9055_/Q VGND VPWR _5692_/A VGND VPWR sky130_fd_sc_hd__or2_2
XFILLER_175_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7430_ _7430_/A VGND VPWR _7430_/X VGND VPWR sky130_fd_sc_hd__buf_6
X_4642_ _4642_/A VGND VPWR _4642_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_175_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7361_ _6577_/Y _7079_/B _6510_/Y _7059_/A VGND VPWR _7361_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4573_ _9749_/Q _4566_/A _5966_/B1 _4566_/Y VGND VPWR _9749_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_6312_ _6310_/Y _6081_/B _6311_/Y _5583_/B VGND VPWR _6312_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_7292_ _4761_/Y _7048_/B _4784_/Y _7077_/A _7291_/X VGND VPWR _7299_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9100_ _9652_/CLK _9100_/D _9647_/SET_B VGND VPWR _9100_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6243_ _9745_/Q VGND VPWR _6243_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9031_ _9039_/CLK _9031_/D VGND VPWR _9031_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_115_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6174_ _6174_/A _6174_/B _6174_/C _6174_/D VGND VPWR _6237_/A VGND VPWR sky130_fd_sc_hd__and4_1
X_5125_ _9630_/Q _5123_/A _5964_/B1 _5123_/Y VGND VPWR _9630_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_84_234 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5056_ _7733_/A _7734_/A _8810_/A VGND VPWR _5062_/A VGND VPWR sky130_fd_sc_hd__a21oi_1
XFILLER_52_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_1_wb_clk_i clkbuf_1_0_1_wb_clk_i/A VGND VPWR clkbuf_2_1_0_wb_clk_i/A VGND
+ VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_40_304 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5958_ _9107_/Q _5951_/A _8930_/A1 _5951_/Y VGND VPWR _9107_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8746_ _8746_/A VGND VPWR _8746_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_52_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_540 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4909_ _9758_/Q VGND VPWR _4909_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_21_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8677_ _8677_/A _8677_/B _8677_/C _8677_/D VGND VPWR _8731_/D VGND VPWR sky130_fd_sc_hd__or4_4
X_5889_ _5889_/A1 _8885_/X _8924_/X _9144_/Q VGND VPWR _9144_/D VGND VPWR sky130_fd_sc_hd__o22a_2
X_7628_ _6801_/Y _7400_/X _6927_/Y _7405_/X _7627_/X VGND VPWR _7644_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_193_397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7559_ _6246_/Y _7427_/X _6320_/Y _5699_/X VGND VPWR _7559_/X VGND VPWR sky130_fd_sc_hd__o22a_1
Xclkbuf_2_2_0_csclk clkbuf_2_3_0_csclk/A VGND VPWR clkbuf_2_2_0_csclk/X VGND VPWR
+ sky130_fd_sc_hd__clkbuf_2
X_9229_ _9440_/CLK _9229_/D _9685_/SET_B VGND VPWR _9229_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_96_25 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_76 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_98 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_540 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_470 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_114 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_484 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_351 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_340 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_384 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_362 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_23 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_5 _7155_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_112_114 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_359 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6930_ _6928_/Y _5671_/B _6929_/Y _5960_/B VGND VPWR _6930_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_6861_ _9741_/Q VGND VPWR _6861_/Y VGND VPWR sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_6_csclk clkbuf_leaf_6_csclk/A VGND VPWR _9440_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_34_131 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5812_ _5812_/A VGND VPWR _5812_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_6792_ _6787_/Y _5355_/B _6788_/Y _5267_/B _6791_/X VGND VPWR _6830_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9580_ _9620_/CLK _9580_/D _9633_/SET_B VGND VPWR _9580_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_8600_ _8600_/A _8600_/B VGND VPWR _8662_/C VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_179_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_8531_ _8607_/A _8531_/B _8734_/D _8614_/D VGND VPWR _8535_/A VGND VPWR sky130_fd_sc_hd__or4_1
Xclkbuf_1_0_0_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/X VGND VPWR clkbuf_1_0_1_mgmt_gpio_in[4]/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_2
X_5743_ _5743_/A VGND VPWR _5744_/A VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_22_348 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_320 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5674_ _9268_/Q _5673_/A _8843_/X _5673_/Y VGND VPWR _9268_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8462_ _7836_/B _8299_/B _7862_/Y _8544_/A _7987_/Y VGND VPWR _8668_/A VGND VPWR
+ sky130_fd_sc_hd__a32o_1
XFILLER_148_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8393_ _8393_/A VGND VPWR _8393_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7413_ _7413_/A _9253_/Q VGND VPWR _7474_/C VGND VPWR sky130_fd_sc_hd__or2_4
X_4625_ _4625_/A VGND VPWR _9720_/D VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_7344_ _6632_/Y _7112_/X _6750_/Y _7077_/B VGND VPWR _7344_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4556_ _4556_/A VGND VPWR _9758_/D VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_143_250 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_592 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7275_ _6126_/Y _7068_/A _6083_/Y _7105_/X VGND VPWR _7275_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4487_ _4661_/C _8938_/X _4801_/C VGND VPWR _4488_/A VGND VPWR sky130_fd_sc_hd__or3_1
X_9014_ _9027_/CLK _9014_/D VGND VPWR _9014_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_6226_ _9768_/Q VGND VPWR _6226_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_103_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6157_ _9652_/Q VGND VPWR _6157_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_106_79 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5108_ _9061_/Q _9062_/Q _9063_/Q _9065_/D VGND VPWR _5108_/X VGND VPWR sky130_fd_sc_hd__or4_2
X_6088_ _6085_/Y _6086_/X _6087_/Y _4870_/X VGND VPWR _6088_/X VGND VPWR sky130_fd_sc_hd__o22a_1
Xrepeater361 _8842_/X VGND VPWR _5964_/B1 VGND VPWR sky130_fd_sc_hd__buf_12
Xrepeater372 _9647_/SET_B VGND VPWR _9528_/SET_B VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_38_492 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5039_ _8974_/X _4551_/B _9680_/Q _5062_/D VGND VPWR _9680_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_13_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9778_ _9785_/CLK _9778_/D _9779_/SET_B VGND VPWR _9778_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_15_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_8729_ _8729_/A VGND VPWR _8729_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_31_42 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_31 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_86 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_442 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_230 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput120 sram_ro_data[5] VGND VPWR _6270_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_102_180 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput142 wb_adr_i[1] VGND VPWR _8394_/C VGND VPWR sky130_fd_sc_hd__buf_4
Xinput153 wb_adr_i[2] VGND VPWR _8379_/B VGND VPWR sky130_fd_sc_hd__buf_4
Xinput131 wb_adr_i[0] VGND VPWR _7839_/A VGND VPWR sky130_fd_sc_hd__clkbuf_4
Xinput164 wb_dat_i[0] VGND VPWR _8961_/A1 VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput175 wb_dat_i[1] VGND VPWR _8962_/A1 VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput186 wb_dat_i[2] VGND VPWR _8963_/A1 VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput197 wb_sel_i[0] VGND VPWR _5059_/B VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_44_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_607 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_170 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_192 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5390_ _9452_/Q _5384_/A _8841_/X _5384_/Y VGND VPWR _9452_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_172_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7060_ _7104_/A _7127_/B _7073_/C VGND VPWR _7061_/A VGND VPWR sky130_fd_sc_hd__or3_1
X_6011_ _9084_/Q _5995_/A _8899_/X _5995_/Y VGND VPWR _9084_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_39_234 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_212 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_267 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7962_ _8528_/A _7960_/Y _8193_/A _8193_/B VGND VPWR _7994_/B VGND VPWR sky130_fd_sc_hd__o22a_1
X_9701_ _4446_/A1 _9701_/D _4984_/X VGND VPWR _9701_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6913_ _9094_/Q VGND VPWR _6913_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_7893_ _8077_/A _8232_/B _8441_/A _7892_/X VGND VPWR _7893_/X VGND VPWR sky130_fd_sc_hd__o211a_1
X_9632_ _9639_/CLK _9632_/D _9633_/SET_B VGND VPWR _9632_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_22_123 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6844_ _9779_/Q VGND VPWR _6844_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_22_156 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9563_ _9617_/CLK _9563_/D _9295_/SET_B VGND VPWR _9563_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6775_ _9108_/Q VGND VPWR _6775_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
XFILLER_50_465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_8514_ _8514_/A _8514_/B _8514_/C VGND VPWR _8605_/B VGND VPWR sky130_fd_sc_hd__or3_1
X_9494_ _9534_/CLK _9494_/D _9647_/SET_B VGND VPWR _9494_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_5726_ _5726_/A VGND VPWR _7127_/C VGND VPWR sky130_fd_sc_hd__buf_4
X_8445_ _8272_/A _8521_/B _8164_/A _8525_/C _8085_/A VGND VPWR _8445_/X VGND VPWR
+ sky130_fd_sc_hd__a311o_1
XFILLER_148_386 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5657_ _9054_/Q _9056_/Q _5724_/B _5647_/X _5656_/Y VGND VPWR _9278_/D VGND VPWR
+ sky130_fd_sc_hd__o311a_2
XFILLER_2_506 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5588_ _9317_/Q _5585_/A _8844_/X _5585_/Y VGND VPWR _9317_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_4608_ _9728_/Q _4604_/A _5965_/B1 _4604_/Y VGND VPWR _9728_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8376_ _8376_/A _8539_/A VGND VPWR _8380_/B VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_190_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_412 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7327_ _6856_/Y _5728_/X _6902_/Y _7040_/A _7326_/X VGND VPWR _7330_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_2
X_4539_ _4539_/A VGND VPWR _9761_/D VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_7258_ _6171_/Y _7118_/X _6205_/Y _7048_/C VGND VPWR _7258_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_131_275 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6209_ _6207_/Y _4822_/X _6208_/Y _4907_/X VGND VPWR _6209_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_7189_ _7189_/A _7189_/B _7189_/C _7189_/D VGND VPWR _7199_/B VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_93_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_203 input83/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_214 _6677_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_186_404 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_73 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_415 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_448 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_583 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_82 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_61 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_215 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_94 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_440 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4890_ _9406_/Q VGND VPWR _4890_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_32_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6560_ _6555_/Y _5518_/B _6556_/Y _5404_/B _6559_/X VGND VPWR _6567_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_5511_ _9370_/Q _5509_/A _8845_/X _5509_/Y VGND VPWR _9370_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_6491_ _9341_/Q VGND VPWR _6491_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_118_537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8230_ _8230_/A _8260_/B VGND VPWR _8573_/B VGND VPWR sky130_fd_sc_hd__nor2_1
X_5442_ _5671_/A _5442_/B VGND VPWR _5443_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_5373_ _9463_/Q _5368_/A _5967_/B1 _5368_/Y VGND VPWR _9463_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8161_ _8554_/A _8378_/B VGND VPWR _8370_/A VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_172_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_540 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8092_ _8093_/B VGND VPWR _8092_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7112_ _7112_/A VGND VPWR _7112_/X VGND VPWR sky130_fd_sc_hd__buf_8
Xclkbuf_leaf_24_csclk clkbuf_2_3_0_csclk/X VGND VPWR _9788_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_141_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_264 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7043_ _7043_/A VGND VPWR _7048_/B VGND VPWR sky130_fd_sc_hd__buf_8
XFILLER_67_351 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_39_csclk clkbuf_2_1_0_csclk/X VGND VPWR _9655_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_82_332 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_546 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8994_ _9562_/Q _8765_/A VGND VPWR mgmt_gpio_out[17] VGND VPWR sky130_fd_sc_hd__ebufn_8
XFILLER_63_18 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7945_ _8077_/A _8188_/B _9068_/Q VGND VPWR _8514_/B VGND VPWR sky130_fd_sc_hd__o21ai_1
X_7876_ _8226_/C _8230_/A VGND VPWR _8232_/B VGND VPWR sky130_fd_sc_hd__or2_2
X_6827_ _6825_/Y _5317_/B _6826_/Y _5412_/B VGND VPWR _6827_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_9615_ _9788_/CLK _9615_/D _9646_/SET_B VGND VPWR _9615_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_50_273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9546_ _9757_/CLK _9546_/D _9757_/SET_B VGND VPWR _9546_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_137_7 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6758_ _6753_/Y _6081_/B _6754_/Y _5905_/B _6757_/X VGND VPWR _6759_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_12_44 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9477_ _9527_/CLK _9477_/D _9685_/SET_B VGND VPWR _9477_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_5709_ _7476_/A _7401_/B VGND VPWR _7472_/A VGND VPWR sky130_fd_sc_hd__or2_4
X_6689_ _6685_/Y _5024_/B _6686_/Y _5507_/B _6688_/X VGND VPWR _6690_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_8428_ _8687_/B _8428_/B VGND VPWR _8430_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_124_518 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8359_ _8359_/A _8359_/B VGND VPWR _8574_/C VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_151_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_540 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_332 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_579 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_432 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_95 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_343 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5991_ _5991_/A VGND VPWR _5991_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_17_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7730_ _7727_/Y _7726_/Y _9700_/Q _7729_/Y VGND VPWR _7730_/Y VGND VPWR sky130_fd_sc_hd__a31oi_1
X_5848__7 _8924_/X VGND VPWR _5892_/A1 VGND VPWR sky130_fd_sc_hd__inv_4
X_4942_ _9090_/Q VGND VPWR _6022_/C VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_17_270 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7661_ _7661_/A _7661_/B _7661_/C _7661_/D VGND VPWR _7662_/D VGND VPWR sky130_fd_sc_hd__and4_2
XFILLER_60_582 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4873_ _4865_/Y _5336_/B _4867_/Y _4868_/X _4872_/X VGND VPWR _4896_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9400_ _9758_/CLK _9400_/D _9633_/SET_B VGND VPWR _9400_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6612_ _9414_/Q VGND VPWR _6612_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_32_295 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7592_ _6091_/Y _7400_/X _6139_/Y _7405_/X _7591_/X VGND VPWR _7608_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9331_ _9771_/CLK _9331_/D _4628_/A VGND VPWR _9331_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6543_ _9461_/Q VGND VPWR _6543_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
X_6474_ _6474_/A _6474_/B _6474_/C _6474_/D VGND VPWR _6475_/D VGND VPWR sky130_fd_sc_hd__and4_1
X_9262_ _9601_/CLK _9262_/D _9295_/SET_B VGND VPWR _9262_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_5425_ _9429_/Q _5422_/A _8844_/X _5422_/Y VGND VPWR _9429_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8213_ _8213_/A _8213_/B VGND VPWR _8311_/B VGND VPWR sky130_fd_sc_hd__or2_1
Xoutput210 _8756_/X VGND VPWR mgmt_gpio_oeb[12] VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_133_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9193_ _9378_/CLK _9193_/D _9646_/SET_B VGND VPWR _9193_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
Xoutput243 _8748_/X VGND VPWR mgmt_gpio_oeb[8] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput221 _8776_/X VGND VPWR mgmt_gpio_oeb[22] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput232 _8796_/X VGND VPWR mgmt_gpio_oeb[32] VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_58_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_8144_ _8144_/A _8362_/A _8575_/A _8627_/B VGND VPWR _8144_/X VGND VPWR sky130_fd_sc_hd__or4_1
Xoutput254 _8838_/X VGND VPWR pad_flash_io0_do VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput265 _9721_/Q VGND VPWR pll_div[0] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput276 _9743_/Q VGND VPWR pll_trim[11] VGND VPWR sky130_fd_sc_hd__buf_2
X_5356_ _5356_/A VGND VPWR _5357_/A VGND VPWR sky130_fd_sc_hd__clkbuf_4
X_5287_ _9521_/Q _5280_/A _8840_/X _5280_/Y VGND VPWR _9521_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8075_ _8585_/B _8075_/B VGND VPWR _8075_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
Xoutput298 _9740_/Q VGND VPWR pll_trim[8] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput287 _9753_/Q VGND VPWR pll_trim[21] VGND VPWR sky130_fd_sc_hd__buf_2
X_7026_ _9250_/Q _9249_/Q VGND VPWR _7027_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_101_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_302 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8977_ _8930_/S _6322_/Y _8977_/S VGND VPWR _8977_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_82_173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_218 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7928_ _8325_/A _7928_/B VGND VPWR _7929_/B VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_11_413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7859_ _8521_/B _8262_/B VGND VPWR _8463_/A VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_109_323 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_87 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_470 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9529_ _9534_/CLK _9529_/D _9647_/SET_B VGND VPWR _9529_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_7_439 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_495 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_402 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_554 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_118 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_354 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_256 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_304 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5210_ _9571_/Q _5203_/Y _8930_/X _5203_/A VGND VPWR _9571_/D VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_43_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6190_ _9422_/Q VGND VPWR _6190_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_170_498 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5141_ _9621_/Q _5136_/A _8929_/A1 _5136_/Y VGND VPWR _9621_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_111_543 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_243 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5072_ _8964_/X _9662_/Q _5078_/S VGND VPWR _5073_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_8900_ _7710_/X _9082_/Q _9051_/Q VGND VPWR _8900_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_25_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8831_ _6544_/Y input2/X input1/X VGND VPWR _8831_/X VGND VPWR sky130_fd_sc_hd__mux2_2
X_8762_ _8762_/A VGND VPWR _8762_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_5974_ _9097_/Q _5970_/A _8925_/A1 _5970_/Y VGND VPWR _9097_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7713_ _9084_/Q _7713_/B _9085_/Q VGND VPWR _7716_/B VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_33_571 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_8693_ _8693_/A _8693_/B _8693_/C _7929_/A VGND VPWR _8696_/B VGND VPWR sky130_fd_sc_hd__or4b_1
X_4925_ _4925_/A _4931_/B VGND VPWR _5366_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_20_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4856_ _4911_/A _4917_/A VGND VPWR _5317_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_7644_ _7644_/A _7644_/B _7644_/C _7644_/D VGND VPWR _7644_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
XFILLER_165_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7575_ _6232_/Y _7419_/X _6189_/Y _7421_/X VGND VPWR _7575_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4787_ _4787_/A _4921_/A VGND VPWR _5488_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_6526_ _6526_/A _6526_/B _6526_/C _6526_/D VGND VPWR _6629_/B VGND VPWR sky130_fd_sc_hd__and4_1
X_9314_ _9534_/CLK _9314_/D _9647_/SET_B VGND VPWR _9314_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_118_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6457_ _9181_/Q VGND VPWR _6457_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_173_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9245_ _9278_/CLK _9245_/D _9633_/SET_B VGND VPWR _9245_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
X_6388_ _6386_/Y _6086_/X _6387_/Y _5336_/B VGND VPWR _6388_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_5408_ _9440_/Q _5406_/A _5964_/B1 _5406_/Y VGND VPWR _9440_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_9176_ _9280_/CLK _9176_/D _9757_/SET_B VGND VPWR _9176_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_102_510 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_12 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_210 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5339_ _9488_/Q _5338_/A _5963_/B1 _5338_/Y VGND VPWR _9488_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8127_ _8354_/A _8127_/B _8571_/A _8683_/B VGND VPWR _8131_/A VGND VPWR sky130_fd_sc_hd__or4_1
XFILLER_125_45 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_89 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_427 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8058_ _8521_/B VGND VPWR _8061_/A VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_75_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_7009_ _9051_/Q _5993_/B _9050_/Q _7008_/X VGND VPWR _9050_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_47_129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_184 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_258 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_112 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_464 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_332 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_268 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4710_ _9281_/Q VGND VPWR _7304_/A VGND VPWR sky130_fd_sc_hd__inv_2
X_5690_ _9053_/Q VGND VPWR _5691_/A VGND VPWR sky130_fd_sc_hd__inv_2
X_4641_ _4994_/A VGND VPWR _4642_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_175_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_4572_ _9750_/Q _4566_/A _5965_/B1 _4566_/Y VGND VPWR _9750_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7360_ _6589_/Y _7095_/X _6477_/Y _7068_/D _7359_/X VGND VPWR _7365_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_6311_ _9317_/Q VGND VPWR _6311_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_155_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7291_ _4677_/Y _7040_/C _4775_/Y _7059_/C VGND VPWR _7291_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_6242_ _6240_/Y _5306_/B _6241_/Y _4491_/B VGND VPWR _6242_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_9030_ _9039_/CLK _9030_/D VGND VPWR _9030_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_130_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_232 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6173_ _6168_/Y _5278_/B _6169_/Y _5306_/B _6172_/X VGND VPWR _6174_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_69_276 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_574 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5124_ _9631_/Q _5123_/A _5963_/B1 _5123_/Y VGND VPWR _9631_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_57_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_246 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5055_ _9667_/Q _5047_/A _8916_/A1 _5047_/Y VGND VPWR _9667_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8814_ _9791_/Q _6251_/Y _8916_/A1 _6251_/A _8939_/X VGND VPWR _9791_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_71_18 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5957_ _9108_/Q _5951_/A _8955_/A1 _5951_/Y VGND VPWR _9108_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8745_ _8745_/A VGND VPWR _8746_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_4908_ _9740_/Q VGND VPWR _4908_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_8676_ _8676_/A _8676_/B VGND VPWR _8677_/B VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_166_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7627_ _6866_/Y _7408_/X _6902_/Y _7410_/X VGND VPWR _7627_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_5888_ _5849_/X _8887_/X _8924_/X _9145_/Q VGND VPWR _9145_/D VGND VPWR sky130_fd_sc_hd__o22a_2
XFILLER_21_552 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4839_ _4831_/Y _4832_/X _4833_/Y _5431_/B _4838_/X VGND VPWR _4864_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_119_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_602 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_218 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_579 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7558_ _6301_/Y _7415_/X _6297_/Y _7417_/X _7557_/X VGND VPWR _7572_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_134_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7489_ _6799_/Y _7430_/X _6860_/Y _7432_/X _7488_/X VGND VPWR _7489_/X VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_6509_ _9323_/Q VGND VPWR _8763_/A VGND VPWR sky130_fd_sc_hd__clkinv_8
X_9228_ _9440_/CLK _9228_/D _9685_/SET_B VGND VPWR _9228_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_121_148 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9159_ _9358_/CLK _9159_/D _9528_/SET_B VGND VPWR _9159_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_0_456 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_30 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_324 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_352 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_330 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_374 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_363 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_524 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_91 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_9 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_6 _7155_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_98_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_126 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_170 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6860_ _9547_/Q VGND VPWR _6860_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_34_110 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6791_ _6789_/Y _4602_/B _6790_/Y _4524_/B VGND VPWR _6791_/X VGND VPWR sky130_fd_sc_hd__o22a_4
X_5811_ _5811_/A VGND VPWR _5812_/A VGND VPWR sky130_fd_sc_hd__clkbuf_2
X_8530_ _8472_/Y _8528_/Y _8518_/X _8459_/C VGND VPWR _8614_/D VGND VPWR sky130_fd_sc_hd__a31o_1
X_5742_ _5960_/A _5742_/B VGND VPWR _5743_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_175_332 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5673_ _5673_/A VGND VPWR _5673_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_8461_ _8461_/A _8627_/A VGND VPWR _8464_/B VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_163_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8392_ _8392_/A VGND VPWR _8708_/A VGND VPWR sky130_fd_sc_hd__inv_2
X_7412_ _4877_/Y _7400_/X _4720_/Y _7405_/X _7411_/X VGND VPWR _7481_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_4624_ _5966_/B1 _9720_/Q _4626_/S VGND VPWR _4625_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_116_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_410 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7343_ _7343_/A _7343_/B _7343_/C _7343_/D VGND VPWR _7353_/B VGND VPWR sky130_fd_sc_hd__and4_1
X_4555_ _5967_/B1 _9758_/Q _4555_/S VGND VPWR _4556_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_9013_ _9039_/CLK _9013_/D VGND VPWR _9013_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_7274_ _6067_/Y _7059_/B _6081_/A _7068_/C _7273_/X VGND VPWR _7277_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_4486_ _4486_/A VGND VPWR _9786_/D VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_6225_ _9430_/Q VGND VPWR _6225_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_6156_ _6151_/Y _5545_/B _6152_/Y _5496_/B _6155_/X VGND VPWR _6174_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_66_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5107_ _9641_/Q _5102_/A _5967_/B1 _5102_/Y VGND VPWR _9641_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_6087_ _6087_/A VGND VPWR _6087_/Y VGND VPWR sky130_fd_sc_hd__inv_2
Xrepeater362 _8842_/X VGND VPWR _8929_/A1 VGND VPWR sky130_fd_sc_hd__buf_12
X_5038_ _8975_/X _4551_/B _9681_/Q _5062_/D VGND VPWR _9681_/D VGND VPWR sky130_fd_sc_hd__a22o_1
Xrepeater373 _9685_/SET_B VGND VPWR _9647_/SET_B VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_167_7 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_9777_ _9777_/CLK _9777_/D _7011_/B VGND VPWR _9777_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_13_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6989_ _8813_/A _8809_/A _6950_/B VGND VPWR _9068_/D VGND VPWR sky130_fd_sc_hd__o21ai_1
X_8728_ _8728_/A VGND VPWR _8728_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_8659_ _8659_/A _8659_/B _8659_/C _7893_/X VGND VPWR _8727_/C VGND VPWR sky130_fd_sc_hd__or4b_1
XFILLER_166_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_218 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_98 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_360 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xinput110 sram_ro_data[25] VGND VPWR _6817_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_76_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput143 wb_adr_i[20] VGND VPWR _7837_/B VGND VPWR sky130_fd_sc_hd__buf_2
Xinput121 sram_ro_data[6] VGND VPWR _6233_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput132 wb_adr_i[10] VGND VPWR _7771_/B VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput154 wb_adr_i[30] VGND VPWR _5931_/B VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_102_192 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xinput165 wb_dat_i[10] VGND VPWR _7741_/B2 VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput176 wb_dat_i[20] VGND VPWR _7744_/B VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput187 wb_dat_i[30] VGND VPWR _7749_/A2 VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput198 wb_sel_i[1] VGND VPWR _5058_/B VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_63_216 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_146 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_160 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_94 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_402 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6010_ _6010_/A VGND VPWR _6010_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_79_371 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_490 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7961_ _7959_/A _8195_/B _7960_/Y VGND VPWR _7979_/A VGND VPWR sky130_fd_sc_hd__a21oi_1
X_7892_ _8515_/B _8305_/A _8496_/A _8305_/B VGND VPWR _7892_/X VGND VPWR sky130_fd_sc_hd__a211o_1
X_6912_ _6908_/Y _5089_/B _6909_/Y _5864_/B _6911_/X VGND VPWR _6925_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9700_ _9709_/CLK _9700_/D _4987_/X VGND VPWR _9700_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_9631_ _9757_/CLK _9631_/D _9757_/SET_B VGND VPWR _9631_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6843_ _9490_/Q VGND VPWR _6843_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_22_135 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6774_ _9629_/Q VGND VPWR _6774_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9562_ _9617_/CLK _9562_/D _9295_/SET_B VGND VPWR _9562_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_9493_ _9493_/CLK _9493_/D _4628_/A VGND VPWR _9493_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_5725_ _9250_/Q _5725_/B VGND VPWR _5726_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_8513_ _8513_/A VGND VPWR _8513_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_50_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_600 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5656_ _5647_/A _5651_/A _5751_/C VGND VPWR _5656_/Y VGND VPWR sky130_fd_sc_hd__o21ai_2
X_8444_ _8444_/A _8444_/B VGND VPWR _8448_/B VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_148_398 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4607_ _9729_/Q _4604_/A _5964_/B1 _4604_/Y VGND VPWR _9729_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_5587_ _9318_/Q _5585_/A _8845_/X _5585_/Y VGND VPWR _9318_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8375_ _8375_/A _8582_/A _8678_/A _8646_/A VGND VPWR _8380_/A VGND VPWR sky130_fd_sc_hd__or4_1
XFILLER_116_273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4538_ _5967_/B1 _9761_/Q _4540_/S VGND VPWR _4539_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_7326_ _7326_/A _7392_/B VGND VPWR _7326_/X VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_117_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4469_ _4456_/Y _8942_/X _8941_/X VGND VPWR _4801_/C VGND VPWR sky130_fd_sc_hd__a21bo_1
X_7257_ _6194_/Y _7040_/D _6154_/Y _7110_/X _7256_/X VGND VPWR _7264_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_104_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6208_ _6208_/A VGND VPWR _6208_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7188_ _8751_/A _7048_/D _6517_/Y _7040_/B _7187_/X VGND VPWR _7189_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_6139_ _9263_/Q VGND VPWR _6139_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_93_38 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_204 input83/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_215 _6679_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_41_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_416 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_64 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_5_csclk clkbuf_2_2_0_csclk/X VGND VPWR _9789_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_49_500 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_574 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_595 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_73 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_536 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5510_ _9371_/Q _5509_/A _8846_/X _5509_/Y VGND VPWR _9371_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_145_313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_172 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6490_ _9096_/Q VGND VPWR _7705_/A VGND VPWR sky130_fd_sc_hd__inv_6
X_5441_ _9416_/Q _5433_/A _8916_/A1 _5433_/Y VGND VPWR _9416_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_172_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5372_ _9464_/Q _5368_/A _5966_/B1 _5368_/Y VGND VPWR _9464_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8160_ _8160_/A _8645_/A VGND VPWR _8162_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_99_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8091_ _8525_/A _8091_/B _8386_/A VGND VPWR _8093_/B VGND VPWR sky130_fd_sc_hd__or3_1
X_7111_ _9246_/Q _9245_/Q _7111_/C _7127_/C VGND VPWR _7112_/A VGND VPWR sky130_fd_sc_hd__or4_2
XFILLER_87_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_552 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_308 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7042_ _7127_/A _7127_/B _7073_/C VGND VPWR _7043_/A VGND VPWR sky130_fd_sc_hd__or3_1
XFILLER_101_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_363 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8993_ _9561_/Q _8763_/A VGND VPWR mgmt_gpio_out[16] VGND VPWR sky130_fd_sc_hd__ebufn_8
XFILLER_82_344 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7944_ _7944_/A VGND VPWR _7944_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_70_528 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_19 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7875_ _8525_/A _7894_/B _7903_/C _8193_/A VGND VPWR _8230_/A VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_23_444 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6826_ _9433_/Q VGND VPWR _6826_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9614_ _9788_/CLK _9614_/D _9295_/SET_B VGND VPWR _9614_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6757_ _6755_/Y _5872_/B _6756_/Y _5526_/B VGND VPWR _6757_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_9545_ _9545_/CLK _9545_/D _4628_/A VGND VPWR _9545_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_11_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5708_ _9251_/Q VGND VPWR _7401_/B VGND VPWR sky130_fd_sc_hd__inv_2
X_9476_ _9527_/CLK _9476_/D _9685_/SET_B VGND VPWR _9476_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6688_ input45/X _8926_/S _6687_/Y _5837_/B VGND VPWR _6688_/X VGND VPWR sky130_fd_sc_hd__o2bb2a_1
XFILLER_12_56 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5639_ _9281_/Q _5634_/A _8839_/X _5634_/Y VGND VPWR _9281_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8427_ _8427_/A _8601_/D VGND VPWR _8428_/B VGND VPWR sky130_fd_sc_hd__or2_1
X_8358_ _8358_/A _8358_/B VGND VPWR _8642_/C VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_2_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7309_ _7309_/A _7309_/B _7309_/C VGND VPWR _7309_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
XFILLER_132_552 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_11 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_8289_ _8625_/A _8340_/B _8340_/C _8288_/X VGND VPWR _8290_/B VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_132_596 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_63 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_63 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_466 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_460 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5990_ _6040_/A VGND VPWR _5991_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_91_196 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4941_ _9091_/Q VGND VPWR _6022_/D VGND VPWR sky130_fd_sc_hd__inv_2
X_5848__8 _8924_/X VGND VPWR _5891_/A1 VGND VPWR sky130_fd_sc_hd__inv_4
XFILLER_17_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7660_ _6750_/Y _7471_/X _7348_/A _7473_/X _7659_/X VGND VPWR _7661_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_4872_ _4869_/Y _4870_/X _4871_/Y _4558_/B VGND VPWR _4872_/X VGND VPWR sky130_fd_sc_hd__o22a_2
X_6611_ _9427_/Q VGND VPWR _8771_/A VGND VPWR sky130_fd_sc_hd__inv_6
XFILLER_20_436 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7591_ _6078_/Y _7408_/X _6059_/Y _7410_/X VGND VPWR _7591_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_9330_ _9776_/CLK _9330_/D _4628_/A VGND VPWR _9330_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6542_ _8799_/A _5507_/B _6530_/X _6536_/X _6541_/X VGND VPWR _6629_/C VGND VPWR
+ sky130_fd_sc_hd__o2111a_1
XFILLER_145_143 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6473_ _6473_/A _6473_/B _6473_/C _6473_/D VGND VPWR _6474_/D VGND VPWR sky130_fd_sc_hd__and4_1
X_9261_ _9601_/CLK _9261_/D _9295_/SET_B VGND VPWR _9261_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_5424_ _9430_/Q _5422_/A _8845_/X _5422_/Y VGND VPWR _9430_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8212_ _8341_/B _8260_/B _8312_/D VGND VPWR _8224_/B VGND VPWR sky130_fd_sc_hd__o21ai_1
X_9192_ _9378_/CLK _9192_/D _9646_/SET_B VGND VPWR _9192_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_133_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8143_ _8164_/A _8551_/A VGND VPWR _8627_/B VGND VPWR sky130_fd_sc_hd__nor2_1
Xoutput244 _8750_/X VGND VPWR mgmt_gpio_oeb[9] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput211 _8758_/X VGND VPWR mgmt_gpio_oeb[13] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput222 _8778_/X VGND VPWR mgmt_gpio_oeb[23] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput233 _8798_/X VGND VPWR mgmt_gpio_oeb[33] VGND VPWR sky130_fd_sc_hd__buf_2
X_5355_ _5545_/A _5355_/B VGND VPWR _5356_/A VGND VPWR sky130_fd_sc_hd__or2_1
Xoutput255 _7014_/A VGND VPWR pad_flash_io0_ieb VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput266 _9722_/Q VGND VPWR pll_div[1] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput277 _9744_/Q VGND VPWR pll_trim[12] VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_114_596 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5286_ _9522_/Q _5280_/A _8955_/A1 _5280_/Y VGND VPWR _9522_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8074_ _8074_/A _8704_/A VGND VPWR _8075_/B VGND VPWR sky130_fd_sc_hd__or2_1
Xoutput299 _9741_/Q VGND VPWR pll_trim[9] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput288 _9754_/Q VGND VPWR pll_trim[22] VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_141_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7025_ _7025_/A VGND VPWR _7079_/B VGND VPWR sky130_fd_sc_hd__buf_8
XFILLER_74_119 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_620 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_322 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8976_ _8926_/S _6322_/Y _8977_/S VGND VPWR _8976_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_7927_ _8615_/A _7927_/B VGND VPWR _7928_/B VGND VPWR sky130_fd_sc_hd__nor2_1
X_7858_ _7858_/A VGND VPWR _8262_/B VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_23_11 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_274 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6809_ _6807_/Y _4481_/B _6808_/Y _4893_/X VGND VPWR _6809_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_11_425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7789_ _7903_/C _7823_/A _8528_/A _8193_/A _7787_/X VGND VPWR _7900_/A VGND VPWR
+ sky130_fd_sc_hd__a32o_1
XFILLER_139_33 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9528_ _9535_/CLK _9528_/D _9528_/SET_B VGND VPWR _9528_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_136_110 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9459_ _9532_/CLK _9459_/D _9647_/SET_B VGND VPWR _9459_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_151_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_31 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_73 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_23_csclk clkbuf_2_3_0_csclk/X VGND VPWR _9617_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_9_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_38_csclk clkbuf_2_1_0_csclk/X VGND VPWR _9757_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_6_451 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5140_ _9622_/Q _5136_/A _8925_/A1 _5136_/Y VGND VPWR _9622_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_123_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_555 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5071_ _5071_/A VGND VPWR _9663_/D VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_84_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8830_ _9593_/Q input91/X _8835_/S VGND VPWR _8830_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_52_303 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5973_ _9098_/Q _5970_/A _8844_/X _5970_/Y VGND VPWR _9098_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8761_ _8761_/A VGND VPWR _8762_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_7712_ _9084_/Q _7713_/B _9084_/Q _7713_/B VGND VPWR _7712_/X VGND VPWR sky130_fd_sc_hd__o2bb2a_1
X_4924_ _9463_/Q VGND VPWR _4924_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_33_550 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_8692_ _8671_/Y _8673_/X _8680_/Y _8682_/X _8691_/Y VGND VPWR _8692_/Y VGND VPWR
+ sky130_fd_sc_hd__o221ai_4
X_4855_ _9494_/Q VGND VPWR _4855_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7643_ _7643_/A _7643_/B _7643_/C _7643_/D VGND VPWR _7644_/D VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_20_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4786_ _9380_/Q VGND VPWR _4786_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7574_ _6152_/Y _7400_/X _6178_/Y _7405_/X _7573_/X VGND VPWR _7590_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_165_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9313_ _9534_/CLK _9313_/D _9647_/SET_B VGND VPWR _9313_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6525_ _8747_/A _5837_/B _6521_/Y _6135_/A _6524_/X VGND VPWR _6526_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_134_614 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_9244_ _9789_/CLK _9244_/D _9685_/SET_B VGND VPWR _9244_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_106_338 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6456_ _9110_/Q VGND VPWR _6456_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_5407_ _9441_/Q _5406_/A _5963_/B1 _5406_/Y VGND VPWR _9441_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_9175_ _9280_/CLK _9175_/D _9757_/SET_B VGND VPWR _9175_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6387_ _9488_/Q VGND VPWR _6387_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
XFILLER_87_200 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_24 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5338_ _5338_/A VGND VPWR _5338_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_8126_ _8164_/A _8130_/B VGND VPWR _8683_/B VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_102_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8057_ _8057_/A _8536_/A VGND VPWR _8062_/A VGND VPWR sky130_fd_sc_hd__nand2_1
X_7008_ _7008_/A _7008_/B VGND VPWR _7008_/X VGND VPWR sky130_fd_sc_hd__or2_1
X_5269_ _5269_/A VGND VPWR _5269_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_75_439 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_163 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_8959_ _7133_/X _4875_/Y _8959_/S VGND VPWR _8959_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_34_54 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_208 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_168 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_371 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_330 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_74 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_374 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_620 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4640_ _9717_/Q _4636_/A _8948_/X _4636_/Y VGND VPWR hold2/A VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_116_603 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4571_ _9751_/Q _4566_/A _5964_/B1 _4566_/Y VGND VPWR _9751_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_6310_ _9395_/Q VGND VPWR _6310_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_183_580 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7290_ _4888_/Y _7082_/X _4865_/Y _7084_/X _7289_/X VGND VPWR _7309_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_6241_ _9783_/Q VGND VPWR _6241_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_131_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6172_ _6170_/Y _5621_/B _6171_/Y _5267_/B VGND VPWR _6172_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_69_244 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5123_ _5123_/A VGND VPWR _5123_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_97_586 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_288 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5054_ _9668_/Q _5047_/A _8930_/A1 _5047_/Y VGND VPWR _9668_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_65_472 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_163 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_8813_ _8813_/A _8813_/B VGND VPWR _9060_/D VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_52_111 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5956_ _9109_/Q _5951_/A _8929_/A1 _5951_/Y VGND VPWR _9109_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8744_ _8744_/A VGND VPWR _8744_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_33_380 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_4907_ _6158_/A _6111_/B VGND VPWR _4907_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_8675_ _8675_/A _8675_/B _8675_/C _8675_/D VGND VPWR _8716_/D VGND VPWR sky130_fd_sc_hd__or4_4
X_5887_ _5849_/X _8889_/X _8924_/X _9146_/Q VGND VPWR _9146_/D VGND VPWR sky130_fd_sc_hd__o22a_2
XFILLER_178_385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4838_ _4835_/Y _4481_/B _4836_/Y _5232_/B VGND VPWR _4838_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_7626_ _7626_/A _7626_/B _7626_/C _7626_/D VGND VPWR _7626_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
X_4769_ _9646_/Q VGND VPWR _4769_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7557_ _6282_/Y _7419_/X _6241_/Y _7421_/X VGND VPWR _7557_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_119_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6508_ _9336_/Q VGND VPWR _6508_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7488_ _6788_/Y _7434_/X _6854_/Y _7436_/X VGND VPWR _7488_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_134_455 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9227_ _9440_/CLK _9227_/D _9685_/SET_B VGND VPWR _9227_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6439_ _9650_/Q VGND VPWR _6439_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
XFILLER_0_413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_263 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9158_ _9695_/CLK _9158_/D _9646_/SET_B VGND VPWR _9158_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_102_330 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_435 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_8109_ _8640_/A VGND VPWR _8110_/C VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_75_203 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9089_ _9089_/CLK _9089_/D _5991_/X VGND VPWR _9089_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_75_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_42 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_336 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_342 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_331 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_320 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_188 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_391 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_386 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_375 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_364 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_52 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_238 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_536 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_400 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_7 _7177_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_125_499 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_406 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_182 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_512 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_291 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6790_ _9763_/Q VGND VPWR _6790_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_5810_ _5960_/A _5810_/B VGND VPWR _5811_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_5741_ _9245_/Q _5713_/A _5738_/B _5724_/B VGND VPWR _9245_/D VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_34_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_188 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_8460_ _8460_/A VGND VPWR _8627_/A VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_30_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_7411_ _4897_/Y _7408_/X _4842_/Y _7410_/X VGND VPWR _7411_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_5672_ _5672_/A VGND VPWR _5673_/A VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_30_394 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4623_ _5259_/A _4623_/B VGND VPWR _4626_/S VGND VPWR sky130_fd_sc_hd__or2_1
X_8391_ _8544_/C VGND VPWR _8401_/B VGND VPWR sky130_fd_sc_hd__clkinv_4
X_4554_ _6158_/A _4925_/A _5259_/A VGND VPWR _4555_/S VGND VPWR sky130_fd_sc_hd__or3_1
X_7342_ _6646_/Y _7048_/D _6745_/Y _7040_/B _7341_/X VGND VPWR _7343_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_116_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7273_ _6103_/Y _7079_/B _6066_/Y _7059_/A VGND VPWR _7273_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_116_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_9012_ _9027_/CLK _9012_/D VGND VPWR _9012_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_4485_ _8840_/X _9786_/Q _6018_/S VGND VPWR _4486_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_6224_ _9131_/Q VGND VPWR _6224_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_131_458 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6155_ _6153_/Y _4870_/X _6154_/Y _5534_/B VGND VPWR _6155_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_85_512 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5106_ _9642_/Q _5102_/A _5966_/B1 _5102_/Y VGND VPWR _9642_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_6086_ _6158_/A _6086_/B VGND VPWR _6086_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_85_578 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5037_ _9049_/Q _5034_/Y _5985_/B _9682_/Q VGND VPWR _9682_/D VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_122_47 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xrepeater374 _4628_/A VGND VPWR _9685_/SET_B VGND VPWR sky130_fd_sc_hd__buf_12
Xrepeater363 _8841_/X VGND VPWR _5965_/B1 VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_82_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9776_ _9776_/CLK _9776_/D _7011_/B VGND VPWR _9776_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_8727_ _8727_/A _8727_/B _8727_/C _8727_/D VGND VPWR _8728_/A VGND VPWR sky130_fd_sc_hd__or4_1
X_6988_ _8812_/A _8809_/A _6962_/B VGND VPWR _9067_/D VGND VPWR sky130_fd_sc_hd__o21ai_1
X_5939_ _5939_/A _5939_/B VGND VPWR _5939_/X VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_21_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_8658_ _8676_/B _8658_/B VGND VPWR _8659_/B VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_154_506 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7609_ _4924_/Y _7408_/X _4692_/A _7410_/X VGND VPWR _7609_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_8589_ _8650_/B _8650_/C _8651_/B _8588_/X VGND VPWR _8589_/X VGND VPWR sky130_fd_sc_hd__or4b_2
XFILLER_134_230 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_350 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xinput100 sram_ro_data[16] VGND VPWR _4840_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput111 sram_ro_data[26] VGND VPWR _6669_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_0_287 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_372 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput144 wb_adr_i[21] VGND VPWR _7832_/A VGND VPWR sky130_fd_sc_hd__buf_2
Xinput122 sram_ro_data[7] VGND VPWR _6075_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput133 wb_adr_i[11] VGND VPWR _7771_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_76_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput155 wb_adr_i[31] VGND VPWR _5931_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput166 wb_dat_i[11] VGND VPWR _7743_/B2 VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput177 wb_dat_i[21] VGND VPWR _7746_/B VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_76_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput199 wb_sel_i[2] VGND VPWR _7733_/A VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
Xinput188 wb_dat_i[31] VGND VPWR _7751_/A2 VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_56_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_80 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_150 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_119 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_194 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_183 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_172 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_182 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_73 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_354 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_6 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_119 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_108 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_383 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7960_ _8193_/B VGND VPWR _7960_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_94_397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6911_ input62/X _4680_/Y _6910_/Y _5045_/B VGND VPWR _6911_/X VGND VPWR sky130_fd_sc_hd__o2bb2a_1
X_7891_ _7896_/A _8305_/B VGND VPWR _8441_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_9630_ _9639_/CLK _9630_/D _9757_/SET_B VGND VPWR _9630_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6842_ _6837_/Y _5121_/B _6838_/Y _5110_/B _6841_/X VGND VPWR _6878_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_50_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_412 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6773_ _9648_/Q VGND VPWR _6773_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9561_ _9788_/CLK _9561_/D _9295_/SET_B VGND VPWR _9561_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_10_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8512_ _8603_/A _8512_/B _8603_/C _8512_/D VGND VPWR _8513_/A VGND VPWR sky130_fd_sc_hd__or4_1
X_5724_ _5725_/B _5724_/B _7041_/A VGND VPWR _5724_/Y VGND VPWR sky130_fd_sc_hd__nor3_1
X_9492_ _9545_/CLK _9492_/D _4628_/A VGND VPWR _9492_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_8443_ _7902_/B _8624_/B _7896_/X VGND VPWR _8444_/B VGND VPWR sky130_fd_sc_hd__o21ai_1
X_5655_ _5649_/B _5647_/X _5651_/A _5654_/X VGND VPWR _9279_/D VGND VPWR sky130_fd_sc_hd__o2bb2a_2
X_4606_ _9730_/Q _4604_/A _5963_/B1 _4604_/Y VGND VPWR _9730_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8374_ _8204_/A _8279_/C _8280_/C VGND VPWR _8646_/A VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_7_90 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5586_ _9319_/Q _5585_/A _8846_/X _5585_/Y VGND VPWR _9319_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7325_ _6929_/Y _7059_/D _6801_/Y _7116_/X _7324_/X VGND VPWR _7330_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_190_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4537_ _5259_/A _4537_/B VGND VPWR _4540_/S VGND VPWR sky130_fd_sc_hd__or2_2
XFILLER_116_285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4468_ _8938_/X VGND VPWR _4665_/B VGND VPWR sky130_fd_sc_hd__inv_2
X_7256_ _6176_/Y _7112_/X _6212_/Y _7077_/B VGND VPWR _7256_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_6207_ _6207_/A VGND VPWR _6207_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7187_ _8753_/A _7068_/A _8785_/A _7105_/X VGND VPWR _7187_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_6138_ _9301_/Q VGND VPWR _7282_/A VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_85_331 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_364 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6069_ _6067_/Y _5621_/B _6068_/Y _5507_/B VGND VPWR _6069_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_58_578 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA_216 _7703_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_205 input83/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_60_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_604 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_66 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_77 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_9759_ _4450_/A1 _9759_/D _6146_/A VGND VPWR _9759_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_9_129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_480 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_388 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_263 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_62 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_375 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_288 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_163 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5440_ _9417_/Q _5433_/A _8840_/X _5433_/Y VGND VPWR _9417_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_5371_ _9465_/Q _5368_/A _5965_/B1 _5368_/Y VGND VPWR _9465_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_99_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_380 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8090_ _8218_/A _8096_/B _7968_/A _8120_/A VGND VPWR _8386_/A VGND VPWR sky130_fd_sc_hd__or4bb_4
X_7110_ _7110_/A VGND VPWR _7110_/X VGND VPWR sky130_fd_sc_hd__buf_8
X_7041_ _7041_/A _7073_/C VGND VPWR _7392_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_113_299 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8992_ _8992_/A _8761_/A VGND VPWR mgmt_gpio_out[15] VGND VPWR sky130_fd_sc_hd__ebufn_2
X_7943_ _8636_/A _7943_/B VGND VPWR _7944_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_7874_ _8238_/A _8226_/C VGND VPWR _8239_/B VGND VPWR sky130_fd_sc_hd__or2_2
X_9613_ _9613_/CLK _9613_/D _9646_/SET_B VGND VPWR _9613_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
Xclkbuf_3_7_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/A VGND VPWR _9664_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_2
X_6825_ _9495_/Q VGND VPWR _6825_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_168_428 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9544_ _9768_/CLK _9544_/D _4628_/A VGND VPWR _9544_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6756_ _9356_/Q VGND VPWR _6756_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_148_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5707_ _9252_/Q VGND VPWR _7476_/A VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_164_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9475_ _9687_/CLK _9475_/D _9528_/SET_B VGND VPWR _9475_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6687_ _9179_/Q VGND VPWR _6687_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_12_68 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5638_ _9282_/Q _5634_/A _8840_/X _5634_/Y VGND VPWR _9282_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8426_ _8476_/A _8539_/A VGND VPWR _8601_/D VGND VPWR sky130_fd_sc_hd__or2_2
XFILLER_117_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5569_ _9330_/Q _5566_/A _5965_/B1 _5566_/Y VGND VPWR _9330_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8357_ _8357_/A _8658_/B VGND VPWR _8573_/C VGND VPWR sky130_fd_sc_hd__or2_1
X_7308_ _7308_/A _7308_/B _7308_/C _7308_/D VGND VPWR _7309_/C VGND VPWR sky130_fd_sc_hd__and4_1
X_8288_ _8340_/C _8390_/B _8340_/B _8287_/X VGND VPWR _8288_/X VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_144_34 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7239_ _6246_/Y _5728_/X _6303_/Y _7040_/A _7238_/X VGND VPWR _7242_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_37_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_272 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_412 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_236 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_75 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_472 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_464 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_143 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_198 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4940_ _9092_/Q VGND VPWR _6022_/A VGND VPWR sky130_fd_sc_hd__inv_2
X_5848__9 _8924_/X VGND VPWR _5890_/A1 VGND VPWR sky130_fd_sc_hd__inv_4
X_4871_ _9756_/Q VGND VPWR _4871_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_60_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7590_ _7590_/A _7590_/B _7590_/C _7590_/D VGND VPWR _7590_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
X_6610_ _9349_/Q VGND VPWR _8765_/A VGND VPWR sky130_fd_sc_hd__clkinv_8
XFILLER_20_448 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6541_ _7703_/A _5949_/B _6538_/Y _5178_/B _6540_/X VGND VPWR _6541_/X VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_118_325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6472_ _6467_/Y _5829_/B _6468_/Y _5872_/B _6471_/X VGND VPWR _6473_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9260_ _9601_/CLK _9260_/D _9295_/SET_B VGND VPWR _9260_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_5423_ _9431_/Q _5422_/A _8846_/X _5422_/Y VGND VPWR _9431_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_9191_ _9378_/CLK _9191_/D _9646_/SET_B VGND VPWR _9191_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_8211_ _8341_/B _8264_/B VGND VPWR _8312_/D VGND VPWR sky130_fd_sc_hd__or2_2
X_5354_ _9476_/Q _5346_/A _8916_/A1 _5346_/Y VGND VPWR _9476_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8142_ _8213_/A _8550_/A VGND VPWR _8575_/A VGND VPWR sky130_fd_sc_hd__nor2_1
Xoutput212 _8760_/X VGND VPWR mgmt_gpio_oeb[14] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput223 _8780_/X VGND VPWR mgmt_gpio_oeb[24] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput234 _8800_/X VGND VPWR mgmt_gpio_oeb[34] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput256 _7014_/Y VGND VPWR pad_flash_io0_oeb VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput267 _9723_/Q VGND VPWR pll_div[2] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput245 _8824_/X VGND VPWR mgmt_gpio_out[0] VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_114_575 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_415 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5285_ _9523_/Q _5280_/A _8842_/X _5280_/Y VGND VPWR _9523_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8073_ _8713_/A _8540_/A VGND VPWR _8704_/A VGND VPWR sky130_fd_sc_hd__or2_1
Xoutput278 _9745_/Q VGND VPWR pll_trim[13] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput289 _9755_/Q VGND VPWR pll_trim[23] VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_101_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7024_ _9246_/Q _9245_/Q _7111_/C _7075_/A VGND VPWR _7025_/A VGND VPWR sky130_fd_sc_hd__or4_1
XFILLER_114_48 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8975_ _8742_/X _8728_/X _8975_/S VGND VPWR _8975_/X VGND VPWR sky130_fd_sc_hd__mux2_2
XFILLER_55_378 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7926_ _8305_/A _8270_/B _7925_/Y VGND VPWR _7927_/B VGND VPWR sky130_fd_sc_hd__o21ai_1
X_7857_ _8496_/A _8260_/A VGND VPWR _7858_/A VGND VPWR sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_4_csclk _9329_/CLK VGND VPWR _9380_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_90_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6808_ _6808_/A VGND VPWR _6808_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_23_23 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7788_ _7903_/C _7823_/A _7787_/X VGND VPWR _8528_/B VGND VPWR sky130_fd_sc_hd__o21ai_2
XFILLER_11_437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6739_ _6737_/Y _5534_/B _6738_/Y _5583_/B VGND VPWR _6739_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_9527_ _9527_/CLK _9527_/D _9528_/SET_B VGND VPWR _9527_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_136_122 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9458_ _9789_/CLK _9458_/D _9647_/SET_B VGND VPWR _9458_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_8409_ _8137_/B _8401_/B _8406_/X _8408_/Y VGND VPWR _8409_/X VGND VPWR sky130_fd_sc_hd__o211a_1
XFILLER_124_339 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_9389_ _9775_/CLK _9389_/D _7011_/B VGND VPWR _9389_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_151_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_542 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_315 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_203 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_264 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_40 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_463 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_147 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_467 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5070_ _8965_/X _9663_/Q _5078_/S VGND VPWR _5071_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_49_161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_131 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5972_ _9099_/Q _5970_/A _8845_/X _5970_/Y VGND VPWR _9099_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8760_ _8760_/A VGND VPWR _8760_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_178_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7711_ _7711_/A VGND VPWR _7713_/B VGND VPWR sky130_fd_sc_hd__inv_2
X_4923_ _4914_/Y _5420_/B _4916_/Y _5382_/B _4922_/X VGND VPWR _4934_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_64_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_8691_ _8713_/A _8689_/X _8635_/Y _8690_/Y VGND VPWR _8691_/Y VGND VPWR sky130_fd_sc_hd__o211ai_2
X_4854_ _4846_/Y _5267_/B _4848_/Y _5442_/B _4853_/X VGND VPWR _4864_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_7642_ _6896_/Y _7471_/X _7326_/A _7473_/X _7641_/X VGND VPWR _7643_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_178_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7573_ _6196_/Y _7408_/X _6230_/Y _7410_/X VGND VPWR _7573_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4785_ _4900_/B _4843_/B VGND VPWR _5941_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_6524_ _6522_/Y _5602_/B _8743_/A _5045_/B VGND VPWR _6524_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_9312_ _9534_/CLK _9312_/D _9647_/SET_B VGND VPWR _9312_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_9243_ _9789_/CLK _9243_/D _9647_/SET_B VGND VPWR _9243_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_146_497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6455_ _6455_/A VGND VPWR _8808_/B VGND VPWR sky130_fd_sc_hd__clkinv_4
X_5406_ _5406_/A VGND VPWR _5406_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_6386_ input7/X VGND VPWR _6386_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9174_ _9280_/CLK _9174_/D _9757_/SET_B VGND VPWR _9174_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_133_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_8125_ _8213_/A _8401_/A VGND VPWR _8571_/A VGND VPWR sky130_fd_sc_hd__nor2_1
X_5337_ _5337_/A VGND VPWR _5338_/A VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_102_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8056_ _8389_/A _8168_/A VGND VPWR _8536_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_5268_ _5268_/A VGND VPWR _5269_/A VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_102_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7007_ _4952_/Y _4953_/Y _6023_/Y _9051_/Q _7008_/A VGND VPWR _9051_/D VGND VPWR
+ sky130_fd_sc_hd__a32o_1
X_5199_ _9580_/Q _5193_/Y _8955_/X _5193_/A VGND VPWR _9580_/D VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_141_46 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_378 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8958_ _9090_/Q _9092_/Q _9091_/Q VGND VPWR _8958_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_188_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7909_ _8077_/A _8239_/B _7877_/X _7907_/X _8303_/A VGND VPWR _7909_/X VGND VPWR
+ sky130_fd_sc_hd__o2111a_1
XFILLER_24_551 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8889_ _8888_/X _9145_/Q _9054_/Q VGND VPWR _8889_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_34_66 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_212 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_515 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_400 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_434 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_136 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_383 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_367 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_510 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_584 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4570_ _9752_/Q _4566_/A _5963_/B1 _4566_/Y VGND VPWR _9752_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_162_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_592 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6240_ _9507_/Q VGND VPWR _6240_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_115_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6171_ _9534_/Q VGND VPWR _6171_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_5122_ _5122_/A VGND VPWR _5123_/A VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_111_364 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_256 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5053_ _9669_/Q _5047_/A _8955_/A1 _5047_/Y VGND VPWR _9669_/D VGND VPWR sky130_fd_sc_hd__a22o_1
Xclkbuf_opt_6_0_csclk clkbuf_2_3_0_csclk/X VGND VPWR clkbuf_opt_6_0_csclk/X VGND VPWR
+ sky130_fd_sc_hd__clkbuf_16
X_8812_ _8812_/A _8813_/B VGND VPWR _9061_/D VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_1_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_326 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5955_ _9110_/Q _5951_/A _8925_/A1 _5951_/Y VGND VPWR _9110_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8743_ _8743_/A VGND VPWR _8744_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_4906_ _4906_/A VGND VPWR _4906_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_5886_ _5849_/X _8891_/X _8924_/X _9147_/Q VGND VPWR _9147_/D VGND VPWR sky130_fd_sc_hd__o22a_2
X_8674_ _8674_/A _8674_/B VGND VPWR _8675_/B VGND VPWR sky130_fd_sc_hd__or2_1
X_4837_ _4919_/A _4911_/A VGND VPWR _5232_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_7625_ _7625_/A _7625_/B _7625_/C _7625_/D VGND VPWR _7626_/D VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_178_397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4768_ _7121_/A _5610_/B _4761_/Y _5829_/B _4767_/X VGND VPWR _4790_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_7556_ _6276_/Y _7400_/X _6309_/Y _7405_/X _7555_/X VGND VPWR _7572_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_119_497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7487_ _6818_/Y _7427_/X _6895_/Y _5699_/X VGND VPWR _7487_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_6507_ _8755_/A _5757_/B _6503_/Y _5488_/B _6506_/X VGND VPWR _6526_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_4699_ _9133_/Q VGND VPWR _4699_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_136_35 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6438_ _6438_/A VGND VPWR _6438_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9226_ _9440_/CLK _9226_/D _9685_/SET_B VGND VPWR _9226_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_161_275 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_467 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9157_ _9378_/CLK _9157_/D _9646_/SET_B VGND VPWR _9157_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_121_128 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6369_ _9202_/Q VGND VPWR _6369_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_8108_ _8108_/A VGND VPWR _8640_/A VGND VPWR sky130_fd_sc_hd__buf_6
Xclkbuf_leaf_22_csclk clkbuf_2_3_0_csclk/X VGND VPWR _9601_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
X_9088_ _9089_/CLK _9088_/D _5998_/X VGND VPWR _9088_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_152_23 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8039_ _8039_/A _8416_/A VGND VPWR _8041_/A VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_75_215 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_37_csclk clkbuf_2_1_0_csclk/X VGND VPWR _9639_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_16_348 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_310 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_106 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_343 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_332 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0_mgmt_gpio_in[4] mgmt_gpio_in[4] VGND VPWR clkbuf_0_mgmt_gpio_in[4]/X VGND
+ VPWR sky130_fd_sc_hd__clkbuf_16
XPHY_376 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_354 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_387 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_548 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_412 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_8 _7243_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_125_434 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_74 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_72 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_524 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_440 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_484 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5740_ _5740_/A VGND VPWR _9246_/D VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_175_301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5671_ _5671_/A _5671_/B VGND VPWR _5672_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_7410_ _7410_/A VGND VPWR _7410_/X VGND VPWR sky130_fd_sc_hd__buf_6
X_4622_ _6158_/A _4917_/A VGND VPWR _4623_/B VGND VPWR sky130_fd_sc_hd__or2_2
X_8390_ _8518_/B _8390_/B VGND VPWR _8544_/C VGND VPWR sky130_fd_sc_hd__or2_1
X_4553_ _4669_/A _8932_/X _8946_/X _4729_/B VGND VPWR _4925_/A VGND VPWR sky130_fd_sc_hd__or4_4
X_7341_ _6640_/Y _7068_/A _6725_/Y _7105_/X VGND VPWR _7341_/X VGND VPWR sky130_fd_sc_hd__o22a_2
XFILLER_116_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4484_ _9787_/Q _4466_/A _8930_/A1 _4466_/Y VGND VPWR _9787_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7272_ _6078_/Y _7095_/X _6122_/Y _7068_/D _7271_/X VGND VPWR _7277_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_116_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6223_ _6218_/Y _5949_/B _6219_/Y _4841_/X _6222_/X VGND VPWR _6236_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9011_ _9590_/Q _8799_/A VGND VPWR mgmt_gpio_out[34] VGND VPWR sky130_fd_sc_hd__ebufn_8
X_6154_ _9352_/Q VGND VPWR _6154_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_85_524 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6085_ _6085_/A VGND VPWR _6085_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_5105_ _9643_/Q _5102_/A _5965_/B1 _5102_/Y VGND VPWR _9643_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_57_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5036_ _5981_/B VGND VPWR _5985_/B VGND VPWR sky130_fd_sc_hd__inv_2
Xrepeater375 _7011_/B VGND VPWR _4628_/A VGND VPWR sky130_fd_sc_hd__buf_12
Xrepeater364 _8841_/X VGND VPWR _8955_/A1 VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_65_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6987_ _8810_/A _8809_/A _6974_/A VGND VPWR _9066_/D VGND VPWR sky130_fd_sc_hd__o21ai_1
X_9775_ _9775_/CLK _9775_/D _7011_/B VGND VPWR _9775_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_5938_ _6147_/B _7001_/B VGND VPWR _5938_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
X_8726_ _8077_/A _8246_/B _8243_/A _8314_/X _8504_/C VGND VPWR _8727_/B VGND VPWR
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_166_312 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5869_ _9161_/Q _5866_/A _8841_/X _5866_/Y VGND VPWR _9161_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8657_ _8657_/A _8657_/B _8657_/C _8657_/D VGND VPWR _8696_/C VGND VPWR sky130_fd_sc_hd__or4_2
X_8588_ _8720_/B _8588_/B _8705_/A _8681_/A VGND VPWR _8588_/X VGND VPWR sky130_fd_sc_hd__or4_1
X_7608_ _7608_/A _7608_/B _7608_/C _7608_/D VGND VPWR _7608_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
XFILLER_154_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7539_ _6463_/Y _7419_/X _6403_/Y _7421_/X VGND VPWR _7539_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_181_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_456 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_9209_ _9652_/CLK _9209_/D _9646_/SET_B VGND VPWR _9209_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_0_244 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xinput101 sram_ro_data[17] VGND VPWR _6806_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_88_384 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput123 sram_ro_data[8] VGND VPWR _4892_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput112 sram_ro_data[27] VGND VPWR _6561_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput134 wb_adr_i[12] VGND VPWR _7771_/D VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput145 wb_adr_i[22] VGND VPWR _7781_/B VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_76_524 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xinput156 wb_adr_i[3] VGND VPWR _8379_/D VGND VPWR sky130_fd_sc_hd__buf_4
Xinput167 wb_dat_i[12] VGND VPWR _7745_/B2 VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput178 wb_dat_i[22] VGND VPWR _7748_/B VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_76_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput189 wb_dat_i[3] VGND VPWR _8964_/A1 VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_56_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_432 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_454 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_251 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_151 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_140 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_63 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_194 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_184 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_195 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_359 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_104 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_278 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6910_ _9668_/Q VGND VPWR _6910_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7890_ _7890_/A VGND VPWR _8305_/B VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_47_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6841_ _6839_/Y _4558_/B _6840_/Y _5450_/B VGND VPWR _6841_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_9560_ _9776_/CLK _9560_/D _4628_/A VGND VPWR _9560_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_167_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6772_ _9116_/Q VGND VPWR _6772_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_8511_ _8282_/C _8566_/B _8587_/A _8673_/A VGND VPWR _8512_/D VGND VPWR sky130_fd_sc_hd__a211o_1
XFILLER_148_301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_9491_ _9493_/CLK _9491_/D _4628_/A VGND VPWR _9491_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_5723_ _7104_/A _7098_/C VGND VPWR _7041_/A VGND VPWR sky130_fd_sc_hd__or2_2
X_8442_ _7896_/A _8498_/A _8624_/B _8013_/B VGND VPWR _8444_/A VGND VPWR sky130_fd_sc_hd__o22ai_1
X_5654_ _5649_/B _5751_/C _5647_/A _5651_/B VGND VPWR _5654_/X VGND VPWR sky130_fd_sc_hd__o31a_1
X_4605_ _9731_/Q _4604_/A _8844_/X _4604_/Y VGND VPWR _9731_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8373_ _8373_/A _8693_/B VGND VPWR _8582_/A VGND VPWR sky130_fd_sc_hd__or2_2
XFILLER_144_540 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5585_ _5585_/A VGND VPWR _5585_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7324_ _6874_/Y _7118_/X _6892_/Y _7048_/C VGND VPWR _7324_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4536_ _6111_/A _4929_/A VGND VPWR _4537_/B VGND VPWR sky130_fd_sc_hd__or2_2
XFILLER_116_297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4467_ _9790_/Q _4466_/A _8845_/X _4466_/Y VGND VPWR _9790_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7255_ _7255_/A _7255_/B _7255_/C _7255_/D VGND VPWR _7265_/B VGND VPWR sky130_fd_sc_hd__and4_1
X_6206_ input9/X VGND VPWR _6206_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7186_ _6582_/Y _7059_/B _8797_/A _7068_/C _7185_/X VGND VPWR _7189_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_2
XFILLER_133_14 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6137_ _6132_/Y _6322_/A _6133_/Y _5545_/B _6136_/Y VGND VPWR _6144_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_2
XFILLER_97_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_376 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_218 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6068_ _9371_/Q VGND VPWR _6068_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_26_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5019_ _9692_/Q _5015_/A _8925_/A1 _5015_/Y VGND VPWR _9692_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XANTENNA_206 input83/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_73_549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA_217 _8916_/A1 VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_53_273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_104 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_616 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9758_ _9758_/CLK _9758_/D _7011_/B VGND VPWR _9758_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_139_312 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_492 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8709_ _8709_/A _8709_/B _8709_/C _8709_/D VGND VPWR _8738_/A VGND VPWR sky130_fd_sc_hd__or4_1
X_9689_ _9695_/CLK _9689_/D _9779_/SET_B VGND VPWR _9689_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_21_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_275 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_223 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_74 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_387 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_170 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5370_ _9466_/Q _5368_/A _5964_/B1 _5368_/Y VGND VPWR _9466_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_113_201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_7040_ _7040_/A _7040_/B _7040_/C _7040_/D VGND VPWR _7079_/C VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_141_587 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8991_ _8991_/A _8759_/A VGND VPWR mgmt_gpio_out[14] VGND VPWR sky130_fd_sc_hd__ebufn_2
XFILLER_67_376 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7942_ _8651_/A _8562_/A _7942_/C VGND VPWR _7943_/B VGND VPWR sky130_fd_sc_hd__or3_1
X_9612_ _9788_/CLK _9612_/D _9646_/SET_B VGND VPWR _9612_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_7873_ _7873_/A VGND VPWR _8238_/A VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_168_407 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6824_ _9485_/Q VGND VPWR _6824_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_6755_ _9153_/Q VGND VPWR _6755_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9543_ _9768_/CLK _9543_/D _4628_/A VGND VPWR _9543_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_11_608 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5706_ _7406_/B _5704_/Y _9055_/Q _5705_/X VGND VPWR _9253_/D VGND VPWR sky130_fd_sc_hd__a31o_1
X_9474_ _9687_/CLK _9474_/D _9528_/SET_B VGND VPWR _9474_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_136_304 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6686_ _9366_/Q VGND VPWR _6686_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_8425_ _8688_/A _8631_/A _8425_/C VGND VPWR _8427_/A VGND VPWR sky130_fd_sc_hd__or3_1
XFILLER_163_123 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5637_ _9283_/Q _5634_/A _8841_/X _5634_/Y VGND VPWR _9283_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_5568_ _9331_/Q _5566_/A _5964_/B1 _5566_/Y VGND VPWR _9331_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8356_ _8356_/A _8356_/B _8571_/C _8677_/A VGND VPWR _8360_/A VGND VPWR sky130_fd_sc_hd__or4_1
XFILLER_117_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4519_ _4931_/A _6158_/A _5259_/A VGND VPWR _4520_/S VGND VPWR sky130_fd_sc_hd__or3_1
X_7307_ _4918_/Y _7124_/X _4763_/Y _7068_/B _7306_/X VGND VPWR _7308_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_8287_ _8713_/A _8287_/B VGND VPWR _8287_/X VGND VPWR sky130_fd_sc_hd__or2_1
X_5499_ _9379_/Q _5498_/A _8846_/X _5498_/Y VGND VPWR _9379_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7238_ _7238_/A _7392_/B VGND VPWR _7238_/X VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_144_46 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7169_ _6687_/Y _7040_/D _6737_/Y _7110_/X _7168_/X VGND VPWR _7176_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_37_11 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_590 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_56 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_346 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_284 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_87 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_248 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_276 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_142 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_112 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_540 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_155 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_188 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_91 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_383 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_4870_ _6158_/A _4900_/B VGND VPWR _4870_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_32_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6540_ _4629_/C _8955_/S _6539_/Y _5941_/B VGND VPWR _6540_/X VGND VPWR sky130_fd_sc_hd__o2bb2a_1
XFILLER_60_596 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6471_ _6469_/Y _4524_/B _6470_/Y _4870_/X VGND VPWR _6471_/X VGND VPWR sky130_fd_sc_hd__o22a_2
X_5422_ _5422_/A VGND VPWR _5422_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9190_ _9352_/CLK _9190_/D _9646_/SET_B VGND VPWR _9190_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_8210_ _8210_/A VGND VPWR _8260_/B VGND VPWR sky130_fd_sc_hd__buf_4
X_5353_ _9477_/Q _5346_/A _8840_/X _5346_/Y VGND VPWR _9477_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8141_ _8550_/A _8378_/B VGND VPWR _8362_/A VGND VPWR sky130_fd_sc_hd__nor2_1
Xoutput213 _8762_/X VGND VPWR mgmt_gpio_oeb[15] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput224 _8782_/X VGND VPWR mgmt_gpio_oeb[25] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput235 _8833_/X VGND VPWR mgmt_gpio_oeb[35] VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_99_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xoutput257 _8816_/X VGND VPWR pad_flash_io1_do VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput268 _9724_/Q VGND VPWR pll_div[3] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput246 _8827_/X VGND VPWR mgmt_gpio_out[1] VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_87_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_427 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5284_ _9524_/Q _5280_/A _8925_/A1 _5280_/Y VGND VPWR _9524_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8072_ _8305_/A _8437_/B VGND VPWR _8540_/A VGND VPWR sky130_fd_sc_hd__nor2_1
Xoutput279 _9746_/Q VGND VPWR pll_trim[14] VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_101_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7023_ _9248_/Q _9247_/Q VGND VPWR _7111_/C VGND VPWR sky130_fd_sc_hd__or2_2
X_8974_ _8725_/Y _8697_/X _8975_/S VGND VPWR _8974_/X VGND VPWR sky130_fd_sc_hd__mux2_2
XFILLER_82_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7925_ _8599_/A _7925_/B VGND VPWR _7925_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
X_7856_ _8525_/A _7894_/B _7959_/A _8528_/A VGND VPWR _8260_/A VGND VPWR sky130_fd_sc_hd__or4_4
X_6807_ _9786_/Q VGND VPWR _6807_/Y VGND VPWR sky130_fd_sc_hd__inv_4
X_9526_ _9527_/CLK _9526_/D _9528_/SET_B VGND VPWR _9526_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_7787_ _7959_/A _7787_/B VGND VPWR _7787_/X VGND VPWR sky130_fd_sc_hd__or2_1
X_4999_ _6040_/A VGND VPWR _5000_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_23_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6738_ _9314_/Q VGND VPWR _6738_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_6669_ _6669_/A VGND VPWR _6669_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9457_ _9483_/CLK _9457_/D _9528_/SET_B VGND VPWR _9457_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_136_167 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_134 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8408_ _8607_/B _8573_/A VGND VPWR _8408_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
X_9388_ _9775_/CLK _9388_/D _7011_/B VGND VPWR _9388_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_105_521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_8339_ _8651_/A _8672_/C VGND VPWR _8705_/A VGND VPWR sky130_fd_sc_hd__or2_2
XFILLER_105_554 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_416 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_419 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_66 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_327 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_215 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_276 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_50 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_159 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_202 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_482 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5971_ _9100_/Q _5970_/A _8846_/X _5970_/Y VGND VPWR _9100_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_18_582 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8690_ _8714_/C VGND VPWR _8690_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7710_ _9083_/Q _9082_/Q _7711_/A VGND VPWR _7710_/X VGND VPWR sky130_fd_sc_hd__o21a_1
X_4922_ _4918_/Y _5480_/B _4920_/Y _5518_/B VGND VPWR _4922_/X VGND VPWR sky130_fd_sc_hd__o22a_2
XFILLER_178_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7641_ _6812_/Y _7475_/X _6928_/Y _7477_/X VGND VPWR _7641_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4853_ _4850_/Y _5355_/B _4852_/Y _4524_/B VGND VPWR _4853_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_165_207 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4784_ _9114_/Q VGND VPWR _4784_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7572_ _7572_/A _7572_/B _7572_/C _7572_/D VGND VPWR _7572_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
XFILLER_193_549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_9311_ _9789_/CLK _9311_/D _9685_/SET_B VGND VPWR _9311_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6523_ _9670_/Q VGND VPWR _8743_/A VGND VPWR sky130_fd_sc_hd__inv_4
Xclkbuf_opt_2_0_csclk clkbuf_2_1_0_csclk/X VGND VPWR clkbuf_opt_2_0_csclk/X VGND VPWR
+ sky130_fd_sc_hd__clkbuf_16
X_9242_ _9789_/CLK _9242_/D _9647_/SET_B VGND VPWR _9242_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6454_ _6449_/Y _4590_/B _6450_/Y _6135_/A _6453_/X VGND VPWR _6473_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_5405_ _5405_/A VGND VPWR _5406_/A VGND VPWR sky130_fd_sc_hd__clkbuf_2
X_6385_ _6385_/A VGND VPWR _6385_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9173_ _9280_/CLK _9173_/D _9757_/SET_B VGND VPWR _9173_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_8124_ _8114_/Y _8115_/Y _8115_/Y _8390_/B _8123_/X VGND VPWR _8127_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_5336_ _5671_/A _5336_/B VGND VPWR _5337_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_102_524 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_8055_ _8055_/A _8708_/C VGND VPWR _8057_/A VGND VPWR sky130_fd_sc_hd__nor2_1
X_5267_ _5545_/A _5267_/B VGND VPWR _5268_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_102_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_19 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7006_ _9708_/Q _5993_/B _9048_/Q _9052_/Q VGND VPWR _9052_/D VGND VPWR sky130_fd_sc_hd__a31o_1
X_5198_ _9581_/Q _5193_/Y _8923_/X _5193_/A VGND VPWR _9581_/D VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_55_154 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8957_ _5007_/S _6022_/B _8957_/S VGND VPWR _8957_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_55_176 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7908_ _8521_/B _8232_/B VGND VPWR _8303_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_34_23 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_8888_ _7309_/Y _9627_/Q _8959_/S VGND VPWR _8888_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_78 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7839_ _7839_/A VGND VPWR _8195_/A VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_184_527 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9509_ _9509_/CLK _9509_/D _9528_/SET_B VGND VPWR _9509_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_109_145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_456 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_302 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_52 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_379 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_91 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_596 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6170_ _9292_/Q VGND VPWR _6170_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_130_129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5121_ _5259_/A _5121_/B VGND VPWR _5122_/A VGND VPWR sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_3_csclk _9329_/CLK VGND VPWR _9771_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_111_376 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5052_ _9670_/Q _5047_/A _8929_/A1 _5047_/Y VGND VPWR _9670_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_92_260 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8811_ _8811_/A _8813_/B VGND VPWR _9062_/D VGND VPWR sky130_fd_sc_hd__nor2_1
X_9791_ _9791_/CLK _9791_/D _9633_/SET_B VGND VPWR _9791_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_80_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8742_ _8729_/Y _8723_/Y _8731_/X _8741_/X VGND VPWR _8742_/X VGND VPWR sky130_fd_sc_hd__a31o_1
X_5954_ _9111_/Q _5951_/A _8844_/X _5951_/Y VGND VPWR _9111_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_80_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_360 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4905_ _4897_/Y _5344_/B _4899_/Y _5404_/B _4904_/X VGND VPWR _4934_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_5885_ _5849_/X _8893_/X _8924_/X _9148_/Q VGND VPWR _9148_/D VGND VPWR sky130_fd_sc_hd__o22a_2
X_8673_ _8673_/A _8706_/A _8673_/C _8707_/B VGND VPWR _8673_/X VGND VPWR sky130_fd_sc_hd__or4_2
XFILLER_178_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7624_ _4699_/Y _7471_/X _7304_/A _7473_/X _7623_/X VGND VPWR _7625_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_4836_ _9554_/Q VGND VPWR _4836_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_33_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7555_ _6290_/Y _7408_/X _6303_/Y _7410_/X VGND VPWR _7555_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_146_240 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_379 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6506_ _6504_/Y _5829_/B _6505_/Y _6134_/A VGND VPWR _6506_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4767_ _4763_/Y _5564_/B _4765_/Y _5960_/B VGND VPWR _4767_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_20_14 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7486_ _6890_/Y _7415_/X _6921_/Y _7417_/X _7485_/X VGND VPWR _7500_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_4698_ _4698_/A VGND VPWR _6165_/A VGND VPWR sky130_fd_sc_hd__buf_12
X_6437_ _6435_/Y _5110_/B _6436_/Y _5507_/B VGND VPWR _6437_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_9225_ _9695_/CLK _9225_/D _9779_/SET_B VGND VPWR _9225_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_20_47 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_47 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6368_ _9235_/Q VGND VPWR _6368_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9156_ _9695_/CLK _9156_/D _9779_/SET_B VGND VPWR _9156_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_96_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5319_ _5319_/A VGND VPWR _5319_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_8107_ _8218_/A _8200_/B _8218_/C VGND VPWR _8108_/A VGND VPWR sky130_fd_sc_hd__or3_1
XFILLER_29_12 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6299_ input49/X _8926_/S _6298_/Y _5818_/B VGND VPWR _6299_/X VGND VPWR sky130_fd_sc_hd__o2bb2a_1
X_9087_ _9089_/CLK _9087_/D _6001_/X VGND VPWR _9087_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_102_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_387 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_8038_ _8521_/A _8552_/A VGND VPWR _8416_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_16_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_400 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_271 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_300 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_322 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_311 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_366 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_355 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_344 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_207 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_555 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_262 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_9 _7265_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_3_264 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_192 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_496 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_516 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5670_ _9269_/Q _5662_/A _8839_/X _5662_/Y VGND VPWR _9269_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_175_313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4621_ _4669_/A _8932_/X _8946_/X _8944_/X VGND VPWR _4917_/A VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_163_519 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7340_ _6707_/Y _7059_/B _6719_/Y _7068_/C _7339_/X VGND VPWR _7343_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_4552_ _7731_/A _5062_/D _9759_/Q _8960_/X _4551_/X VGND VPWR _9759_/D VGND VPWR
+ sky130_fd_sc_hd__a32o_1
X_7271_ _6110_/Y _7097_/X _6079_/Y _7099_/X VGND VPWR _7271_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4483_ _4483_/A VGND VPWR _9788_/D VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_131_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_468 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6222_ _6220_/Y _4564_/B _6221_/Y _4893_/X VGND VPWR _6222_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_9010_ _9010_/A _8797_/A VGND VPWR mgmt_gpio_out[33] VGND VPWR sky130_fd_sc_hd__ebufn_8
X_6153_ _6153_/A VGND VPWR _6153_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_6084_ _9739_/Q VGND VPWR _6084_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_5104_ _9644_/Q _5102_/A _5964_/B1 _5102_/Y VGND VPWR _9644_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_85_536 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5035_ _9048_/Q _9050_/Q _9051_/Q VGND VPWR _5981_/B VGND VPWR sky130_fd_sc_hd__or3_1
Xrepeater376 _9757_/SET_B VGND VPWR _9633_/SET_B VGND VPWR sky130_fd_sc_hd__buf_12
Xrepeater365 _8840_/X VGND VPWR _5966_/B1 VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_65_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_271 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6986_ _8811_/A _8809_/A _5939_/X VGND VPWR _9064_/D VGND VPWR sky130_fd_sc_hd__o21ai_1
X_9774_ _9774_/CLK _9774_/D _7011_/B VGND VPWR _9774_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_8725_ _8702_/Y _8733_/A _8712_/Y _8739_/A _8724_/Y VGND VPWR _8725_/Y VGND VPWR
+ sky130_fd_sc_hd__o221ai_1
X_5937_ _9059_/Q _5939_/B VGND VPWR _7001_/B VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_41_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_8656_ _7836_/B _7862_/Y _8518_/A _8367_/B VGND VPWR _8657_/B VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_166_324 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5868_ _9162_/Q _5866_/A _8842_/X _5866_/Y VGND VPWR _9162_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7607_ _7607_/A _7607_/B _7607_/C _7607_/D VGND VPWR _7608_/D VGND VPWR sky130_fd_sc_hd__and4_1
X_4819_ _4816_/Y _5393_/B _4818_/Y _4623_/B VGND VPWR _4819_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_8587_ _8587_/A _8606_/B VGND VPWR _8681_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_5799_ _5799_/A VGND VPWR _5799_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_31_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7538_ _6421_/Y _7400_/X _6371_/Y _7405_/X _7537_/X VGND VPWR _7554_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_181_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7469_ _4716_/Y _7461_/X _4910_/Y _7463_/X _7468_/X VGND VPWR _7480_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_107_468 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9208_ _9788_/CLK _9208_/D _9647_/SET_B VGND VPWR _9208_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_0_201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_330 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9139_ _9278_/CLK _9139_/D _9633_/SET_B VGND VPWR _9139_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
Xinput102 sram_ro_data[18] VGND VPWR _6744_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_193_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xinput124 sram_ro_data[9] VGND VPWR _6808_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput113 sram_ro_data[28] VGND VPWR _6444_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput135 wb_adr_i[13] VGND VPWR _7771_/C VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_48_227 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput157 wb_adr_i[4] VGND VPWR _7894_/B VGND VPWR sky130_fd_sc_hd__buf_4
Xinput146 wb_adr_i[23] VGND VPWR _7781_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput168 wb_dat_i[13] VGND VPWR _7747_/B2 VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_91_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput179 wb_dat_i[23] VGND VPWR _7750_/B VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_189_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_263 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_151 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_152 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_130 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_324 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_163 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_368 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_196 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_606 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_438 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_90 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_116 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_344 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_528 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6840_ _9407_/Q VGND VPWR _6840_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_6771_ _6766_/Y _4907_/X _6767_/Y _5458_/B _6770_/X VGND VPWR _6783_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_23_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_8510_ _8510_/A _8660_/B _8660_/C VGND VPWR _8603_/C VGND VPWR sky130_fd_sc_hd__nor3_1
X_5722_ _7037_/A _7056_/B VGND VPWR _7098_/C VGND VPWR sky130_fd_sc_hd__or2_2
X_9490_ _9545_/CLK _9490_/D _4628_/A VGND VPWR _9490_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_21_csclk clkbuf_2_3_0_csclk/X VGND VPWR _9371_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
X_5653_ _5649_/B _5647_/X _5649_/A _5651_/X _5652_/Y VGND VPWR _9280_/D VGND VPWR
+ sky130_fd_sc_hd__o311a_2
X_8441_ _8441_/A _8441_/B VGND VPWR _8449_/A VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_136_508 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_8372_ _8372_/A _8645_/C _8579_/C _8715_/C VGND VPWR _8375_/A VGND VPWR sky130_fd_sc_hd__or4_4
X_4604_ _4604_/A VGND VPWR _4604_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_5584_ _5584_/A VGND VPWR _5585_/A VGND VPWR sky130_fd_sc_hd__clkbuf_4
X_4535_ _8946_/X _8944_/X _8934_/X _4729_/D VGND VPWR _4929_/A VGND VPWR sky130_fd_sc_hd__or4_4
X_7323_ _6909_/Y _7040_/D _6898_/Y _7110_/X _7322_/X VGND VPWR _7330_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_2
Xclkbuf_leaf_36_csclk clkbuf_2_1_0_csclk/X VGND VPWR _9791_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_144_552 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7254_ _6184_/Y _7048_/D _6157_/Y _7040_/B _7253_/X VGND VPWR _7255_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_4466_ _4466_/A VGND VPWR _4466_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_171_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7185_ _8795_/A _7079_/B _8759_/A _7059_/A VGND VPWR _7185_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_6205_ _9370_/Q VGND VPWR _6205_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
XFILLER_97_160 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6136_ input42/X _8930_/S input51/X _8926_/S VGND VPWR _6136_/Y VGND VPWR sky130_fd_sc_hd__a22oi_1
XFILLER_97_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_48 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_26 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_344 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6067_ _9293_/Q VGND VPWR _6067_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_85_388 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5018_ _9693_/Q _5015_/A _8844_/X _5015_/Y VGND VPWR _9693_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XANTENNA_207 input83/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_218 _8822_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_81_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_296 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9757_ _9757_/CLK _9757_/D _9757_/SET_B VGND VPWR _9757_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6969_ _6629_/Y _6964_/A _9023_/Q _6964_/Y VGND VPWR _9023_/D VGND VPWR sky130_fd_sc_hd__o22a_1
X_8708_ _8708_/A _8708_/B _8708_/C _8708_/D VGND VPWR _8709_/B VGND VPWR sky130_fd_sc_hd__or4_1
X_9688_ _9695_/CLK _9688_/D _9779_/SET_B VGND VPWR _9688_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_8639_ _8115_/Y _8390_/B _8595_/C _8356_/A _8572_/C VGND VPWR _8677_/D VGND VPWR
+ sky130_fd_sc_hd__a2111o_1
XFILLER_21_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_348 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_574 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_235 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_28 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_108 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_31 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_399 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_583 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_182 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_179 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_596 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_311 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8990_ _8990_/A _8757_/A VGND VPWR mgmt_gpio_out[13] VGND VPWR sky130_fd_sc_hd__ebufn_8
XFILLER_94_130 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7941_ _8587_/A _7941_/B VGND VPWR _7942_/C VGND VPWR sky130_fd_sc_hd__or2_1
X_7872_ _8583_/A _8189_/A _7959_/A _8528_/A VGND VPWR _7873_/A VGND VPWR sky130_fd_sc_hd__or4_4
X_9611_ _9613_/CLK _9611_/D _9646_/SET_B VGND VPWR _9611_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6823_ _9071_/Q VGND VPWR _6823_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
X_9542_ _9545_/CLK _9542_/D _4628_/A VGND VPWR _9542_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6754_ _9127_/Q VGND VPWR _6754_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_148_110 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5705_ _5724_/B _7462_/A _5692_/A _9253_/Q VGND VPWR _5705_/X VGND VPWR sky130_fd_sc_hd__o211a_1
X_9473_ _9687_/CLK _9473_/D _9528_/SET_B VGND VPWR _9473_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_6685_ _9685_/Q VGND VPWR _6685_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
X_5636_ _9284_/Q _5634_/A _8842_/X _5634_/Y VGND VPWR _9284_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8424_ _8168_/A _8401_/B _8423_/X VGND VPWR _8425_/C VGND VPWR sky130_fd_sc_hd__o21bai_1
XFILLER_163_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5567_ _9332_/Q _5566_/A _5963_/B1 _5566_/Y VGND VPWR _9332_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8355_ _8683_/B _8499_/B VGND VPWR _8677_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_88_19 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5498_ _5498_/A VGND VPWR _5498_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7306_ _4882_/Y _7126_/X _4809_/Y _7128_/X VGND VPWR _7306_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_8286_ _8585_/B _8721_/A _8286_/C VGND VPWR _8287_/B VGND VPWR sky130_fd_sc_hd__or3_1
X_4518_ _9771_/Q _4517_/Y _5967_/B1 _4517_/A _8939_/X VGND VPWR _9771_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_7237_ _6315_/Y _7059_/D _6276_/Y _7116_/X _7236_/X VGND VPWR _7242_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_4449_ _9577_/Q user_clock _9786_/Q VGND VPWR _8992_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_7168_ _6661_/Y _7112_/X _6755_/Y _7077_/B VGND VPWR _7168_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_6119_ _6119_/A _6119_/B _6119_/C _6119_/D VGND VPWR _6145_/C VGND VPWR sky130_fd_sc_hd__and4_1
X_7099_ _7099_/A VGND VPWR _7099_/X VGND VPWR sky130_fd_sc_hd__buf_8
XFILLER_100_496 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_68 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_33 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_296 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_44 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_124 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_411 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_444 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_146 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_574 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_352 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_290 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_303 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_244 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6470_ _6470_/A VGND VPWR _6470_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_161_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5421_ _5421_/A VGND VPWR _5422_/A VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_173_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5352_ _9478_/Q _5346_/A _8841_/X _5346_/Y VGND VPWR _9478_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8140_ _8140_/A _8574_/A _8361_/A _8730_/A VGND VPWR _8144_/A VGND VPWR sky130_fd_sc_hd__or4_1
Xoutput203 _8806_/X VGND VPWR debug_in VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput214 _8764_/X VGND VPWR mgmt_gpio_oeb[16] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput225 _8784_/X VGND VPWR mgmt_gpio_oeb[26] VGND VPWR sky130_fd_sc_hd__buf_2
X_8071_ _8202_/A _8077_/A VGND VPWR _8713_/A VGND VPWR sky130_fd_sc_hd__nor2_4
Xoutput258 _7017_/Y VGND VPWR pad_flash_io1_ieb VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput247 _8828_/X VGND VPWR mgmt_gpio_out[35] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput236 _8834_/X VGND VPWR mgmt_gpio_oeb[36] VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_141_363 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5283_ _9525_/Q _5280_/A _8844_/X _5280_/Y VGND VPWR _9525_/D VGND VPWR sky130_fd_sc_hd__a22o_1
Xoutput269 _9725_/Q VGND VPWR pll_div[4] VGND VPWR sky130_fd_sc_hd__buf_2
X_7022_ _7022_/A _7022_/B VGND VPWR _7022_/Y VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_87_439 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8973_ _8692_/Y _8664_/X _8975_/S VGND VPWR _8973_/X VGND VPWR sky130_fd_sc_hd__mux2_2
X_7924_ _8463_/A _7924_/B VGND VPWR _7925_/B VGND VPWR sky130_fd_sc_hd__or2_1
X_7855_ _8077_/A _8270_/B VGND VPWR _8599_/A VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_11_406 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_255 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6806_ _6806_/A VGND VPWR _6806_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_23_288 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7786_ _7787_/B VGND VPWR _7823_/A VGND VPWR sky130_fd_sc_hd__inv_2
X_9525_ _9684_/CLK _9525_/D _9685_/SET_B VGND VPWR _9525_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_4998_ _6050_/A VGND VPWR _6040_/A VGND VPWR sky130_fd_sc_hd__buf_8
XFILLER_23_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6737_ _9348_/Q VGND VPWR _6737_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_128_7 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6668_ _9382_/Q VGND VPWR _6668_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9456_ _9509_/CLK _9456_/D _9528_/SET_B VGND VPWR _9456_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_8407_ _8407_/A VGND VPWR _8607_/B VGND VPWR sky130_fd_sc_hd__inv_2
X_6599_ _9729_/Q VGND VPWR _6599_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_5619_ _9295_/Q _5612_/A _8840_/X _5612_/Y VGND VPWR _9295_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_9387_ _9775_/CLK _9387_/D _7011_/B VGND VPWR _9387_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_136_179 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_8338_ _8338_/A VGND VPWR _8338_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_117_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_68 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_352 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_8269_ _8269_/A _8579_/B VGND VPWR _8271_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_171_78 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_163 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_222 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_98 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_260 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_135 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_80 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_91 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_84 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_90 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_6 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_214 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_431 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5970_ _5970_/A VGND VPWR _5970_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_4921_ _4921_/A _4931_/B VGND VPWR _5518_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_178_525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4852_ _9762_/Q VGND VPWR _4852_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7640_ _6909_/Y _7461_/X _6845_/Y _7463_/X _7639_/X VGND VPWR _7643_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_60_383 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_219 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7571_ _7571_/A _7571_/B _7571_/C _7571_/D VGND VPWR _7572_/D VGND VPWR sky130_fd_sc_hd__and4_2
X_4783_ _4783_/A VGND VPWR _6322_/A VGND VPWR sky130_fd_sc_hd__buf_12
X_9310_ _9789_/CLK _9310_/D _9647_/SET_B VGND VPWR _9310_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6522_ _9305_/Q VGND VPWR _6522_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_9_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6453_ _6451_/Y _4861_/X _6452_/Y _4602_/B VGND VPWR _6453_/X VGND VPWR sky130_fd_sc_hd__o22a_2
X_9241_ _9789_/CLK _9241_/D _9647_/SET_B VGND VPWR _9241_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_133_105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_9172_ _9203_/CLK _9172_/D _9757_/SET_B VGND VPWR _9172_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_5404_ _5671_/A _5404_/B VGND VPWR _5405_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_133_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6384_ _9752_/Q VGND VPWR _6384_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_8123_ _8394_/C _7839_/A _8393_/A _8118_/X _8122_/X VGND VPWR _8123_/X VGND VPWR
+ sky130_fd_sc_hd__a41o_2
X_5335_ _9489_/Q _5330_/A _5967_/B1 _5330_/Y VGND VPWR _9489_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_87_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5266_ _9536_/Q _5261_/A _5967_/B1 _5261_/Y VGND VPWR _9536_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8054_ _8624_/B _8168_/A VGND VPWR _8708_/C VGND VPWR sky130_fd_sc_hd__nor2_1
X_7005_ _7005_/A VGND VPWR _9048_/D VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_18_25 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5197_ _9582_/Q _5193_/Y _8920_/X _5193_/A VGND VPWR _9582_/D VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_55_133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_26 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_144 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_8956_ _8955_/S _6322_/Y _8977_/S VGND VPWR _8956_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_7907_ _7864_/X _8230_/A _7887_/Y _7893_/X _7906_/X VGND VPWR _7907_/X VGND VPWR
+ sky130_fd_sc_hd__o2111a_2
X_8887_ _8886_/X _9144_/Q _9054_/Q VGND VPWR _8887_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_51_372 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7838_ _8379_/D _7838_/B _8394_/D _7879_/A VGND VPWR _8298_/A VGND VPWR sky130_fd_sc_hd__or4_1
X_7769_ _8528_/A VGND VPWR _8193_/A VGND VPWR sky130_fd_sc_hd__clkinv_4
XFILLER_11_269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_9508_ _9508_/CLK _9508_/D _9528_/SET_B VGND VPWR _9508_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_9439_ _9440_/CLK _9439_/D _9685_/SET_B VGND VPWR _9439_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_125_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_171 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_88 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_280 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_556 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_411 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_190 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5120_ _9632_/Q _5112_/A _5967_/B1 _5112_/Y VGND VPWR _9632_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_69_214 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_491 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5051_ _9671_/Q _5047_/A _8925_/A1 _5047_/Y VGND VPWR _9671_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_111_388 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_50 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8810_ _8810_/A _8813_/B VGND VPWR _9063_/D VGND VPWR sky130_fd_sc_hd__nor2_1
X_9790_ _9790_/CLK _9790_/D _9757_/SET_B VGND VPWR _9790_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_8741_ _8732_/Y _8733_/Y _8735_/X _8740_/X VGND VPWR _8741_/X VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_92_272 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5953_ _9112_/Q _5951_/A _8845_/X _5951_/Y VGND VPWR _9112_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_80_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8672_ _8703_/B _8672_/B _8672_/C VGND VPWR _8673_/C VGND VPWR sky130_fd_sc_hd__or3_1
X_4904_ _6158_/A _4927_/A _4901_/Y _4902_/Y _5412_/B VGND VPWR _4904_/X VGND VPWR
+ sky130_fd_sc_hd__o32a_1
X_5884_ _5849_/X _8895_/X _8924_/X _9149_/Q VGND VPWR _9149_/D VGND VPWR sky130_fd_sc_hd__o22a_2
XFILLER_33_372 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7623_ _4882_/Y _7475_/X _4706_/Y _7477_/X VGND VPWR _7623_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4835_ _9081_/Q VGND VPWR _4835_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
X_4766_ _6111_/B _4843_/B VGND VPWR _5960_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_7554_ _7554_/A _7554_/B _7554_/C _7554_/D VGND VPWR _7554_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
X_6505_ _6505_/A VGND VPWR _6505_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_107_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7485_ _6910_/Y _7419_/X _6844_/Y _7421_/X VGND VPWR _7485_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4697_ _4787_/A _4903_/B VGND VPWR _4698_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_161_211 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6436_ _9368_/Q VGND VPWR _6436_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9224_ _9695_/CLK _9224_/D _9779_/SET_B VGND VPWR _9224_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_136_59 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9155_ _9695_/CLK _9155_/D _9646_/SET_B VGND VPWR _9155_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6367_ _9208_/Q VGND VPWR _6367_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
XFILLER_0_427 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_8106_ _8200_/C VGND VPWR _8218_/C VGND VPWR sky130_fd_sc_hd__inv_2
X_5318_ _5318_/A VGND VPWR _5319_/A VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_114_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_24 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6298_ _9195_/Q VGND VPWR _6298_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9086_ _9089_/CLK _9086_/D _6004_/X VGND VPWR _9086_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_29_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5249_ _9547_/Q _5242_/A _5966_/B1 _5242_/Y VGND VPWR _9547_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8037_ _8544_/A _7987_/Y _8036_/Y VGND VPWR _8039_/A VGND VPWR sky130_fd_sc_hd__a21oi_1
XFILLER_29_79 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_412 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_8939_ _9710_/Q _9759_/Q _9587_/Q VGND VPWR _8939_/X VGND VPWR sky130_fd_sc_hd__mux2_8
XPHY_334 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_323 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_312 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_322 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_367 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_356 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_33 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_219 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_378 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_274 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_276 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_96 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_604 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_372 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_163 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_528 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4620_ _9721_/Q _4615_/A _5967_/B1 _4615_/Y VGND VPWR _9721_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_187_196 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4551_ _9065_/Q _4551_/B VGND VPWR _4551_/X VGND VPWR sky130_fd_sc_hd__or2_1
X_7270_ _6140_/Y _7048_/B _6120_/Y _7077_/A _7269_/X VGND VPWR _7277_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_4482_ _8955_/A1 _9788_/Q _6018_/S VGND VPWR _4483_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_6221_ _6221_/A VGND VPWR _6221_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_103_108 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6152_ _9378_/Q VGND VPWR _6152_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_106_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5103_ _9645_/Q _5102_/A _5963_/B1 _5102_/Y VGND VPWR _9645_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_6083_ _9553_/Q VGND VPWR _6083_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
X_5034_ _9052_/Q VGND VPWR _5034_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_72_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xrepeater377 _7011_/B VGND VPWR _9757_/SET_B VGND VPWR sky130_fd_sc_hd__buf_12
Xrepeater366 _8840_/X VGND VPWR _8930_/A1 VGND VPWR sky130_fd_sc_hd__buf_12
X_6985_ _9710_/Q _9569_/Q _8977_/S VGND VPWR _8809_/A VGND VPWR sky130_fd_sc_hd__o21ai_4
X_9773_ _9775_/CLK _9773_/D _7011_/B VGND VPWR _9773_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_25_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_264 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8724_ _8729_/A _8731_/C _8723_/Y VGND VPWR _8724_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
X_5936_ _5936_/A _5936_/B _5936_/C _5936_/D VGND VPWR _5939_/B VGND VPWR sky130_fd_sc_hd__or4_2
XFILLER_178_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8655_ _8655_/A VGND VPWR _8655_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_5867_ _9163_/Q _5866_/A _8843_/X _5866_/Y VGND VPWR _9163_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7606_ _6128_/Y _7471_/X _7282_/A _7473_/X _7605_/X VGND VPWR _7607_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_166_336 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_386 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8586_ _8586_/A _8646_/B _8678_/B _8721_/B VGND VPWR _8588_/B VGND VPWR sky130_fd_sc_hd__or4_1
X_4818_ _9719_/Q VGND VPWR _4818_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_5798_ _5798_/A VGND VPWR _5799_/A VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_193_155 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7537_ _6396_/Y _7408_/X _6334_/Y _7410_/X VGND VPWR _7537_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4749_ _9302_/Q VGND VPWR _4749_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_110_7 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7468_ _4734_/Y _7465_/X _4855_/Y _7467_/X VGND VPWR _7468_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_134_244 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9207_ _9788_/CLK _9207_/D _9647_/SET_B VGND VPWR _9207_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_6419_ _6417_/Y _5412_/B _6418_/Y _5024_/B VGND VPWR _6419_/X VGND VPWR sky130_fd_sc_hd__o22a_2
XFILLER_134_288 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7399_ _7476_/A _9251_/Q _7456_/A _7474_/D VGND VPWR _7400_/A VGND VPWR sky130_fd_sc_hd__or4_1
X_9138_ _9203_/CLK _9138_/D _9633_/SET_B VGND VPWR _9138_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_88_342 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9069_ _9790_/CLK _9069_/D _9757_/SET_B VGND VPWR _9069_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
Xinput125 trap VGND VPWR _4901_/A VGND VPWR sky130_fd_sc_hd__buf_6
Xinput103 sram_ro_data[19] VGND VPWR _6558_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput114 sram_ro_data[29] VGND VPWR _6249_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput136 wb_adr_i[14] VGND VPWR _7770_/B VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_48_239 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput158 wb_adr_i[5] VGND VPWR _8525_/A VGND VPWR sky130_fd_sc_hd__buf_6
Xinput147 wb_adr_i[24] VGND VPWR _5925_/C VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput169 wb_dat_i[14] VGND VPWR _7749_/B2 VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_17_604 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_570 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_77 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_294 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_275 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_10 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_32 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_106 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_142 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_120 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_175 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_2_csclk clkbuf_leaf_2_csclk/A VGND VPWR _9514_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XPHY_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_186 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_111 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_299 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_128 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_574 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_0 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6770_ _6768_/Y _4564_/B _6769_/Y _6086_/X VGND VPWR _6770_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_62_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5721_ _9247_/Q VGND VPWR _7056_/B VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_176_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8440_ _7864_/X _8230_/A _8544_/A _8115_/Y VGND VPWR _8665_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_1
X_5652_ _5649_/B _5647_/X _5649_/A VGND VPWR _5652_/Y VGND VPWR sky130_fd_sc_hd__o21ai_2
XFILLER_129_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_572 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8371_ _8708_/D _8506_/B VGND VPWR _8715_/C VGND VPWR sky130_fd_sc_hd__or2_1
X_5583_ _6052_/A _5583_/B VGND VPWR _5584_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_4603_ _4603_/A VGND VPWR _4604_/A VGND VPWR sky130_fd_sc_hd__buf_2
X_4534_ _9762_/Q _4526_/A _5967_/B1 _4526_/Y VGND VPWR _9762_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7322_ _6938_/Y _7112_/X _6896_/Y _7077_/B VGND VPWR _7322_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_144_564 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7253_ _6182_/Y _7068_/A _6199_/Y _7105_/X VGND VPWR _7253_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4465_ _4465_/A VGND VPWR _4466_/A VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_131_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6204_ _6199_/Y _5240_/B _6200_/Y _5393_/B _6203_/X VGND VPWR _6211_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_7184_ _8775_/A _7095_/X _8755_/A _7068_/D _7183_/X VGND VPWR _7189_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_112_450 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6135_ _6135_/A VGND VPWR _8926_/S VGND VPWR sky130_fd_sc_hd__clkinv_8
X_6066_ _9276_/Q VGND VPWR _6066_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_5017_ _9694_/Q _5015_/A _8845_/X _5015_/Y VGND VPWR _9694_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_26_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_412 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_220 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_208 input83/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_26_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9756_ _9757_/CLK _9756_/D _9757_/SET_B VGND VPWR _9756_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_81_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6968_ _6475_/Y _6964_/A _9024_/Q _6964_/Y VGND VPWR _9024_/D VGND VPWR sky130_fd_sc_hd__o22a_2
X_8707_ _8707_/A _8707_/B _8707_/C VGND VPWR _8733_/A VGND VPWR sky130_fd_sc_hd__or3_2
X_5919_ _9124_/Q _5918_/A _5963_/B1 _5918_/Y VGND VPWR _9124_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_6899_ _6897_/Y _5810_/B _6898_/Y _5556_/B VGND VPWR _6899_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_9687_ _9687_/CLK _9687_/D _9685_/SET_B VGND VPWR _9687_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_8638_ _8721_/B VGND VPWR _8638_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_8569_ _8640_/A _8568_/X _8223_/A _8352_/C VGND VPWR _8719_/A VGND VPWR sky130_fd_sc_hd__o211ai_4
XFILLER_181_103 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_586 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_150 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_43 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_304 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_100 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_90 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_19 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_7940_ _8202_/A _8341_/A _7939_/X VGND VPWR _7941_/B VGND VPWR sky130_fd_sc_hd__o21ai_1
X_7871_ _8515_/B _8246_/B VGND VPWR _8734_/A VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_94_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6822_ _6817_/Y _4832_/X _6818_/Y _5393_/B _6821_/X VGND VPWR _6829_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9610_ _9613_/CLK _9610_/D _9646_/SET_B VGND VPWR _9610_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6753_ _9392_/Q VGND VPWR _6753_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9541_ _9545_/CLK _9541_/D _4628_/A VGND VPWR _9541_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_148_122 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5704_ _7462_/A VGND VPWR _5704_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_6684_ _6679_/Y _4861_/X _6680_/Y _6322_/A _6683_/X VGND VPWR _6690_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9472_ _9684_/CLK _9472_/D _9685_/SET_B VGND VPWR _9472_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_176_453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5635_ _9285_/Q _5634_/A _8843_/X _5634_/Y VGND VPWR _9285_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8423_ _8708_/A _8708_/B _8422_/X VGND VPWR _8423_/X VGND VPWR sky130_fd_sc_hd__or3b_1
X_5566_ _5566_/A VGND VPWR _5566_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_8354_ _8354_/A _8595_/B VGND VPWR _8571_/C VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_132_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4517_ _4517_/A VGND VPWR _4517_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7305_ _4858_/Y _5728_/X _4692_/A _7040_/A _7304_/X VGND VPWR _7308_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_2
X_8285_ _8476_/B _8285_/B VGND VPWR _8286_/C VGND VPWR sky130_fd_sc_hd__or2_1
X_5497_ _5497_/A VGND VPWR _5498_/A VGND VPWR sky130_fd_sc_hd__clkbuf_4
X_7236_ _6275_/Y _7118_/X _6321_/Y _7048_/C VGND VPWR _7236_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4448_ _9584_/Q input77/X _8801_/B VGND VPWR _8983_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_86_621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7167_ _7167_/A _7167_/B _7167_/C _7167_/D VGND VPWR _7177_/B VGND VPWR sky130_fd_sc_hd__and4_1
X_7098_ _9246_/Q _9245_/Q _7098_/C _7127_/C VGND VPWR _7099_/A VGND VPWR sky130_fd_sc_hd__or4_1
X_6118_ _6113_/Y _5382_/B _6114_/Y _5355_/B _6117_/X VGND VPWR _6119_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_6049_ _6049_/A VGND VPWR _6049_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_18_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_46 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_304 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_79 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_9739_ _9774_/CLK _9739_/D _9757_/SET_B VGND VPWR _9739_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_127_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_158 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_136 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_456 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_88 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_60 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_331 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_20_csclk clkbuf_2_3_0_csclk/X VGND VPWR _9596_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_134_70 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_96 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_156 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_35_csclk clkbuf_opt_4_0_csclk/X VGND VPWR _9790_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_177_217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_470 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_103 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5420_ _5545_/A _5420_/B VGND VPWR _5421_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_126_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_512 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5351_ _9479_/Q _5346_/A _8842_/X _5346_/Y VGND VPWR _9479_/D VGND VPWR sky130_fd_sc_hd__a22o_1
Xoutput204 _9771_/Q VGND VPWR irq[0] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput215 _8766_/X VGND VPWR mgmt_gpio_oeb[17] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput226 _8786_/X VGND VPWR mgmt_gpio_oeb[27] VGND VPWR sky130_fd_sc_hd__buf_2
X_5282_ _9526_/Q _5280_/A _8845_/X _5280_/Y VGND VPWR _9526_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8070_ _8515_/A _8305_/A _8069_/Y VGND VPWR _8074_/A VGND VPWR sky130_fd_sc_hd__o21bai_1
Xoutput259 _7017_/A VGND VPWR pad_flash_io1_oeb VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput237 _8835_/X VGND VPWR mgmt_gpio_oeb[37] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput248 _8829_/X VGND VPWR mgmt_gpio_out[36] VGND VPWR sky130_fd_sc_hd__buf_2
X_7021_ _7021_/A VGND VPWR _7021_/X VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_141_375 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_518 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_8972_ _8655_/Y _8604_/X _8975_/S VGND VPWR _8972_/X VGND VPWR sky130_fd_sc_hd__mux2_2
XFILLER_55_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_348 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_495 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7923_ _8667_/A _7923_/B VGND VPWR _7924_/B VGND VPWR sky130_fd_sc_hd__or2_1
X_7854_ _8515_/B _8270_/B VGND VPWR _8615_/A VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_51_532 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7785_ _8583_/A _8189_/A _7791_/B VGND VPWR _7787_/B VGND VPWR sky130_fd_sc_hd__or3_1
X_6805_ _9555_/Q VGND VPWR _6805_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_9524_ _9527_/CLK _9524_/D _9528_/SET_B VGND VPWR _9524_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6736_ _9478_/Q VGND VPWR _6736_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
X_4997_ _4997_/A VGND VPWR _9699_/D VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_176_283 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6667_ _9669_/Q VGND VPWR _6667_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9455_ _9483_/CLK _9455_/D _9528_/SET_B VGND VPWR _9455_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6598_ _9549_/Q VGND VPWR _8785_/A VGND VPWR sky130_fd_sc_hd__inv_8
X_5618_ _9296_/Q _5612_/A _8955_/A1 _5612_/Y VGND VPWR _9296_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8406_ _8130_/B _8401_/B _8402_/X _8405_/Y VGND VPWR _8406_/X VGND VPWR sky130_fd_sc_hd__o211a_1
X_9386_ _9777_/CLK _9386_/D _7011_/B VGND VPWR _9386_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_124_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8337_ _8636_/A _8650_/B _8337_/C VGND VPWR _8338_/A VGND VPWR sky130_fd_sc_hd__or3_1
X_5549_ _9344_/Q _5547_/A _8845_/X _5547_/Y VGND VPWR _9344_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_3_606 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_320 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_191 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_504 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_8268_ _8660_/A _8270_/B VGND VPWR _8579_/B VGND VPWR sky130_fd_sc_hd__nor2_1
X_8199_ _8213_/B VGND VPWR _8340_/B VGND VPWR sky130_fd_sc_hd__clkinvlp_2
X_7219_ _6328_/Y _7124_/X _6410_/Y _7068_/B _7218_/X VGND VPWR _7220_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_58_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_326 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_123 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_451 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_272 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_434 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_147 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_92 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_96 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_6_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/A VGND VPWR _4450_/A1 VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_1_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_186 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4920_ _9359_/Q VGND VPWR _4920_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_4851_ _4911_/A _4898_/A VGND VPWR _5355_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_60_395 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7570_ _6302_/Y _7471_/X _7238_/A _7473_/X _7569_/X VGND VPWR _7571_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_4782_ _4787_/A _4898_/A VGND VPWR _4783_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_118_103 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6521_ _6521_/A VGND VPWR _6521_/Y VGND VPWR sky130_fd_sc_hd__inv_4
XFILLER_173_220 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_456 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_147 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6452_ _9730_/Q VGND VPWR _6452_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9240_ _9789_/CLK _9240_/D _9647_/SET_B VGND VPWR _9240_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_106_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5403_ _9442_/Q _5395_/A _8916_/A1 _5395_/Y VGND VPWR _9442_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_9171_ _9280_/CLK _9171_/D _9757_/SET_B VGND VPWR _9171_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_8122_ _7886_/B _8566_/A _8546_/A _8121_/Y VGND VPWR _8122_/X VGND VPWR sky130_fd_sc_hd__o31a_1
X_6383_ _6367_/Y _5797_/B _6370_/X _6376_/X _6382_/X VGND VPWR _6475_/C VGND VPWR
+ sky130_fd_sc_hd__o2111a_1
X_5334_ _9490_/Q _5330_/A _5966_/B1 _5330_/Y VGND VPWR _9490_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_114_375 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5265_ _9537_/Q _5261_/A _5966_/B1 _5261_/Y VGND VPWR _9537_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8053_ _8053_/A _8392_/A VGND VPWR _8055_/A VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_87_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5196_ _9583_/Q _5193_/Y _8915_/X _5193_/A VGND VPWR _9583_/D VGND VPWR sky130_fd_sc_hd__o22a_1
X_7004_ _4964_/B _7008_/A _7008_/B _6022_/B _7003_/X VGND VPWR _7005_/A VGND VPWR
+ sky130_fd_sc_hd__o32a_1
XFILLER_28_304 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8955_ _9620_/Q _8955_/A1 _8955_/S VGND VPWR _8955_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_83_487 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7906_ _7864_/X _7885_/B _7896_/X _7902_/X _7905_/X VGND VPWR _7906_/X VGND VPWR
+ sky130_fd_sc_hd__o2111a_1
X_8886_ _7287_/Y _9639_/Q _8959_/S VGND VPWR _8886_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_70_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_148 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7837_ _7837_/A _7837_/B _7837_/C VGND VPWR _7879_/A VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_140_7 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_384 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7768_ _7768_/A _7768_/B _7768_/C _7768_/D VGND VPWR _7966_/A VGND VPWR sky130_fd_sc_hd__nand4_1
XFILLER_50_24 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_9507_ _9509_/CLK _9507_/D _9528_/SET_B VGND VPWR _9507_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6719_ _9408_/Q VGND VPWR _6719_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_7699_ _7699_/A VGND VPWR _7700_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_164_220 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_46 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9438_ _9514_/CLK _9438_/D _9685_/SET_B VGND VPWR _9438_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_152_415 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_9369_ _9371_/CLK _9369_/D _9295_/SET_B VGND VPWR _9369_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_132_183 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_440 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_292 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_270 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_318 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_340 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_323 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_524 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_568 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_459 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_194 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5050_ _9672_/Q _5047_/A _8844_/X _5047_/Y VGND VPWR _9672_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_77_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5952_ _9113_/Q _5951_/A _8846_/X _5951_/Y VGND VPWR _9113_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8740_ _8712_/B _8737_/Y _8689_/A _8738_/Y _8739_/Y VGND VPWR _8740_/X VGND VPWR
+ sky130_fd_sc_hd__o311a_1
X_4903_ _4911_/A _4903_/B VGND VPWR _5412_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_8671_ _8735_/D _8699_/D _8671_/C _8703_/A VGND VPWR _8671_/Y VGND VPWR sky130_fd_sc_hd__nor4_2
X_5883_ _5849_/X _8897_/X _8924_/X _9150_/Q VGND VPWR _9150_/D VGND VPWR sky130_fd_sc_hd__o22a_2
XFILLER_60_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4834_ _4911_/A _4876_/B VGND VPWR _5431_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_7622_ _4694_/Y _7461_/X _4883_/Y _7463_/X _7621_/X VGND VPWR _7625_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_138_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7553_ _7553_/A _7553_/B _7553_/C _7553_/D VGND VPWR _7554_/D VGND VPWR sky130_fd_sc_hd__and4_1
X_4765_ _9101_/Q VGND VPWR _4765_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_193_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_592 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6504_ _9188_/Q VGND VPWR _6504_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
X_4696_ _8805_/A VGND VPWR _4696_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7484_ _6859_/Y _7400_/X _6891_/Y _7405_/X _7483_/X VGND VPWR _7500_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9223_ _9695_/CLK _9223_/D _9646_/SET_B VGND VPWR _9223_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_174_584 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6435_ _9636_/Q VGND VPWR _6435_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_6366_ _6353_/Y _5818_/B _6355_/X _6359_/X _6365_/X VGND VPWR _6475_/B VGND VPWR
+ sky130_fd_sc_hd__o2111a_2
X_9154_ _9695_/CLK _9154_/D _9779_/SET_B VGND VPWR _9154_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_0_406 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_8105_ _7756_/B _8103_/Y _7837_/B _8103_/A VGND VPWR _8200_/C VGND VPWR sky130_fd_sc_hd__o22a_1
X_9085_ _9089_/CLK _9085_/D _6007_/X VGND VPWR _9085_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_5317_ _5545_/A _5317_/B VGND VPWR _5318_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_102_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8036_ _8389_/A _8551_/A _8035_/X VGND VPWR _8036_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
X_6297_ _9693_/Q VGND VPWR _6297_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_5248_ _9548_/Q _5242_/A _5965_/B1 _5242_/Y VGND VPWR _9548_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_29_36 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5179_ _5179_/A VGND VPWR _5180_/A VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_71_424 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8938_ _8937_/X _9680_/Q _9587_/Q VGND VPWR _8938_/X VGND VPWR sky130_fd_sc_hd__mux2_2
XFILLER_43_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_52 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_324 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_302 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_8869_ _8868_/X _9173_/Q _9054_/Q VGND VPWR _8869_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XPHY_368 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_346 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_335 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_379 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_326 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_45 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_200 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_299 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_590 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_384 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_242 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4550_ _4551_/B VGND VPWR _5062_/D VGND VPWR sky130_fd_sc_hd__inv_6
XFILLER_183_370 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4481_ _5259_/A _4481_/B VGND VPWR _6018_/S VGND VPWR sky130_fd_sc_hd__or2_2
XFILLER_7_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6220_ _9754_/Q VGND VPWR _6220_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_6151_ _9344_/Q VGND VPWR _6151_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_5102_ _5102_/A VGND VPWR _5102_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_85_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6082_ _6078_/Y _5344_/B _6079_/Y _5278_/B _6081_/X VGND VPWR _6096_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_2
XFILLER_57_218 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5033_ _5033_/A VGND VPWR _5033_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_122_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xrepeater367 _8839_/X VGND VPWR _5967_/B1 VGND VPWR sky130_fd_sc_hd__buf_12
X_6984_ _4936_/Y _6976_/A _9012_/Q _6976_/Y VGND VPWR _9012_/D VGND VPWR sky130_fd_sc_hd__o22a_1
X_9772_ _9790_/CLK _9772_/D _9757_/SET_B VGND VPWR _9772_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_5935_ _7837_/C _5935_/B _5935_/C _5934_/X VGND VPWR _5936_/D VGND VPWR sky130_fd_sc_hd__or4b_1
X_8723_ _8723_/A _8723_/B _8723_/C VGND VPWR _8723_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_33_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5866_ _5866_/A VGND VPWR _5866_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_8654_ _8705_/A _8707_/B _8620_/Y _8637_/X _8653_/X VGND VPWR _8655_/A VGND VPWR
+ sky130_fd_sc_hd__o311a_1
XFILLER_178_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_7605_ _6104_/Y _7475_/X _6066_/Y _7477_/X VGND VPWR _7605_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4817_ _4911_/A _4927_/A VGND VPWR _5393_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_166_348 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5797_ _6052_/A _5797_/B VGND VPWR _5798_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_8585_ _8585_/A _8585_/B VGND VPWR _8721_/B VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_147_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4748_ _4726_/Y _5660_/B _4731_/X _4736_/X _4747_/X VGND VPWR _4791_/C VGND VPWR
+ sky130_fd_sc_hd__o2111a_1
X_7536_ _7536_/A _7536_/B _7536_/C _7536_/D VGND VPWR _7536_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
X_4679_ _4787_/A _4925_/A VGND VPWR _5178_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_7467_ _7467_/A VGND VPWR _7467_/X VGND VPWR sky130_fd_sc_hd__buf_8
XFILLER_162_565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_9206_ _9652_/CLK _9206_/D _9647_/SET_B VGND VPWR _9206_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6418_ _9687_/Q VGND VPWR _6418_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
X_7398_ _7456_/A _7462_/A _9255_/Q VGND VPWR _8978_/S VGND VPWR sky130_fd_sc_hd__nor3_4
X_9137_ _9354_/CLK _9137_/D _9685_/SET_B VGND VPWR _9137_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6349_ _9524_/Q VGND VPWR _6349_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
XFILLER_0_258 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9068_ _4450_/A1 _9068_/D _6146_/A VGND VPWR _9068_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
Xinput126 uart_enabled VGND VPWR _8801_/B VGND VPWR sky130_fd_sc_hd__buf_4
Xinput104 sram_ro_data[1] VGND VPWR _6820_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput115 sram_ro_data[2] VGND VPWR _6679_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_102_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8019_ _8612_/A _8016_/X _8019_/C _8441_/B VGND VPWR _8019_/X VGND VPWR sky130_fd_sc_hd__and4bb_1
Xinput159 wb_adr_i[6] VGND VPWR _7903_/C VGND VPWR sky130_fd_sc_hd__buf_4
Xinput137 wb_adr_i[15] VGND VPWR _7770_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput148 wb_adr_i[25] VGND VPWR input148/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_84_582 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_446 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_143 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_110 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_22 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_176 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_154 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_198 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_187 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_134 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_123 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_348 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_508 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_552 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_608 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5720_ _9248_/Q VGND VPWR _7037_/A VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_62_298 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_490 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5651_ _5651_/A _5651_/B VGND VPWR _5651_/X VGND VPWR sky130_fd_sc_hd__or2_2
X_5582_ _9320_/Q _5574_/A _8916_/A1 _5574_/Y VGND VPWR _9320_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_4602_ _5960_/A _4602_/B VGND VPWR _4603_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_8370_ _8370_/A _8599_/B VGND VPWR _8579_/C VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_7_72 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_584 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4533_ _9763_/Q _4526_/A _5966_/B1 _4526_/Y VGND VPWR _9763_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7321_ _7321_/A _7321_/B _7321_/C _7321_/D VGND VPWR _7331_/B VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_190_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_7252_ _6170_/Y _7059_/B _6201_/Y _7068_/C _7251_/X VGND VPWR _7255_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_171_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_576 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6203_ _6201_/Y _6081_/B _6202_/Y _4590_/B VGND VPWR _6203_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4464_ _5960_/A _6251_/A VGND VPWR _4465_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_7183_ _8777_/A _7097_/X _8787_/A _7099_/X VGND VPWR _7183_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_112_462 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6134_ _6134_/A VGND VPWR _8930_/S VGND VPWR sky130_fd_sc_hd__clkinv_8
XFILLER_133_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6065_ _9184_/Q VGND VPWR _6065_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_5016_ _9695_/Q _5015_/A _8846_/X _5015_/Y VGND VPWR _9695_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_38_240 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_209 input83/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_9755_ _9755_/CLK _9755_/D _9757_/SET_B VGND VPWR _9755_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6967_ _6326_/Y _6964_/A _9025_/Q _6964_/Y VGND VPWR _9025_/D VGND VPWR sky130_fd_sc_hd__o22a_1
X_5918_ _5918_/A VGND VPWR _5918_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_8706_ _8706_/A _8706_/B _8706_/C _8706_/D VGND VPWR _8707_/C VGND VPWR sky130_fd_sc_hd__or4_1
XFILLER_41_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6898_ _9334_/Q VGND VPWR _6898_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_139_304 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9686_ _9687_/CLK _9686_/D _9685_/SET_B VGND VPWR _9686_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_158_36 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8637_ _8621_/Y _8633_/Y _8635_/Y _8714_/C VGND VPWR _8637_/X VGND VPWR sky130_fd_sc_hd__a31o_1
X_5849_ _5849_/A VGND VPWR _5849_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_166_156 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_359 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8568_ _8213_/A _8640_/C _8215_/X VGND VPWR _8568_/X VGND VPWR sky130_fd_sc_hd__o21a_1
XFILLER_5_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7519_ _8767_/A _7400_/X _8757_/A _7405_/X VGND VPWR _7519_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_181_159 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_8499_ _8571_/B _8499_/B VGND VPWR _8659_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_135_598 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_11 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_316 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_298 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_432 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7870_ _7870_/A VGND VPWR _8246_/B VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_23_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6821_ _6819_/Y _5431_/B _6820_/Y _4861_/X VGND VPWR _6821_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_9540_ _9768_/CLK _9540_/D _4628_/A VGND VPWR _9540_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_16_490 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6752_ _6748_/Y _5621_/B _6749_/Y _6052_/C _6751_/X VGND VPWR _6759_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_176_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_460 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5703_ _9253_/Q VGND VPWR _7406_/B VGND VPWR sky130_fd_sc_hd__inv_2
X_6683_ _6681_/Y _5013_/B _6682_/Y _5829_/B VGND VPWR _6683_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_9471_ _9687_/CLK _9471_/D _9685_/SET_B VGND VPWR _9471_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_5634_ _5634_/A VGND VPWR _5634_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_8422_ _8554_/A _8401_/B _8419_/X _8421_/Y VGND VPWR _8422_/X VGND VPWR sky130_fd_sc_hd__o211a_1
X_8353_ _8164_/A _8117_/A _8343_/Y _8223_/X _8352_/X VGND VPWR _8356_/B VGND VPWR
+ sky130_fd_sc_hd__o2111ai_4
X_7304_ _7304_/A _7392_/B VGND VPWR _7304_/X VGND VPWR sky130_fd_sc_hd__or2_1
X_5565_ _5565_/A VGND VPWR _5566_/A VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_132_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4516_ _4898_/A _6158_/A VGND VPWR _4517_/A VGND VPWR sky130_fd_sc_hd__or2_2
X_5496_ _5545_/A _5496_/B VGND VPWR _5497_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_8284_ _8539_/A _8284_/B VGND VPWR _8285_/B VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_171_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7235_ _6284_/Y _7040_/D _6277_/Y _7110_/X _7234_/X VGND VPWR _7242_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_4447_ _9570_/Q _4629_/C _9080_/Q VGND VPWR _8985_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_132_568 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7166_ _6637_/Y _7048_/D _6773_/Y _7040_/B _7165_/X VGND VPWR _7167_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_6117_ _6115_/Y _4564_/B _6116_/Y _4491_/B VGND VPWR _6117_/X VGND VPWR sky130_fd_sc_hd__o22a_2
Xclkbuf_leaf_1_csclk _9329_/CLK VGND VPWR _9493_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_100_432 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_335 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7097_ _7097_/A VGND VPWR _7097_/X VGND VPWR sky130_fd_sc_hd__buf_8
X_6048_ _6050_/A VGND VPWR _6049_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_26_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_13 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7999_ _8116_/B _8050_/B VGND VPWR _8000_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_9738_ _9774_/CLK _9738_/D _9757_/SET_B VGND VPWR _9738_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_179_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9669_ _9674_/CLK _9669_/D _9633_/SET_B VGND VPWR _9669_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_10_622 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_424 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_351 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_343 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_568 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_0_0_mgmt_gpio_in[4] clkbuf_2_1_0_mgmt_gpio_in[4]/A VGND VPWR _8837_/A1 VGND
+ VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_49_302 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_482 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_431 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5350_ _9480_/Q _5346_/A _8925_/A1 _5346_/Y VGND VPWR _9480_/D VGND VPWR sky130_fd_sc_hd__a22o_1
Xoutput205 _8807_/Y VGND VPWR irq[1] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput216 _8768_/X VGND VPWR mgmt_gpio_oeb[18] VGND VPWR sky130_fd_sc_hd__buf_2
X_5281_ _9527_/Q _5280_/A _8846_/X _5280_/Y VGND VPWR _9527_/D VGND VPWR sky130_fd_sc_hd__a22o_1
Xoutput238 _7706_/X VGND VPWR mgmt_gpio_oeb[3] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput227 _8788_/X VGND VPWR mgmt_gpio_oeb[28] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput249 _8830_/X VGND VPWR mgmt_gpio_out[37] VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_99_268 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7020_ _9586_/Q _7020_/B VGND VPWR _7021_/A VGND VPWR sky130_fd_sc_hd__and2b_1
XFILLER_68_622 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_132 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_19 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_603 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8971_ _8590_/Y _8513_/X _8975_/S VGND VPWR _8971_/X VGND VPWR sky130_fd_sc_hd__mux2_4
X_7922_ _7836_/B _8299_/B _7862_/Y _7921_/Y VGND VPWR _7923_/B VGND VPWR sky130_fd_sc_hd__a31o_1
X_7853_ _8521_/B _8270_/B VGND VPWR _8325_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_168_207 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6804_ _6799_/Y _5905_/B _6800_/Y _5941_/B _6803_/X VGND VPWR _6830_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_4996_ _8901_/X _9699_/Q _5001_/S VGND VPWR _4997_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_7784_ _7897_/A _7898_/B VGND VPWR _8084_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_9523_ _9684_/CLK _9523_/D _9685_/SET_B VGND VPWR _9523_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_6735_ _9522_/Q VGND VPWR _6735_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_23_38 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9454_ _9483_/CLK _9454_/D _9528_/SET_B VGND VPWR _9454_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_164_424 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6666_ _6661_/Y _5572_/B _6662_/Y _5556_/B _6665_/X VGND VPWR _6691_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_164_435 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_8405_ _8405_/A VGND VPWR _8405_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_5617_ _9297_/Q _5612_/A _8842_/X _5612_/Y VGND VPWR _9297_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_9385_ _9775_/CLK _9385_/D _7011_/B VGND VPWR _9385_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6597_ _9557_/Q VGND VPWR _6597_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_155_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5548_ _9345_/Q _5547_/A _8846_/X _5547_/Y VGND VPWR _9345_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8336_ _8673_/A _8336_/B VGND VPWR _8337_/C VGND VPWR sky130_fd_sc_hd__or2_1
X_8267_ _8267_/A _8599_/B VGND VPWR _8269_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_132_332 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7218_ _6430_/Y _7126_/X _6403_/Y _7128_/X VGND VPWR _7218_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_5479_ _9390_/Q _5471_/A _8916_/A1 _5471_/Y VGND VPWR _9390_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_132_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8198_ _8525_/A _8583_/B _8583_/C VGND VPWR _8213_/B VGND VPWR sky130_fd_sc_hd__or3_1
X_7149_ _6919_/Y _7059_/D _6859_/Y _7116_/X _7148_/X VGND VPWR _7154_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_58_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_316 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_135 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_338 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_34 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_126 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_276 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_340 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_159 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_198 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_91 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4850_ _9468_/Q VGND VPWR _4850_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_33_599 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4781_ _4781_/A VGND VPWR _4781_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_6520_ _9180_/Q VGND VPWR _8747_/A VGND VPWR sky130_fd_sc_hd__clkinv_4
XFILLER_118_115 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_19 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6451_ _6451_/A VGND VPWR _6451_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_9_272 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_159 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_468 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5402_ _9443_/Q _5395_/A _8930_/A1 _5395_/Y VGND VPWR _9443_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_6382_ _6377_/Y _5660_/B _7392_/A _5632_/B _6381_/X VGND VPWR _6382_/X VGND VPWR
+ sky130_fd_sc_hd__o221a_2
X_9170_ _9203_/CLK _9170_/D _9633_/SET_B VGND VPWR _9170_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_173_298 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5333_ _9491_/Q _5330_/A _5965_/B1 _5330_/Y VGND VPWR _9491_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8121_ _8397_/A _8397_/B _8098_/A VGND VPWR _8121_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
X_5264_ _9538_/Q _5261_/A _5965_/B1 _5261_/Y VGND VPWR _9538_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8052_ _8521_/A _8168_/A VGND VPWR _8392_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_5195_ _9584_/Q _5193_/Y _8904_/X _5193_/A VGND VPWR _9584_/D VGND VPWR sky130_fd_sc_hd__o22a_1
X_7003_ _4951_/B _4958_/Y _7003_/C _8958_/X VGND VPWR _7003_/X VGND VPWR sky130_fd_sc_hd__and4bb_1
XFILLER_18_16 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_8954_ _7707_/Y _5214_/A _9050_/Q VGND VPWR _9058_/D VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_70_105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7905_ _8496_/A _8077_/A _8341_/B _7896_/A _8498_/A VGND VPWR _7905_/X VGND VPWR
+ sky130_fd_sc_hd__o32a_1
X_8885_ _8884_/X _9143_/Q _9054_/Q VGND VPWR _8885_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_169_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_382 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_330 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7836_ _7836_/A _7836_/B _7836_/C VGND VPWR _8662_/A VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_149_240 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4979_ _9703_/Q _4966_/A _9702_/Q _4966_/Y VGND VPWR _9703_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7767_ _8394_/A _8394_/B _7767_/C VGND VPWR _7791_/B VGND VPWR sky130_fd_sc_hd__or3_2
X_6718_ _9361_/Q VGND VPWR _6718_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7698_ _7698_/A _7698_/B _7698_/C _7698_/D VGND VPWR _7698_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
X_9506_ _9527_/CLK _9506_/D _9528_/SET_B VGND VPWR _9506_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_50_58 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6649_ _6649_/A _6649_/B _6649_/C VGND VPWR _6785_/A VGND VPWR sky130_fd_sc_hd__and3_1
X_9437_ _9514_/CLK _9437_/D _4628_/A VGND VPWR _9437_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_166_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9368_ _9508_/CLK _9368_/D _9295_/SET_B VGND VPWR _9368_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_34_csclk clkbuf_2_1_0_csclk/X VGND VPWR _9620_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_3_415 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_8319_ _8319_/A _8498_/B VGND VPWR _8493_/C VGND VPWR sky130_fd_sc_hd__nor2_1
X_9299_ _9371_/CLK _9299_/D _9295_/SET_B VGND VPWR _9299_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_78_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_49_csclk _9329_/CLK VGND VPWR _9769_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_74_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_168 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_330 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_352 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_346 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_374 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_582 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_530 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_424 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_275 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_514 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_324 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_488 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5951_ _5951_/A VGND VPWR _5951_/Y VGND VPWR sky130_fd_sc_hd__inv_2
Xclkbuf_1_0_1_mgmt_gpio_in[4] clkbuf_1_0_1_mgmt_gpio_in[4]/A VGND VPWR clkbuf_2_1_0_mgmt_gpio_in[4]/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_2
X_4902_ _9432_/Q VGND VPWR _4902_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_8670_ _8703_/C _8705_/D _8670_/C _8707_/A VGND VPWR _8671_/C VGND VPWR sky130_fd_sc_hd__or4_1
X_5882_ _9151_/Q _5874_/A _8916_/A1 _5874_/Y VGND VPWR _9151_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7621_ _4685_/Y _7465_/X _4888_/Y _7467_/X VGND VPWR _7621_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4833_ _9416_/Q VGND VPWR _4833_/Y VGND VPWR sky130_fd_sc_hd__inv_4
XFILLER_60_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_402 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7552_ _6468_/Y _7471_/X _7216_/A _7473_/X _7551_/X VGND VPWR _7553_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_4764_ _4787_/A _6111_/B VGND VPWR _5564_/B VGND VPWR sky130_fd_sc_hd__or2_2
X_6503_ _9383_/Q VGND VPWR _6503_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7483_ _6865_/Y _7408_/X _6913_/Y _7410_/X VGND VPWR _7483_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_6434_ _9163_/Q VGND VPWR _6434_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_4695_ _4903_/B _4843_/B VGND VPWR _5864_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_9222_ _9695_/CLK _9222_/D _9779_/SET_B VGND VPWR _9222_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6365_ _6360_/Y _5572_/B _6361_/Y _5594_/B _6364_/X VGND VPWR _6365_/X VGND VPWR
+ sky130_fd_sc_hd__o221a_2
X_9153_ _9352_/CLK _9153_/D _9646_/SET_B VGND VPWR _9153_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6296_ _9291_/Q VGND VPWR _6296_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_8104_ _7832_/A _8103_/A _7969_/A _8103_/Y VGND VPWR _8200_/B VGND VPWR sky130_fd_sc_hd__a22o_1
X_5316_ _9502_/Q _5308_/A _8916_/A1 _5308_/Y VGND VPWR _9502_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_9084_ _8837_/A1 _9084_/D _6010_/X VGND VPWR _9084_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_5247_ _9549_/Q _5242_/A _5964_/B1 _5242_/Y VGND VPWR _9549_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8035_ _8035_/A _8460_/A VGND VPWR _8035_/X VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_102_357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_379 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_282 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5178_ _5960_/A _5178_/B VGND VPWR _5179_/A VGND VPWR sky130_fd_sc_hd__or2_2
XFILLER_56_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_179 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8937_ _9087_/Q _9086_/Q _9051_/Q VGND VPWR _8937_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_71_436 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_314 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_303 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_302 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_31 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_190 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8868_ _7662_/Y _9629_/Q _8978_/S VGND VPWR _8868_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XPHY_358 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_347 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_336 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_7819_ _7819_/A VGND VPWR _8660_/B VGND VPWR sky130_fd_sc_hd__clkbuf_4
X_8799_ _8799_/A VGND VPWR _8800_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XPHY_369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_13 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_338 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_254 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_235 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_212 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_514 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_208 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_403 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_322 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_382 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4480_ _6111_/A _4931_/A VGND VPWR _4481_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_143_268 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6150_ _6145_/Y _6149_/A _9043_/Q _6149_/Y VGND VPWR _9043_/D VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_97_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5101_ _5101_/A VGND VPWR _5102_/A VGND VPWR sky130_fd_sc_hd__clkbuf_2
X_6081_ _6081_/A _6081_/B VGND VPWR _6081_/X VGND VPWR sky130_fd_sc_hd__or2_1
X_5032_ _6040_/A VGND VPWR _5033_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xrepeater368 _8839_/X VGND VPWR _8916_/A1 VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_38_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6983_ _6946_/Y _6976_/A _9013_/Q _6976_/Y VGND VPWR _9013_/D VGND VPWR sky130_fd_sc_hd__o22a_1
X_9771_ _9771_/CLK _9771_/D _4628_/A VGND VPWR _9771_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_8722_ _8722_/A _8722_/B _8722_/C VGND VPWR _8723_/B VGND VPWR sky130_fd_sc_hd__or3_1
X_5934_ _7837_/A _7756_/B VGND VPWR _5934_/X VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_80_288 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_8653_ _8638_/Y _8647_/Y _8649_/Y _8652_/X VGND VPWR _8653_/X VGND VPWR sky130_fd_sc_hd__a31o_1
X_5865_ _5865_/A VGND VPWR _5866_/A VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_80_299 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7604_ _6065_/Y _7461_/X _6079_/Y _7463_/X _7603_/X VGND VPWR _7607_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_4816_ _9442_/Q VGND VPWR _4816_/Y VGND VPWR sky130_fd_sc_hd__inv_4
X_5796_ _9212_/Q _5791_/A _5967_/B1 _5791_/Y VGND VPWR _9212_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8584_ _8340_/C _8544_/B _8583_/Y _8330_/B _8380_/B VGND VPWR _8678_/B VGND VPWR
+ sky130_fd_sc_hd__a311o_1
XFILLER_147_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4747_ _4737_/Y _6134_/A _4740_/Y _5818_/B _4746_/X VGND VPWR _4747_/X VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_7535_ _7535_/A _7535_/B _7535_/C _7535_/D VGND VPWR _7536_/D VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_147_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_319 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_371 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7466_ _7466_/A _7476_/C _7474_/D VGND VPWR _7467_/A VGND VPWR sky130_fd_sc_hd__or3_1
X_4678_ _4921_/A _4843_/B VGND VPWR _5080_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_6417_ _9436_/Q VGND VPWR _6417_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9205_ _9613_/CLK _9205_/D _9646_/SET_B VGND VPWR _9205_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_7397_ _7397_/A _7397_/B _7397_/C VGND VPWR _7397_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
XFILLER_122_408 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9136_ _9354_/CLK _9136_/D _9685_/SET_B VGND VPWR _9136_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6348_ _9441_/Q VGND VPWR _6348_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_0_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_290 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_208 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9067_ _4450_/A1 _9067_/D _6146_/A VGND VPWR _9067_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_6279_ _6274_/Y _5382_/B _6275_/Y _5267_/B _6278_/X VGND VPWR _6280_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_2
Xinput105 sram_ro_data[20] VGND VPWR _6438_/A VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
Xinput116 sram_ro_data[30] VGND VPWR _6227_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput127 usr1_vcc_pwrgood VGND VPWR _6593_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_130_496 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_400 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8018_ _8624_/B _8401_/A VGND VPWR _8441_/B VGND VPWR sky130_fd_sc_hd__or2_1
Xinput138 wb_adr_i[16] VGND VPWR _7768_/B VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput149 wb_adr_i[26] VGND VPWR input149/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_17_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_100 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_119 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_300 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_166 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_78 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_199 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_596 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_60 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_238 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_550 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_564 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_244 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5650_ _9054_/Q _6997_/C _9056_/Q VGND VPWR _5651_/B VGND VPWR sky130_fd_sc_hd__a21o_1
XFILLER_87_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4601_ _6111_/A _4921_/A VGND VPWR _4602_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_5581_ _9321_/Q _5574_/A _8930_/A1 _5574_/Y VGND VPWR _9321_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_156_360 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_596 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_62 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4532_ _9764_/Q _4526_/A _5965_/B1 _4526_/Y VGND VPWR _9764_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7320_ _6897_/Y _7048_/D _6833_/Y _7040_/B _7319_/X VGND VPWR _7321_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_183_190 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7251_ _6190_/Y _7079_/B _6179_/Y _7059_/A VGND VPWR _7251_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4463_ _6111_/A _4919_/A VGND VPWR _6251_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_89_108 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_19 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6202_ _9738_/Q VGND VPWR _6202_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_171_385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7182_ _8749_/A _7048_/B _8745_/A _7077_/A _7181_/X VGND VPWR _7189_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_58_506 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6133_ _9345_/Q VGND VPWR _6133_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_58_528 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6064_ _6059_/Y _5968_/B _8807_/B _6165_/A _6063_/X VGND VPWR _6071_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_5015_ _5015_/A VGND VPWR _5015_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_81_553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_9754_ _9755_/CLK _9754_/D _9757_/SET_B VGND VPWR _9754_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6966_ _6237_/Y _6964_/A _9026_/Q _6964_/Y VGND VPWR _9026_/D VGND VPWR sky130_fd_sc_hd__o22a_1
X_8705_ _8705_/A _8705_/B _8705_/C _8705_/D VGND VPWR _8706_/D VGND VPWR sky130_fd_sc_hd__or4_1
X_5917_ _5917_/A VGND VPWR _5918_/A VGND VPWR sky130_fd_sc_hd__clkbuf_2
X_9685_ _9687_/CLK _9685_/D _9685_/SET_B VGND VPWR _9685_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6897_ _9199_/Q VGND VPWR _6897_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_8636_ _8636_/A _8636_/B _8636_/C _8636_/D VGND VPWR _8714_/C VGND VPWR sky130_fd_sc_hd__or4_2
XFILLER_139_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5779_ _9225_/Q _5778_/A _8846_/X _5778_/Y VGND VPWR _9225_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8567_ _8640_/A _8566_/Y _8352_/A VGND VPWR _8641_/B VGND VPWR sky130_fd_sc_hd__o21ai_2
XFILLER_166_168 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7518_ _7518_/A _7518_/B _7518_/C _7518_/D VGND VPWR _7518_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
XFILLER_174_14 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8498_ _8498_/A _8498_/B VGND VPWR _8695_/A VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_150_503 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7449_ _4779_/Y _7441_/X _4850_/Y _7443_/X _7448_/X VGND VPWR _7480_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9119_ _4450_/A1 _9119_/D _6146_/A VGND VPWR _9119_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_76_303 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_474 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_358 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_403 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_414 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_288 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_88 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_439 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_71 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_444 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6820_ _6820_/A VGND VPWR _6820_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_50_203 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6751_ input37/X _8930_/S _6750_/Y _5897_/B VGND VPWR _6751_/X VGND VPWR sky130_fd_sc_hd__o2bb2a_1
XFILLER_176_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5702_ _5696_/Y _5701_/X _5692_/A VGND VPWR _9254_/D VGND VPWR sky130_fd_sc_hd__o21a_1
X_9470_ _9687_/CLK _9470_/D _9528_/SET_B VGND VPWR _9470_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
Xclkbuf_1_1_0_wb_clk_i clkbuf_0_wb_clk_i/X VGND VPWR clkbuf_1_1_1_wb_clk_i/A VGND
+ VPWR sky130_fd_sc_hd__clkbuf_2
X_6682_ _9187_/Q VGND VPWR _6682_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
XFILLER_31_472 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8421_ _8630_/C VGND VPWR _8421_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_5633_ _5633_/A VGND VPWR _5634_/A VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_12_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8352_ _8352_/A _8352_/B _8352_/C VGND VPWR _8352_/X VGND VPWR sky130_fd_sc_hd__and3_1
X_5564_ _5671_/A _5564_/B VGND VPWR _5565_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_128_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7303_ _4765_/Y _7059_/D _4920_/Y _7116_/X _7302_/X VGND VPWR _7308_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_4515_ _4515_/A VGND VPWR _6158_/A VGND VPWR sky130_fd_sc_hd__buf_8
X_5495_ _9380_/Q _5490_/A _5967_/B1 _5490_/Y VGND VPWR _9380_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8283_ _8283_/A _8330_/B VGND VPWR _8284_/B VGND VPWR sky130_fd_sc_hd__or2_1
X_7234_ _6320_/Y _7112_/X _6302_/Y _7077_/B VGND VPWR _7234_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4446_ _9571_/Q _4446_/A1 _9682_/Q VGND VPWR _8986_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_7165_ _6639_/Y _7068_/A _6761_/Y _7105_/X VGND VPWR _7165_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_98_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6116_ _9785_/Q VGND VPWR _6116_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_58_347 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7096_ _7127_/C _7096_/B VGND VPWR _7097_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_39_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6047_ _6047_/A VGND VPWR _6047_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_85_199 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7998_ _7998_/A VGND VPWR _8401_/A VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_53_25 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6949_ _9063_/Q VGND VPWR _6950_/B VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_169_14 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9737_ _9774_/CLK _9737_/D _9757_/SET_B VGND VPWR _9737_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_139_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_271 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9668_ _9674_/CLK _9668_/D _9779_/SET_B VGND VPWR _9668_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_179_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_124 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_8619_ _8619_/A _8707_/A _8706_/B _8619_/D VGND VPWR _8620_/D VGND VPWR sky130_fd_sc_hd__or4_1
XFILLER_155_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_9599_ _9601_/CLK _9599_/D _9528_/SET_B VGND VPWR _9599_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_185_35 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_612 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_271 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_94 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_103 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_60 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_400 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_443 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_494 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xoutput206 _8808_/Y VGND VPWR irq[2] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput217 _8770_/X VGND VPWR mgmt_gpio_oeb[19] VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_114_525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5280_ _5280_/A VGND VPWR _5280_/Y VGND VPWR sky130_fd_sc_hd__inv_2
Xoutput239 _7704_/X VGND VPWR mgmt_gpio_oeb[4] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput228 _8790_/X VGND VPWR mgmt_gpio_oeb[29] VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_141_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_464 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8970_ _8488_/X _8338_/X _8975_/S VGND VPWR _8970_/X VGND VPWR sky130_fd_sc_hd__mux2_4
X_7921_ _8077_/A _8262_/B _7920_/X VGND VPWR _7921_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_70_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_19 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7852_ _7852_/A VGND VPWR _8270_/B VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_90_191 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7783_ _7969_/A _7777_/Y _7832_/A _7777_/A _8218_/A VGND VPWR _7898_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_6803_ _6801_/Y _5518_/B _6802_/Y _5602_/B _6158_/X VGND VPWR _6803_/X VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_4995_ _4995_/A VGND VPWR _4995_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_23_247 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6734_ _6729_/Y _5366_/B _6730_/Y _5298_/B _6733_/X VGND VPWR _6741_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9522_ _9527_/CLK _9522_/D _9528_/SET_B VGND VPWR _9522_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_9453_ _9483_/CLK _9453_/D _9528_/SET_B VGND VPWR _9453_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6665_ _7348_/A _5632_/B _6664_/Y _5679_/B VGND VPWR _6665_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_8404_ _8665_/B _8571_/A VGND VPWR _8405_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_5616_ _9298_/Q _5612_/A _8925_/A1 _5612_/Y VGND VPWR _9298_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_6596_ _6591_/Y _4564_/B _6592_/Y _6086_/X _6595_/X VGND VPWR _6596_/X VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9384_ _9771_/CLK _9384_/D _4628_/A VGND VPWR _9384_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_5547_ _5547_/A VGND VPWR _5547_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_8335_ _8335_/A _8334_/X VGND VPWR _8336_/B VGND VPWR sky130_fd_sc_hd__or2b_1
XFILLER_155_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5478_ _9391_/Q _5471_/A _8840_/X _5471_/Y VGND VPWR _9391_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8266_ _8510_/A _8270_/B VGND VPWR _8599_/B VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_132_344 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7217_ _6422_/Y _5728_/X _6334_/Y _7040_/A _7216_/X VGND VPWR _7220_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_132_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8197_ _8346_/A _8346_/B _8196_/X VGND VPWR _8583_/C VGND VPWR sky130_fd_sc_hd__o21ai_2
X_7148_ _6788_/Y _7118_/X _6915_/Y _7048_/C VGND VPWR _7148_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_100_230 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_464 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7079_ _7127_/C _7079_/B _7079_/C _7079_/D VGND VPWR _7080_/A VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_73_147 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_350 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_67 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_160 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_322 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_355 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_442 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4780_ _6086_/B _4780_/B VGND VPWR _5757_/B VGND VPWR sky130_fd_sc_hd__or2_4
Xclkbuf_leaf_0_csclk _9329_/CLK VGND VPWR _9545_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_146_425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_262 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_127 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6450_ _6450_/A VGND VPWR _6450_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
X_5401_ _9444_/Q _5395_/A _5965_/B1 _5395_/Y VGND VPWR _9444_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_6381_ _6379_/Y _5671_/B _7216_/A _5610_/B VGND VPWR _6381_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_173_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_119 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_439 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5332_ _9492_/Q _5330_/A _5964_/B1 _5330_/Y VGND VPWR _9492_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8120_ _8120_/A _8120_/B VGND VPWR _8397_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_141_130 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5263_ _9539_/Q _5261_/A _5964_/B1 _5261_/Y VGND VPWR _9539_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8051_ _8051_/A VGND VPWR _8168_/A VGND VPWR sky130_fd_sc_hd__buf_2
X_5194_ _9585_/Q _5193_/Y _8914_/X _5193_/A VGND VPWR _9585_/D VGND VPWR sky130_fd_sc_hd__o22a_1
X_7002_ _7002_/A VGND VPWR _9059_/D VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_83_434 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8953_ _9717_/Q _6145_/Y _8957_/S VGND VPWR _8953_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_70_117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_512 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8884_ _7265_/Y _9638_/Q _8959_/S VGND VPWR _8884_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_7904_ _7904_/A VGND VPWR _8498_/A VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_36_394 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7835_ _8496_/A VGND VPWR _7836_/B VGND VPWR sky130_fd_sc_hd__inv_4
XFILLER_169_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7766_ _7838_/B VGND VPWR _7767_/C VGND VPWR sky130_fd_sc_hd__inv_2
X_9505_ _9527_/CLK _9505_/D _9528_/SET_B VGND VPWR _9505_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_4978_ _4978_/A VGND VPWR _4978_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_149_252 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7697_ _7697_/A _7697_/B _7697_/C _7697_/D VGND VPWR _7698_/D VGND VPWR sky130_fd_sc_hd__and4_1
X_6717_ _9496_/Q VGND VPWR _6717_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_192_520 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6648_ _6643_/Y _5757_/B _6644_/Y _5818_/B _6647_/X VGND VPWR _6649_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9436_ _9440_/CLK _9436_/D _4628_/A VGND VPWR _9436_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_125_609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_9367_ _9371_/CLK _9367_/D _9295_/SET_B VGND VPWR _9367_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_8318_ _8318_/A _8490_/C _8597_/C VGND VPWR _8318_/X VGND VPWR sky130_fd_sc_hd__or3_1
X_6579_ _6574_/Y _5298_/B _8767_/A _5496_/B _6578_/X VGND VPWR _6586_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9298_ _9788_/CLK _9298_/D _9295_/SET_B VGND VPWR _9298_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_160_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8249_ _8510_/A _8254_/B VGND VPWR _8250_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_120_347 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_114 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_78 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_40 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_73 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_77 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_211 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_436 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_287 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_526 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_103 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_404 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5950_ _5950_/A VGND VPWR _5951_/A VGND VPWR sky130_fd_sc_hd__clkbuf_4
X_4901_ _4901_/A VGND VPWR _4901_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_5881_ _9152_/Q _5874_/A _8930_/A1 _5874_/Y VGND VPWR _9152_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7620_ _4761_/Y _7451_/X _4899_/Y _7453_/X _7619_/X VGND VPWR _7625_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_4832_ _6111_/A _6086_/B VGND VPWR _4832_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA_190 _7021_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_193_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_4763_ _9328_/Q VGND VPWR _4763_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7551_ _6430_/Y _7475_/X _6377_/Y _7477_/X VGND VPWR _7551_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_6502_ _9234_/Q VGND VPWR _8755_/A VGND VPWR sky130_fd_sc_hd__inv_6
X_4694_ _9159_/Q VGND VPWR _4694_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
X_7482_ _7482_/A VGND VPWR _7482_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_6433_ _6433_/A _6433_/B _6433_/C _6433_/D VGND VPWR _6474_/B VGND VPWR sky130_fd_sc_hd__and4_1
X_9221_ _9695_/CLK _9221_/D _9779_/SET_B VGND VPWR _9221_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_106_119 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_108 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9152_ _9352_/CLK _9152_/D _9646_/SET_B VGND VPWR _9152_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6364_ _6362_/Y _5742_/B _6363_/Y _5556_/B VGND VPWR _6364_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_114_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8103_ _8103_/A VGND VPWR _8103_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_5315_ _9503_/Q _5308_/A _8840_/X _5308_/Y VGND VPWR _9503_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_6295_ _6287_/Y _5545_/B _6288_/Y _5797_/B _6294_/X VGND VPWR _6307_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9083_ _9709_/CLK _9083_/D _6013_/X VGND VPWR _9083_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_114_185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5246_ _9550_/Q _5242_/A _5963_/B1 _5242_/Y VGND VPWR _9550_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8034_ _8624_/B _8551_/A VGND VPWR _8460_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_5177_ _9594_/Q _5169_/A _8916_/A1 _5169_/Y VGND VPWR _9594_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_28_147 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_8936_ _8935_/X _9679_/Q _9587_/Q VGND VPWR _8936_/X VGND VPWR sky130_fd_sc_hd__mux2_2
XFILLER_16_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_315 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_304 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_43 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_8867_ _8866_/X _9172_/Q _9054_/Q VGND VPWR _8867_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XPHY_359 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_348 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_326 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_7818_ _7903_/C _8528_/A _8583_/A _7894_/B VGND VPWR _7819_/A VGND VPWR sky130_fd_sc_hd__or4_1
X_8798_ _8798_/A VGND VPWR _8798_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_177_25 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7749_ _9068_/Q _7749_/A2 _9067_/Q _7749_/B2 _7748_/X VGND VPWR _7749_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_61_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_9419_ _9684_/CLK _9419_/D _9685_/SET_B VGND VPWR _9419_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_180_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_247 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_130 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_40 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_612 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_526 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_291 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_456 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_61 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_211 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_203 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_491 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_472 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5100_ _5259_/A _5100_/B VGND VPWR _5101_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_6080_ _9397_/Q VGND VPWR _6081_/A VGND VPWR sky130_fd_sc_hd__clkinv_2
X_5031_ _9683_/Q _5026_/A _8839_/X _5026_/Y VGND VPWR _9683_/D VGND VPWR sky130_fd_sc_hd__a22o_1
Xrepeater369 _9779_/SET_B VGND VPWR _9646_/SET_B VGND VPWR sky130_fd_sc_hd__buf_12
X_9770_ _9770_/CLK _9770_/D _7011_/B VGND VPWR _9770_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_8721_ _8721_/A _8721_/B _8721_/C _8721_/D VGND VPWR _8722_/C VGND VPWR sky130_fd_sc_hd__or4_1
X_6982_ _6785_/Y _6976_/A _9014_/Q _6976_/Y VGND VPWR _9014_/D VGND VPWR sky130_fd_sc_hd__o22a_1
X_5933_ _7837_/B VGND VPWR _7756_/B VGND VPWR sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_33_csclk clkbuf_2_1_0_csclk/X VGND VPWR _9674_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_178_133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8652_ _8681_/A _8722_/B _8681_/C VGND VPWR _8652_/X VGND VPWR sky130_fd_sc_hd__or3_1
X_5864_ _5960_/A _5864_/B VGND VPWR _5865_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_8583_ _8583_/A _8583_/B _8583_/C VGND VPWR _8583_/Y VGND VPWR sky130_fd_sc_hd__nor3_1
X_7603_ _6121_/Y _7465_/X _6073_/Y _7467_/X VGND VPWR _7603_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4815_ _4911_/A _6158_/B VGND VPWR _6027_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_31_17 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_380 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5795_ _9213_/Q _5791_/A _8930_/A1 _5791_/Y VGND VPWR _9213_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7534_ _7699_/A _7471_/X _8761_/A _7473_/X _7533_/X VGND VPWR _7535_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_4746_ _4742_/Y _5572_/B _4744_/Y _6081_/B VGND VPWR _4746_/X VGND VPWR sky130_fd_sc_hd__o22a_1
Xclkbuf_leaf_48_csclk _9329_/CLK VGND VPWR _9774_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_174_350 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_383 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7465_ _7465_/A VGND VPWR _7465_/X VGND VPWR sky130_fd_sc_hd__buf_8
X_4677_ _9654_/Q VGND VPWR _4677_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_6416_ _9118_/Q VGND VPWR _6416_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9204_ _9652_/CLK _9204_/D _9647_/SET_B VGND VPWR _9204_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_7396_ _7396_/A _7396_/B _7396_/C _7396_/D VGND VPWR _7397_/C VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_162_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_9135_ _9354_/CLK _9135_/D _9685_/SET_B VGND VPWR _9135_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6347_ _9493_/Q VGND VPWR _6347_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_0_216 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_38 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_144 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6278_ _6276_/Y _5496_/B _6277_/Y _5534_/B VGND VPWR _6278_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_9066_ _4450_/A1 _9066_/D _6146_/A VGND VPWR _9066_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
Xinput106 sram_ro_data[21] VGND VPWR _6252_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput117 sram_ro_data[31] VGND VPWR _6097_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_130_464 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_412 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8017_ _8521_/A _8401_/A VGND VPWR _8019_/C VGND VPWR sky130_fd_sc_hd__or2_1
X_5229_ _5229_/A VGND VPWR _9560_/D VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput139 wb_adr_i[17] VGND VPWR _7768_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput128 usr1_vdd_pwrgood VGND VPWR _6847_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_29_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8919_ _9603_/Q _8840_/X _8926_/S VGND VPWR _8919_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XPHY_134 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_167 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_575 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_90 _4450_/A1 VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_21_72 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_72 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_3_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A VGND VPWR clkbuf_3_7_0_wb_clk_i/A VGND
+ VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_121_431 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_87 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_576 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_470 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_194 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4600_ _9732_/Q _4592_/A _5967_/B1 _4592_/Y VGND VPWR _9732_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_5580_ _9322_/Q _5574_/A _8955_/A1 _5574_/Y VGND VPWR _9322_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_175_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4531_ _9765_/Q _4526_/A _5964_/B1 _4526_/Y VGND VPWR _9765_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7250_ _6196_/Y _7095_/X _6183_/Y _7068_/D _7249_/X VGND VPWR _7255_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_4462_ _4729_/A _4729_/B _8934_/X _8932_/X VGND VPWR _4919_/A VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_144_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6201_ _9396_/Q VGND VPWR _6201_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
X_7181_ _8743_/A _7040_/C _7701_/A _7059_/C VGND VPWR _7181_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_6132_ _6132_/A VGND VPWR _6132_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_97_131 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_518 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6063_ _6061_/Y _5583_/B _6062_/Y _5089_/B VGND VPWR _6063_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_5014_ _5014_/A VGND VPWR _5015_/A VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_38_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_448 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9753_ _9755_/CLK _9753_/D _9757_/SET_B VGND VPWR _9753_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6965_ _6145_/Y _6964_/A _9027_/Q _6964_/Y VGND VPWR _9027_/D VGND VPWR sky130_fd_sc_hd__o22a_1
X_9684_ _9684_/CLK _9684_/D _9685_/SET_B VGND VPWR _9684_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_5916_ _5960_/A _5916_/B VGND VPWR _5917_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_8704_ _8704_/A _8704_/B VGND VPWR _8705_/C VGND VPWR sky130_fd_sc_hd__or2_1
X_8635_ _8713_/B _8714_/A VGND VPWR _8635_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
X_6896_ _9134_/Q VGND VPWR _6896_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_21_142 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5847_ _9177_/Q _5839_/A _8916_/A1 _5839_/Y VGND VPWR _9177_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_166_147 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8566_ _8566_/A _8566_/B VGND VPWR _8566_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
X_5778_ _5778_/A VGND VPWR _5778_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_154_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_618 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4729_ _4729_/A _4729_/B _8934_/X _4729_/D VGND VPWR _4900_/B VGND VPWR sky130_fd_sc_hd__or4_4
X_7517_ _7517_/A _7517_/B _7517_/C _7517_/D VGND VPWR _7518_/D VGND VPWR sky130_fd_sc_hd__and4_2
X_8497_ _8497_/A _8395_/X VGND VPWR _8501_/C VGND VPWR sky130_fd_sc_hd__or2b_1
XFILLER_107_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7448_ _4914_/Y _7445_/X _4928_/Y _7447_/X VGND VPWR _7448_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_174_37 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_515 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7379_ _6464_/Y _7040_/C _6331_/Y _7059_/C VGND VPWR _7379_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_1_536 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9118_ _9779_/CLK _9118_/D _9779_/SET_B VGND VPWR _9118_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_103_486 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_9049_ _9709_/CLK _9049_/D _6049_/X VGND VPWR _9049_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_83_23 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_223 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_74 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_426 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_451 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_512 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_71 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_180 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_9 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_567 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_291 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_576 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6750_ _9135_/Q VGND VPWR _6750_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_5701_ _9253_/Q _7462_/A _5724_/B _9254_/Q VGND VPWR _5701_/X VGND VPWR sky130_fd_sc_hd__o31a_1
X_6681_ _9690_/Q VGND VPWR _6681_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_31_484 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_8420_ _8615_/B _8578_/A VGND VPWR _8630_/C VGND VPWR sky130_fd_sc_hd__or2_1
X_5632_ _5671_/A _5632_/B VGND VPWR _5633_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_136_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_19 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_8351_ _8640_/A _8378_/B _8640_/C VGND VPWR _8352_/C VGND VPWR sky130_fd_sc_hd__or3_1
X_5563_ _9333_/Q _5558_/A _8839_/X _5558_/Y VGND VPWR _9333_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_12_19 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_512 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7302_ _4800_/Y _7118_/X _4786_/Y _7048_/C VGND VPWR _7302_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4514_ _8936_/X _8938_/X _4665_/C VGND VPWR _4515_/A VGND VPWR sky130_fd_sc_hd__or3_1
X_5494_ _9381_/Q _5490_/A _5966_/B1 _5490_/Y VGND VPWR _9381_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8282_ _8625_/A _8282_/B _8282_/C VGND VPWR _8330_/B VGND VPWR sky130_fd_sc_hd__and3_1
X_7233_ _7233_/A _7233_/B _7233_/C _7233_/D VGND VPWR _7243_/B VGND VPWR sky130_fd_sc_hd__and4_1
X_4445_ _9572_/Q _4949_/A _9682_/Q VGND VPWR _8987_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_7164_ _6748_/Y _7059_/B _6753_/Y _7068_/C _7163_/X VGND VPWR _7167_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_58_304 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_451 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6115_ _9755_/Q VGND VPWR _6115_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_85_123 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7095_ _7095_/A VGND VPWR _7095_/X VGND VPWR sky130_fd_sc_hd__buf_8
XFILLER_58_359 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6046_ _6050_/A VGND VPWR _6047_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_37_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_543 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_256 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7997_ _8116_/B _7997_/B VGND VPWR _7998_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_156_7 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_26 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9736_ _9774_/CLK _9736_/D _9757_/SET_B VGND VPWR _9736_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6948_ _4936_/Y _6149_/A _9036_/Q _6149_/Y VGND VPWR _9036_/D VGND VPWR sky130_fd_sc_hd__o22a_1
X_6879_ _9205_/Q VGND VPWR _6879_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9667_ _9674_/CLK _9667_/D _9779_/SET_B VGND VPWR _9667_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_167_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_8618_ _8515_/A _8305_/A _8521_/A _8515_/A VGND VPWR _8706_/B VGND VPWR sky130_fd_sc_hd__o22ai_2
X_9598_ _9601_/CLK _9598_/D _9528_/SET_B VGND VPWR _9598_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_139_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_8549_ _8130_/B _8554_/B _8137_/B _8554_/B _8548_/X VGND VPWR _8553_/A VGND VPWR
+ sky130_fd_sc_hd__o221ai_1
XFILLER_185_47 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_526 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_375 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_52 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_311 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_234 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xoutput207 _8831_/X VGND VPWR mgmt_gpio_oeb[0] VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_141_301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput218 _8832_/X VGND VPWR mgmt_gpio_oeb[1] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput229 _8744_/X VGND VPWR mgmt_gpio_oeb[2] VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_99_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_443 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_476 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_104 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7920_ _7864_/X _8319_/A _7917_/Y _8492_/A _8320_/A VGND VPWR _7920_/X VGND VPWR
+ sky130_fd_sc_hd__o2111a_1
X_7851_ _8324_/A _8496_/A VGND VPWR _7852_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_6802_ _9303_/Q VGND VPWR _6802_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_7782_ _7832_/A _7837_/B _7781_/Y _7837_/C _5934_/X VGND VPWR _8218_/A VGND VPWR
+ sky130_fd_sc_hd__a32o_2
X_4994_ _4994_/A VGND VPWR _4995_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_51_568 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6733_ _6731_/Y _5960_/B _6732_/Y _5080_/B VGND VPWR _6733_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_9521_ _9684_/CLK _9521_/D _9685_/SET_B VGND VPWR _9521_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_9452_ _9483_/CLK _9452_/D _9685_/SET_B VGND VPWR _9452_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6664_ _9258_/Q VGND VPWR _6664_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
XFILLER_31_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8403_ _8403_/A VGND VPWR _8665_/B VGND VPWR sky130_fd_sc_hd__inv_2
X_5615_ _9299_/Q _5612_/A _8844_/X _5612_/Y VGND VPWR _9299_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_6595_ _6593_/Y _4868_/X _8795_/A _5431_/B VGND VPWR _6595_/X VGND VPWR sky130_fd_sc_hd__o22a_4
X_9383_ _9771_/CLK _9383_/D _4628_/A VGND VPWR _9383_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_191_256 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_8334_ _8202_/A _8510_/A _8660_/A _8202_/A VGND VPWR _8334_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_5546_ _5546_/A VGND VPWR _5547_/A VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_151_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_108 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5477_ _9392_/Q _5471_/A _8841_/X _5471_/Y VGND VPWR _9392_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8265_ _8265_/A _8645_/B VGND VPWR _8267_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_7216_ _7216_/A _7392_/B VGND VPWR _7216_/X VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_132_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_602 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8196_ _7903_/C _8195_/Y _7839_/A _7960_/Y VGND VPWR _8196_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_1
XFILLER_86_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7147_ _6920_/Y _7040_/D _6793_/Y _7110_/X _7146_/X VGND VPWR _7154_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_100_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_242 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7078_ _7078_/A _7078_/B _7078_/C _7078_/D VGND VPWR _7079_/D VGND VPWR sky130_fd_sc_hd__and4_1
X_6029_ _6029_/A VGND VPWR _6029_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_73_159 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_340 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9719_ _9770_/CLK _9719_/D _7011_/B VGND VPWR _9719_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_120_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_33 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_402 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_318 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_404 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5400_ _9445_/Q _5395_/A _5964_/B1 _5395_/Y VGND VPWR _9445_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_6380_ _9298_/Q VGND VPWR _7216_/A VGND VPWR sky130_fd_sc_hd__inv_4
XFILLER_161_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5331_ _9493_/Q _5330_/A _5963_/B1 _5330_/Y VGND VPWR _9493_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_154_492 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_8050_ _8096_/B _8050_/B VGND VPWR _8051_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_5262_ _9540_/Q _5261_/A _5963_/B1 _5261_/Y VGND VPWR _9540_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7001_ _9065_/Q _7001_/B VGND VPWR _7002_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_5193_ _5193_/A VGND VPWR _5193_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_95_262 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8952_ _9711_/Q _6946_/Y _8957_/S VGND VPWR _8952_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_36_351 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_7903_ _8583_/A _8189_/A _7903_/C _8193_/A VGND VPWR _7904_/A VGND VPWR sky130_fd_sc_hd__or4_1
X_8883_ _8882_/X _9142_/Q _9054_/Q VGND VPWR _8883_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_63_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7834_ _8226_/C VGND VPWR _8496_/A VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_24_524 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7765_ _7894_/B VGND VPWR _8189_/A VGND VPWR sky130_fd_sc_hd__inv_6
X_6716_ _6716_/A _6716_/B _6716_/C _6716_/D VGND VPWR _6784_/A VGND VPWR sky130_fd_sc_hd__and4_1
X_9504_ _9508_/CLK _9504_/D _9528_/SET_B VGND VPWR _9504_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_4977_ _4994_/A VGND VPWR _4978_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_149_264 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7696_ _6441_/Y _7471_/X _7392_/A _7473_/X _7695_/X VGND VPWR _7697_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_177_595 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6647_ _6645_/Y _5742_/B _6646_/Y _5810_/B VGND VPWR _6647_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_9435_ _9440_/CLK _9435_/D _4628_/A VGND VPWR _9435_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6578_ _8779_/A _5267_/B _6577_/Y _5412_/B VGND VPWR _6578_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_9366_ _9508_/CLK _9366_/D _9647_/SET_B VGND VPWR _9366_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_117_161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5529_ _9358_/Q _5528_/A _8843_/X _5528_/Y VGND VPWR _9358_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8317_ _8317_/A _8317_/B VGND VPWR _8597_/C VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_117_194 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9297_ _9788_/CLK _9297_/D _9295_/SET_B VGND VPWR _9297_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_120_304 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8248_ _8248_/A _8490_/B _8317_/B VGND VPWR _8251_/A VGND VPWR sky130_fd_sc_hd__or3_1
XFILLER_132_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_8179_ _8379_/B _8431_/A _8178_/X VGND VPWR _8179_/X VGND VPWR sky130_fd_sc_hd__a21o_1
XFILLER_120_359 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_24 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_402 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_262 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_52 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_448 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_295 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_299 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_538 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_6 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_402 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_416 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_90 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5880_ _9153_/Q _5874_/A _8955_/A1 _5874_/Y VGND VPWR _9153_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_4900_ _4931_/B _4900_/B VGND VPWR _5404_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_4831_ _4831_/A VGND VPWR _4831_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_21_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_191 _7021_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_180 _6785_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_4762_ _4891_/A _4843_/B VGND VPWR _5829_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_7550_ _6457_/Y _7461_/X _6349_/Y _7463_/X _7549_/X VGND VPWR _7553_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_4693_ _4685_/Y _5810_/B _4687_/Y _5949_/B _4692_/X VGND VPWR _4705_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_6501_ _6501_/A _6501_/B _6501_/C _6501_/D VGND VPWR _6629_/A VGND VPWR sky130_fd_sc_hd__and4_1
X_7481_ _7481_/A _7481_/B _7481_/C _7481_/D VGND VPWR _7482_/A VGND VPWR sky130_fd_sc_hd__and4_2
XFILLER_146_256 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6432_ _6427_/Y _5317_/B _6428_/Y _5431_/B _6431_/X VGND VPWR _6433_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9220_ _9695_/CLK _9220_/D _9779_/SET_B VGND VPWR _9220_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_146_267 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_9151_ _9378_/CLK _9151_/D _9646_/SET_B VGND VPWR _9151_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_161_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6363_ _9337_/Q VGND VPWR _6363_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_136_19 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_8102_ _8195_/A _8102_/B VGND VPWR _8103_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_5314_ _9504_/Q _5308_/A _8955_/A1 _5308_/Y VGND VPWR _9504_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_6294_ _6289_/Y _4564_/B _6290_/Y _5344_/B _6293_/X VGND VPWR _6294_/X VGND VPWR
+ sky130_fd_sc_hd__o221a_4
X_9082_ _9709_/CLK _9082_/D _6016_/X VGND VPWR _9082_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_130_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_164 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5245_ _9551_/Q _5242_/A _8844_/X _5242_/Y VGND VPWR _9551_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8033_ _8033_/A _8614_/B VGND VPWR _8035_/A VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_152_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5176_ _9595_/Q _5169_/A _8840_/X _5169_/Y VGND VPWR _9595_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_28_159 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8935_ _9086_/Q _9085_/Q _9051_/Q VGND VPWR _8935_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_71_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_316 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_332 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8866_ _7644_/Y _9628_/Q _8978_/S VGND VPWR _8866_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xclkbuf_3_5_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/A VGND VPWR _9039_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_169_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_338 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_327 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_151 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7817_ _8341_/A VGND VPWR _7836_/C VGND VPWR sky130_fd_sc_hd__inv_2
X_8797_ _8797_/A VGND VPWR _8798_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_7748_ _9066_/Q _7748_/B VGND VPWR _7748_/X VGND VPWR sky130_fd_sc_hd__and2_1
X_7679_ _7679_/A _7679_/B _7679_/C _7679_/D VGND VPWR _7680_/D VGND VPWR sky130_fd_sc_hd__and4_2
X_9418_ _9687_/CLK _9418_/D _9685_/SET_B VGND VPWR _9418_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_3_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_9349_ _9613_/CLK _9349_/D _9646_/SET_B VGND VPWR _9349_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_10_52 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_484 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_74 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_295 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_73 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_416 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_215 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_568 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_291 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_91 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_368 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5030_ _9684_/Q _5026_/A _8840_/X _5026_/Y VGND VPWR _9684_/D VGND VPWR sky130_fd_sc_hd__a22o_1
Xrepeater359 _8843_/X VGND VPWR _5963_/B1 VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_38_468 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6981_ _6629_/Y _6976_/A _9015_/Q _6976_/Y VGND VPWR _9015_/D VGND VPWR sky130_fd_sc_hd__o22a_1
X_5932_ _7832_/A VGND VPWR _7837_/A VGND VPWR sky130_fd_sc_hd__inv_2
X_8720_ _8720_/A _8720_/B _8720_/C VGND VPWR _8721_/D VGND VPWR sky130_fd_sc_hd__or3_1
XFILLER_18_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_123 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5863_ _8924_/X _6997_/A _5862_/Y _5863_/B1 _9164_/Q VGND VPWR _9164_/D VGND VPWR
+ sky130_fd_sc_hd__a32o_2
X_8651_ _8651_/A _8651_/B VGND VPWR _8681_/C VGND VPWR sky130_fd_sc_hd__or2_1
X_5794_ _9214_/Q _5791_/A _5965_/B1 _5791_/Y VGND VPWR _9214_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7602_ _6140_/Y _7451_/X _6113_/Y _7453_/X _7601_/X VGND VPWR _7607_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_8582_ _8582_/A _8582_/B VGND VPWR _8646_/B VGND VPWR sky130_fd_sc_hd__or2_1
X_4814_ _9070_/Q VGND VPWR _4814_/Y VGND VPWR sky130_fd_sc_hd__inv_6
X_7533_ _8783_/A _7475_/X _8759_/A _7477_/X VGND VPWR _7533_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4745_ _4787_/A _4805_/A VGND VPWR _6081_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_119_245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7464_ _7476_/A _9251_/Q _7474_/C _9255_/Q VGND VPWR _7465_/A VGND VPWR sky130_fd_sc_hd__or4_1
X_4676_ _4787_/A _6158_/B VGND VPWR _5507_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_7395_ _6404_/Y _7124_/X _6343_/Y _7068_/B _7394_/X VGND VPWR _7396_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9203_ _9203_/CLK _9203_/D _9633_/SET_B VGND VPWR _9203_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6415_ _9454_/Q VGND VPWR _6415_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
X_6346_ _9532_/Q VGND VPWR _6346_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9134_ _9358_/CLK _9134_/D _9685_/SET_B VGND VPWR _9134_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_9065_ _9664_/CLK _9065_/D _6146_/A VGND VPWR _9065_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6277_ _9351_/Q VGND VPWR _6277_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_8016_ _8016_/A _8016_/B _8016_/C _8016_/D VGND VPWR _8016_/X VGND VPWR sky130_fd_sc_hd__or4_1
Xinput118 sram_ro_data[3] VGND VPWR _6564_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput107 sram_ro_data[22] VGND VPWR _6219_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_102_156 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5228_ _5966_/B1 _9560_/Q _5230_/S VGND VPWR _5229_/A VGND VPWR sky130_fd_sc_hd__mux2_1
Xinput129 usr2_vcc_pwrgood VGND VPWR _6676_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_29_424 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5159_ _9609_/Q _5158_/A _8846_/X _5158_/Y VGND VPWR _9609_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_112_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_8918_ _9608_/Q _8845_/X _8926_/S VGND VPWR _8918_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XPHY_124 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_102 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_8849_ _9618_/Q _8916_/A1 _8955_/S VGND VPWR _8849_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xclkbuf_2_1_0_csclk clkbuf_2_1_0_csclk/A VGND VPWR clkbuf_2_1_0_csclk/X VGND VPWR
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_72_47 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_179 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_168 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_510 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_91 _6326_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_80 _7308_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_180_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_84 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_218 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_443 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_99 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_232 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_276 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_279 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_4 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_482 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_159 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4530_ _9766_/Q _4526_/A _5963_/B1 _4526_/Y VGND VPWR _9766_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_116_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_4461_ _8944_/X VGND VPWR _4729_/B VGND VPWR sky130_fd_sc_hd__clkinv_2
X_6200_ _9448_/Q VGND VPWR _6200_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7180_ _8789_/A _7082_/X _8791_/A _7084_/X _7179_/X VGND VPWR _7199_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_2
X_6131_ _6126_/Y _5776_/B _6127_/Y _5949_/B _6130_/X VGND VPWR _6144_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_112_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6062_ _9653_/Q VGND VPWR _6062_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_5013_ _5960_/A _5013_/B VGND VPWR _5014_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_38_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6964_ _6964_/A VGND VPWR _6964_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9752_ _9755_/CLK _9752_/D _9757_/SET_B VGND VPWR _9752_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_81_599 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5915_ _9125_/Q _5907_/A _8916_/A1 _5907_/Y VGND VPWR _9125_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8703_ _8703_/A _8703_/B _8703_/C _8703_/D VGND VPWR _8706_/C VGND VPWR sky130_fd_sc_hd__or4_1
X_9683_ _9684_/CLK _9683_/D _9685_/SET_B VGND VPWR _9683_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6895_ _9321_/Q VGND VPWR _6895_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_5846_ _9178_/Q _5839_/A _8930_/A1 _5839_/Y VGND VPWR _9178_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8634_ _8544_/A _8092_/Y _8587_/A _8431_/A VGND VPWR _8714_/A VGND VPWR sky130_fd_sc_hd__a211o_1
XFILLER_21_154 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_104 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_8565_ _8565_/A _8640_/B VGND VPWR _8720_/B VGND VPWR sky130_fd_sc_hd__nor2_1
X_5777_ _5777_/A VGND VPWR _5778_/A VGND VPWR sky130_fd_sc_hd__clkbuf_4
X_4728_ _9240_/Q VGND VPWR _4731_/A VGND VPWR sky130_fd_sc_hd__inv_2
X_7516_ _6755_/Y _7471_/X _7172_/A _7473_/X _7515_/X VGND VPWR _7517_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_8496_ _8496_/A _8496_/B VGND VPWR _8695_/C VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_174_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7447_ _7447_/A VGND VPWR _7447_/X VGND VPWR sky130_fd_sc_hd__buf_8
X_4659_ _7003_/C VGND VPWR _8957_/S VGND VPWR sky130_fd_sc_hd__clkinv_4
XFILLER_162_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_7 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_527 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_49 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_526 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7378_ _6397_/Y _7082_/X _6387_/Y _7084_/X _7377_/X VGND VPWR _7397_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_88_110 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_548 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_590 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_9117_ _9785_/CLK _9117_/D _9779_/SET_B VGND VPWR _9117_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6329_ _9506_/Q VGND VPWR _6329_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
XFILLER_130_240 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9048_ _9709_/CLK _9048_/D _6051_/X VGND VPWR _9048_/Q VGND VPWR sky130_fd_sc_hd__dfstp_4
XFILLER_123_31 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_35 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_235 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_110 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_463 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_524 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_579 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_192 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_32_csclk clkbuf_opt_3_0_csclk/X VGND VPWR _9695_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_164_71 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_262 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_240 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_154 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_592 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_47_csclk _9329_/CLK VGND VPWR _9776_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_57_91 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_330 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_588 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5700_ _9255_/Q _5692_/Y _5696_/Y _5724_/B _5699_/X VGND VPWR _9255_/D VGND VPWR
+ sky130_fd_sc_hd__o32a_1
X_6680_ _6680_/A VGND VPWR _6680_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
X_5631_ _9286_/Q _5623_/A _8916_/A1 _5623_/Y VGND VPWR _9286_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_31_496 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5562_ _9334_/Q _5558_/A _8930_/A1 _5558_/Y VGND VPWR _9334_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8350_ _8583_/A _8583_/B _8350_/C VGND VPWR _8640_/C VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_117_524 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4513_ _4669_/A _8932_/X _4729_/A _8944_/X VGND VPWR _4898_/A VGND VPWR sky130_fd_sc_hd__or4_4
X_7301_ _4694_/Y _7040_/D _4660_/Y _7110_/X _7300_/X VGND VPWR _7308_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_2
X_8281_ _8678_/A _8281_/B VGND VPWR _8283_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_5493_ _9382_/Q _5490_/A _5965_/B1 _5490_/Y VGND VPWR _9382_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7232_ _6288_/Y _7048_/D _6314_/Y _7040_/B _7231_/X VGND VPWR _7233_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_144_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4444_ _9589_/Q input78/X _8833_/S VGND VPWR _9010_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_7163_ _6720_/Y _7079_/B _6633_/Y _7059_/A VGND VPWR _7163_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_7094_ _7127_/C _7094_/B VGND VPWR _7095_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_6114_ _9475_/Q VGND VPWR _6114_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
XFILLER_112_273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6045_ _6045_/A VGND VPWR _6045_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_100_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_179 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_555 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9735_ _9774_/CLK _9735_/D _9757_/SET_B VGND VPWR _9735_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_7996_ _7996_/A VGND VPWR _8130_/B VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_81_385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6947_ _6149_/A _6946_/Y _9037_/Q _6149_/Y VGND VPWR _9037_/D VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_149_7 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6878_ _6878_/A _6878_/B _6878_/C _6878_/D VGND VPWR _6946_/B VGND VPWR sky130_fd_sc_hd__and4_1
X_9666_ _4450_/A1 _9666_/D _6146_/A VGND VPWR _9666_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_9597_ _9601_/CLK _9597_/D _9528_/SET_B VGND VPWR _9597_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_5829_ _5960_/A _5829_/B VGND VPWR _5830_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_8617_ _8617_/A _8617_/B VGND VPWR _8707_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_8548_ _8393_/Y _8554_/B _8401_/A _8554_/B _8547_/X VGND VPWR _8548_/X VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_5_106 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8479_ _8704_/B _8479_/B VGND VPWR _8481_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_123_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_538 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_323 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_327 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_12 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_67 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_330 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_50 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_8 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_71 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_343 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xoutput208 _8752_/X VGND VPWR mgmt_gpio_oeb[10] VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_126_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput219 _8772_/X VGND VPWR mgmt_gpio_oeb[20] VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_4_43 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_590 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_116 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_500 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7850_ _7850_/A VGND VPWR _8521_/B VGND VPWR sky130_fd_sc_hd__buf_12
X_6801_ _9360_/Q VGND VPWR _6801_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_23_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_547 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7781_ _7781_/A _7781_/B VGND VPWR _7781_/Y VGND VPWR sky130_fd_sc_hd__nand2_1
X_4993_ _4993_/A VGND VPWR _9700_/D VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_6732_ _9656_/Q VGND VPWR _6732_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9520_ _9527_/CLK _9520_/D _9528_/SET_B VGND VPWR _9520_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6663_ _9283_/Q VGND VPWR _7348_/A VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_139_19 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9451_ _9483_/CLK _9451_/D _9685_/SET_B VGND VPWR _9451_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_31_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5614_ _9300_/Q _5612_/A _8845_/X _5612_/Y VGND VPWR _9300_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8402_ _8213_/A _8117_/A _8019_/C _8400_/X _8401_/X VGND VPWR _8402_/X VGND VPWR
+ sky130_fd_sc_hd__o2111a_1
X_9382_ _9771_/CLK _9382_/D _4628_/A VGND VPWR _9382_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6594_ _9419_/Q VGND VPWR _8795_/A VGND VPWR sky130_fd_sc_hd__inv_6
X_8333_ _8720_/A _8713_/A _8333_/C VGND VPWR _8335_/A VGND VPWR sky130_fd_sc_hd__or3_1
X_5545_ _5545_/A _5545_/B VGND VPWR _5546_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_5476_ _9393_/Q _5471_/A _8842_/X _5471_/Y VGND VPWR _9393_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8264_ _8324_/A _8264_/B VGND VPWR _8645_/B VGND VPWR sky130_fd_sc_hd__nor2_1
X_8195_ _8195_/A _8195_/B VGND VPWR _8195_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
X_7215_ _6456_/Y _7059_/D _6421_/Y _7116_/X _7214_/X VGND VPWR _7220_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_7146_ _6895_/Y _7112_/X _6889_/Y _7077_/B VGND VPWR _7146_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_86_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7077_ _7077_/A _7077_/B _7077_/C _7077_/D VGND VPWR _7078_/D VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_100_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6028_ _6028_/A VGND VPWR _6029_/A VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_39_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_588 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_7979_ _7979_/A VGND VPWR _7994_/A VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_42_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9718_ _8837_/A1 _9718_/D _4994_/A VGND VPWR _9718_/Q VGND VPWR sky130_fd_sc_hd__dfrtn_1
X_9649_ _9652_/CLK _9649_/D _9646_/SET_B VGND VPWR _9649_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_155_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_118 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_63 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_519 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_120 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_606 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_179 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_71 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_414 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_80 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_438 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_302 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5330_ _5330_/A VGND VPWR _5330_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_5_481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5261_ _5261_/A VGND VPWR _5261_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7000_ _9056_/Q _5753_/B _6996_/Y _7000_/B2 VGND VPWR _9056_/D VGND VPWR sky130_fd_sc_hd__a22o_2
X_5192_ _6322_/A _6165_/A _5259_/A _8956_/X VGND VPWR _5193_/A VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_68_455 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_274 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8951_ _9712_/Q _6785_/Y _8957_/S VGND VPWR _8951_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_56_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_596 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7902_ _8077_/A _7902_/B VGND VPWR _7902_/X VGND VPWR sky130_fd_sc_hd__or2_1
X_8882_ _7243_/Y _9637_/Q _8959_/S VGND VPWR _8882_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_7833_ _7833_/A VGND VPWR _8226_/C VGND VPWR sky130_fd_sc_hd__buf_8
X_7764_ _7764_/A VGND VPWR _8510_/A VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_149_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_4976_ _9704_/Q _4966_/A _9703_/Q _4966_/Y VGND VPWR _9704_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_9503_ _9527_/CLK _9503_/D _9528_/SET_B VGND VPWR _9503_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6715_ _6710_/Y _5420_/B _6711_/Y _5259_/B _6714_/X VGND VPWR _6716_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_7695_ _6429_/Y _7475_/X _6379_/Y _7477_/X VGND VPWR _7695_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_149_276 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_298 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6646_ _9200_/Q VGND VPWR _6646_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_192_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9434_ _9440_/CLK _9434_/D _4628_/A VGND VPWR _9434_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_192_544 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6577_ _9435_/Q VGND VPWR _6577_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9365_ _9508_/CLK _9365_/D _9647_/SET_B VGND VPWR _9365_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_133_611 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5528_ _5528_/A VGND VPWR _5528_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_8316_ _8316_/A _8498_/B VGND VPWR _8490_/C VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_132_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_9296_ _9788_/CLK _9296_/D _9295_/SET_B VGND VPWR _9296_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_8247_ _8319_/A _8264_/B VGND VPWR _8317_/B VGND VPWR sky130_fd_sc_hd__nor2_1
X_5459_ _5459_/A VGND VPWR _5460_/A VGND VPWR sky130_fd_sc_hd__clkbuf_4
X_8178_ _8703_/A _8178_/B VGND VPWR _8178_/X VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_101_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7129_ _4814_/Y _7126_/X _4857_/Y _7128_/X VGND VPWR _7129_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_75_36 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_574 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_76 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_98 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_108 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_64 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_514 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_522 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_460 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_61 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_176 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_60 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_414 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_222 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_4830_ _4830_/A _4830_/B _4830_/C _4830_/D VGND VPWR _4935_/A VGND VPWR sky130_fd_sc_hd__and4_1
XANTENNA_170 _6902_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_21_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA_192 _7021_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_181 _4901_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_60_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4761_ _9185_/Q VGND VPWR _4761_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_6500_ _7370_/A _5632_/B _7701_/A _5905_/B _6499_/X VGND VPWR _6501_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_7480_ _7480_/A _7480_/B _7480_/C _7480_/D VGND VPWR _7481_/D VGND VPWR sky130_fd_sc_hd__and4_1
X_4692_ _4692_/A _5024_/B VGND VPWR _4692_/X VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_174_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6431_ _6429_/Y _4504_/B _6430_/Y _6027_/B VGND VPWR _6431_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_6362_ _9244_/Q VGND VPWR _6362_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9150_ _9280_/CLK _9150_/D _9757_/SET_B VGND VPWR _9150_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_5313_ _9505_/Q _5308_/A _8842_/X _5308_/Y VGND VPWR _9505_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8101_ _8213_/A VGND VPWR _8625_/A VGND VPWR sky130_fd_sc_hd__clkinv_2
X_6293_ _6291_/Y _6027_/B _6292_/Y _4893_/X VGND VPWR _6293_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_9081_ _9788_/CLK _9081_/D _9646_/SET_B VGND VPWR _9081_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_88_528 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_176 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5244_ _9552_/Q _5242_/A _8845_/X _5242_/Y VGND VPWR _9552_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8032_ _8521_/A _8551_/A VGND VPWR _8614_/B VGND VPWR sky130_fd_sc_hd__nor2_1
X_5175_ _9596_/Q _5169_/A _8841_/X _5169_/Y VGND VPWR _9596_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_110_360 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_211 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_127 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_458 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8934_ _8933_/X _9678_/Q _9587_/Q VGND VPWR _8934_/X VGND VPWR sky130_fd_sc_hd__mux2_4
XFILLER_83_288 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_8865_ _8864_/X _9171_/Q _9054_/Q VGND VPWR _8865_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_344 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_306 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_7816_ _8202_/A _8097_/B VGND VPWR _8094_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_51_163 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_339 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_328 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_8796_ _8796_/A VGND VPWR _8796_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_24_355 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_399 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7747_ _9068_/Q _7747_/A2 _9067_/Q _7747_/B2 _7746_/X VGND VPWR _7747_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_4959_ _9048_/Q VGND VPWR _6022_/B VGND VPWR sky130_fd_sc_hd__clkinv_4
XFILLER_131_7 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_371 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7678_ _6528_/Y _7471_/X _7370_/A _7473_/X _7677_/X VGND VPWR _7679_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_177_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9417_ _9684_/CLK _9417_/D _9685_/SET_B VGND VPWR _9417_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6629_ _6629_/A _6629_/B _6629_/C _6629_/D VGND VPWR _6629_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
X_9348_ _9352_/CLK _9348_/D _9646_/SET_B VGND VPWR _9348_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_133_430 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_64 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9279_ _9280_/CLK _9279_/D _9633_/SET_B VGND VPWR _9279_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_133_474 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_496 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_152 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_235 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_576 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_550 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_146 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6980_ _6475_/Y _6976_/A _9016_/Q _6976_/Y VGND VPWR _9016_/D VGND VPWR sky130_fd_sc_hd__o22a_2
XFILLER_80_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5931_ _5931_/A _5931_/B input163/X input201/X VGND VPWR _5935_/C VGND VPWR sky130_fd_sc_hd__or4bb_1
X_5862_ _8978_/X VGND VPWR _5862_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_8650_ _8672_/C _8650_/B _8650_/C VGND VPWR _8722_/B VGND VPWR sky130_fd_sc_hd__or3_1
X_4813_ _9761_/Q VGND VPWR _4813_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_5793_ _9215_/Q _5791_/A _5964_/B1 _5791_/Y VGND VPWR _9215_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8581_ _8005_/A _8279_/C _8280_/B VGND VPWR _8582_/B VGND VPWR sky130_fd_sc_hd__o21ai_1
X_7601_ _6098_/Y _7455_/X _6062_/Y _7457_/X VGND VPWR _7601_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_21_325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4744_ _9390_/Q VGND VPWR _4744_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7532_ _8747_/A _7461_/X _8787_/A _7463_/X _7531_/X VGND VPWR _7535_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_119_257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_9202_ _9440_/CLK _9202_/D _4628_/A VGND VPWR _9202_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_7463_ _7463_/A VGND VPWR _7463_/X VGND VPWR sky130_fd_sc_hd__buf_8
X_4675_ _9364_/Q VGND VPWR _4675_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_7394_ _6429_/Y _7126_/X _6341_/Y _7128_/X VGND VPWR _7394_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_6414_ _6409_/Y _5442_/B _6410_/Y _5583_/B _6413_/X VGND VPWR _6433_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_127_290 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6345_ _6340_/Y _5259_/B _6341_/Y _5251_/B _6344_/X VGND VPWR _6352_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9133_ _9354_/CLK _9133_/D _9685_/SET_B VGND VPWR _9133_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6276_ _9377_/Q VGND VPWR _6276_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9064_ _4450_/A1 _9064_/D _6146_/A VGND VPWR _9064_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_102_124 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8015_ _7902_/B _8013_/B _8093_/A VGND VPWR _8016_/D VGND VPWR sky130_fd_sc_hd__a21oi_1
X_5227_ _5259_/A _5227_/B VGND VPWR _5230_/S VGND VPWR sky130_fd_sc_hd__or2_1
Xinput108 sram_ro_data[23] VGND VPWR _6100_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_102_168 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xinput119 sram_ro_data[4] VGND VPWR _6451_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_29_436 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5158_ _5158_/A VGND VPWR _5158_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_5089_ _5545_/A _5089_/B VGND VPWR _5090_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_8917_ _9609_/Q _8846_/X _8926_/S VGND VPWR _8917_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XPHY_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_103 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8848_ _9602_/Q _8916_/A1 _8926_/S VGND VPWR _8848_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_130 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_158 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_136 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_8779_ _8779_/A VGND VPWR _8780_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XPHY_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_347 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA_81 _7330_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_70 _6727_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_92 _9571_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_192_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_96 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_45 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_466 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_95 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_266 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_512 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_299 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_5 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_144 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_555 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_514 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4460_ _8946_/X VGND VPWR _4729_/A VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_116_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6130_ _6128_/Y _5872_/B _6129_/Y _5045_/B VGND VPWR _6130_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_112_411 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_306 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6061_ _9319_/Q VGND VPWR _6061_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_5012_ _9048_/Q _8957_/S _4949_/A _9696_/Q _5011_/X VGND VPWR _9696_/D VGND VPWR
+ sky130_fd_sc_hd__a32o_1
XFILLER_38_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9751_ _9755_/CLK _9751_/D _9757_/SET_B VGND VPWR _9751_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6963_ _6963_/A VGND VPWR _6964_/A VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_38_299 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_400 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5914_ _9126_/Q _5907_/A _8930_/A1 _5907_/Y VGND VPWR _9126_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8702_ _8732_/A _8735_/C VGND VPWR _8702_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
X_9682_ _9709_/CLK _9682_/D _5033_/X VGND VPWR _9682_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_6894_ _6889_/Y _5872_/B _6890_/Y _5776_/B _6893_/X VGND VPWR _6901_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_5845_ _9179_/Q _5839_/A _8955_/A1 _5839_/Y VGND VPWR _9179_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8633_ _8633_/A _8709_/C _8688_/C _8687_/C VGND VPWR _8633_/Y VGND VPWR sky130_fd_sc_hd__nor4_1
XFILLER_167_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_18 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_8564_ _8636_/A _8636_/B _8636_/C _8563_/X VGND VPWR _8564_/X VGND VPWR sky130_fd_sc_hd__or4b_1
X_5776_ _6052_/A _5776_/B VGND VPWR _5777_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_7515_ _6650_/Y _7475_/X _6633_/Y _7477_/X VGND VPWR _7515_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_8495_ _8341_/A _8498_/A _8189_/A _7885_/X VGND VPWR _8496_/B VGND VPWR sky130_fd_sc_hd__o22a_1
X_4727_ _4898_/A _4780_/B VGND VPWR _5660_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_7446_ _7456_/A _7472_/A _7474_/D VGND VPWR _7447_/A VGND VPWR sky130_fd_sc_hd__or3_1
X_4658_ _9091_/Q _9090_/Q _9092_/Q VGND VPWR _7003_/C VGND VPWR sky130_fd_sc_hd__or3_2
XFILLER_174_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput90 spimemio_flash_io2_oeb VGND VPWR input90/X VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_162_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9116_ _9779_/CLK _9116_/D _9779_/SET_B VGND VPWR _9116_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_4589_ _6158_/A _4903_/B VGND VPWR _4590_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_7377_ _6362_/Y _7077_/C _6440_/Y _7077_/D _7376_/X VGND VPWR _7377_/X VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_1_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_122 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_411 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6328_ _9402_/Q VGND VPWR _6328_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_130_230 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_99 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6259_ input8/X VGND VPWR _6259_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9047_ _9790_/CLK _9047_/D VGND VPWR _9047_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_190_49 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_200 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_188 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_43 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_247 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_383 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_612 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_116 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_119 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_311 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_344 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_274 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_342 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_420 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5630_ _9287_/Q _5623_/A _8840_/X _5623_/Y VGND VPWR _9287_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_5561_ _9335_/Q _5558_/A _8841_/X _5558_/Y VGND VPWR _9335_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_117_536 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5492_ _9383_/Q _5490_/A _5964_/B1 _5490_/Y VGND VPWR _9383_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8280_ _8275_/X _8280_/B _8280_/C VGND VPWR _8281_/B VGND VPWR sky130_fd_sc_hd__nand3b_1
X_7300_ _4718_/Y _7112_/X _4699_/Y _7077_/B VGND VPWR _7300_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4512_ _9772_/Q _4466_/A _5963_/B1 _4466_/Y VGND VPWR _9772_/D VGND VPWR sky130_fd_sc_hd__a22o_2
XFILLER_156_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_322 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7231_ _6301_/Y _7068_/A _6263_/Y _7105_/X VGND VPWR _7231_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_144_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4443_ _9588_/Q input80/X _8833_/S VGND VPWR _9009_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_7162_ _6736_/Y _7095_/X _6643_/Y _7068_/D _7161_/X VGND VPWR _7167_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_6113_ _9457_/Q VGND VPWR _6113_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7093_ _4740_/Y _7048_/B _4701_/Y _7077_/A _7092_/X VGND VPWR _7108_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_112_285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_414 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6044_ _6050_/A VGND VPWR _6045_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_85_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_19 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7995_ _8116_/B _7995_/B VGND VPWR _7996_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_54_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_567 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9734_ _9774_/CLK _9734_/D _9757_/SET_B VGND VPWR _9734_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6946_ _6946_/A _6946_/B _6946_/C VGND VPWR _6946_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
XFILLER_81_397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6877_ _6877_/A _6877_/B _6877_/C _6877_/D VGND VPWR _6878_/D VGND VPWR sky130_fd_sc_hd__and4_1
X_9665_ _4450_/A1 _9665_/D _6146_/A VGND VPWR _9665_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_5828_ _9190_/Q _5820_/A _8916_/A1 _5820_/Y VGND VPWR _9190_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8616_ _8735_/A _8616_/B _8668_/D _8699_/C VGND VPWR _8619_/A VGND VPWR sky130_fd_sc_hd__or4_2
X_9596_ _9596_/CLK _9596_/D _9528_/SET_B VGND VPWR _9596_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_5759_ _5759_/A VGND VPWR _5759_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_8547_ _8098_/A _8546_/Y _8398_/Y VGND VPWR _8547_/X VGND VPWR sky130_fd_sc_hd__o21a_1
X_8478_ _8703_/D _8478_/B VGND VPWR _8479_/B VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_123_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7429_ _7476_/A _9251_/Q _7470_/B _9255_/Q VGND VPWR _7430_/A VGND VPWR sky130_fd_sc_hd__or4_1
XFILLER_78_47 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_24 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_342 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_258 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_61 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_402 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_255 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_266 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_479 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput209 _8754_/X VGND VPWR mgmt_gpio_oeb[11] VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_141_325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_55 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_158 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_512 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_128 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_191 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6800_ _9115_/Q VGND VPWR _6800_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_36_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7780_ _8218_/B VGND VPWR _7969_/A VGND VPWR sky130_fd_sc_hd__inv_2
X_4992_ _8909_/X _9700_/Q _5001_/S VGND VPWR _4993_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_6731_ _9103_/Q VGND VPWR _6731_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_31_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9450_ _9483_/CLK _9450_/D _9528_/SET_B VGND VPWR _9450_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6662_ _9335_/Q VGND VPWR _6662_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_5613_ _9301_/Q _5612_/A _8846_/X _5612_/Y VGND VPWR _9301_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_9381_ _9771_/CLK _9381_/D _4628_/A VGND VPWR _9381_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_8401_ _8401_/A _8401_/B VGND VPWR _8401_/X VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_129_160 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_8332_ _8299_/A _8282_/C _8282_/B _8331_/X VGND VPWR _8333_/C VGND VPWR sky130_fd_sc_hd__a31o_1
X_6593_ _6593_/A VGND VPWR _6593_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_144_130 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5544_ _9346_/Q _5536_/A _8916_/A1 _5536_/Y VGND VPWR _9346_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_144_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5475_ _9394_/Q _5471_/A _8925_/A1 _5471_/Y VGND VPWR _9394_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8263_ _8263_/A _8369_/B VGND VPWR _8265_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_105_528 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8194_ _8204_/A VGND VPWR _8346_/B VGND VPWR sky130_fd_sc_hd__inv_2
X_7214_ _6346_/Y _7118_/X _6436_/Y _7048_/C VGND VPWR _7214_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_132_358 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7145_ _7145_/A _7145_/B _7145_/C _7145_/D VGND VPWR _7155_/B VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_113_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7076_ _7076_/A VGND VPWR _7077_/D VGND VPWR sky130_fd_sc_hd__buf_8
XFILLER_86_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6027_ _6052_/A _6027_/B VGND VPWR _6028_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_64_16 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_320 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7978_ _8096_/A _8098_/A VGND VPWR _7995_/B VGND VPWR sky130_fd_sc_hd__or2_1
X_6929_ _9102_/Q VGND VPWR _6929_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9717_ _9709_/CLK hold2/X _4639_/X VGND VPWR _9717_/Q VGND VPWR sky130_fd_sc_hd__dfrtn_1
Xclkbuf_leaf_31_csclk clkbuf_opt_2_0_csclk/X VGND VPWR _9379_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_81_194 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9648_ _9652_/CLK _9648_/D _9646_/SET_B VGND VPWR _9648_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_9579_ _9674_/CLK _9579_/D _9633_/SET_B VGND VPWR _9579_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_129_75 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_46_csclk _9329_/CLK VGND VPWR _9775_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_108_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_622 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_132 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0_wb_clk_i clkbuf_0_wb_clk_i/X VGND VPWR clkbuf_1_0_1_wb_clk_i/A VGND
+ VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_49_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_456 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_183 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_250 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5260_ _5260_/A VGND VPWR _5261_/A VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_141_144 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5191_ _9052_/Q _5985_/B _9586_/Q VGND VPWR _9586_/D VGND VPWR sky130_fd_sc_hd__a21o_1
XFILLER_83_415 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8950_ _9714_/Q _6475_/Y _8957_/S VGND VPWR _8950_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_7901_ _8472_/A _8517_/A VGND VPWR _7902_/B VGND VPWR sky130_fd_sc_hd__or2_1
X_8881_ _8880_/X _9141_/Q _9054_/Q VGND VPWR _8881_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_7832_ _7832_/A _7837_/B _7837_/C VGND VPWR _7833_/A VGND VPWR sky130_fd_sc_hd__or3_1
X_7763_ _8394_/A _8379_/B _7838_/B VGND VPWR _7764_/A VGND VPWR sky130_fd_sc_hd__or3_1
X_4975_ _4975_/A VGND VPWR _4975_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_9502_ _9527_/CLK _9502_/D _9528_/SET_B VGND VPWR _9502_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6714_ _6712_/Y _5374_/B _6713_/Y _5382_/B VGND VPWR _6714_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_7694_ _6434_/Y _7461_/X _6340_/Y _7463_/X _7693_/X VGND VPWR _7697_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9433_ _9440_/CLK _9433_/D _4628_/A VGND VPWR _9433_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_192_512 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6645_ _9242_/Q VGND VPWR _6645_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_192_556 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9364_ _9508_/CLK _9364_/D _9647_/SET_B VGND VPWR _9364_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6576_ _9531_/Q VGND VPWR _8779_/A VGND VPWR sky130_fd_sc_hd__clkinv_8
XFILLER_192_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9295_ _9371_/CLK _9295_/D _9295_/SET_B VGND VPWR _9295_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_8315_ _8238_/A _8498_/B _8304_/Y _8313_/X _8314_/X VGND VPWR _8318_/A VGND VPWR
+ sky130_fd_sc_hd__o2111ai_1
X_5527_ _5527_/A VGND VPWR _5528_/A VGND VPWR sky130_fd_sc_hd__clkbuf_2
X_8246_ _8341_/A _8246_/B VGND VPWR _8490_/B VGND VPWR sky130_fd_sc_hd__nor2_1
X_5458_ _5545_/A _5458_/B VGND VPWR _5459_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_8177_ _8720_/A _8560_/A _8177_/C VGND VPWR _8178_/B VGND VPWR sky130_fd_sc_hd__or3_1
X_5389_ _9453_/Q _5384_/A _8842_/X _5384_/Y VGND VPWR _9453_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7128_ _7128_/A VGND VPWR _7128_/X VGND VPWR sky130_fd_sc_hd__buf_8
XFILLER_101_553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7059_ _7059_/A _7059_/B _7059_/C _7059_/D VGND VPWR _7078_/B VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_15_526 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_36 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_306 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_570 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_202 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_472 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_73 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_420 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_426 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_160 _6027_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_182 _8801_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_171 _6929_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_193 _7021_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_60_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4760_ _4927_/A _4780_/B VGND VPWR _5610_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_4691_ _4919_/A _4843_/B VGND VPWR _5024_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_174_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6430_ _9074_/Q VGND VPWR _6430_/Y VGND VPWR sky130_fd_sc_hd__inv_4
XFILLER_127_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6361_ _9311_/Q VGND VPWR _6361_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_5312_ _9506_/Q _5308_/A _8925_/A1 _5308_/Y VGND VPWR _9506_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8100_ _8100_/A VGND VPWR _8213_/A VGND VPWR sky130_fd_sc_hd__buf_12
X_9080_ _9709_/CLK _9080_/D _6021_/X VGND VPWR _9080_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_6292_ _6292_/A VGND VPWR _6292_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_142_464 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5243_ _9553_/Q _5242_/A _8846_/X _5242_/Y VGND VPWR _9553_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8031_ _8097_/B _8550_/A _8030_/X VGND VPWR _8033_/A VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_142_497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5174_ _9597_/Q _5169_/A _8842_/X _5169_/Y VGND VPWR _9597_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8933_ _9085_/Q _9084_/Q _9051_/Q VGND VPWR _8933_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_8864_ _7626_/Y _9627_/Q _8978_/S VGND VPWR _8864_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XPHY_307 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_183 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_7815_ _7815_/A VGND VPWR _8097_/B VGND VPWR sky130_fd_sc_hd__buf_12
XPHY_329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_318 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_507 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_518 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8795_ _8795_/A VGND VPWR _8796_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_101_68 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_79 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4958_ _9091_/Q _6022_/C VGND VPWR _4958_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
X_7746_ _9066_/Q _7746_/B VGND VPWR _7746_/X VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_184_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7677_ _6549_/Y _7475_/X _6510_/Y _7477_/X VGND VPWR _7677_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4889_ _4911_/A _4900_/B VGND VPWR _5298_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_20_584 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_7 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9416_ _9684_/CLK _9416_/D _9685_/SET_B VGND VPWR _9416_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6628_ _6628_/A _6628_/B _6628_/C _6628_/D VGND VPWR _6629_/D VGND VPWR sky130_fd_sc_hd__and4_2
XFILLER_106_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_450 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9347_ _9352_/CLK _9347_/D _9646_/SET_B VGND VPWR _9347_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_192_397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6559_ _6557_/Y _5450_/B _6558_/Y _4841_/X VGND VPWR _6559_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_10_32 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_442 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_122 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9278_ _9278_/CLK _9278_/D _9633_/SET_B VGND VPWR _9278_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_126_43 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8229_ _8510_/A _8232_/B VGND VPWR _8658_/B VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_59_220 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_158 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_30 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_604 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_312 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_304 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_158 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_448 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_470 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5930_ _5930_/A _5930_/B input149/X input152/X VGND VPWR _5935_/B VGND VPWR sky130_fd_sc_hd__or4bb_1
X_7600_ _6122_/Y _7441_/X _6114_/Y _7443_/X _7599_/X VGND VPWR _7607_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_5861_ _5849_/X _8851_/X _8924_/X _9165_/Q VGND VPWR _9165_/D VGND VPWR sky130_fd_sc_hd__o22a_2
XFILLER_21_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5792_ _9216_/Q _5791_/A _5963_/B1 _5791_/Y VGND VPWR _9216_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_4812_ _4800_/Y _5290_/B _4804_/Y _5534_/B _4811_/X VGND VPWR _4830_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_8580_ _8580_/A _8675_/C _8645_/D _8716_/A VGND VPWR _8586_/A VGND VPWR sky130_fd_sc_hd__or4_4
X_7531_ _8751_/A _7465_/X _8789_/A _7467_/X VGND VPWR _7531_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4743_ _4876_/B _4780_/B VGND VPWR _5572_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_7462_ _7462_/A _7476_/C _7474_/D VGND VPWR _7463_/A VGND VPWR sky130_fd_sc_hd__or3_1
X_4674_ _4660_/Y _5556_/B _4664_/Y _5905_/B _4673_/X VGND VPWR _4705_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_6413_ _6411_/Y _4822_/X _6412_/Y _5232_/B VGND VPWR _6413_/X VGND VPWR sky130_fd_sc_hd__o22a_2
X_9201_ _9789_/CLK _9201_/D _4628_/A VGND VPWR _9201_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_7393_ _6391_/Y _5728_/X _6418_/Y _7040_/A _7392_/X VGND VPWR _7396_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_6344_ _6342_/Y _4613_/B _6343_/Y _5564_/B VGND VPWR _6344_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_9132_ _9379_/CLK _9132_/D _9779_/SET_B VGND VPWR _9132_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_0_208 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6275_ _9533_/Q VGND VPWR _6275_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9063_ _4450_/A1 _9063_/D _6146_/A VGND VPWR _9063_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_8014_ _8521_/A _8117_/A _8013_/X VGND VPWR _8016_/C VGND VPWR sky130_fd_sc_hd__o21ai_1
X_5226_ _9561_/Q _5218_/Y _8848_/X _5218_/A VGND VPWR _9561_/D VGND VPWR sky130_fd_sc_hd__o22a_1
Xinput109 sram_ro_data[24] VGND VPWR _4831_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_130_456 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5157_ _5157_/A VGND VPWR _5158_/A VGND VPWR sky130_fd_sc_hd__clkbuf_4
X_5088_ _5133_/A VGND VPWR _5545_/A VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_71_204 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8916_ _9610_/Q _8916_/A1 _8930_/S VGND VPWR _8916_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XPHY_115 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_104 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_8847_ _7022_/Y _9640_/Q _9587_/Q VGND VPWR _8847_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_52_440 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_148 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_175 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8778_ _8778_/A VGND VPWR _8778_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_12_359 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_159 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7729_ _7727_/Y _7726_/Y _9700_/Q VGND VPWR _7729_/Y VGND VPWR sky130_fd_sc_hd__a21oi_1
XFILLER_24_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_364 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_556 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA_93 _8831_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_82 _7482_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_60 _6280_/D VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_71 _6759_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_180_301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_478 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_30 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_587 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_524 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_6 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_167 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_71 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_323 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_526 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5658__14 _5651_/A VGND VPWR _5659_/B2 VGND VPWR sky130_fd_sc_hd__inv_2
X_6060_ _6060_/A VGND VPWR _8807_/B VGND VPWR sky130_fd_sc_hd__inv_4
XFILLER_112_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5011_ _6022_/B _7003_/C VGND VPWR _5011_/X VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_66_521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9750_ _9755_/CLK _9750_/D _9757_/SET_B VGND VPWR _9750_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6962_ _6974_/B _6962_/B VGND VPWR _6963_/A VGND VPWR sky130_fd_sc_hd__or2_2
XFILLER_179_412 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_440 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6893_ _6891_/Y _5679_/B _6892_/Y _5488_/B VGND VPWR _6893_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_5913_ _9127_/Q _5907_/A _8955_/A1 _5907_/Y VGND VPWR _9127_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8701_ _8064_/C _8700_/Y _8016_/C _8527_/C _8613_/B VGND VPWR _8735_/C VGND VPWR
+ sky130_fd_sc_hd__a2111o_2
X_9681_ _9681_/CLK _9681_/D _6146_/A VGND VPWR _9681_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_179_456 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5844_ _9180_/Q _5839_/A _8929_/A1 _5839_/Y VGND VPWR _9180_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8632_ _8632_/A _8632_/B VGND VPWR _8687_/C VGND VPWR sky130_fd_sc_hd__nor2_1
X_8563_ _8563_/A _8713_/D _8713_/B _8636_/D VGND VPWR _8563_/X VGND VPWR sky130_fd_sc_hd__or4_1
XFILLER_166_117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5775_ _9226_/Q _5770_/A _5967_/B1 _5770_/Y VGND VPWR _9226_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7514_ _6687_/Y _7461_/X _6735_/Y _7463_/X _7513_/X VGND VPWR _7517_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_159_191 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8494_ _8515_/B _8305_/A _8660_/A _8496_/A _8341_/B VGND VPWR _8594_/A VGND VPWR
+ sky130_fd_sc_hd__a311oi_2
X_4726_ _9269_/Q VGND VPWR _4726_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_135_537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7445_ _7445_/A VGND VPWR _7445_/X VGND VPWR sky130_fd_sc_hd__buf_8
X_4657_ _4657_/A VGND VPWR _4657_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_162_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7376_ _6348_/Y _7086_/X _6409_/Y _7088_/X VGND VPWR _7376_/X VGND VPWR sky130_fd_sc_hd__o22a_1
Xinput80 spi_sck VGND VPWR input80/X VGND VPWR sky130_fd_sc_hd__buf_6
Xinput91 spimemio_flash_io3_do VGND VPWR input91/X VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_162_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_12 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6327_ _6149_/A _6326_/Y _9041_/Q _6149_/Y VGND VPWR _9041_/D VGND VPWR sky130_fd_sc_hd__o22a_1
X_4588_ _4669_/A _4729_/D _8946_/X _4729_/B VGND VPWR _4903_/B VGND VPWR sky130_fd_sc_hd__or4_4
X_9115_ _9129_/CLK _9115_/D _9779_/SET_B VGND VPWR _9115_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_130_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_134 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6258_ _9737_/Q VGND VPWR _6258_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9046_ _9790_/CLK _9046_/D VGND VPWR _9046_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_29_212 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6189_ _9784_/Q VGND VPWR _6189_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_5209_ _9572_/Q _5203_/Y _8905_/X _5203_/A VGND VPWR _9572_/D VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_29_267 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_410 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_470 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_344 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_543 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_82 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_432 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5560_ _9336_/Q _5558_/A _8842_/X _5558_/Y VGND VPWR _9336_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_156_161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5491_ _9384_/Q _5490_/A _5963_/B1 _5490_/Y VGND VPWR _9384_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_4511_ _9773_/Q _4506_/A _5967_/B1 _4506_/Y VGND VPWR _9773_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_144_334 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_548 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7230_ _6296_/Y _7059_/B _6310_/Y _7068_/C _7229_/X VGND VPWR _7233_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_7_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7161_ _6760_/Y _7097_/X _6735_/Y _7099_/X VGND VPWR _7161_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_7092_ _4773_/Y _7040_/C _4664_/Y _7059_/C VGND VPWR _7092_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_6112_ _6109_/Y _5267_/B _6110_/Y _5306_/B _6111_/X VGND VPWR _6119_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_140_584 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6043_ _6043_/A VGND VPWR _6043_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_85_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7994_ _7994_/A _7994_/B VGND VPWR _8116_/B VGND VPWR sky130_fd_sc_hd__nand2_4
X_9733_ _9774_/CLK _9733_/D _9757_/SET_B VGND VPWR _9733_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6945_ _6945_/A _6945_/B _6945_/C VGND VPWR _6946_/C VGND VPWR sky130_fd_sc_hd__and3_2
XFILLER_54_579 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_2_2_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A VGND VPWR clkbuf_3_5_0_wb_clk_i/A VGND
+ VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_22_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6876_ _6871_/Y _5458_/B _6872_/Y _5480_/B _6875_/X VGND VPWR _6877_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9664_ _9664_/CLK _9664_/D _6146_/A VGND VPWR _9664_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_5827_ _9191_/Q _5820_/A _8930_/A1 _5820_/Y VGND VPWR _9191_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8615_ _8615_/A _8615_/B _8615_/C _8615_/D VGND VPWR _8699_/C VGND VPWR sky130_fd_sc_hd__or4_1
X_9595_ _9596_/CLK _9595_/D _9528_/SET_B VGND VPWR _9595_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_8546_ _8546_/A _8566_/B VGND VPWR _8546_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
X_5758_ _5758_/A VGND VPWR _5759_/A VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_135_301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4709_ _4929_/A _4780_/B VGND VPWR _5776_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_8477_ _8477_/A _8721_/C VGND VPWR _8478_/B VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_175_481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_492 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7428_ _4816_/Y _7427_/X _4742_/Y _5699_/X VGND VPWR _7428_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_5689_ _9256_/Q _5681_/A _8916_/A1 _5681_/Y VGND VPWR _9256_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_162_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7359_ _6604_/Y _7097_/X _6550_/Y _7099_/X VGND VPWR _7359_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_78_59 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_104 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9029_ _9039_/CLK _9029_/D VGND VPWR _9029_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_1_369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_354 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_75 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_415 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_67 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_524 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4991_ _4991_/A _8957_/X VGND VPWR _5001_/S VGND VPWR sky130_fd_sc_hd__or2b_1
X_6730_ _9512_/Q VGND VPWR _6730_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_189_551 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6661_ _9322_/Q VGND VPWR _6661_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_6592_ input6/X VGND VPWR _6592_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_8400_ _8521_/A _8117_/A _8393_/Y _8401_/B _8399_/X VGND VPWR _8400_/X VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9380_ _9380_/CLK _9380_/D _4628_/A VGND VPWR _9380_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_5612_ _5612_/A VGND VPWR _5612_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_5543_ _9347_/Q _5536_/A _8930_/A1 _5536_/Y VGND VPWR _9347_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8331_ _8331_/A _8331_/B VGND VPWR _8331_/X VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_129_183 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5474_ _9395_/Q _5471_/A _8844_/X _5471_/Y VGND VPWR _9395_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8262_ _8341_/A _8262_/B VGND VPWR _8369_/B VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_144_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7213_ _6457_/Y _7040_/D _6398_/Y _7110_/X _7212_/X VGND VPWR _7220_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_8193_ _8193_/A _8193_/B _8195_/A VGND VPWR _8204_/A VGND VPWR sky130_fd_sc_hd__or3_2
X_7144_ _6879_/Y _7048_/D _6908_/Y _7040_/B _7143_/X VGND VPWR _7145_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_48_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_18 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_7075_ _7075_/A _7123_/B VGND VPWR _7076_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_39_351 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6026_ _9078_/Q _4466_/A _8955_/A1 _4466_/Y VGND VPWR _9078_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_104_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_332 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7977_ _8091_/B _7988_/A VGND VPWR _8096_/A VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_154_7 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9716_ _9089_/CLK _9716_/D _4642_/X VGND VPWR hold1/A VGND VPWR sky130_fd_sc_hd__dfrtn_1
X_6928_ _9265_/Q VGND VPWR _6928_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_6859_ _9373_/Q VGND VPWR _6859_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9647_ _9652_/CLK _9647_/D _9647_/SET_B VGND VPWR _9647_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_10_413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_571 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_9578_ _9674_/CLK _9578_/D _9633_/SET_B VGND VPWR _9578_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_8529_ _8523_/Y _8528_/Y _8518_/X _8455_/B VGND VPWR _8734_/D VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_135_142 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_356 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_107 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_50 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_262 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_3_0_mgmt_gpio_in[4] clkbuf_2_3_0_mgmt_gpio_in[4]/A VGND VPWR _4446_/A1 VGND
+ VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_173_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5190_ _5190_/A VGND VPWR _5190_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_83_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7900_ _7900_/A _8528_/B VGND VPWR _8517_/A VGND VPWR sky130_fd_sc_hd__or2b_2
X_8880_ _7221_/Y _9636_/Q _8959_/S VGND VPWR _8880_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_91_471 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7831_ _8324_/A VGND VPWR _7831_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_36_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7762_ _8379_/D VGND VPWR _8394_/A VGND VPWR sky130_fd_sc_hd__clkinv_4
X_4974_ _4994_/A VGND VPWR _4975_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_6713_ _9452_/Q VGND VPWR _6713_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7693_ _6369_/Y _7465_/X _6397_/Y _7467_/X VGND VPWR _7693_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_9501_ _9501_/CLK _9501_/D _9647_/SET_B VGND VPWR _9501_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6644_ _9192_/Q VGND VPWR _6644_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9432_ _9440_/CLK _9432_/D _4628_/A VGND VPWR _9432_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_109_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_19 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9363_ _9771_/CLK _9363_/D _4628_/A VGND VPWR _9363_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6575_ _9375_/Q VGND VPWR _8767_/A VGND VPWR sky130_fd_sc_hd__clkinv_8
XFILLER_192_579 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_568 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9294_ _9371_/CLK _9294_/D _9295_/SET_B VGND VPWR _9294_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_8314_ _8316_/A _8264_/B _8454_/A VGND VPWR _8314_/X VGND VPWR sky130_fd_sc_hd__o21a_1
X_5526_ _5671_/A _5526_/B VGND VPWR _5527_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_145_484 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_8245_ _8245_/A _8362_/B _8575_/B VGND VPWR _8248_/A VGND VPWR sky130_fd_sc_hd__or3_1
X_5457_ _9406_/Q _5452_/A _5967_/B1 _5452_/Y VGND VPWR _9406_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_105_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_318 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_582 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5388_ _9454_/Q _5384_/A _8925_/A1 _5384_/Y VGND VPWR _9454_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8176_ _8521_/A _8515_/A _8175_/Y VGND VPWR _8177_/C VGND VPWR sky130_fd_sc_hd__o21bai_1
X_7127_ _7127_/A _7127_/B _7127_/C VGND VPWR _7128_/A VGND VPWR sky130_fd_sc_hd__or3_1
X_7058_ _7058_/A VGND VPWR _7059_/D VGND VPWR sky130_fd_sc_hd__buf_8
XFILLER_47_608 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_587 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6009_ _6040_/A VGND VPWR _6010_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_15_549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_48 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_232 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_568 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_443 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_438 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_471 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_151 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_302 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_110 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_150 _5259_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_161 _6251_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_183 _8801_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_172 _7343_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_194 _7021_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_159_554 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4690_ _9683_/Q VGND VPWR _4692_/A VGND VPWR sky130_fd_sc_hd__clkinv_4
XFILLER_174_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6360_ _9324_/Q VGND VPWR _6360_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
XFILLER_127_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5311_ _9507_/Q _5308_/A _8844_/X _5308_/Y VGND VPWR _9507_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_114_134 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8030_ _8389_/A _8550_/A _8027_/X _8410_/A _8029_/X VGND VPWR _8030_/X VGND VPWR
+ sky130_fd_sc_hd__o2111a_1
X_6291_ _9075_/Q VGND VPWR _6291_/Y VGND VPWR sky130_fd_sc_hd__inv_6
X_5242_ _5242_/A VGND VPWR _5242_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_5173_ _9598_/Q _5169_/A _8925_/A1 _5169_/Y VGND VPWR _9598_/D VGND VPWR sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_30_csclk clkbuf_2_1_0_csclk/X VGND VPWR _9129_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_96_596 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xinput1 debug_mode VGND VPWR input1/X VGND VPWR sky130_fd_sc_hd__buf_4
X_8932_ _8931_/X _9677_/Q _9587_/Q VGND VPWR _8932_/X VGND VPWR sky130_fd_sc_hd__mux2_4
Xclkbuf_leaf_45_csclk _9329_/CLK VGND VPWR _9777_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
X_8863_ _8862_/X _9170_/Q _9054_/Q VGND VPWR _8863_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_52_622 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_7814_ _8379_/C _7839_/A _8394_/A _8394_/B VGND VPWR _7815_/A VGND VPWR sky130_fd_sc_hd__or4_1
XPHY_319 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_308 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_368 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8794_ _8794_/A VGND VPWR _8794_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_7745_ _9068_/Q _7745_/A2 _9067_/Q _7745_/B2 _7744_/X VGND VPWR _7745_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_4957_ _4957_/A VGND VPWR _4957_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_4888_ _9510_/Q VGND VPWR _4888_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7676_ _6486_/Y _7461_/X _6550_/Y _7463_/X _7675_/X VGND VPWR _7679_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_137_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6627_ _6627_/A _6627_/B _6627_/C _6627_/D VGND VPWR _6628_/D VGND VPWR sky130_fd_sc_hd__and4_1
X_9415_ _9514_/CLK _9415_/D _4628_/A VGND VPWR _9415_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_192_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_7 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9346_ _9352_/CLK _9346_/D _9646_/SET_B VGND VPWR _9346_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6558_ _6558_/A VGND VPWR _6558_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_5509_ _5509_/A VGND VPWR _5509_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_145_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9277_ _9278_/CLK _9277_/D _9757_/SET_B VGND VPWR _9277_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_6489_ _9393_/Q VGND VPWR _8797_/A VGND VPWR sky130_fd_sc_hd__inv_4
XFILLER_126_55 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8228_ _8230_/A _8264_/B VGND VPWR _8676_/B VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_86_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8159_ _8554_/A _8640_/B VGND VPWR _8645_/A VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_101_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_42 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_140 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_30 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_324 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_616 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_316 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_395 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_40 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_596 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_126 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_104 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_235 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_544 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_460 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5860_ _5849_/X _8853_/X _8924_/X _9166_/Q VGND VPWR _9166_/D VGND VPWR sky130_fd_sc_hd__o22a_2
XFILLER_92_80 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4811_ _4931_/A _6158_/A _4808_/Y _4809_/Y _5251_/B VGND VPWR _4811_/X VGND VPWR
+ sky130_fd_sc_hd__o32a_1
X_5791_ _5791_/A VGND VPWR _5791_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_21_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4742_ _9320_/Q VGND VPWR _4742_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_178_159 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7530_ _8749_/A _7451_/X _8773_/A _7453_/X _7529_/X VGND VPWR _7535_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_4673_ _4668_/Y _5872_/B _4671_/Y _5526_/B VGND VPWR _4673_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_7461_ _7461_/A VGND VPWR _7461_/X VGND VPWR sky130_fd_sc_hd__buf_8
X_6412_ _9558_/Q VGND VPWR _6412_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9200_ _9789_/CLK _9200_/D _4628_/A VGND VPWR _9200_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_174_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_218 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7392_ _7392_/A _7392_/B VGND VPWR _7392_/X VGND VPWR sky130_fd_sc_hd__or2_1
Xclkbuf_opt_5_0_csclk clkbuf_2_2_0_csclk/X VGND VPWR clkbuf_leaf_6_csclk/A VGND VPWR
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_127_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6343_ _9332_/Q VGND VPWR _6343_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9131_ _9379_/CLK _9131_/D _9779_/SET_B VGND VPWR _9131_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_88_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_476 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9062_ _4450_/A1 _9062_/D _6146_/A VGND VPWR _9062_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6274_ _9455_/Q VGND VPWR _6274_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
X_5225_ _9562_/Q _5218_/Y _8919_/X _5218_/A VGND VPWR _9562_/D VGND VPWR sky130_fd_sc_hd__o22a_1
X_8013_ _8097_/B _8013_/B VGND VPWR _8013_/X VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_130_446 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5156_ _6135_/A _5156_/B VGND VPWR _5157_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_84_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5087_ _9654_/Q _5082_/A _5967_/B1 _5082_/Y VGND VPWR _9654_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8915_ _9623_/Q _8844_/X _8955_/S VGND VPWR _8915_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_71_216 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_116 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_8846_ _9707_/Q _9666_/Q _9587_/Q VGND VPWR _8846_/X VGND VPWR sky130_fd_sc_hd__mux2_8
XPHY_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_127 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_463 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5989_ _6022_/C _5985_/B _5985_/Y VGND VPWR _9090_/D VGND VPWR sky130_fd_sc_hd__a21oi_1
X_8777_ _8777_/A VGND VPWR _8778_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_24_187 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7728_ _7727_/Y _7726_/Y _9699_/Q _9698_/Q VGND VPWR _7728_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_177_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_50 _6119_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_7659_ _6652_/Y _7475_/X _6634_/Y _7477_/X VGND VPWR _7659_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XANTENNA_83 _7649_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_72 _6784_/D VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_61 _6291_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_165_376 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_94 _8824_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_106_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9329_ _9329_/CLK _9329_/D _4628_/A VGND VPWR _9329_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_97_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_599 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_62 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_7 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_154 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_107 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_124 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_179 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_331 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_78 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_3_4_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/A VGND VPWR _9027_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_97_146 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5010_ _5010_/A VGND VPWR _5010_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_85_319 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_330 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6961_ _9062_/Q VGND VPWR _6962_/B VGND VPWR sky130_fd_sc_hd__inv_2
X_8700_ _8515_/B _8305_/A _8341_/B VGND VPWR _8700_/Y VGND VPWR sky130_fd_sc_hd__a21oi_1
X_5912_ _9128_/Q _5907_/A _8929_/A1 _5907_/Y VGND VPWR _9128_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_9680_ _9681_/CLK _9680_/D _6146_/A VGND VPWR _9680_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6892_ _9381_/Q VGND VPWR _6892_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_53_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_424 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5843_ _9181_/Q _5839_/A _8925_/A1 _5839_/Y VGND VPWR _9181_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8631_ _8631_/A _8631_/B VGND VPWR _8688_/C VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_21_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_468 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8562_ _8562_/A _8672_/C _8673_/A VGND VPWR _8636_/D VGND VPWR sky130_fd_sc_hd__or3_1
X_5774_ _9227_/Q _5770_/A _5966_/B1 _5770_/Y VGND VPWR _9227_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7513_ _6637_/Y _7465_/X _6717_/Y _7467_/X VGND VPWR _7513_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_8493_ _8614_/A _8493_/B _8493_/C VGND VPWR _8657_/C VGND VPWR sky130_fd_sc_hd__or3_1
X_4725_ _4716_/Y _5837_/B _4718_/Y _5594_/B _4724_/X VGND VPWR _4791_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_107_218 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7444_ _7462_/A _7470_/B _7474_/D VGND VPWR _7445_/A VGND VPWR sky130_fd_sc_hd__or3_1
X_4656_ _4994_/A VGND VPWR _4657_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_4587_ _9740_/Q _4579_/A _5967_/B1 _4579_/Y VGND VPWR _9740_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7375_ _7375_/A _7375_/B _7375_/C VGND VPWR _7375_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
Xinput81 spi_sdo VGND VPWR input81/X VGND VPWR sky130_fd_sc_hd__buf_6
Xinput70 mgmt_gpio_in[7] VGND VPWR _6060_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_162_357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6326_ _6326_/A _6326_/B _6326_/C _6326_/D VGND VPWR _6326_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
X_9114_ _9779_/CLK _9114_/D _9779_/SET_B VGND VPWR _9114_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
Xinput92 spimemio_flash_io3_oeb VGND VPWR input92/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_130_210 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_24 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6257_ _6257_/A VGND VPWR _6257_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9045_ _9790_/CLK _9045_/D VGND VPWR _9045_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_130_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5208_ _9573_/Q _5203_/Y _8929_/X _5203_/A VGND VPWR _9573_/D VGND VPWR sky130_fd_sc_hd__o22a_1
X_6188_ _9076_/Q VGND VPWR _6188_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
XFILLER_69_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5139_ _9623_/Q _5136_/A _8844_/X _5136_/Y VGND VPWR _9623_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_57_555 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8829_ _9592_/Q input89/X _8835_/S VGND VPWR _8829_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_185_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_146 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_611 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_590 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_508 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_560 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_124 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_63 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_96 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_584 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_555 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_452 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_444 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_460 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_150 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_302 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5490_ _5490_/A VGND VPWR _5490_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_4510_ _9774_/Q _4506_/A _5966_/B1 _4506_/Y VGND VPWR _9774_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_156_173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_346 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7160_ _6644_/Y _7048_/B _6681_/Y _7077_/A _7159_/X VGND VPWR _7167_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_6111_ _6111_/A _6111_/B _9769_/Q VGND VPWR _6111_/X VGND VPWR sky130_fd_sc_hd__or3b_4
XFILLER_112_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7091_ _4855_/Y _7082_/X _4850_/Y _7084_/X _7090_/X VGND VPWR _7132_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_98_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6042_ _6050_/A VGND VPWR _6043_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_85_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7993_ _7993_/A VGND VPWR _8137_/B VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_81_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_355 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9732_ _9774_/CLK _9732_/D _9757_/SET_B VGND VPWR _9732_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6944_ _6944_/A _6944_/B _6944_/C VGND VPWR _6945_/C VGND VPWR sky130_fd_sc_hd__and3_1
X_9663_ _9664_/CLK _9663_/D _6146_/A VGND VPWR _9663_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_167_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_271 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6875_ _6873_/Y _5404_/B _6874_/Y _5290_/B VGND VPWR _6875_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_8614_ _8614_/A _8614_/B _8614_/C _8614_/D VGND VPWR _8668_/D VGND VPWR sky130_fd_sc_hd__or4_1
XFILLER_22_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5826_ _9192_/Q _5820_/A _8955_/A1 _5820_/Y VGND VPWR _9192_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_9594_ _9596_/CLK _9594_/D _9528_/SET_B VGND VPWR _9594_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_5757_ _6052_/A _5757_/B VGND VPWR _5758_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_8545_ _8625_/B VGND VPWR _8554_/B VGND VPWR sky130_fd_sc_hd__clkinv_4
X_4708_ _9218_/Q VGND VPWR _4708_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_8476_ _8476_/A _8476_/B VGND VPWR _8721_/C VGND VPWR sky130_fd_sc_hd__or2_2
XFILLER_135_313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5688_ _9257_/Q _5681_/A _8840_/X _5681_/Y VGND VPWR _9257_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7427_ _7427_/A VGND VPWR _7427_/X VGND VPWR sky130_fd_sc_hd__buf_8
X_4639_ _4639_/A VGND VPWR _4639_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_78_38 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7358_ _6504_/Y _7048_/B _6539_/Y _7077_/A _7357_/X VGND VPWR _7365_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_2
XFILLER_89_400 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6309_ _9261_/Q VGND VPWR _6309_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_131_552 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7289_ _4731_/A _7077_/C _4671_/Y _7077_/D _7288_/X VGND VPWR _7289_/X VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_76_116 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9028_ _9039_/CLK _9028_/D VGND VPWR _9028_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_77_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_55 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_190 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_539 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_271 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_95 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_186 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_79 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_92 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4990_ _7008_/A _5992_/B _4966_/A _6022_/B _4989_/X VGND VPWR _4991_/A VGND VPWR
+ sky130_fd_sc_hd__o32a_1
XFILLER_149_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6660_ _6656_/Y _4524_/B _6657_/Y _5412_/B _6659_/X VGND VPWR _6691_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_6591_ _9751_/Q VGND VPWR _6591_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_5611_ _5611_/A VGND VPWR _5612_/A VGND VPWR sky130_fd_sc_hd__clkbuf_4
X_5542_ _9348_/Q _5536_/A _8955_/A1 _5536_/Y VGND VPWR _9348_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8330_ _8376_/A _8330_/B VGND VPWR _8331_/B VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_129_195 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5473_ _9396_/Q _5471_/A _8845_/X _5471_/Y VGND VPWR _9396_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8261_ _8261_/A _8578_/B VGND VPWR _8263_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_7212_ _6360_/Y _7112_/X _6468_/Y _7077_/B VGND VPWR _7212_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_8192_ _8195_/A _8193_/B _8193_/A VGND VPWR _8346_/A VGND VPWR sky130_fd_sc_hd__o21a_1
X_7143_ _6890_/Y _7068_/A _6860_/Y _7105_/X VGND VPWR _7143_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_140_360 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7074_ _7074_/A VGND VPWR _7077_/C VGND VPWR sky130_fd_sc_hd__buf_8
XFILLER_113_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6025_ _9079_/Q _4466_/A _8844_/X _4466_/Y VGND VPWR _9079_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_39_374 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7976_ _8583_/A _7966_/B _8195_/B VGND VPWR _7988_/A VGND VPWR sky130_fd_sc_hd__a21bo_1
X_9715_ _9089_/CLK _9715_/D _4645_/X VGND VPWR _9715_/Q VGND VPWR sky130_fd_sc_hd__dfrtn_1
X_6927_ _9241_/Q VGND VPWR _6927_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9646_ _9652_/CLK _9646_/D _9646_/SET_B VGND VPWR _9646_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6858_ _6853_/Y _5382_/B _6854_/Y _5306_/B _6857_/X VGND VPWR _6877_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_2
X_5809_ _9053_/Q _9791_/Q _5643_/Y _5808_/X VGND VPWR _9203_/D VGND VPWR sky130_fd_sc_hd__a31o_1
X_9577_ _9788_/CLK _9577_/D _9295_/SET_B VGND VPWR _9577_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6789_ _9727_/Q VGND VPWR _6789_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_8528_ _8528_/A _8528_/B VGND VPWR _8528_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
X_8459_ _8459_/A _8734_/C _8459_/C _8614_/C VGND VPWR _8464_/A VGND VPWR sky130_fd_sc_hd__or4_1
XFILLER_131_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_620 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_439 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_119 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_274 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_316 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_92 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7830_ _7903_/C _8528_/A _8583_/A _8189_/A VGND VPWR _8324_/A VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_91_483 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_539 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4973_ _9705_/Q _4966_/A _9704_/Q _4966_/Y VGND VPWR _9705_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7761_ _8299_/A _8282_/C _7836_/A VGND VPWR _8636_/A VGND VPWR sky130_fd_sc_hd__and3_2
X_6712_ _9460_/Q VGND VPWR _6712_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_149_213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7692_ _6467_/Y _7451_/X _6348_/Y _7453_/X _7691_/X VGND VPWR _7697_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9500_ _9501_/CLK _9500_/D _9647_/SET_B VGND VPWR _9500_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_32_583 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_9431_ _9508_/CLK _9431_/D _9295_/SET_B VGND VPWR _9431_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6643_ _9233_/Q VGND VPWR _6643_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_6574_ _9513_/Q VGND VPWR _6574_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9362_ _9514_/CLK _9362_/D _4628_/A VGND VPWR _9362_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_145_441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5525_ _9359_/Q _5520_/A _5967_/B1 _5520_/Y VGND VPWR _9359_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8313_ _8496_/A _8306_/X _8230_/A _8498_/B _8312_/X VGND VPWR _8313_/X VGND VPWR
+ sky130_fd_sc_hd__o221a_2
X_9293_ _9596_/CLK _9293_/D _9528_/SET_B VGND VPWR _9293_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_105_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_411 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5456_ _9407_/Q _5452_/A _5966_/B1 _5452_/Y VGND VPWR _9407_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8244_ _8316_/A _8260_/B VGND VPWR _8575_/B VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_105_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_496 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5387_ _9455_/Q _5384_/A _8844_/X _5384_/Y VGND VPWR _9455_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8175_ _8175_/A _8175_/B VGND VPWR _8175_/Y VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_101_500 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_594 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_382 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7126_ _7126_/A VGND VPWR _7126_/X VGND VPWR sky130_fd_sc_hd__buf_8
XFILLER_140_190 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7057_ _7073_/C _7087_/B VGND VPWR _7058_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_74_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_599 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6008_ _9085_/Q _5995_/A _8910_/X _5995_/Y VGND VPWR _9085_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_54_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7959_ _7959_/A _8583_/A _7966_/B VGND VPWR _8193_/B VGND VPWR sky130_fd_sc_hd__or3_2
XFILLER_24_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_9629_ _9757_/CLK _9629_/D _9757_/SET_B VGND VPWR _9629_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_10_244 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_222 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_226 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_400 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_271 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_360 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_14 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_163 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_483 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_122 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_314 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_151 _4590_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_140 _7199_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_162 _6264_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_184 input2/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_173 _7343_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_195 _7021_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_5310_ _9508_/Q _5308_/A _8845_/X _5308_/Y VGND VPWR _9508_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_6290_ _9481_/Q VGND VPWR _6290_/Y VGND VPWR sky130_fd_sc_hd__inv_6
XFILLER_5_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5241_ _5241_/A VGND VPWR _5242_/A VGND VPWR sky130_fd_sc_hd__clkbuf_4
X_5172_ _9599_/Q _5169_/A _8844_/X _5169_/Y VGND VPWR _9599_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_96_553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_190 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_406 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_8931_ _9084_/Q _9083_/Q _9051_/Q VGND VPWR _8931_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xinput2 debug_oeb VGND VPWR input2/X VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_83_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_opt_1_0_csclk _9329_/CLK VGND VPWR clkbuf_leaf_2_csclk/A VGND VPWR sky130_fd_sc_hd__clkbuf_16
X_8862_ _7608_/Y _9639_/Q _8978_/S VGND VPWR _8862_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_7813_ _7813_/A VGND VPWR _8341_/A VGND VPWR sky130_fd_sc_hd__clkbuf_16
X_8793_ _8793_/A VGND VPWR _8794_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XPHY_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_7744_ _9066_/Q _7744_/B VGND VPWR _7744_/X VGND VPWR sky130_fd_sc_hd__and2_1
X_4956_ _4994_/A VGND VPWR _4957_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_4887_ _9732_/Q VGND VPWR _4887_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7675_ _6498_/Y _7465_/X _6574_/Y _7467_/X VGND VPWR _7675_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_6626_ _6621_/Y _4524_/B _8787_/A _5278_/B _6625_/X VGND VPWR _6627_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9414_ _9514_/CLK _9414_/D _9685_/SET_B VGND VPWR _9414_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_192_344 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6557_ _9409_/Q VGND VPWR _6557_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9345_ _9371_/CLK _9345_/D _9295_/SET_B VGND VPWR _9345_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_192_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5508_ _5508_/A VGND VPWR _5509_/A VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_105_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6488_ _8761_/A _5610_/B _6484_/Y _5594_/B _6487_/X VGND VPWR _6501_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9276_ _9596_/CLK _9276_/D _9528_/SET_B VGND VPWR _9276_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_160_241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_466 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5439_ _9418_/Q _5433_/A _8841_/X _5433_/Y VGND VPWR _9418_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8227_ _8595_/B _8227_/B _8571_/B _8499_/B VGND VPWR _8231_/A VGND VPWR sky130_fd_sc_hd__or4_1
Xoutput350 _9042_/Q VGND VPWR wb_dat_o[30] VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_126_67 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_8158_ _8158_/A _8630_/B VGND VPWR _8160_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_7109_ _7127_/C _7109_/B VGND VPWR _7110_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_19_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_8089_ _8218_/B _7837_/A _8102_/B VGND VPWR _8120_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_101_385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_152 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_494 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_42 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_352 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_52 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_96 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_474 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_203 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_247 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4810_ _4891_/A _4931_/B VGND VPWR _5251_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_21_306 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_155 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5790_ _5790_/A VGND VPWR _5791_/A VGND VPWR sky130_fd_sc_hd__clkbuf_2
X_4741_ _4805_/A _4780_/B VGND VPWR _5818_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_119_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_300 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7460_ _7462_/A _7474_/C _9255_/Q VGND VPWR _7461_/A VGND VPWR sky130_fd_sc_hd__or3_1
X_4672_ _4919_/A _4787_/A VGND VPWR _5526_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_6411_ _6411_/A VGND VPWR _6411_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_7391_ _6458_/Y _7059_/D _6424_/Y _7116_/X _7390_/X VGND VPWR _7396_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9130_ _9379_/CLK _9130_/D _9779_/SET_B VGND VPWR _9130_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_155_591 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6342_ _9725_/Q VGND VPWR _6342_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_170_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6273_ _6268_/Y _4524_/B _6269_/Y _5458_/B _6272_/X VGND VPWR _6280_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9061_ _4450_/A1 _9061_/D _6146_/A VGND VPWR _9061_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_5224_ _9563_/Q _5218_/Y _8922_/X _5218_/A VGND VPWR _9563_/D VGND VPWR sky130_fd_sc_hd__o22a_1
X_8012_ _8523_/A _8517_/A VGND VPWR _8013_/B VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_69_575 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5155_ _9610_/Q _5147_/A _8916_/A1 _5147_/Y VGND VPWR _9610_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_5086_ _9655_/Q _5082_/A _8930_/A1 _5082_/Y VGND VPWR _9655_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_37_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8914_ _9625_/Q _8846_/X _8955_/S VGND VPWR _8914_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_56_269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_239 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8845_ _9706_/Q _9665_/Q _9587_/Q VGND VPWR _8845_/X VGND VPWR sky130_fd_sc_hd__mux2_8
XPHY_106 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_139 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5988_ _5988_/A VGND VPWR _5988_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_8776_ _8776_/A VGND VPWR _8776_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_7727_ _9699_/Q VGND VPWR _7727_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_4939_ _4939_/A VGND VPWR _4939_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_7658_ _6674_/Y _7461_/X _6711_/Y _7463_/X _7657_/X VGND VPWR _7661_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XANTENNA_40 _5968_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_21_11 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6609_ _9544_/Q VGND VPWR _6609_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XANTENNA_62 _6291_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_73 _6784_/D VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_51 _6107_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_84 _8375_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_165_388 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7589_ _7589_/A _7589_/B _7589_/C _7589_/D VGND VPWR _7590_/D VGND VPWR sky130_fd_sc_hd__and4_1
XANTENNA_95 _7019_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_4_527 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9328_ _9380_/CLK _9328_/D _4628_/A VGND VPWR _9328_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_97_37 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9259_ _9601_/CLK _9259_/D _9295_/SET_B VGND VPWR _9259_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_106_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_494 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_74 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_8 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_44_csclk _9329_/CLK VGND VPWR _9755_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_100_609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6960_ _4936_/Y _6952_/A _9028_/Q _6952_/Y VGND VPWR _9028_/D VGND VPWR sky130_fd_sc_hd__o22a_1
X_5911_ _9129_/Q _5907_/A _8925_/A1 _5907_/Y VGND VPWR _9129_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_6891_ _9257_/Q VGND VPWR _6891_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
XFILLER_61_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5842_ _9182_/Q _5839_/A _8844_/X _5839_/Y VGND VPWR _9182_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8630_ _8630_/A _8630_/B _8630_/C _8630_/D VGND VPWR _8709_/C VGND VPWR sky130_fd_sc_hd__or4_2
X_5773_ _9228_/Q _5770_/A _5965_/B1 _5770_/Y VGND VPWR _9228_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8561_ _8624_/B _8632_/B VGND VPWR _8713_/B VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_21_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4724_ _4720_/Y _5679_/B _4722_/Y _5768_/B VGND VPWR _4724_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_7512_ _6644_/Y _7451_/X _6713_/Y _7453_/X _7511_/X VGND VPWR _7517_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_8492_ _8492_/A VGND VPWR _8614_/A VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_190_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4655_ _9712_/Q _4636_/A _8952_/X _4636_/Y VGND VPWR _9712_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7443_ _7443_/A VGND VPWR _7443_/X VGND VPWR sky130_fd_sc_hd__buf_8
XFILLER_128_580 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4586_ _9741_/Q _4579_/A _5966_/B1 _4579_/Y VGND VPWR _9741_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7374_ _7374_/A _7374_/B _7374_/C _7374_/D VGND VPWR _7375_/C VGND VPWR sky130_fd_sc_hd__and4_1
Xinput71 mgmt_gpio_in[8] VGND VPWR _4737_/A VGND VPWR sky130_fd_sc_hd__clkbuf_2
Xinput82 spi_sdoenb VGND VPWR input82/X VGND VPWR sky130_fd_sc_hd__buf_4
Xinput60 mgmt_gpio_in[31] VGND VPWR _6132_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_6325_ _6325_/A _6325_/B _6325_/C VGND VPWR _6326_/D VGND VPWR sky130_fd_sc_hd__and3_2
X_9113_ _9378_/CLK _9113_/D _9646_/SET_B VGND VPWR _9113_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
Xinput93 sram_ro_data[0] VGND VPWR _4860_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_1_519 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9044_ _9790_/CLK _9044_/D VGND VPWR _9044_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_103_436 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_222 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6256_ _9473_/Q VGND VPWR _6256_/Y VGND VPWR sky130_fd_sc_hd__inv_4
XFILLER_76_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5207_ _9574_/Q _5203_/Y _8906_/X _5203_/A VGND VPWR _9574_/D VGND VPWR sky130_fd_sc_hd__o22a_1
X_6187_ _6187_/A _6187_/B _6187_/C VGND VPWR _6237_/B VGND VPWR sky130_fd_sc_hd__and3_1
X_5138_ _9624_/Q _5136_/A _8845_/X _5136_/Y VGND VPWR _9624_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_123_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_11 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5069_ _5069_/A VGND VPWR _9664_/D VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_8828_ _9591_/Q input81/X _8833_/S VGND VPWR _8828_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_12_136 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_88 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8759_ _8759_/A VGND VPWR _8760_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_12_158 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_54 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_572 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_136 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_567 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_464 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_412 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_266 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_472 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_122 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_162 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_358 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_550 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6110_ _9509_/Q VGND VPWR _6110_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_140_520 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7090_ _4720_/Y _7077_/C _4751_/Y _7077_/D _7089_/X VGND VPWR _7090_/X VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_58_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6041_ _6041_/A VGND VPWR _6041_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_39_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_7992_ _8116_/A _7992_/B VGND VPWR _7993_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_6943_ _6938_/Y _5594_/B _6939_/Y _5757_/B _6942_/X VGND VPWR _6944_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9731_ _9774_/CLK _9731_/D _7011_/B VGND VPWR _9731_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6874_ _9516_/Q VGND VPWR _6874_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9662_ _9664_/CLK _9662_/D _6146_/A VGND VPWR _9662_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_81_367 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_8613_ _8666_/C _8613_/B _8666_/D VGND VPWR _8616_/B VGND VPWR sky130_fd_sc_hd__or3_1
X_5825_ _9193_/Q _5820_/A _8929_/A1 _5820_/Y VGND VPWR _9193_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_167_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9593_ _9601_/CLK _9593_/D _9295_/SET_B VGND VPWR _9593_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_22_467 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5756_ _5713_/Y _5750_/Y _5755_/Y _9239_/Q _5755_/A VGND VPWR _9239_/D VGND VPWR
+ sky130_fd_sc_hd__a32o_2
X_8544_ _8544_/A _8544_/B _8544_/C VGND VPWR _8625_/B VGND VPWR sky130_fd_sc_hd__or3_2
X_8475_ _8703_/C _8617_/A _8475_/C VGND VPWR _8477_/A VGND VPWR sky130_fd_sc_hd__or3_1
X_5687_ _9258_/Q _5681_/A _8955_/A1 _5681_/Y VGND VPWR _9258_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_4707_ _4925_/A _4780_/B VGND VPWR _5671_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_7426_ _7472_/A _7476_/C _7474_/D VGND VPWR _7427_/A VGND VPWR sky130_fd_sc_hd__or3_1
X_4638_ _4994_/A VGND VPWR _4639_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_162_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_572 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7357_ _6533_/Y _7040_/C _6479_/Y _7059_/C VGND VPWR _7357_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4569_ _9753_/Q _4566_/A _8844_/X _4566_/Y VGND VPWR _9753_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7288_ _4899_/Y _7086_/X _4848_/Y _7088_/X VGND VPWR _7288_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_6308_ _9236_/Q VGND VPWR _6308_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_6239_ _9429_/Q VGND VPWR _6239_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9027_ _9027_/CLK _9027_/D VGND VPWR _9027_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_76_128 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_331 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_38 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_42 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_564 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6590_ _8777_/A _5306_/B _6589_/Y _5366_/B VGND VPWR _6590_/X VGND VPWR sky130_fd_sc_hd__o22a_2
X_5610_ _6052_/A _5610_/B VGND VPWR _5611_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_129_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5541_ _9349_/Q _5536_/A _8929_/A1 _5536_/Y VGND VPWR _9349_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_144_111 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8260_ _8260_/A _8260_/B VGND VPWR _8578_/B VGND VPWR sky130_fd_sc_hd__nor2_1
X_5472_ _9397_/Q _5471_/A _8846_/X _5471_/Y VGND VPWR _9397_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7211_ _7211_/A _7211_/B _7211_/C _7211_/D VGND VPWR _7221_/B VGND VPWR sky130_fd_sc_hd__and4_1
X_8191_ _8345_/A VGND VPWR _8583_/B VGND VPWR sky130_fd_sc_hd__inv_2
X_7142_ _6914_/Y _7059_/B _6905_/Y _7068_/C _7141_/X VGND VPWR _7145_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_86_404 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7073_ _7098_/C _7127_/A _7073_/C VGND VPWR _7074_/A VGND VPWR sky130_fd_sc_hd__or3_1
XFILLER_98_297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6024_ _9709_/Q _6023_/Y _9080_/Q _6023_/A VGND VPWR _9080_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_66_161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_386 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7975_ _7975_/A VGND VPWR _8389_/A VGND VPWR sky130_fd_sc_hd__buf_8
X_6926_ _9270_/Q VGND VPWR _6926_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9714_ _9089_/CLK _9714_/D _4648_/X VGND VPWR _9714_/Q VGND VPWR sky130_fd_sc_hd__dfrtn_1
XFILLER_14_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_9645_ _9774_/CLK _9645_/D _7011_/B VGND VPWR _9645_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6857_ _6855_/Y _5420_/B _6856_/Y _5374_/B VGND VPWR _6857_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_167_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6788_ _9529_/Q VGND VPWR _6788_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_5808_ _9056_/Q _5691_/A _5643_/Y _5753_/B _9203_/Q VGND VPWR _5808_/X VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9576_ _9788_/CLK _9576_/D _9646_/SET_B VGND VPWR _9576_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_136_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8527_ _8612_/B _8527_/B _8527_/C _8666_/A VGND VPWR _8531_/B VGND VPWR sky130_fd_sc_hd__or4_1
X_5739_ _9055_/Q _7125_/A _7127_/A _5737_/A _5713_/Y VGND VPWR _5740_/A VGND VPWR
+ sky130_fd_sc_hd__a32o_1
X_8458_ _7864_/X _8319_/A _8097_/B _8550_/A VGND VPWR _8614_/C VGND VPWR sky130_fd_sc_hd__o22ai_1
X_8389_ _8389_/A VGND VPWR _8518_/B VGND VPWR sky130_fd_sc_hd__inv_2
X_7409_ _7456_/A _7472_/A _9255_/Q VGND VPWR _7410_/A VGND VPWR sky130_fd_sc_hd__or3_1
XFILLER_38_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_540 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_584 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_246 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_328 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_6 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_183 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_7760_ _8394_/D VGND VPWR _7836_/A VGND VPWR sky130_fd_sc_hd__inv_2
X_4972_ _4972_/A VGND VPWR _4972_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_51_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_495 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_7691_ _6363_/Y _7455_/X _6445_/Y _7457_/X VGND VPWR _7691_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_6711_ _9538_/Q VGND VPWR _6711_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
X_6642_ _6637_/Y _5797_/B _6638_/Y _5768_/B _6641_/X VGND VPWR _6649_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9430_ _9508_/CLK _9430_/D _9295_/SET_B VGND VPWR _9430_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_9361_ _9545_/CLK _9361_/D _4628_/A VGND VPWR _9361_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_118_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6573_ _8789_/A _5317_/B _6569_/Y _4590_/B _6572_/X VGND VPWR _6586_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_8312_ _8310_/X _8676_/B _8592_/A _8312_/D VGND VPWR _8312_/X VGND VPWR sky130_fd_sc_hd__and4bb_1
X_5524_ _9360_/Q _5520_/A _5966_/B1 _5520_/Y VGND VPWR _9360_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_9292_ _9596_/CLK _9292_/D _9528_/SET_B VGND VPWR _9292_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
Xclkbuf_1_1_0_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/X VGND VPWR clkbuf_1_1_1_mgmt_gpio_in[4]/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_105_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8243_ _8243_/A VGND VPWR _8362_/B VGND VPWR sky130_fd_sc_hd__inv_2
X_5455_ _9408_/Q _5452_/A _5965_/B1 _5452_/Y VGND VPWR _9408_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8174_ _8376_/A _8174_/B VGND VPWR _8175_/B VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_132_147 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7125_ _7125_/A _7127_/B _7127_/C VGND VPWR _7126_/A VGND VPWR sky130_fd_sc_hd__or3_1
X_5386_ _9456_/Q _5384_/A _8845_/X _5384_/Y VGND VPWR _9456_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_86_234 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7056_ _9248_/Q _7056_/B _9246_/Q _9245_/Q VGND VPWR _7087_/B VGND VPWR sky130_fd_sc_hd__or4_1
XFILLER_55_610 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6007_ _6007_/A VGND VPWR _6007_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_39_194 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_484 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7958_ _8189_/A _8099_/B VGND VPWR _7966_/B VGND VPWR sky130_fd_sc_hd__or2_1
X_7889_ _8525_/A _8189_/A _7903_/C _8193_/A VGND VPWR _7890_/A VGND VPWR sky130_fd_sc_hd__or4_1
X_6909_ _9160_/Q VGND VPWR _6909_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
X_9628_ _9639_/CLK _9628_/D _9757_/SET_B VGND VPWR _9628_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_168_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_9559_ _9776_/CLK _9559_/D _4628_/A VGND VPWR _9559_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_108_133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_412 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_467 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_499 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_26 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_440 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA_130 _8816_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_141 _7199_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_152 _4602_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_178_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_134 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_163 _6264_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_174 _8632_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_185 input201/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_196 _7021_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_127_497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5240_ _5545_/A _5240_/B VGND VPWR _5241_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_102_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5171_ _9600_/Q _5169_/A _8845_/X _5169_/Y VGND VPWR _9600_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_96_565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_8930_ _9611_/Q _8930_/A1 _8930_/S VGND VPWR _8930_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_83_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput3 debug_out VGND VPWR input3/X VGND VPWR sky130_fd_sc_hd__buf_4
X_8861_ _8860_/X _9169_/Q _9054_/Q VGND VPWR _8861_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_304 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7812_ _8379_/D _8379_/B _7838_/B VGND VPWR _7813_/A VGND VPWR sky130_fd_sc_hd__or3_1
X_8792_ _8792_/A VGND VPWR _8792_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_36_175 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7743_ _9068_/Q _7743_/A2 _9067_/Q _7743_/B2 _7742_/X VGND VPWR _7743_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_4955_ _4949_/Y _4951_/Y _4952_/Y _4954_/X VGND VPWR _9709_/D VGND VPWR sky130_fd_sc_hd__o22ai_1
XFILLER_36_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4886_ _4882_/Y _4504_/B _4883_/Y _5259_/B _4885_/X VGND VPWR _4896_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_7674_ _6504_/Y _7451_/X _6556_/Y _7453_/X _7673_/X VGND VPWR _7679_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_137_206 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_543 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_386 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6625_ _8781_/A _4491_/B _6624_/Y _4822_/X VGND VPWR _6625_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_9413_ _9514_/CLK _9413_/D _9685_/SET_B VGND VPWR _9413_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_20_598 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_9344_ _9344_/CLK _9344_/D _9295_/SET_B VGND VPWR _9344_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6556_ _9440_/Q VGND VPWR _6556_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_192_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9275_ _9371_/CLK _9275_/D _9295_/SET_B VGND VPWR _9275_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_5507_ _5545_/A _5507_/B VGND VPWR _5508_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_6487_ _6485_/Y _5583_/B _6486_/Y _5864_/B VGND VPWR _6487_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_8226_ _8341_/A _8305_/B _8226_/C VGND VPWR _8499_/B VGND VPWR sky130_fd_sc_hd__nor3_1
XFILLER_105_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5438_ _9419_/Q _5433_/A _8842_/X _5433_/Y VGND VPWR _9419_/D VGND VPWR sky130_fd_sc_hd__a22o_1
Xoutput340 _9033_/Q VGND VPWR wb_dat_o[21] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput351 _9043_/Q VGND VPWR wb_dat_o[31] VGND VPWR sky130_fd_sc_hd__buf_2
X_5369_ _9467_/Q _5368_/A _5963_/B1 _5368_/Y VGND VPWR _9467_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8157_ _8164_/A _8554_/A VGND VPWR _8630_/B VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_86_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_320 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8088_ _8188_/B _8389_/A VGND VPWR _8433_/B VGND VPWR sky130_fd_sc_hd__nor2_1
X_7108_ _7108_/A _7108_/B _7108_/C _7108_/D VGND VPWR _7132_/B VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_87_598 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_267 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7039_ _7039_/A VGND VPWR _7040_/D VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_74_248 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_164 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_106 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_375 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_64 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_31 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_75 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_318 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_61 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_215 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_259 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_440 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_71 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_292 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_320 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4740_ _9190_/Q VGND VPWR _4740_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_119_217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4671_ _9354_/Q VGND VPWR _4671_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7390_ _6330_/Y _7118_/X _6335_/Y _7048_/C VGND VPWR _7390_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_6410_ _9316_/Q VGND VPWR _6410_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_6341_ _9545_/Q VGND VPWR _6341_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_115_412 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6272_ _6270_/Y _4861_/X _6271_/Y _5278_/B VGND VPWR _6272_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_9060_ _4450_/A1 _9060_/D _6146_/A VGND VPWR _9065_/D VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_115_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_404 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_318 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5223_ _9564_/Q _5218_/Y _8926_/X _5218_/A VGND VPWR _9564_/D VGND VPWR sky130_fd_sc_hd__o22a_1
X_8011_ _8583_/A _8538_/B _8525_/C VGND VPWR _8523_/A VGND VPWR sky130_fd_sc_hd__or3_2
X_5154_ _9611_/Q _5147_/A _8930_/A1 _5147_/Y VGND VPWR _9611_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_69_587 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5085_ _9656_/Q _5082_/A _5965_/B1 _5082_/Y VGND VPWR _9656_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_112_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8913_ _7723_/X _9087_/Q _9051_/Q VGND VPWR _8913_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_64_270 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8844_ _9705_/Q _9664_/Q _9587_/Q VGND VPWR _8844_/X VGND VPWR sky130_fd_sc_hd__mux2_8
XPHY_107 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_118 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_139 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5987_ _6040_/A VGND VPWR _5988_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_8775_ _8775_/A VGND VPWR _8776_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_7726_ _9698_/Q VGND VPWR _7726_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
X_4938_ _4994_/A VGND VPWR _4939_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_4869_ input4/X VGND VPWR _4869_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7657_ _6646_/Y _7465_/X _6730_/Y _7467_/X VGND VPWR _7657_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XANTENNA_30 _4681_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_41 _5355_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_20_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6608_ _8775_/A _5344_/B _6604_/Y _5328_/B _6607_/X VGND VPWR _6627_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XANTENNA_74 _6829_/D VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_52 _6111_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_63 _6294_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_192_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_518 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7588_ _6212_/Y _7471_/X _7260_/A _7473_/X _7587_/X VGND VPWR _7589_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XANTENNA_96 _7019_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_85 _8586_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_137_34 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6539_ _9117_/Q VGND VPWR _6539_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_192_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9327_ _9352_/CLK _9327_/D _9646_/SET_B VGND VPWR _9327_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_133_220 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9258_ _9601_/CLK _9258_/D _9295_/SET_B VGND VPWR _9258_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_106_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9189_ _9655_/CLK _9189_/D _9633_/SET_B VGND VPWR _9189_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_8209_ _8660_/A _8226_/C VGND VPWR _8210_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_153_88 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_9 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_150 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_362 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_204 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_470 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_579 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_354 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_462 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5910_ _9130_/Q _5907_/A _8844_/X _5907_/Y VGND VPWR _9130_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_6890_ _9219_/Q VGND VPWR _6890_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_34_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5841_ _9183_/Q _5839_/A _8845_/X _5839_/Y VGND VPWR _9183_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_34_454 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5772_ _9229_/Q _5770_/A _5964_/B1 _5770_/Y VGND VPWR _9229_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8560_ _8560_/A _8560_/B VGND VPWR _8713_/D VGND VPWR sky130_fd_sc_hd__or2_2
X_7511_ _6737_/Y _7455_/X _6773_/Y _7457_/X VGND VPWR _7511_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_8491_ _7862_/Y _8302_/Y _8667_/A _8369_/B VGND VPWR _8599_/D VGND VPWR sky130_fd_sc_hd__a211o_1
X_4723_ _6111_/B _4780_/B VGND VPWR _5768_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_187_481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7442_ _7476_/A _9251_/Q _7476_/C _7474_/D VGND VPWR _7443_/A VGND VPWR sky130_fd_sc_hd__or4_1
X_4654_ _4654_/A VGND VPWR _4654_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_147_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4585_ _9742_/Q _4579_/A _5965_/B1 _4579_/Y VGND VPWR _9742_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7373_ _6587_/Y _7124_/X _6480_/Y _7068_/B _7372_/X VGND VPWR _7374_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
Xinput50 mgmt_gpio_in[22] VGND VPWR input50/X VGND VPWR sky130_fd_sc_hd__clkbuf_4
Xinput61 mgmt_gpio_in[32] VGND VPWR input61/X VGND VPWR sky130_fd_sc_hd__clkbuf_4
Xinput72 mgmt_gpio_in[9] VGND VPWR _6941_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_6324_ _6320_/Y _5572_/B _6321_/Y _5507_/B _6323_/Y VGND VPWR _6325_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9112_ _9379_/CLK _9112_/D _9779_/SET_B VGND VPWR _9112_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
Xinput94 sram_ro_data[10] VGND VPWR _6778_/A VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
Xinput83 spimemio_flash_clk VGND VPWR input83/X VGND VPWR sky130_fd_sc_hd__buf_6
X_9043_ _9664_/CLK _9043_/D VGND VPWR _9043_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_6255_ _6239_/Y _5420_/B _6242_/X _6248_/X _6254_/X VGND VPWR _6326_/A VGND VPWR
+ sky130_fd_sc_hd__o2111a_1
XFILLER_67_19 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_286 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5206_ _9575_/Q _5203_/Y _8928_/X _5203_/A VGND VPWR _9575_/D VGND VPWR sky130_fd_sc_hd__o22a_1
X_6186_ _7260_/A _5610_/B _6182_/Y _5776_/B _6185_/X VGND VPWR _6187_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_130_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5137_ _9625_/Q _5136_/A _8846_/X _5136_/Y VGND VPWR _9625_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_5068_ _8966_/X _9664_/Q _5078_/S VGND VPWR _5069_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_72_516 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_23 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_410 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8827_ _8826_/X _7020_/B _9586_/Q VGND VPWR _8827_/X VGND VPWR sky130_fd_sc_hd__mux2_4
XFILLER_16_45 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_8758_ _8758_/A VGND VPWR _8758_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_7709_ _9083_/Q _9082_/Q VGND VPWR _7711_/A VGND VPWR sky130_fd_sc_hd__nand2_1
X_8689_ _8689_/A _8709_/D _8713_/C _8714_/D VGND VPWR _8689_/X VGND VPWR sky130_fd_sc_hd__or4_1
XFILLER_193_440 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_358 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_584 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_520 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_608 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_579 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_292 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_7 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_134 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_510 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_554 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6040_ _6040_/A VGND VPWR _6041_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_66_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7991_ _7991_/A VGND VPWR _8550_/A VGND VPWR sky130_fd_sc_hd__clkbuf_4
X_6942_ _6940_/Y _5080_/B _6941_/Y _6134_/A VGND VPWR _6942_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_9730_ _9774_/CLK _9730_/D _7011_/B VGND VPWR _9730_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
X_9661_ _9664_/CLK _9661_/D _6146_/A VGND VPWR _9661_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6873_ _9438_/Q VGND VPWR _6873_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_179_245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5824_ _9194_/Q _5820_/A _8925_/A1 _5820_/Y VGND VPWR _9194_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8612_ _8612_/A _8612_/B VGND VPWR _8666_/D VGND VPWR sky130_fd_sc_hd__or2_1
X_9592_ _9617_/CLK _9592_/D _9295_/SET_B VGND VPWR _9592_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_8543_ _8543_/A VGND VPWR _8543_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_5755_ _5755_/A VGND VPWR _5755_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_147_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5686_ _9259_/Q _5681_/A _8842_/X _5681_/Y VGND VPWR _9259_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8474_ _8474_/A _8474_/B VGND VPWR _8475_/C VGND VPWR sky130_fd_sc_hd__or2_1
X_4706_ _9264_/Q VGND VPWR _4706_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_163_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_175 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_14 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4637_ _9718_/Q _4636_/A _8953_/X _4636_/Y VGND VPWR _9718_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7425_ _7425_/A VGND VPWR _7425_/X VGND VPWR sky130_fd_sc_hd__buf_8
XFILLER_162_123 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4568_ _9754_/Q _4566_/A _8845_/X _4566_/Y VGND VPWR _9754_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7356_ _6574_/Y _7082_/X _6615_/Y _7084_/X _7355_/X VGND VPWR _7375_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_116_584 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_212 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4499_ _9780_/Q _4493_/A _5965_/B1 _4493_/Y VGND VPWR _9780_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7287_ _7287_/A _7287_/B _7287_/C VGND VPWR _7287_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
X_6307_ _6307_/A _6307_/B _6307_/C _6307_/D VGND VPWR _6326_/C VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_134_24 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_9026_ _9027_/CLK _9026_/D VGND VPWR _9026_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_6238_ _6149_/A _6237_/Y _9042_/Q _6149_/Y VGND VPWR _9042_/D VGND VPWR sky130_fd_sc_hd__o22a_1
X_6169_ _9508_/Q VGND VPWR _6169_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_57_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_43_csclk _9329_/CLK VGND VPWR _9758_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_13_413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_402 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_98 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_166 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_63 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_372 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_350 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_416 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_346 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_576 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_248 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_276 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_290 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5540_ _9350_/Q _5536_/A _8925_/A1 _5536_/Y VGND VPWR _9350_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_157_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5471_ _5471_/A VGND VPWR _5471_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_117_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7210_ _6367_/Y _7048_/D _6439_/Y _7040_/B _7209_/X VGND VPWR _7211_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_8190_ _8189_/A _8213_/A _8189_/Y VGND VPWR _8345_/A VGND VPWR sky130_fd_sc_hd__a21oi_1
XFILLER_125_370 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7141_ _6819_/Y _7079_/B _6926_/Y _7059_/A VGND VPWR _7141_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_7072_ _7072_/A VGND VPWR _7077_/B VGND VPWR sky130_fd_sc_hd__buf_8
XFILLER_98_276 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_416 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6023_ _6023_/A VGND VPWR _6023_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_39_343 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_471 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_516 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7974_ _8379_/B _8093_/A VGND VPWR _7975_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_27_549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9713_ _9089_/CLK _9713_/D _4651_/X VGND VPWR _9713_/Q VGND VPWR sky130_fd_sc_hd__dfrtn_1
X_6925_ _6925_/A _6925_/B _6925_/C _6925_/D VGND VPWR _6945_/B VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_120_48 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_37 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_9644_ _9776_/CLK _9644_/D _4628_/A VGND VPWR _9644_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6856_ _9459_/Q VGND VPWR _6856_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_22_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5807_ _9204_/Q _5799_/A _8916_/A1 _5799_/Y VGND VPWR _9204_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_9575_ _9613_/CLK _9575_/D _9646_/SET_B VGND VPWR _9575_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6787_ _9469_/Q VGND VPWR _6787_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
XFILLER_167_248 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8526_ _8525_/Y _8517_/Y _8518_/X _8449_/A VGND VPWR _8666_/A VGND VPWR sky130_fd_sc_hd__a31o_1
X_5738_ _9246_/Q _5738_/B VGND VPWR _7127_/A VGND VPWR sky130_fd_sc_hd__or2_2
XFILLER_136_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5669_ _9270_/Q _5662_/A _8840_/X _5662_/Y VGND VPWR _9270_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8457_ _8521_/B _8246_/B _8029_/X VGND VPWR _8459_/C VGND VPWR sky130_fd_sc_hd__o21ai_2
X_8388_ _8098_/B _8397_/B _8171_/X VGND VPWR _8631_/A VGND VPWR sky130_fd_sc_hd__o21ai_1
X_7408_ _7408_/A VGND VPWR _7408_/X VGND VPWR sky130_fd_sc_hd__buf_6
XFILLER_150_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_210 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7339_ _6657_/Y _7079_/B _6634_/Y _7059_/A VGND VPWR _7339_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_77_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_384 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9009_ _9009_/A _8795_/A VGND VPWR mgmt_gpio_out[32] VGND VPWR sky130_fd_sc_hd__ebufn_8
XFILLER_57_151 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_324 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_379 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_64 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_552 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_596 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_579 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_9 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_159 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_2_1_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A VGND VPWR clkbuf_3_3_0_wb_clk_i/A VGND
+ VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_0_180 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_246 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4971_ _4994_/A VGND VPWR _4972_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_6710_ _9426_/Q VGND VPWR _6710_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7690_ _6374_/Y _7441_/X _6387_/Y _7443_/X _7689_/X VGND VPWR _7697_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_6641_ _6639_/Y _5776_/B _6640_/Y _5789_/B VGND VPWR _6641_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_177_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_568 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_9360_ _9771_/CLK _9360_/D _4628_/A VGND VPWR _9360_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_118_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6572_ _6570_/Y _4907_/X _8773_/A _5382_/B VGND VPWR _6572_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_8311_ _8640_/A _8311_/B VGND VPWR _8592_/A VGND VPWR sky130_fd_sc_hd__or2_2
X_5523_ _9361_/Q _5520_/A _5965_/B1 _5520_/Y VGND VPWR _9361_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_9291_ _9596_/CLK _9291_/D _9528_/SET_B VGND VPWR _9291_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_5454_ _9409_/Q _5452_/A _5964_/B1 _5452_/Y VGND VPWR _9409_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8242_ _8510_/A _8246_/B VGND VPWR _8243_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_132_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5385_ _9457_/Q _5384_/A _8846_/X _5384_/Y VGND VPWR _9457_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8173_ _8688_/A _8173_/B VGND VPWR _8174_/B VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_132_159 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_552 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7124_ _7124_/A VGND VPWR _7124_/X VGND VPWR sky130_fd_sc_hd__buf_8
X_7055_ _7055_/A VGND VPWR _7059_/C VGND VPWR sky130_fd_sc_hd__buf_6
X_6006_ _6040_/A VGND VPWR _6007_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_54_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_452 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_603 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_496 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7957_ _8583_/A _8189_/A _8099_/B VGND VPWR _8195_/B VGND VPWR sky130_fd_sc_hd__or3_1
X_6908_ _9647_/Q VGND VPWR _6908_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7888_ _8496_/A _8521_/B VGND VPWR _7896_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_6839_ _9757_/Q VGND VPWR _6839_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_168_546 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9627_ _9757_/CLK _9627_/D _9757_/SET_B VGND VPWR _9627_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_24_89 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_596 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9558_ _9758_/CLK _9558_/D _9633_/SET_B VGND VPWR _9558_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_136_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_239 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8509_ _8509_/A _8693_/A _8600_/B _8662_/B VGND VPWR _8512_/B VGND VPWR sky130_fd_sc_hd__or4_1
X_9489_ _9493_/CLK _9489_/D _4628_/A VGND VPWR _9489_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_108_178 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_479 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_38 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_302 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_52 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_120 input86/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_131 _7015_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_142 _7221_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_153 _5013_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_164 _6461_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_175 _8098_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_197 input78/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_186 input201/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_186_376 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5170_ _9601_/Q _5169_/A _8846_/X _5169_/Y VGND VPWR _9601_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_110_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_387 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_471 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput4 mask_rev_in[0] VGND VPWR input4/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_8860_ _7590_/Y _9638_/Q _8978_/S VGND VPWR _8860_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_7811_ _7811_/A VGND VPWR _8202_/A VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_8791_ _8791_/A VGND VPWR _8792_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_51_102 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4954_ _4953_/Y _7008_/A _9092_/Q _9048_/Q _9091_/Q VGND VPWR _4954_/X VGND VPWR
+ sky130_fd_sc_hd__o2111a_1
X_7742_ _9066_/Q _7742_/B VGND VPWR _7742_/X VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_189_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7673_ _6508_/Y _7455_/X _6551_/Y _7457_/X VGND VPWR _7673_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4885_ _6158_/A _6086_/B input34/X VGND VPWR _4885_/X VGND VPWR sky130_fd_sc_hd__or3b_1
X_9412_ _9493_/CLK _9412_/D _4628_/A VGND VPWR _9412_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_165_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6624_ _6624_/A VGND VPWR _6624_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_9343_ _9344_/CLK _9343_/D _9295_/SET_B VGND VPWR _9343_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6555_ _9362_/Q VGND VPWR _6555_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_180_519 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5506_ _9372_/Q _5498_/A _8916_/A1 _5498_/Y VGND VPWR _9372_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_9274_ _9371_/CLK _9274_/D _9295_/SET_B VGND VPWR _9274_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_10_25 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6486_ _9162_/Q VGND VPWR _6486_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_8225_ _8305_/B _8260_/B VGND VPWR _8571_/B VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_105_159 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5437_ _9420_/Q _5433_/A _8925_/A1 _5433_/Y VGND VPWR _9420_/D VGND VPWR sky130_fd_sc_hd__a22o_1
Xoutput352 _9023_/Q VGND VPWR wb_dat_o[3] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput330 _9016_/Q VGND VPWR wb_dat_o[12] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput341 _9034_/Q VGND VPWR wb_dat_o[22] VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_120_118 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5368_ _5368_/A VGND VPWR _5368_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_8156_ _8156_/A _8578_/A VGND VPWR _8158_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_113_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7107_ _4734_/Y _7048_/D _4769_/Y _7040_/B _7106_/X VGND VPWR _7108_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_8087_ _8514_/B _8086_/Y VGND VPWR _8296_/A VGND VPWR sky130_fd_sc_hd__or2b_1
X_5299_ _5299_/A VGND VPWR _5300_/A VGND VPWR sky130_fd_sc_hd__clkbuf_2
X_7038_ _9246_/Q _9245_/Q _7127_/B _7073_/C VGND VPWR _7039_/A VGND VPWR sky130_fd_sc_hd__or4_1
X_8989_ _9574_/Q _8755_/A VGND VPWR mgmt_gpio_out[12] VGND VPWR sky130_fd_sc_hd__ebufn_8
XFILLER_70_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_43 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_240 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_242 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_8 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_452 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_332 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4670_ _4927_/A _4843_/B VGND VPWR _5872_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_147_549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6340_ _9540_/Q VGND VPWR _6340_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_6_581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_424 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6271_ _9525_/Q VGND VPWR _6271_/Y VGND VPWR sky130_fd_sc_hd__inv_6
XFILLER_130_416 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_8010_ _7864_/X _8085_/A _8009_/X VGND VPWR _8016_/B VGND VPWR sky130_fd_sc_hd__o21ai_1
X_5222_ _9565_/Q _5218_/Y _8925_/X _5218_/A VGND VPWR _9565_/D VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_130_438 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5153_ _9612_/Q _5147_/A _8955_/A1 _5147_/Y VGND VPWR _9612_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_69_599 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5084_ _9657_/Q _5082_/A _5964_/B1 _5082_/Y VGND VPWR _9657_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8912_ _7720_/X _9086_/Q _9051_/Q VGND VPWR _8912_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_37_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8843_ _9704_/Q _9663_/Q _9587_/Q VGND VPWR _8843_/X VGND VPWR sky130_fd_sc_hd__mux2_8
XFILLER_25_603 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_282 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_580 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_119 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_108 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5986_ _9091_/Q _5985_/Y _5981_/X VGND VPWR _9091_/D VGND VPWR sky130_fd_sc_hd__o21ba_1
X_8774_ _8774_/A VGND VPWR _8774_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_4937_ _4636_/Y _8957_/S _4936_/Y _9711_/Q _4636_/A VGND VPWR _9711_/D VGND VPWR
+ sky130_fd_sc_hd__a32o_1
X_7725_ _9088_/Q _7722_/B _7724_/Y _9089_/Q _7722_/Y VGND VPWR _7725_/X VGND VPWR
+ sky130_fd_sc_hd__a32o_1
X_4868_ _6111_/A _4898_/A VGND VPWR _4868_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_7656_ _6682_/Y _7451_/X _6723_/Y _7453_/X _7655_/X VGND VPWR _7661_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XANTENNA_31 _4681_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_20 _7518_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_6607_ _8769_/A _5458_/B _6606_/Y _5290_/B VGND VPWR _6607_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XANTENNA_75 _6832_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_64 _6446_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_53 _6117_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_42 _5355_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_4_507 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7587_ _6188_/Y _7475_/X _6179_/Y _7477_/X VGND VPWR _7587_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4799_ _4792_/Y _4564_/B _4793_/Y _5240_/B _4798_/X VGND VPWR _4830_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9326_ _9352_/CLK _9326_/D _9646_/SET_B VGND VPWR _9326_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XANTENNA_97 _7019_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_86 _8586_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_20_385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_7 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_46 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6538_ _6538_/A VGND VPWR _6538_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
XFILLER_106_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6469_ _9766_/Q VGND VPWR _6469_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9257_ _9601_/CLK _9257_/D _9295_/SET_B VGND VPWR _9257_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_133_276 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_308 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8208_ _8305_/B _8264_/B VGND VPWR _8595_/C VGND VPWR sky130_fd_sc_hd__nor2_1
X_9188_ _9758_/CLK _9188_/D _9633_/SET_B VGND VPWR _9188_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_121_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_8139_ _8550_/A _8640_/B VGND VPWR _8730_/A VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_101_173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_514 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_32 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_591 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_116 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_216 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_300 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_388 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_208 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_474 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_260 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5840_ _9184_/Q _5839_/A _8846_/X _5839_/Y VGND VPWR _9184_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_5771_ _9230_/Q _5770_/A _5963_/B1 _5770_/Y VGND VPWR _9230_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_4722_ _9226_/Q VGND VPWR _4722_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_8490_ _8734_/A _8490_/B _8490_/C VGND VPWR _8597_/D VGND VPWR sky130_fd_sc_hd__or3_1
X_7510_ _6643_/Y _7441_/X _6704_/Y _7443_/X _7509_/X VGND VPWR _7517_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_187_493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7441_ _7441_/A VGND VPWR _7441_/X VGND VPWR sky130_fd_sc_hd__buf_8
X_4653_ _4994_/A VGND VPWR _4654_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput40 mgmt_gpio_in[13] VGND VPWR _6317_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_7372_ _6549_/Y _7126_/X _6609_/Y _7128_/X VGND VPWR _7372_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4584_ _9743_/Q _4579_/A _5964_/B1 _4579_/Y VGND VPWR _9743_/D VGND VPWR sky130_fd_sc_hd__a22o_1
Xinput51 mgmt_gpio_in[23] VGND VPWR input51/X VGND VPWR sky130_fd_sc_hd__clkbuf_2
Xinput62 mgmt_gpio_in[33] VGND VPWR input62/X VGND VPWR sky130_fd_sc_hd__clkbuf_4
Xinput73 pad_flash_io0_di VGND VPWR _7018_/B VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_143_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_232 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6323_ _8818_/A _4680_/Y input57/X _6322_/Y VGND VPWR _6323_/Y VGND VPWR sky130_fd_sc_hd__a22oi_4
X_9111_ _9379_/CLK _9111_/D _9646_/SET_B VGND VPWR _9111_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
Xinput84 spimemio_flash_csb VGND VPWR input84/X VGND VPWR sky130_fd_sc_hd__buf_4
Xinput95 sram_ro_data[11] VGND VPWR _6552_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_89_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_9042_ _9664_/CLK _9042_/D VGND VPWR _9042_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_6254_ _6249_/Y _4832_/X _6250_/Y _5110_/B _6253_/X VGND VPWR _6254_/X VGND VPWR
+ sky130_fd_sc_hd__o221a_2
XFILLER_170_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5205_ _9576_/Q _5203_/Y _8927_/X _5203_/A VGND VPWR _9576_/D VGND VPWR sky130_fd_sc_hd__o22a_1
X_6185_ _6183_/Y _5757_/B _6184_/Y _5797_/B VGND VPWR _6185_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_69_341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5136_ _5136_/A VGND VPWR _5136_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_84_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5067_ _5067_/A VGND VPWR _9665_/D VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_72_528 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_422 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_8826_ _8825_/X _6505_/A _9682_/Q VGND VPWR _8826_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_13_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5969_ _5969_/A VGND VPWR _5970_/A VGND VPWR sky130_fd_sc_hd__clkbuf_4
X_8757_ _8757_/A VGND VPWR _8758_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_178_460 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7708_ _9082_/Q VGND VPWR _7708_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_8688_ _8688_/A _8688_/B _8688_/C VGND VPWR _8714_/D VGND VPWR sky130_fd_sc_hd__or3_1
X_7639_ _6897_/Y _7465_/X _6848_/Y _7467_/X VGND VPWR _7639_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_4_304 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9309_ _9789_/CLK _9309_/D _9647_/SET_B VGND VPWR _9309_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_106_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_108 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_598 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_303 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_366 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_400 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_572 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_621 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_530 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_146 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_506 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7990_ _8050_/B _7992_/B VGND VPWR _7991_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_6941_ _6941_/A VGND VPWR _6941_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9660_ _9664_/CLK _9660_/D _6146_/A VGND VPWR _9660_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6872_ _9386_/Q VGND VPWR _6872_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_34_285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5823_ _9195_/Q _5820_/A _8844_/X _5820_/Y VGND VPWR _9195_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8611_ _8064_/C _8610_/Y _8016_/A _8527_/B VGND VPWR _8613_/B VGND VPWR sky130_fd_sc_hd__a211o_1
X_9591_ _9601_/CLK _9591_/D _9295_/SET_B VGND VPWR _9591_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_179_257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_8542_ _8703_/B _8605_/A _8705_/A _8541_/Y VGND VPWR _8543_/A VGND VPWR sky130_fd_sc_hd__or4b_1
X_5754_ _6997_/A _5643_/Y _5713_/Y _5753_/X VGND VPWR _5755_/A VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_175_441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5685_ _9260_/Q _5681_/A _8925_/A1 _5681_/Y VGND VPWR _9260_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8473_ _8471_/Y _8472_/Y _8061_/A _8708_/C VGND VPWR _8474_/B VGND VPWR sky130_fd_sc_hd__a31o_1
X_4705_ _4705_/A _4705_/B _4705_/C _4705_/D VGND VPWR _4936_/A VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_147_187 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_519 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4636_ _4636_/A VGND VPWR _4636_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7424_ _7462_/A _7470_/B _9255_/Q VGND VPWR _7425_/A VGND VPWR sky130_fd_sc_hd__or3_1
XFILLER_162_135 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7355_ _6497_/Y _7077_/C _6583_/Y _7077_/D _7354_/X VGND VPWR _7355_/X VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_150_319 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4567_ _9755_/Q _4566_/A _8846_/X _4566_/Y VGND VPWR _9755_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_6306_ _6301_/Y _5776_/B _6302_/Y _5872_/B _6305_/X VGND VPWR _6307_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_143_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4498_ _9781_/Q _4493_/A _5964_/B1 _4493_/Y VGND VPWR _9781_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7286_ _7286_/A _7286_/B _7286_/C _7286_/D VGND VPWR _7287_/C VGND VPWR sky130_fd_sc_hd__and4_1
X_9025_ _9027_/CLK _9025_/D VGND VPWR _9025_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_6237_ _6237_/A _6237_/B _6237_/C _6237_/D VGND VPWR _6237_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
X_6168_ _9526_/Q VGND VPWR _6168_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_5119_ _9633_/Q _5112_/A _5966_/B1 _5112_/Y VGND VPWR _9633_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_6099_ _6099_/A VGND VPWR _6099_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
Xclkbuf_3_3_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/A VGND VPWR _9278_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_53_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_8809_ _8809_/A VGND VPWR _8813_/B VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_185_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_458 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9789_ _9789_/CLK _9789_/D _9685_/SET_B VGND VPWR _9789_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_138_132 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_187 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_428 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_300 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_122 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_358 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_230 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_588 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_291 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_280 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5470_ _5470_/A VGND VPWR _5471_/A VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_117_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_606 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_466 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_511 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7140_ _6865_/Y _7095_/X _6939_/Y _7068_/D _7139_/X VGND VPWR _7145_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_140_330 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_7071_ _7096_/B _7073_/C VGND VPWR _7072_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_39_300 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6022_ _6022_/A _6022_/B _6022_/C _6022_/D VGND VPWR _6023_/A VGND VPWR sky130_fd_sc_hd__or4_1
XFILLER_82_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_130 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7973_ _7973_/A VGND VPWR _8554_/A VGND VPWR sky130_fd_sc_hd__clkbuf_4
X_9712_ _9089_/CLK _9712_/D _4654_/X VGND VPWR _9712_/Q VGND VPWR sky130_fd_sc_hd__dfrtn_1
X_6924_ _6919_/Y _5949_/B _6920_/Y _5837_/B _6923_/X VGND VPWR _6925_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9643_ _9776_/CLK _9643_/D _7011_/B VGND VPWR _9643_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_167_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6855_ _9425_/Q VGND VPWR _6855_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_22_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5806_ _9205_/Q _5799_/A _8930_/A1 _5799_/Y VGND VPWR _9205_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_6786_ _6149_/A _6785_/Y _9038_/Q _6149_/Y VGND VPWR _9038_/D VGND VPWR sky130_fd_sc_hd__o22a_1
X_9574_ _9788_/CLK _9574_/D _9646_/SET_B VGND VPWR _9574_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_8525_ _8525_/A _8538_/B _8525_/C VGND VPWR _8525_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
X_5737_ _5737_/A _9245_/Q VGND VPWR _7125_/A VGND VPWR sky130_fd_sc_hd__or2_2
X_8456_ _7864_/X _8316_/A _8097_/B _8137_/B VGND VPWR _8734_/C VGND VPWR sky130_fd_sc_hd__o22ai_1
XFILLER_135_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5668_ _9271_/Q _5662_/A _8841_/X _5662_/Y VGND VPWR _9271_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7407_ _7476_/A _9251_/Q _7470_/B _7474_/D VGND VPWR _7408_/A VGND VPWR sky130_fd_sc_hd__or4_1
XFILLER_151_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5599_ _9309_/Q _5596_/A _8841_/X _5596_/Y VGND VPWR _9309_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_4619_ _9722_/Q _4615_/A _5966_/B1 _4615_/Y VGND VPWR _9722_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8387_ _8389_/A _8632_/B VGND VPWR _8687_/B VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_150_105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_24 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7338_ _6729_/Y _7095_/X _6638_/Y _7068_/D _7337_/X VGND VPWR _7343_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_104_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7269_ _6129_/Y _7040_/C _6123_/Y _7059_/C VGND VPWR _7269_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_9008_ _9601_/Q _8793_/A VGND VPWR mgmt_gpio_out[31] VGND VPWR sky130_fd_sc_hd__ebufn_8
XFILLER_57_130 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_163 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_76 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_20 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_208 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_135 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_91 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_382 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4970_ _9706_/Q _4966_/A _9705_/Q _4966_/Y VGND VPWR _9706_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_177_525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6640_ _9214_/Q VGND VPWR _6640_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_6571_ _9453_/Q VGND VPWR _8773_/A VGND VPWR sky130_fd_sc_hd__inv_6
XFILLER_145_400 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5522_ _9362_/Q _5520_/A _5964_/B1 _5520_/Y VGND VPWR _9362_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8310_ _8571_/B _8310_/B _8497_/A _8309_/X VGND VPWR _8310_/X VGND VPWR sky130_fd_sc_hd__or4b_1
XFILLER_117_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9290_ _9483_/CLK _9290_/D _9528_/SET_B VGND VPWR _9290_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_133_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5453_ _9410_/Q _5452_/A _5963_/B1 _5452_/Y VGND VPWR _9410_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8241_ _8241_/A _8574_/B _8361_/B _8730_/B VGND VPWR _8245_/A VGND VPWR sky130_fd_sc_hd__or4_1
X_5384_ _5384_/A VGND VPWR _5384_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_8172_ _8172_/A _8373_/A _8171_/X VGND VPWR _8173_/B VGND VPWR sky130_fd_sc_hd__or3b_1
X_7123_ _7127_/C _7123_/B VGND VPWR _7124_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_5848__10 _8924_/X VGND VPWR _5889_/A1 VGND VPWR sky130_fd_sc_hd__inv_4
XFILLER_5_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_428 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7054_ _7094_/B _7073_/C VGND VPWR _7055_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_67_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6005_ _9086_/Q _5995_/A _8911_/X _5995_/Y VGND VPWR _9086_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_67_494 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_464 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7956_ _8379_/C _8394_/A _8394_/B VGND VPWR _8099_/B VGND VPWR sky130_fd_sc_hd__or3_1
XFILLER_70_615 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6907_ _6902_/Y _5024_/B _6903_/Y _6135_/A _6906_/X VGND VPWR _6925_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_7887_ _7836_/B _7879_/Y _7886_/X VGND VPWR _7887_/Y VGND VPWR sky130_fd_sc_hd__o21ai_2
X_6838_ _9633_/Q VGND VPWR _6838_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9626_ _8837_/A1 _9626_/D _5130_/X VGND VPWR _9626_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_9557_ _9755_/CLK _9557_/D _9633_/SET_B VGND VPWR _9557_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6769_ input5/X VGND VPWR _6769_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_8508_ _8282_/C _7831_/Y _8394_/A _7767_/C _8331_/B VGND VPWR _8662_/B VGND VPWR
+ sky130_fd_sc_hd__a41o_1
X_9488_ _9777_/CLK _9488_/D _9757_/SET_B VGND VPWR _9488_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_191_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_45 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_8439_ _8518_/A _8064_/B _8061_/C _8062_/B VGND VPWR _8617_/A VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_77_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_450 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_121 input86/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_132 _7015_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_143 _7536_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_110 input77/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_154 _5960_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_165 _6549_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_176 _8647_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_186_322 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_350 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA_198 input83/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_187 _8807_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_186_388 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_506 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_90 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_422 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_572 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_116 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_490 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_399 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xinput5 mask_rev_in[10] VGND VPWR input5/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_49_483 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7810_ _8660_/C _7878_/A VGND VPWR _7811_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_91_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8790_ _8790_/A VGND VPWR _8790_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_4953_ _9708_/Q VGND VPWR _4953_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7741_ _9068_/Q _7741_/A2 _9067_/Q _7741_/B2 _7740_/X VGND VPWR _7741_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_51_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7672_ _6477_/Y _7441_/X _6615_/Y _7443_/X _7671_/X VGND VPWR _7679_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_177_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4884_ _4911_/A _6111_/B VGND VPWR _5259_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_9411_ _9514_/CLK _9411_/D _9685_/SET_B VGND VPWR _9411_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6623_ _9781_/Q VGND VPWR _8781_/A VGND VPWR sky130_fd_sc_hd__inv_6
XFILLER_165_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_580 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6554_ _6549_/Y _4504_/B _6550_/Y _5259_/B _6553_/X VGND VPWR _6567_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9342_ _9508_/CLK _9342_/D _9647_/SET_B VGND VPWR _9342_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_173_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5505_ _9373_/Q _5498_/A _8930_/A1 _5498_/Y VGND VPWR _9373_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_9273_ _9535_/CLK _9273_/D _9528_/SET_B VGND VPWR _9273_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6485_ _9315_/Q VGND VPWR _6485_/Y VGND VPWR sky130_fd_sc_hd__inv_4
XFILLER_118_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5436_ _9421_/Q _5433_/A _8844_/X _5433_/Y VGND VPWR _9421_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8224_ _8595_/C _8224_/B _8224_/C _8223_/X VGND VPWR _8227_/B VGND VPWR sky130_fd_sc_hd__or4b_2
Xoutput320 _9766_/Q VGND VPWR sram_ro_addr[4] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput353 _9024_/Q VGND VPWR wb_dat_o[4] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput331 _9017_/Q VGND VPWR wb_dat_o[13] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput342 _9035_/Q VGND VPWR wb_dat_o[23] VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_99_372 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8155_ _8213_/A _8552_/A VGND VPWR _8578_/A VGND VPWR sky130_fd_sc_hd__nor2_1
X_5367_ _5367_/A VGND VPWR _5368_/A VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_141_491 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7106_ _4708_/Y _7068_/A _4793_/Y _7105_/X VGND VPWR _7106_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_5298_ _5671_/A _5298_/B VGND VPWR _5299_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_8086_ _8086_/A _8086_/B VGND VPWR _8086_/Y VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_59_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_578 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7037_ _7037_/A _9247_/Q VGND VPWR _7127_/B VGND VPWR sky130_fd_sc_hd__or2_2
XFILLER_19_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_306 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_8988_ _9573_/Q _8753_/A VGND VPWR mgmt_gpio_out[11] VGND VPWR sky130_fd_sc_hd__ebufn_8
XFILLER_42_136 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7939_ _8202_/A _8510_/A _7938_/Y VGND VPWR _7939_/X VGND VPWR sky130_fd_sc_hd__o21ba_1
XFILLER_11_523 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9609_ _9617_/CLK _9609_/D _9295_/SET_B VGND VPWR _9609_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_109_444 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_358 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_512 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_171 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_280 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_155 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_434 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_174 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_436 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6270_ _6270_/A VGND VPWR _6270_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_5221_ _9566_/Q _5218_/Y _8921_/X _5218_/A VGND VPWR _9566_/D VGND VPWR sky130_fd_sc_hd__o22a_1
X_5152_ _9613_/Q _5147_/A _8929_/A1 _5147_/Y VGND VPWR _9613_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_96_331 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5083_ _9658_/Q _5082_/A _5963_/B1 _5082_/Y VGND VPWR _9658_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_110_185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_8911_ _7717_/X _9085_/Q _9051_/Q VGND VPWR _8911_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_8842_ _9703_/Q _9662_/Q _9587_/Q VGND VPWR _8842_/X VGND VPWR sky130_fd_sc_hd__mux2_8
XFILLER_37_497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8773_ _8773_/A VGND VPWR _8774_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_24_114 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7724_ _9089_/Q VGND VPWR _7724_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_5985_ _6022_/C _5985_/B VGND VPWR _5985_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_52_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4936_ _4936_/A _4936_/B _4936_/C VGND VPWR _4936_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
X_7655_ _6662_/Y _7455_/X _6745_/Y _7457_/X VGND VPWR _7655_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4867_ _4867_/A VGND VPWR _4867_/Y VGND VPWR sky130_fd_sc_hd__inv_4
XANTENNA_21 _7608_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_10 _7265_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_32 _4681_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_192_111 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_314 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_196 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7586_ _6194_/Y _7461_/X _6168_/Y _7463_/X _7585_/X VGND VPWR _7589_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_6606_ _9518_/Q VGND VPWR _6606_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XANTENNA_65 _6595_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_43 _4858_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_54 _6153_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_4798_ _4795_/Y _5121_/B _4797_/Y _4613_/B VGND VPWR _4798_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_9325_ _9613_/CLK _9325_/D _9646_/SET_B VGND VPWR _9325_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6537_ _9109_/Q VGND VPWR _7703_/A VGND VPWR sky130_fd_sc_hd__clkinv_4
XANTENNA_76 _6847_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_87 _8753_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_98 _7019_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_192_166 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_18 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6468_ _9155_/Q VGND VPWR _6468_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9256_ _9601_/CLK _9256_/D _9528_/SET_B VGND VPWR _9256_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_106_469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6399_ _9467_/Q VGND VPWR _6399_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_5419_ _9432_/Q _5414_/A _5967_/B1 _5414_/Y VGND VPWR _9432_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_9187_ _9757_/CLK _9187_/D _9633_/SET_B VGND VPWR _9187_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_8207_ _8207_/A VGND VPWR _8264_/B VGND VPWR sky130_fd_sc_hd__buf_6
X_8138_ _8164_/A _8550_/A VGND VPWR _8361_/A VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_87_342 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_79 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_375 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_526 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8069_ _8069_/A _8203_/A VGND VPWR _8069_/Y VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_101_185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_220 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_336 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_16 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_274 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_520 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_139 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_228 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_486 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5770_ _5770_/A VGND VPWR _5770_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_175_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4721_ _4917_/A _4780_/B VGND VPWR _5679_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_174_100 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7440_ _7462_/A _7476_/C _9255_/Q VGND VPWR _7441_/A VGND VPWR sky130_fd_sc_hd__or3_1
X_4652_ _9713_/Q _4636_/A _8951_/X _4636_/Y VGND VPWR _9713_/D VGND VPWR sky130_fd_sc_hd__a22o_1
Xinput30 mask_rev_in[4] VGND VPWR _6470_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_4583_ _9744_/Q _4579_/A _5963_/B1 _4579_/Y VGND VPWR _9744_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7371_ _6543_/Y _5728_/X _6529_/Y _7040_/A _7370_/X VGND VPWR _7374_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9110_ _9695_/CLK _9110_/D _9779_/SET_B VGND VPWR _9110_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
Xinput41 mgmt_gpio_in[14] VGND VPWR input41/X VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
Xinput63 mgmt_gpio_in[34] VGND VPWR _8803_/A VGND VPWR sky130_fd_sc_hd__buf_6
Xinput52 mgmt_gpio_in[24] VGND VPWR _4781_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_155_380 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput74 pad_flash_io1_di VGND VPWR _7020_/B VGND VPWR sky130_fd_sc_hd__buf_2
Xinput85 spimemio_flash_io0_do VGND VPWR input85/X VGND VPWR sky130_fd_sc_hd__buf_4
X_6322_ _6322_/A VGND VPWR _6322_/Y VGND VPWR sky130_fd_sc_hd__inv_6
Xinput96 sram_ro_data[12] VGND VPWR _6336_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_115_244 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_9041_ _9664_/CLK _9041_/D VGND VPWR _9041_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_6253_ _8822_/X _6251_/Y _6252_/Y _4841_/X VGND VPWR _6253_/X VGND VPWR sky130_fd_sc_hd__o2bb2a_1
XFILLER_89_607 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_428 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5204_ _9577_/Q _5203_/Y _8898_/X _5203_/A VGND VPWR _9577_/D VGND VPWR sky130_fd_sc_hd__o22a_1
X_6184_ _9210_/Q VGND VPWR _6184_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_111_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5135_ _5135_/A VGND VPWR _5136_/A VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_111_483 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5066_ _8967_/X _9665_/Q _5078_/S VGND VPWR _5067_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_25_434 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_231 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8825_ _9579_/Q _9718_/Q _8977_/S VGND VPWR _8825_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_52_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5968_ _6052_/A _5968_/B VGND VPWR _5969_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_8756_ _8756_/A VGND VPWR _8756_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_166_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7707_ _9049_/Q _9052_/Q VGND VPWR _7707_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
X_4919_ _4919_/A _4931_/B VGND VPWR _5480_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_178_472 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_35 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5899_ _5899_/A VGND VPWR _5899_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_8687_ _8720_/A _8687_/B _8687_/C VGND VPWR _8713_/C VGND VPWR sky130_fd_sc_hd__or3_1
X_7638_ _6883_/Y _7451_/X _6873_/Y _7453_/X _7637_/X VGND VPWR _7643_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_193_486 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7569_ _6291_/Y _7475_/X _6316_/Y _7477_/X VGND VPWR _7569_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_180_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_211 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9308_ _9789_/CLK _9308_/D _9647_/SET_B VGND VPWR _9308_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_161_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_106 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_9239_ _9278_/CLK _9239_/D _9757_/SET_B VGND VPWR _9239_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_0_555 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_504 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_570 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_584 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_604 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_61 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_158 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_372 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6940_ _9655_/Q VGND VPWR _6940_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_66_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_203 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6871_ _9399_/Q VGND VPWR _6871_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
X_5822_ _9196_/Q _5820_/A _8845_/X _5820_/Y VGND VPWR _9196_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8610_ _8189_/A _7885_/X _7881_/A VGND VPWR _8610_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
X_9590_ _9601_/CLK _9590_/D _9295_/SET_B VGND VPWR _9590_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_148_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5753_ _9056_/Q _5753_/B _5787_/A VGND VPWR _5753_/X VGND VPWR sky130_fd_sc_hd__and3_1
X_8541_ _8541_/A _8617_/B _8705_/D _8619_/D VGND VPWR _8541_/Y VGND VPWR sky130_fd_sc_hd__nor4_1
XFILLER_34_297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4704_ _4694_/Y _5864_/B _4696_/Y _6165_/A _4703_/X VGND VPWR _4705_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_5684_ _9261_/Q _5681_/A _8844_/X _5681_/Y VGND VPWR _9261_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8472_ _8472_/A VGND VPWR _8472_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_175_475 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_7423_ _4708_/Y _7415_/X _4701_/Y _7417_/X _7422_/X VGND VPWR _7481_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_4635_ _4635_/A VGND VPWR _4636_/A VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_147_199 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_328 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7354_ _6556_/Y _7086_/X _6612_/Y _7088_/X VGND VPWR _7354_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4566_ _4566_/A VGND VPWR _4566_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_150_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6305_ _6303_/Y _5968_/B _6304_/Y _5905_/B VGND VPWR _6305_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4497_ _9782_/Q _4493_/A _5963_/B1 _4493_/Y VGND VPWR _9782_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_9024_ _9027_/CLK _9024_/D VGND VPWR _9024_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_7285_ _6090_/Y _7124_/X _6061_/Y _7068_/B _7284_/X VGND VPWR _7286_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_103_247 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6236_ _6236_/A _6236_/B _6236_/C _6236_/D VGND VPWR _6237_/D VGND VPWR sky130_fd_sc_hd__and4_2
X_6167_ _6163_/Y _5583_/B _6164_/Y _5458_/B _6166_/Y VGND VPWR _6174_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_5118_ _9634_/Q _5112_/A _5965_/B1 _5112_/Y VGND VPWR _9634_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_6098_ _9353_/Q VGND VPWR _6098_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_45_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5049_ _9673_/Q _5047_/A _8845_/X _5047_/Y VGND VPWR _9673_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8808_ _8808_/A _8808_/B VGND VPWR _8808_/Y VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_80_392 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9788_ _9788_/CLK _9788_/D _9646_/SET_B VGND VPWR _9788_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_8739_ _8739_/A VGND VPWR _8739_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_153_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_74 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_134 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_242 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_270 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_292 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_103 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_618 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_523 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7070_ _7070_/A VGND VPWR _7077_/A VGND VPWR sky130_fd_sc_hd__buf_8
XFILLER_100_206 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6021_ _6021_/A VGND VPWR _6021_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_1_csclk clkbuf_1_1_1_csclk/A VGND VPWR clkbuf_2_3_0_csclk/A VGND VPWR
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_39_312 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_484 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7972_ _8096_/B _8116_/A VGND VPWR _7973_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_6923_ _6921_/Y _5013_/B _6922_/Y _5916_/B VGND VPWR _6923_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_9711_ _9709_/CLK _9711_/D _4657_/X VGND VPWR _9711_/Q VGND VPWR sky130_fd_sc_hd__dfrtn_1
XFILLER_66_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9642_ _9776_/CLK _9642_/D _4628_/A VGND VPWR _9642_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6854_ _9503_/Q VGND VPWR _6854_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_13_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5805_ _9206_/Q _5799_/A _8955_/A1 _5799_/Y VGND VPWR _9206_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_6785_ _6785_/A _6785_/B _6785_/C VGND VPWR _6785_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
X_9573_ _9613_/CLK _9573_/D _9646_/SET_B VGND VPWR _9573_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_129_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8524_ _8523_/Y _8517_/Y _8518_/X _8444_/A VGND VPWR _8527_/C VGND VPWR sky130_fd_sc_hd__a31o_1
X_5736_ _5724_/B _7104_/A _7056_/B _5692_/A _5735_/X VGND VPWR _9247_/D VGND VPWR
+ sky130_fd_sc_hd__o311a_1
XFILLER_148_453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5667_ _9272_/Q _5662_/A _8929_/A1 _5662_/Y VGND VPWR _9272_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8455_ _8455_/A _8455_/B VGND VPWR _8459_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_135_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4618_ _9723_/Q _4615_/A _5965_/B1 _4615_/Y VGND VPWR _9723_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7406_ _9254_/Q _7406_/B VGND VPWR _7470_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_135_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_231 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5598_ _9310_/Q _5596_/A _8842_/X _5596_/Y VGND VPWR _9310_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8386_ _8386_/A _8386_/B VGND VPWR _8632_/B VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_190_297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_36 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_512 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7337_ _6780_/Y _7097_/X _6711_/Y _7099_/X VGND VPWR _7337_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4549_ _8811_/A _8975_/S VGND VPWR _4551_/B VGND VPWR sky130_fd_sc_hd__nand2_8
XFILLER_145_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7268_ _6073_/Y _7082_/X _6114_/Y _7084_/X _7267_/X VGND VPWR _7287_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_104_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9007_ _9600_/Q _8791_/A VGND VPWR mgmt_gpio_out[30] VGND VPWR sky130_fd_sc_hd__ebufn_8
X_6219_ _6219_/A VGND VPWR _6219_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_7199_ _7199_/A _7199_/B _7199_/C VGND VPWR _7199_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
XFILLER_161_79 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_50 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_220 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_320 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_228 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_386 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6570_ _6570_/A VGND VPWR _6570_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_5521_ _9363_/Q _5520_/A _5963_/B1 _5520_/Y VGND VPWR _9363_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_117_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8240_ _8316_/A _8264_/B VGND VPWR _8730_/B VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_172_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_231 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5452_ _5452_/A VGND VPWR _5452_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_117_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_8171_ _8396_/A _8397_/B VGND VPWR _8171_/X VGND VPWR sky130_fd_sc_hd__or2_1
X_5383_ _5383_/A VGND VPWR _5384_/A VGND VPWR sky130_fd_sc_hd__clkbuf_4
X_7122_ _4816_/Y _5728_/X _4842_/Y _7040_/A _7121_/X VGND VPWR _7131_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_5848__11 _8924_/X VGND VPWR _5863_/B1 VGND VPWR sky130_fd_sc_hd__inv_4
XFILLER_86_204 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_150 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7053_ _7053_/A VGND VPWR _7059_/B VGND VPWR sky130_fd_sc_hd__buf_8
X_6004_ _6004_/A VGND VPWR _6004_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_27_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_318 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7955_ _8437_/B _8164_/A VGND VPWR _8585_/B VGND VPWR sky130_fd_sc_hd__nor2_2
X_7886_ _8566_/A _7886_/B _7879_/B _7885_/X VGND VPWR _7886_/X VGND VPWR sky130_fd_sc_hd__or4bb_1
X_6906_ _6904_/Y _5526_/B _6905_/Y _6081_/B VGND VPWR _6906_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_6837_ _9628_/Q VGND VPWR _6837_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9625_ _9674_/CLK _9625_/D _9633_/SET_B VGND VPWR _9625_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_9556_ _9777_/CLK _9556_/D _9633_/SET_B VGND VPWR _9556_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6768_ _9750_/Q VGND VPWR _6768_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_8507_ _7879_/A _7881_/A _7848_/A _8300_/B _7931_/A VGND VPWR _8600_/B VGND VPWR
+ sky130_fd_sc_hd__o221ai_2
X_6699_ _9742_/Q VGND VPWR _6699_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_5719_ _5737_/A _5738_/B VGND VPWR _7104_/A VGND VPWR sky130_fd_sc_hd__or2_2
X_9487_ _9777_/CLK _9487_/D _7011_/B VGND VPWR _9487_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_163_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_8438_ _8515_/A _8521_/B VGND VPWR _8703_/D VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_156_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8369_ _8630_/B _8369_/B VGND VPWR _8645_/C VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_151_459 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_12 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_150 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_100 _7019_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_122 input86/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_111 input80/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_133 _7015_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_33_329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_144 _7626_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_166 _6590_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_155 _5960_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_81_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA_199 input83/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_188 _8808_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_177 _8761_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_186_334 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_518 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_434 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_584 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xinput6 mask_rev_in[11] VGND VPWR input6/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_64_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_240 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_19 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4952_ _9709_/Q VGND VPWR _4952_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7740_ _9066_/Q _7740_/B VGND VPWR _7740_/X VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_177_301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4883_ _9536_/Q VGND VPWR _4883_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7671_ _6612_/Y _7445_/X _6587_/Y _7447_/X VGND VPWR _7671_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_20_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6622_ _9523_/Q VGND VPWR _8787_/A VGND VPWR sky130_fd_sc_hd__inv_8
X_9410_ _9514_/CLK _9410_/D _4628_/A VGND VPWR _9410_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_165_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_580 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_412 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6553_ _6551_/Y _5100_/B _6552_/Y _4893_/X VGND VPWR _6553_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_9341_ _9344_/CLK _9341_/D _9295_/SET_B VGND VPWR _9341_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6484_ _9310_/Q VGND VPWR _6484_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_5504_ _9374_/Q _5498_/A _8955_/A1 _5498_/Y VGND VPWR _9374_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_9272_ _9344_/CLK _9272_/D _9295_/SET_B VGND VPWR _9272_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_118_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5435_ _9422_/Q _5433_/A _8845_/X _5433_/Y VGND VPWR _9422_/D VGND VPWR sky130_fd_sc_hd__a22o_1
Xoutput310 _8821_/X VGND VPWR serial_resetn VGND VPWR sky130_fd_sc_hd__buf_2
X_8223_ _8223_/A _8223_/B VGND VPWR _8223_/X VGND VPWR sky130_fd_sc_hd__and2_1
Xoutput321 _9767_/Q VGND VPWR sram_ro_addr[5] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput332 _9018_/Q VGND VPWR wb_dat_o[14] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput343 _9036_/Q VGND VPWR wb_dat_o[24] VGND VPWR sky130_fd_sc_hd__buf_2
X_8154_ _8154_/A _8367_/A VGND VPWR _8156_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_5366_ _5671_/A _5366_/B VGND VPWR _5367_/A VGND VPWR sky130_fd_sc_hd__or2_1
Xoutput354 _9025_/Q VGND VPWR wb_dat_o[5] VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_99_384 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5297_ _9515_/Q _5292_/A _5967_/B1 _5292_/Y VGND VPWR _9515_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8085_ _8085_/A _8538_/D VGND VPWR _8086_/B VGND VPWR sky130_fd_sc_hd__or2_1
X_7105_ _7105_/A VGND VPWR _7105_/X VGND VPWR sky130_fd_sc_hd__buf_8
XFILLER_142_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7036_ _7036_/A VGND VPWR _7040_/C VGND VPWR sky130_fd_sc_hd__buf_6
XFILLER_142_37 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8987_ _8987_/A _8751_/A VGND VPWR mgmt_gpio_out[10] VGND VPWR sky130_fd_sc_hd__ebufn_8
XFILLER_43_605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7938_ _8094_/A _7938_/B VGND VPWR _7938_/Y VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_168_301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_9608_ _9617_/CLK _9608_/D _9295_/SET_B VGND VPWR _9608_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_7869_ _8226_/C _8316_/A VGND VPWR _7870_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_11_535 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_423 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9539_ _9768_/CLK _9539_/D _4628_/A VGND VPWR _9539_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_93_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_292 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_70 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_41_csclk clkbuf_2_1_0_csclk/X VGND VPWR _9779_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_33_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_90 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_186 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5220_ _9567_/Q _5218_/Y _8918_/X _5218_/A VGND VPWR _9567_/D VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_102_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_278 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5151_ _9614_/Q _5147_/A _8925_/A1 _5147_/Y VGND VPWR _9614_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_5082_ _5082_/A VGND VPWR _5082_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_96_354 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8910_ _7715_/Y _9084_/Q _9051_/Q VGND VPWR _8910_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_110_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8841_ _9702_/Q _9661_/Q _9587_/Q VGND VPWR _8841_/X VGND VPWR sky130_fd_sc_hd__mux2_8
XFILLER_52_413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8772_ _8772_/A VGND VPWR _8772_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_24_148 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_7723_ _9088_/Q _7722_/B _7722_/Y VGND VPWR _7723_/X VGND VPWR sky130_fd_sc_hd__o21a_1
X_5984_ _5984_/A VGND VPWR _5984_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_4935_ _4935_/A _4935_/B _4935_/C _4935_/D VGND VPWR _4936_/C VGND VPWR sky130_fd_sc_hd__and4_2
XFILLER_177_142 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4866_ _4911_/A _4925_/A VGND VPWR _5336_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_7654_ _6638_/Y _7441_/X _6705_/Y _7443_/X _7653_/X VGND VPWR _7661_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XANTENNA_22 _7608_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_11 _7287_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_165_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4797_ _9721_/Q VGND VPWR _4797_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_6605_ _9401_/Q VGND VPWR _8769_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_165_326 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7585_ _6184_/Y _7465_/X _6160_/Y _7467_/X VGND VPWR _7585_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XANTENNA_44 _4867_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_66 _6676_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_55 _6205_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_33 _4681_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_192_123 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_398 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6536_ _6531_/Y _6322_/A _7699_/A _5872_/B _6535_/X VGND VPWR _6536_/X VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9324_ _9352_/CLK _9324_/D _9646_/SET_B VGND VPWR _9324_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XANTENNA_88 _8783_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_77 _6877_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_99 _7019_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_118_275 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_178 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6467_ _9189_/Q VGND VPWR _6467_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9255_ _9278_/CLK _9255_/D _9779_/SET_B VGND VPWR _9255_/Q VGND VPWR sky130_fd_sc_hd__dfstp_4
X_6398_ _9350_/Q VGND VPWR _6398_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_5418_ _9433_/Q _5414_/A _5966_/B1 _5414_/Y VGND VPWR _9433_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_9186_ _9758_/CLK _9186_/D _9633_/SET_B VGND VPWR _9186_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_8206_ _8272_/A _8226_/C VGND VPWR _8207_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_133_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5349_ _9481_/Q _5346_/A _8844_/X _5346_/Y VGND VPWR _9481_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8137_ _8213_/A _8137_/B VGND VPWR _8574_/A VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_153_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_8068_ _8515_/A _8164_/A VGND VPWR _8203_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_46_12 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_538 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_432 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7019_ _7019_/A VGND VPWR _7019_/X VGND VPWR sky130_fd_sc_hd__buf_6
XFILLER_15_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_77 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_186 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_220 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_348 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_70 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_387 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_498 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4720_ _9256_/Q VGND VPWR _4720_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
XFILLER_175_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_112 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4651_ _4651_/A VGND VPWR _4651_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_147_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xinput31 mask_rev_in[5] VGND VPWR _6257_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput20 mask_rev_in[24] VGND VPWR _4821_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_4582_ _9745_/Q _4579_/A _8844_/X _4579_/Y VGND VPWR _9745_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7370_ _7370_/A _7392_/B VGND VPWR _7370_/X VGND VPWR sky130_fd_sc_hd__or2_1
Xinput53 mgmt_gpio_in[25] VGND VPWR input53/X VGND VPWR sky130_fd_sc_hd__clkbuf_4
Xinput42 mgmt_gpio_in[15] VGND VPWR input42/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput64 mgmt_gpio_in[35] VGND VPWR _6538_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_115_212 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput86 spimemio_flash_io0_oeb VGND VPWR input86/X VGND VPWR sky130_fd_sc_hd__buf_6
Xinput75 porb VGND VPWR _7011_/B VGND VPWR sky130_fd_sc_hd__buf_12
X_6321_ _9369_/Q VGND VPWR _6321_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
Xinput97 sram_ro_data[13] VGND VPWR _6292_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_170_351 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_256 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9040_ _9664_/CLK _9040_/D VGND VPWR _9040_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_6252_ _6252_/A VGND VPWR _6252_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_5203_ _5203_/A VGND VPWR _5203_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_6183_ _9237_/Q VGND VPWR _6183_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_5134_ _6165_/A _5156_/B VGND VPWR _5135_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_57_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_495 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5065_ _5065_/A VGND VPWR _9666_/D VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_8824_ _9578_/Q input3/X input1/X VGND VPWR _8824_/X VGND VPWR sky130_fd_sc_hd__mux2_2
XFILLER_16_59 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_427 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5967_ _9101_/Q _5962_/A _5967_/B1 _5962_/Y VGND VPWR _9101_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8755_ _8755_/A VGND VPWR _8756_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_8686_ _8686_/A _8686_/B _8686_/C _8686_/D VGND VPWR _8709_/D VGND VPWR sky130_fd_sc_hd__or4_2
X_4918_ _9385_/Q VGND VPWR _4918_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_7706_ _7706_/A VGND VPWR _7706_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_166_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_25 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_47 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7637_ _6898_/Y _7455_/X _6833_/Y _7457_/X VGND VPWR _7637_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_5898_ _5898_/A VGND VPWR _5899_/A VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_120_7 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4849_ _6111_/B _4931_/B VGND VPWR _5442_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_7568_ _6284_/Y _7461_/X _6271_/Y _7463_/X _7567_/X VGND VPWR _7571_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_180_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6519_ _8749_/A _5818_/B _8759_/A _5660_/B _6518_/X VGND VPWR _6526_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_7499_ _7499_/A _7499_/B _7499_/C _7499_/D VGND VPWR _7500_/D VGND VPWR sky130_fd_sc_hd__and4_1
X_9307_ _9789_/CLK _9307_/D _9685_/SET_B VGND VPWR _9307_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_134_554 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_9238_ _9371_/CLK _9238_/D _9295_/SET_B VGND VPWR _9238_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_161_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9169_ _9203_/CLK _9169_/D _9633_/SET_B VGND VPWR _9169_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_87_140 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_22 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_516 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_240 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_72 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_582 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_232 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_94 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_616 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_350 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_73 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_251 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6870_ _6865_/Y _5344_/B _6866_/Y _5366_/B _6869_/X VGND VPWR _6877_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_179_215 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5821_ _9197_/Q _5820_/A _8846_/X _5820_/Y VGND VPWR _9197_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_5752_ _9280_/Q _9279_/Q _9278_/Q VGND VPWR _5787_/A VGND VPWR sky130_fd_sc_hd__or3_1
X_8540_ _8540_/A _8704_/B VGND VPWR _8619_/D VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_148_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4703_ _4699_/Y _5897_/B _4701_/Y _5013_/B VGND VPWR _4703_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_5683_ _9262_/Q _5681_/A _8845_/X _5681_/Y VGND VPWR _9262_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8471_ _8538_/C VGND VPWR _8471_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_190_413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_104 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7422_ _4773_/Y _7419_/X _4857_/Y _7421_/X VGND VPWR _7422_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4634_ _5214_/A _4964_/B VGND VPWR _4635_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_7353_ _7353_/A _7353_/B _7353_/C VGND VPWR _7353_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
X_4565_ _4565_/A VGND VPWR _4566_/A VGND VPWR sky130_fd_sc_hd__buf_2
X_6304_ _9130_/Q VGND VPWR _6304_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7284_ _6104_/Y _7126_/X _6116_/Y _7128_/X VGND VPWR _7284_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4496_ _9783_/Q _4493_/A _8844_/X _4493_/Y VGND VPWR _9783_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_9023_ _9027_/CLK _9023_/D VGND VPWR _9023_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_89_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6235_ _6230_/Y _5968_/B _6231_/Y _5110_/B _6234_/X VGND VPWR _6236_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_6166_ input69/X _8955_/S input50/X _8926_/S VGND VPWR _6166_/Y VGND VPWR sky130_fd_sc_hd__a22oi_1
XFILLER_57_302 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5117_ _9635_/Q _5112_/A _5964_/B1 _5112_/Y VGND VPWR _9635_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_6097_ _6097_/A VGND VPWR _6097_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_27_14 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5048_ _9674_/Q _5047_/A _8846_/X _5047_/Y VGND VPWR _9674_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_150_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9787_ _9790_/CLK _9787_/D _9757_/SET_B VGND VPWR _9787_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_8807_ _8807_/A _8807_/B VGND VPWR _8807_/Y VGND VPWR sky130_fd_sc_hd__nor2_2
X_8738_ _8738_/A VGND VPWR _8738_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_40_268 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_246 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8669_ _8713_/A _8703_/D _8706_/B VGND VPWR _8670_/C VGND VPWR sky130_fd_sc_hd__or3_1
XFILLER_4_114 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_89 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_18 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_20 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_260 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_270 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_282 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_271 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6020_ _6040_/A VGND VPWR _6021_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_100_218 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_482 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_496 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7971_ _7971_/A _8098_/A VGND VPWR _8116_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_9710_ _9709_/CLK _9710_/D _4939_/X VGND VPWR _9710_/Q VGND VPWR sky130_fd_sc_hd__dfrtn_1
X_6922_ _9121_/Q VGND VPWR _6922_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_6853_ _9451_/Q VGND VPWR _6853_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9641_ _9774_/CLK _9641_/D _7011_/B VGND VPWR _9641_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_50_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5804_ _9207_/Q _5799_/A _8842_/X _5799_/Y VGND VPWR _9207_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_50_522 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_246 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6784_ _6784_/A _6784_/B _6784_/C _6784_/D VGND VPWR _6785_/C VGND VPWR sky130_fd_sc_hd__and4_1
X_9572_ _9788_/CLK _9572_/D _9646_/SET_B VGND VPWR _9572_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_148_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8523_ _8523_/A VGND VPWR _8523_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_5735_ _9246_/Q _9245_/Q _9055_/Q _9247_/Q VGND VPWR _5735_/X VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_129_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5666_ _9273_/Q _5662_/A _8925_/A1 _5662_/Y VGND VPWR _9273_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8454_ _8454_/A _8454_/B VGND VPWR _8455_/B VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_163_413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4617_ _9724_/Q _4615_/A _5964_/B1 _4615_/Y VGND VPWR _9724_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7405_ _7405_/A VGND VPWR _7405_/X VGND VPWR sky130_fd_sc_hd__buf_6
X_5597_ _9311_/Q _5596_/A _8843_/X _5596_/Y VGND VPWR _9311_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8385_ _8650_/C _8385_/B VGND VPWR _8436_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_190_287 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7336_ _6682_/Y _7048_/B _6772_/Y _7077_/A _7335_/X VGND VPWR _7343_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_2
X_4548_ _4548_/A VGND VPWR _8975_/S VGND VPWR sky130_fd_sc_hd__buf_12
X_7267_ _6139_/Y _7077_/C _6133_/Y _7077_/D _7266_/X VGND VPWR _7267_/X VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_4479_ _4729_/A _4729_/B _4669_/A _8932_/X VGND VPWR _4931_/A VGND VPWR sky130_fd_sc_hd__or4_4
X_9006_ _9599_/Q _8789_/A VGND VPWR mgmt_gpio_out[29] VGND VPWR sky130_fd_sc_hd__ebufn_8
X_6218_ _9112_/Q VGND VPWR _6218_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
X_7198_ _7198_/A _7198_/B _7198_/C _7198_/D VGND VPWR _7199_/C VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_97_290 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6149_ _6149_/A VGND VPWR _6149_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_26_596 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_511 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_382 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_95 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_118 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_63 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_102 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_319 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_354 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_332 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5520_ _5520_/A VGND VPWR _5520_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_157_262 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_104 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_243 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5451_ _5451_/A VGND VPWR _5452_/A VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_172_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8170_ _8170_/A _8389_/A VGND VPWR _8396_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_5382_ _5545_/A _5382_/B VGND VPWR _5383_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_160_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7121_ _7121_/A _7392_/B VGND VPWR _7121_/X VGND VPWR sky130_fd_sc_hd__or2_1
X_5848__12 _8924_/X VGND VPWR _5849_/A VGND VPWR sky130_fd_sc_hd__inv_4
XFILLER_101_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7052_ _7075_/A _7085_/B VGND VPWR _7053_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_140_162 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6003_ _6040_/A VGND VPWR _6004_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_67_430 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_143 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_7954_ _7954_/A VGND VPWR _8164_/A VGND VPWR sky130_fd_sc_hd__buf_12
X_6905_ _9391_/Q VGND VPWR _6905_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_24_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7885_ _8515_/B _7885_/B VGND VPWR _7885_/X VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_35_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6836_ _6831_/Y _4822_/X _6832_/Y _5278_/B _6835_/X VGND VPWR _6878_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9624_ _9674_/CLK _9624_/D _9633_/SET_B VGND VPWR _9624_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_9555_ _9758_/CLK _9555_/D _7011_/B VGND VPWR _9555_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6767_ _9400_/Q VGND VPWR _6767_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
XFILLER_148_240 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_560 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5718_ _9245_/Q VGND VPWR _5738_/B VGND VPWR sky130_fd_sc_hd__inv_2
X_8506_ _8615_/A _8506_/B _8506_/C VGND VPWR _8693_/A VGND VPWR sky130_fd_sc_hd__or3_2
X_9486_ _9777_/CLK _9486_/D _7011_/B VGND VPWR _9486_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6698_ _9078_/Q VGND VPWR _6698_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_5649_ _5649_/A _5649_/B _9278_/Q _9277_/Q VGND VPWR _6997_/C VGND VPWR sky130_fd_sc_hd__or4_1
X_8437_ _8632_/A _8437_/B VGND VPWR _8704_/B VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_156_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8368_ _8368_/A _8577_/C _8675_/A _8578_/C VGND VPWR _8372_/A VGND VPWR sky130_fd_sc_hd__or4_2
XFILLER_49_12 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_298 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7319_ _6932_/Y _7068_/A _6805_/Y _7105_/X VGND VPWR _7319_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_104_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8299_ _8299_/A _8299_/B VGND VPWR _8300_/B VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_172_24 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_89 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_162 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_387 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_84 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_123 input86/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_101 _8805_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_112 input81/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_134 _7015_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_61_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA_145 _7626_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_167 _6807_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_156 _5960_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_14_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_189 _7021_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_178 _8765_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_186_346 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_87 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_0_csclk clkbuf_0_csclk/X VGND VPWR clkbuf_1_1_1_csclk/A VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_60_9 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_302 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xinput7 mask_rev_in[12] VGND VPWR input7/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_64_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_168 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_319 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4951_ _9048_/Q _4951_/B VGND VPWR _4951_/Y VGND VPWR sky130_fd_sc_hd__nand2_1
X_4882_ _9773_/Q VGND VPWR _4882_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7670_ _6516_/Y _7425_/X _7667_/X _7669_/X VGND VPWR _7680_/C VGND VPWR sky130_fd_sc_hd__o211a_1
XFILLER_17_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6621_ _9765_/Q VGND VPWR _6621_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_20_525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_9340_ _9535_/CLK _9340_/D _9528_/SET_B VGND VPWR _9340_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6552_ _6552_/A VGND VPWR _6552_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_145_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5503_ _9375_/Q _5498_/A _8929_/A1 _5498_/Y VGND VPWR _9375_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_9271_ _9535_/CLK _9271_/D _9528_/SET_B VGND VPWR _9271_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6483_ _9297_/Q VGND VPWR _8761_/A VGND VPWR sky130_fd_sc_hd__inv_6
XFILLER_9_592 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_276 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_468 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_8222_ _8341_/A _8498_/A _8640_/A VGND VPWR _8223_/B VGND VPWR sky130_fd_sc_hd__or3_1
X_5434_ _9423_/Q _5433_/A _8846_/X _5433_/Y VGND VPWR _9423_/D VGND VPWR sky130_fd_sc_hd__a22o_1
Xoutput300 _9044_/Q VGND VPWR pwr_ctrl_out[0] VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_133_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_8153_ _8552_/A _8378_/B VGND VPWR _8367_/A VGND VPWR sky130_fd_sc_hd__nor2_1
Xoutput322 _9768_/Q VGND VPWR sram_ro_addr[6] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput311 _8804_/X VGND VPWR spi_sdi VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput333 _9019_/Q VGND VPWR wb_dat_o[15] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput344 _9037_/Q VGND VPWR wb_dat_o[25] VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_160_279 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7104_ _7104_/A _7127_/B _7127_/C VGND VPWR _7105_/A VGND VPWR sky130_fd_sc_hd__or3_1
X_5365_ _9468_/Q _5357_/A _8839_/X _5357_/Y VGND VPWR _9468_/D VGND VPWR sky130_fd_sc_hd__a22o_1
Xoutput355 _9026_/Q VGND VPWR wb_dat_o[6] VGND VPWR sky130_fd_sc_hd__buf_2
X_5296_ _9516_/Q _5292_/A _5966_/B1 _5292_/Y VGND VPWR _9516_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8084_ _8084_/A _8521_/B VGND VPWR _8538_/D VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_87_547 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7035_ _7115_/B _7073_/C VGND VPWR _7036_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_67_260 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_49 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_400 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_8986_ _8986_/A _8749_/A VGND VPWR mgmt_gpio_out[9] VGND VPWR sky130_fd_sc_hd__ebufn_2
XFILLER_43_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7937_ _8282_/C _7836_/C _8282_/B _8703_/A _7936_/X VGND VPWR _7938_/B VGND VPWR
+ sky130_fd_sc_hd__a311oi_1
Xclkbuf_2_0_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A VGND VPWR clkbuf_3_1_0_wb_clk_i/A VGND
+ VPWR sky130_fd_sc_hd__clkbuf_2
X_7868_ _7868_/A VGND VPWR _8316_/A VGND VPWR sky130_fd_sc_hd__clkbuf_4
X_9607_ _9617_/CLK _9607_/D _9295_/SET_B VGND VPWR _9607_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6819_ _9417_/Q VGND VPWR _6819_/Y VGND VPWR sky130_fd_sc_hd__inv_4
XFILLER_11_547 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7799_ _8394_/C VGND VPWR _8379_/C VGND VPWR sky130_fd_sc_hd__inv_6
XFILLER_51_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_402 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9538_ _9768_/CLK _9538_/D _4628_/A VGND VPWR _9538_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_167_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9469_ _9684_/CLK _9469_/D _9685_/SET_B VGND VPWR _9469_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_191_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_490 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_67 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_536 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_528 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_411 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_263 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8815__378 VGND VGND VPWR VPWR _9057_/D _8815__378/LO sky130_fd_sc_hd__conb_1
XFILLER_61_469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_91 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_80 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_338 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_536 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5150_ _9615_/Q _5147_/A _8844_/X _5147_/Y VGND VPWR _9615_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_123_493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5081_ _5081_/A VGND VPWR _5082_/A VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_96_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8840_ _9701_/Q _9660_/Q _9587_/Q VGND VPWR _8840_/X VGND VPWR sky130_fd_sc_hd__mux2_8
XFILLER_64_230 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5983_ _6040_/A VGND VPWR _5984_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_8771_ _8771_/A VGND VPWR _8772_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_4934_ _4934_/A _4934_/B _4934_/C _4934_/D VGND VPWR _4935_/D VGND VPWR sky130_fd_sc_hd__and4_1
X_7722_ _9088_/Q _7722_/B VGND VPWR _7722_/Y VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_32_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_182 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_154 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7653_ _6695_/Y _7445_/X _6700_/Y _7447_/X VGND VPWR _7653_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4865_ _9484_/Q VGND VPWR _4865_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
XANTENNA_23 _7662_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_12 _7287_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_4796_ _6111_/A _4903_/B VGND VPWR _5121_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_7584_ _6175_/Y _7451_/X _6159_/Y _7453_/X _7583_/X VGND VPWR _7589_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_6604_ _9492_/Q VGND VPWR _6604_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XANTENNA_45 _4890_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_56 _6211_/D VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_34 _4777_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_192_135 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_232 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6535_ _6533_/Y _5080_/B _6534_/Y _6052_/C VGND VPWR _6535_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_9323_ _9613_/CLK _9323_/D _9646_/SET_B VGND VPWR _9323_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA_89 _8791_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_67 _6680_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_78 _6910_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_9254_ _9681_/CLK _9254_/D _9633_/SET_B VGND VPWR _9254_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_173_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_287 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_596 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6466_ _6461_/Y _5545_/B _6462_/Y _5013_/B _6465_/X VGND VPWR _6473_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_8205_ _8510_/A _8305_/B _8226_/C VGND VPWR _8595_/B VGND VPWR sky130_fd_sc_hd__nor3_2
X_6397_ _9514_/Q VGND VPWR _6397_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_5417_ _9434_/Q _5414_/A _5965_/B1 _5414_/Y VGND VPWR _9434_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_9185_ _9655_/CLK _9185_/D _9633_/SET_B VGND VPWR _9185_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_121_419 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5348_ _9482_/Q _5346_/A _8845_/X _5346_/Y VGND VPWR _9482_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8136_ _8136_/A _8358_/A _8642_/A _8359_/A VGND VPWR _8140_/A VGND VPWR sky130_fd_sc_hd__or4_1
X_8067_ _8067_/A _8539_/A VGND VPWR _8069_/A VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_87_388 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_7018_ _9626_/Q _7018_/B VGND VPWR _7019_/A VGND VPWR sky130_fd_sc_hd__and2b_1
X_5279_ _5279_/A VGND VPWR _5280_/A VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_46_24 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8969_ _8296_/Y _7944_/X _8975_/S VGND VPWR _8969_/X VGND VPWR sky130_fd_sc_hd__mux2_4
XFILLER_102_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_182 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_316 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_298 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_554 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_460 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_86 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_347 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_414 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_108 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_132 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4650_ _4994_/A VGND VPWR _4651_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_174_124 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput10 mask_rev_in[15] VGND VPWR _6085_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput21 mask_rev_in[25] VGND VPWR _6831_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_4581_ _9746_/Q _4579_/A _8845_/X _4579_/Y VGND VPWR _9746_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_6320_ _9325_/Q VGND VPWR _6320_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
Xinput32 mask_rev_in[6] VGND VPWR _6153_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput43 mgmt_gpio_in[16] VGND VPWR _4754_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput54 mgmt_gpio_in[26] VGND VPWR _6680_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_155_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_202 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xinput76 qspi_enabled VGND VPWR _8835_/S VGND VPWR sky130_fd_sc_hd__buf_6
Xinput87 spimemio_flash_io1_do VGND VPWR _8816_/A VGND VPWR sky130_fd_sc_hd__buf_6
Xinput65 mgmt_gpio_in[36] VGND VPWR _8817_/A VGND VPWR sky130_fd_sc_hd__buf_4
Xinput98 sram_ro_data[14] VGND VPWR _6221_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_6251_ _6251_/A VGND VPWR _6251_/Y VGND VPWR sky130_fd_sc_hd__inv_4
XFILLER_115_268 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5202_ _6134_/A _6322_/A _5259_/A _8977_/X VGND VPWR _5203_/A VGND VPWR sky130_fd_sc_hd__a211o_4
X_6182_ _9224_/Q VGND VPWR _6182_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_5133_ _5133_/A _8977_/S VGND VPWR _5156_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_57_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5064_ _8968_/X _9666_/Q _5078_/S VGND VPWR _5065_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_84_358 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_594 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_8823_ _9150_/Q _9790_/Q _9787_/Q VGND VPWR _8823_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_5966_ _9102_/Q _5962_/A _5966_/B1 _5962_/Y VGND VPWR _9102_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8754_ _8754_/A VGND VPWR _8754_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_40_439 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_430 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4917_ _4917_/A _4931_/B VGND VPWR _5382_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_8685_ _8685_/A _8685_/B VGND VPWR _8686_/B VGND VPWR sky130_fd_sc_hd__or2_1
X_5897_ _5960_/A _5897_/B VGND VPWR _5898_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_7705_ _7705_/A VGND VPWR _7706_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_193_411 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7636_ _6935_/Y _7441_/X _6824_/Y _7443_/X _7635_/X VGND VPWR _7643_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_4848_ _9411_/Q VGND VPWR _4848_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_165_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_59 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_9306_ _9440_/CLK _9306_/D _9685_/SET_B VGND VPWR _9306_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_7567_ _6288_/Y _7465_/X _6244_/Y _7467_/X VGND VPWR _7567_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4779_ _9231_/Q VGND VPWR _4779_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_134_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6518_ _6516_/Y _5960_/B _6517_/Y _5089_/B VGND VPWR _6518_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_7498_ _6889_/Y _7471_/X _7150_/A _7473_/X _7497_/X VGND VPWR _7499_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9237_ _9596_/CLK _9237_/D _9528_/SET_B VGND VPWR _9237_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6449_ _9736_/Q VGND VPWR _6449_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_0_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_279 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_599 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9168_ _9203_/CLK _9168_/D _9633_/SET_B VGND VPWR _9168_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_40_csclk clkbuf_2_1_0_csclk/X VGND VPWR _9785_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
X_8119_ _8119_/A VGND VPWR _8546_/A VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_57_12 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_152 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_34 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9099_ _9344_/CLK _9099_/D _9647_/SET_B VGND VPWR _9099_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
Xclkbuf_2_0_0_csclk clkbuf_2_1_0_csclk/A VGND VPWR _9329_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_48_528 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_347 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_200 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_84 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_255 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_88 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_99 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_588 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_439 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_80 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_271 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_282 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_572 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_274 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5820_ _5820_/A VGND VPWR _5820_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_5751_ _9280_/Q _9279_/Q _5751_/C _9277_/Q VGND VPWR _5753_/B VGND VPWR sky130_fd_sc_hd__or4_2
XFILLER_187_260 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8470_ _8470_/A _8470_/B _8698_/A VGND VPWR _8474_/A VGND VPWR sky130_fd_sc_hd__or3_1
X_4702_ _4917_/A _4843_/B VGND VPWR _5013_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_147_124 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5682_ _9263_/Q _5681_/A _8846_/X _5681_/Y VGND VPWR _9263_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7421_ _7421_/A VGND VPWR _7421_/X VGND VPWR sky130_fd_sc_hd__buf_6
XFILLER_163_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4633_ _9050_/Q VGND VPWR _4964_/B VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_118_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7352_ _7352_/A _7352_/B _7352_/C _7352_/D VGND VPWR _7353_/C VGND VPWR sky130_fd_sc_hd__and4_1
X_4564_ _5960_/A _4564_/B VGND VPWR _4565_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_116_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_330 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7283_ _6072_/Y _5728_/X _6059_/Y _7040_/A _7282_/X VGND VPWR _7286_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_6303_ _9098_/Q VGND VPWR _6303_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_6234_ _6232_/Y _5045_/B _6233_/Y _4861_/X VGND VPWR _6234_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4495_ _9784_/Q _4493_/A _8845_/X _4493_/Y VGND VPWR _9784_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_9022_ _9027_/CLK _9022_/D VGND VPWR _9022_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_6165_ _6165_/A VGND VPWR _8955_/S VGND VPWR sky130_fd_sc_hd__clkinv_8
X_5116_ _9636_/Q _5112_/A _5963_/B1 _5112_/Y VGND VPWR _9636_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_6096_ _6096_/A _6096_/B _6096_/C _6096_/D VGND VPWR _6145_/B VGND VPWR sky130_fd_sc_hd__and4_2
XFILLER_111_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5047_ _5047_/A VGND VPWR _5047_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_84_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6998_ _5691_/A _6991_/Y _6996_/Y _6997_/X VGND VPWR _9055_/D VGND VPWR sky130_fd_sc_hd__o22ai_2
X_9786_ _9788_/CLK _9786_/D _9295_/SET_B VGND VPWR _9786_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_8806_ _8806_/A VGND VPWR _8806_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_159_14 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8737_ _8137_/B _8554_/B _8736_/X _8628_/X VGND VPWR _8737_/Y VGND VPWR sky130_fd_sc_hd__o211ai_4
X_5949_ _6052_/A _5949_/B VGND VPWR _5950_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_159_36 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_260 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8668_ _8668_/A _8668_/B _8668_/C _8668_/D VGND VPWR _8699_/D VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_166_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7619_ _4660_/Y _7455_/X _4823_/Y _7457_/X VGND VPWR _7619_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_8599_ _8599_/A _8599_/B _8599_/C _8599_/D VGND VPWR _8696_/A VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_181_414 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_382 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_514 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_343 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_77 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xinput200 wb_sel_i[3] VGND VPWR _7734_/B VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_191_78 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_50 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_372 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_203 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_250 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_294 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_283 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_272 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_236 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_547 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_494 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7970_ _7970_/A VGND VPWR _8098_/A VGND VPWR sky130_fd_sc_hd__buf_6
X_6921_ _9689_/Q VGND VPWR _6921_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_66_188 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6852_ _6843_/Y _5328_/B _6846_/X _6851_/X VGND VPWR _6878_/C VGND VPWR sky130_fd_sc_hd__o211a_1
X_9640_ _4450_/A1 _9640_/D _6146_/A VGND VPWR _9640_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_5803_ _9208_/Q _5799_/A _8925_/A1 _5799_/Y VGND VPWR _9208_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_9571_ _9613_/CLK _9571_/D _9646_/SET_B VGND VPWR _9571_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_50_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8522_ _8064_/C _8064_/B _8521_/Y _8016_/B VGND VPWR _8527_/B VGND VPWR sky130_fd_sc_hd__a31o_1
X_6783_ _6783_/A _6783_/B _6783_/C _6783_/D VGND VPWR _6784_/D VGND VPWR sky130_fd_sc_hd__and4_2
XFILLER_148_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5734_ _7037_/A _5731_/Y _5724_/B _7096_/B VGND VPWR _9248_/D VGND VPWR sky130_fd_sc_hd__o22ai_1
XFILLER_129_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5665_ _9274_/Q _5662_/A _8844_/X _5662_/Y VGND VPWR _9274_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8453_ _8665_/A _8453_/B _8453_/C _8607_/C VGND VPWR _8455_/A VGND VPWR sky130_fd_sc_hd__or4_1
XFILLER_30_291 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7404_ _7466_/A _7476_/C _9255_/Q VGND VPWR _7405_/A VGND VPWR sky130_fd_sc_hd__or3_1
X_4616_ _9725_/Q _4615_/A _5963_/B1 _4615_/Y VGND VPWR _9725_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8384_ _8384_/A _8651_/B VGND VPWR _8385_/B VGND VPWR sky130_fd_sc_hd__nor2_1
X_5596_ _5596_/A VGND VPWR _5596_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7335_ _6732_/Y _7040_/C _6743_/Y _7059_/C VGND VPWR _7335_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_116_374 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4547_ _8810_/A _8812_/A _8813_/A VGND VPWR _4548_/A VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_89_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7266_ _6113_/Y _7086_/X _6074_/Y _7088_/X VGND VPWR _7266_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4478_ _4478_/A VGND VPWR _9789_/D VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_131_344 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6217_ _6212_/Y _5872_/B _6213_/Y _6251_/A _6216_/X VGND VPWR _6236_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_7197_ _8769_/A _7124_/X _6485_/Y _7068_/B _7196_/X VGND VPWR _7198_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9005_ _9598_/Q _8787_/A VGND VPWR mgmt_gpio_out[28] VGND VPWR sky130_fd_sc_hd__ebufn_8
X_6148_ _6148_/A VGND VPWR _6149_/A VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_161_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_604 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6079_ _9527_/Q VGND VPWR _6079_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_53_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_523 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_214 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_191 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_9769_ _9769_/CLK _9769_/D _4628_/A VGND VPWR _9769_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_110_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_67 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_45 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_322 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_160 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_206 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_31 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_75 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_300 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_372 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5450_ _5671_/A _5450_/B VGND VPWR _5451_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_117_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5381_ _9458_/Q _5376_/A _8839_/X _5376_/Y VGND VPWR _9458_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_113_311 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_160 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7120_ _4687_/Y _7059_/D _4877_/Y _7116_/X _7119_/X VGND VPWR _7131_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
Xclkbuf_3_2_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/A VGND VPWR _9280_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_140_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_344 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_19 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7051_ _9248_/Q _7056_/B _7127_/A VGND VPWR _7085_/B VGND VPWR sky130_fd_sc_hd__or3_1
XFILLER_101_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6002_ _9087_/Q _5995_/A _8912_/X _5995_/Y VGND VPWR _9087_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_27_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_155 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7953_ _8195_/A _8632_/A VGND VPWR _7954_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_6904_ _9355_/Q VGND VPWR _6904_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
X_7884_ _7903_/C _8193_/A _8583_/A VGND VPWR _7885_/B VGND VPWR sky130_fd_sc_hd__or3_2
X_6835_ _6833_/Y _5100_/B _6834_/Y _4590_/B VGND VPWR _6835_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_9623_ _9674_/CLK _9623_/D _9633_/SET_B VGND VPWR _9623_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6766_ _6766_/A VGND VPWR _6766_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9554_ _9755_/CLK _9554_/D _9633_/SET_B VGND VPWR _9554_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_148_230 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5717_ _9246_/Q VGND VPWR _5737_/A VGND VPWR sky130_fd_sc_hd__inv_2
X_8505_ _8597_/D _8599_/D _8657_/C _8504_/X VGND VPWR _8509_/A VGND VPWR sky130_fd_sc_hd__or4b_4
XFILLER_136_403 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6697_ _6692_/Y _4491_/B _6693_/Y _5545_/B _6696_/X VGND VPWR _6716_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9485_ _9774_/CLK _9485_/D _7011_/B VGND VPWR _9485_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_40_37 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5648_ _9280_/Q VGND VPWR _5649_/A VGND VPWR sky130_fd_sc_hd__inv_2
X_8436_ _8436_/A _8436_/B VGND VPWR _8487_/A VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_156_37 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5579_ _9323_/Q _5574_/A _8929_/A1 _5574_/Y VGND VPWR _9323_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8367_ _8367_/A _8367_/B VGND VPWR _8578_/C VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_2_427 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_416 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_8298_ _8298_/A VGND VPWR _8600_/A VGND VPWR sky130_fd_sc_hd__inv_2
X_7318_ _6802_/Y _7059_/B _6840_/Y _7068_/C _7317_/X VGND VPWR _7321_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_49_24 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_7249_ _6169_/Y _7097_/X _6168_/Y _7099_/X VGND VPWR _7249_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_104_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_23 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_102 _8805_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_113 input82/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_124 input86/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_14_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_135 _7015_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_157 _5121_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_146 _7626_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_14_523 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_33 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_168 _6819_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_179 _9404_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_14_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_358 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_210 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xinput8 mask_rev_in[13] VGND VPWR input8/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_24_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4950_ _9092_/Q _9091_/Q _6022_/C VGND VPWR _4951_/B VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_51_139 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4881_ _4874_/Y _4602_/B _4875_/Y _5110_/B _4880_/X VGND VPWR _4896_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_32_342 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6620_ _6615_/Y _5336_/B _8793_/A _5393_/B _6619_/X VGND VPWR _6627_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_6551_ _9644_/Q VGND VPWR _6551_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_5502_ _9376_/Q _5498_/A _8925_/A1 _5498_/Y VGND VPWR _9376_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_9270_ _9535_/CLK _9270_/D _9528_/SET_B VGND VPWR _9270_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6482_ _6477_/Y _5768_/B _8757_/A _5679_/B _6481_/X VGND VPWR _6501_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_133_406 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5433_ _5433_/A VGND VPWR _5433_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_8221_ _8510_/A _8498_/A _8640_/A VGND VPWR _8223_/A VGND VPWR sky130_fd_sc_hd__or3_1
Xoutput301 _9045_/Q VGND VPWR pwr_ctrl_out[1] VGND VPWR sky130_fd_sc_hd__buf_2
X_5364_ _9469_/Q _5357_/A _8840_/X _5357_/Y VGND VPWR _9469_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8152_ _8152_/A _8674_/A VGND VPWR _8154_/A VGND VPWR sky130_fd_sc_hd__or2_1
Xoutput323 _9769_/Q VGND VPWR sram_ro_addr[7] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput334 _9028_/Q VGND VPWR wb_dat_o[16] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput312 _7019_/X VGND VPWR spimemio_flash_io0_di VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_126_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7103_ _4732_/Y _7059_/B _4744_/Y _7068_/C _7102_/X VGND VPWR _7108_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
Xoutput356 _9027_/Q VGND VPWR wb_dat_o[7] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput345 _9038_/Q VGND VPWR wb_dat_o[26] VGND VPWR sky130_fd_sc_hd__buf_2
X_5295_ _9517_/Q _5292_/A _5965_/B1 _5292_/Y VGND VPWR _9517_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8083_ _8185_/A _8187_/A _8083_/C VGND VPWR _8086_/A VGND VPWR sky130_fd_sc_hd__and3_1
X_7034_ _7125_/A _7111_/C VGND VPWR _7115_/B VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_95_581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_8985_ _8985_/A _8747_/A VGND VPWR mgmt_gpio_out[8] VGND VPWR sky130_fd_sc_hd__ebufn_8
XFILLER_55_478 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7936_ _8476_/A _7936_/B VGND VPWR _7936_/X VGND VPWR sky130_fd_sc_hd__or2_1
X_7867_ _7959_/A _8528_/A _8583_/A _7894_/B VGND VPWR _7868_/A VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_143_7 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_375 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9606_ _9617_/CLK _9606_/D _9295_/SET_B VGND VPWR _9606_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6818_ _9443_/Q VGND VPWR _6818_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
X_7798_ _8510_/A _8188_/B VGND VPWR _8651_/A VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_149_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9537_ _9768_/CLK _9537_/D _4628_/A VGND VPWR _9537_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6749_ _9046_/Q VGND VPWR _6749_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
XFILLER_167_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9468_ _9535_/CLK _9468_/D _9528_/SET_B VGND VPWR _9468_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_164_575 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_406 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8419_ _8552_/A _8401_/B _8415_/X _8418_/Y VGND VPWR _8419_/X VGND VPWR sky130_fd_sc_hd__o211a_1
X_9399_ _9758_/CLK _9399_/D _7011_/B VGND VPWR _9399_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_183_79 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_275 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_426 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_106 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_320 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_92 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_70 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_100 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_531 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_91 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_6 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_548 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5080_ _5259_/A _5080_/B VGND VPWR _5081_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_96_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_250 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_423 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_63 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5982_ _9092_/Q _5981_/X _7008_/A _5985_/B VGND VPWR _9092_/D VGND VPWR sky130_fd_sc_hd__o22a_1
X_8770_ _8770_/A VGND VPWR _8770_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_7721_ _7721_/A VGND VPWR _7722_/B VGND VPWR sky130_fd_sc_hd__inv_2
X_4933_ _4924_/Y _5366_/B _4926_/Y _5306_/B _4932_/X VGND VPWR _4934_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_20_301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7652_ _6731_/Y _7425_/X _7649_/X _7651_/X VGND VPWR _7662_/C VGND VPWR sky130_fd_sc_hd__o211a_1
X_4864_ _4864_/A _4864_/B _4864_/C _4864_/D VGND VPWR _4935_/B VGND VPWR sky130_fd_sc_hd__and4_1
XANTENNA_13 _7287_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_4795_ _9627_/Q VGND VPWR _4795_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7583_ _6154_/Y _7455_/X _6157_/Y _7457_/X VGND VPWR _7583_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_6603_ _9479_/Q VGND VPWR _8775_/A VGND VPWR sky130_fd_sc_hd__clkinv_8
XANTENNA_24 _7680_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_46 _4910_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_57 _6252_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_35 _4788_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_6534_ _9047_/Q VGND VPWR _6534_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9322_ _9352_/CLK _9322_/D _9646_/SET_B VGND VPWR _9322_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XANTENNA_79 _7133_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_68 _6716_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_180_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_244 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6465_ _6463_/Y _5045_/B _6464_/Y _5080_/B VGND VPWR _6465_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_9253_ _9681_/CLK _9253_/D _9633_/SET_B VGND VPWR _9253_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_133_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_299 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5416_ _9435_/Q _5414_/A _5964_/B1 _5414_/Y VGND VPWR _9435_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8204_ _8204_/A _8640_/A VGND VPWR _8678_/A VGND VPWR sky130_fd_sc_hd__nor2_1
X_9184_ _9613_/CLK _9184_/D _9646_/SET_B VGND VPWR _9184_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6396_ _9480_/Q VGND VPWR _6396_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
XFILLER_161_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5347_ _9483_/Q _5346_/A _8846_/X _5346_/Y VGND VPWR _9483_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8135_ _8137_/B _8378_/B VGND VPWR _8359_/A VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_87_323 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8066_ _8282_/B _8518_/A _8282_/C VGND VPWR _8539_/A VGND VPWR sky130_fd_sc_hd__and3_1
X_5278_ _5545_/A _5278_/B VGND VPWR _5279_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_7017_ _7017_/A VGND VPWR _7017_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_87_356 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_8968_ _7751_/X _8968_/A1 _8975_/S VGND VPWR _8968_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_43_437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7919_ _8521_/B _8254_/B VGND VPWR _8320_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_102_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_8899_ _7712_/X _9083_/Q _9051_/Q VGND VPWR _8899_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_168_133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_103 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_328 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_244 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_50 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_434 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_144 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_136 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4580_ _9747_/Q _4579_/A _8846_/X _4579_/Y VGND VPWR _9747_/D VGND VPWR sky130_fd_sc_hd__a22o_1
Xinput11 mask_rev_in[16] VGND VPWR _4906_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput22 mask_rev_in[26] VGND VPWR _6726_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_162_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xinput33 mask_rev_in[7] VGND VPWR _6087_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput44 mgmt_gpio_in[17] VGND VPWR _6903_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput55 mgmt_gpio_in[27] VGND VPWR _6531_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput88 spimemio_flash_io1_oeb VGND VPWR _7015_/B VGND VPWR sky130_fd_sc_hd__buf_6
Xinput77 ser_tx VGND VPWR input77/X VGND VPWR sky130_fd_sc_hd__buf_4
Xinput66 mgmt_gpio_in[37] VGND VPWR _8818_/A VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_115_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6250_ _9637_/Q VGND VPWR _6250_/Y VGND VPWR sky130_fd_sc_hd__inv_2
Xinput99 sram_ro_data[15] VGND VPWR _6099_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_6181_ _9300_/Q VGND VPWR _7260_/A VGND VPWR sky130_fd_sc_hd__inv_2
X_5201_ _9578_/Q _5193_/Y _8849_/X _5193_/A VGND VPWR _9578_/D VGND VPWR sky130_fd_sc_hd__o22a_1
X_5132_ _7022_/B VGND VPWR _8977_/S VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_123_19 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5063_ _5063_/A VGND VPWR _5078_/S VGND VPWR sky130_fd_sc_hd__clkbuf_4
X_8822_ _9176_/Q _9079_/Q _9787_/Q VGND VPWR _8822_/X VGND VPWR sky130_fd_sc_hd__mux2_4
X_5965_ _9103_/Q _5962_/A _5965_/B1 _5962_/Y VGND VPWR _9103_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8753_ _8753_/A VGND VPWR _8754_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_52_278 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_610 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4916_ _9450_/Q VGND VPWR _4916_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_8684_ _8115_/Y _8625_/B _8405_/A _8683_/X _8629_/B VGND VPWR _8689_/A VGND VPWR
+ sky130_fd_sc_hd__a2111o_2
X_5896_ _8924_/X _6997_/A _5895_/Y _5896_/B1 _9138_/Q VGND VPWR _9138_/D VGND VPWR
+ sky130_fd_sc_hd__a32o_2
X_7704_ _7704_/A VGND VPWR _7704_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_7635_ _6867_/Y _7445_/X _6872_/Y _7447_/X VGND VPWR _7635_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4847_ _4876_/B _4931_/B VGND VPWR _5267_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_20_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9305_ _9440_/CLK _9305_/D _9685_/SET_B VGND VPWR _9305_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_7566_ _6298_/Y _7451_/X _6274_/Y _7453_/X _7565_/X VGND VPWR _7571_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_4778_ _4769_/Y _5089_/B _4771_/Y _5583_/B _4777_/X VGND VPWR _4790_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_134_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6517_ _9649_/Q VGND VPWR _6517_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7497_ _6823_/Y _7475_/X _6926_/Y _7477_/X VGND VPWR _7497_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_164_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_320 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6448_ _6434_/Y _5864_/B _6437_/X _6443_/X _6447_/X VGND VPWR _6474_/C VGND VPWR
+ sky130_fd_sc_hd__o2111a_1
X_9236_ _9371_/CLK _9236_/D _9295_/SET_B VGND VPWR _9236_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_9167_ _9203_/CLK _9167_/D _9633_/SET_B VGND VPWR _9167_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6379_ _9268_/Q VGND VPWR _6379_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_121_228 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8118_ _8394_/A _8379_/B _8117_/A VGND VPWR _8118_/X VGND VPWR sky130_fd_sc_hd__or3b_1
XFILLER_0_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_9098_ _9344_/CLK _9098_/D _9647_/SET_B VGND VPWR _9098_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_87_164 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_486 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8049_ _8097_/B _8554_/A _8048_/Y VGND VPWR _8053_/A VGND VPWR sky130_fd_sc_hd__o21ba_1
XFILLER_57_46 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_415 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_318 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_67 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_102 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_330 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_239 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_294 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_307 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_584 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_554 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5750_ _9056_/Q _8819_/X VGND VPWR _5750_/Y VGND VPWR sky130_fd_sc_hd__nor2_2
X_4701_ _9688_/Q VGND VPWR _4701_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_5681_ _5681_/A VGND VPWR _5681_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_175_423 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_294 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4632_ _9697_/Q VGND VPWR _5214_/A VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_187_272 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7420_ _7474_/C _7466_/A _7474_/D VGND VPWR _7421_/A VGND VPWR sky130_fd_sc_hd__or3_1
XFILLER_175_456 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_467 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4563_ _4891_/A _6158_/A VGND VPWR _4564_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_7351_ _6700_/Y _7124_/X _6701_/Y _7068_/B _7350_/X VGND VPWR _7352_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_2
XFILLER_116_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4494_ _9785_/Q _4493_/A _8846_/X _4493_/Y VGND VPWR _9785_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7282_ _7282_/A _7392_/B VGND VPWR _7282_/X VGND VPWR sky130_fd_sc_hd__or2_1
X_6302_ _9156_/Q VGND VPWR _6302_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_9021_ _9027_/CLK _9021_/D VGND VPWR _9021_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_6233_ _6233_/A VGND VPWR _6233_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
X_6164_ _9404_/Q VGND VPWR _6164_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_111_250 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5115_ _9637_/Q _5112_/A _8844_/X _5112_/Y VGND VPWR _9637_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_6095_ _6090_/Y _5458_/B _6091_/Y _5496_/B _6094_/X VGND VPWR _6096_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_57_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5046_ _5046_/A VGND VPWR _5047_/A VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_27_38 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_510 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6997_ _6997_/A _8819_/X _6997_/C VGND VPWR _6997_/X VGND VPWR sky130_fd_sc_hd__or3_2
X_9785_ _9785_/CLK _9785_/D _9779_/SET_B VGND VPWR _9785_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_8805_ _8805_/A input1/X VGND VPWR _8806_/A VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_43_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_215 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5948_ _9114_/Q _5943_/A _5967_/B1 _5943_/Y VGND VPWR _9114_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8736_ _8164_/A _8550_/A _8029_/X _8411_/Y VGND VPWR _8736_/X VGND VPWR sky130_fd_sc_hd__o211a_1
XFILLER_166_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_272 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5879_ _9154_/Q _5874_/A _8929_/A1 _5874_/Y VGND VPWR _9154_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8667_ _8667_/A _8667_/B VGND VPWR _8668_/B VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_166_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7618_ _4722_/Y _7441_/X _4865_/Y _7443_/X _7617_/X VGND VPWR _7625_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_8598_ _8695_/D _8659_/C _8727_/A _8657_/D VGND VPWR _8601_/A VGND VPWR sky130_fd_sc_hd__or4_2
XFILLER_181_426 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7549_ _6367_/Y _7465_/X _6427_/Y _7467_/X VGND VPWR _7549_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_5_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_52 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9219_ _9695_/CLK _9219_/D _9779_/SET_B VGND VPWR _9219_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_108_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_526 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_322 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xinput201 wb_stb_i VGND VPWR input201/X VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_191_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_399 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_62 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_148 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_215 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_384 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_251 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_240 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_295 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_284 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_262 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_70 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6920_ _9178_/Q VGND VPWR _6920_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_6851_ _6847_/Y _4868_/X _6848_/Y _5298_/B _6850_/X VGND VPWR _6851_/X VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_50_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5802_ _9209_/Q _5799_/A _8844_/X _5799_/Y VGND VPWR _9209_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_9570_ _9613_/CLK _9570_/D _9646_/SET_B VGND VPWR _9570_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_22_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6782_ _6778_/Y _4893_/X _4949_/Y _6165_/A _6781_/X VGND VPWR _6783_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_8521_ _8521_/A _8521_/B VGND VPWR _8521_/Y VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_188_581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5733_ _9248_/Q _7056_/B _7104_/A VGND VPWR _7096_/B VGND VPWR sky130_fd_sc_hd__or3_2
XFILLER_148_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5664_ _9275_/Q _5662_/A _8845_/X _5662_/Y VGND VPWR _9275_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8452_ _8238_/A _7864_/X _8097_/B _8130_/B VGND VPWR _8607_/C VGND VPWR sky130_fd_sc_hd__o22ai_1
XFILLER_148_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4615_ _4615_/A VGND VPWR _4615_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7403_ _7413_/A _7406_/B VGND VPWR _7476_/C VGND VPWR sky130_fd_sc_hd__or2_4
X_8383_ _8636_/A _8514_/A VGND VPWR _8651_/B VGND VPWR sky130_fd_sc_hd__or2_1
X_5595_ _5595_/A VGND VPWR _5596_/A VGND VPWR sky130_fd_sc_hd__clkbuf_2
X_4546_ _9068_/Q VGND VPWR _8813_/A VGND VPWR sky130_fd_sc_hd__inv_2
X_7334_ _6730_/Y _7082_/X _6705_/Y _7084_/X _7333_/X VGND VPWR _7353_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_190_267 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_386 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7265_ _7265_/A _7265_/B _7265_/C VGND VPWR _7265_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
X_4477_ _8839_/X _9789_/Q _4477_/S VGND VPWR _4478_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_7196_ _8783_/A _7126_/X _8781_/A _7128_/X VGND VPWR _7196_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_6216_ _6214_/Y _4577_/B _6215_/Y _5013_/B VGND VPWR _6216_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_9004_ _9597_/Q _8785_/A VGND VPWR mgmt_gpio_out[27] VGND VPWR sky130_fd_sc_hd__ebufn_8
X_6147_ _6974_/B _6147_/B VGND VPWR _6148_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_85_443 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6078_ _9483_/Q VGND VPWR _6078_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
XFILLER_72_126 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5029_ _9685_/Q _5026_/A _8841_/X _5026_/Y VGND VPWR _9685_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_186_518 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_9768_ _9768_/CLK _9768_/D _4628_/A VGND VPWR _9768_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_8719_ _8719_/A _8719_/B _8719_/C VGND VPWR _8731_/C VGND VPWR sky130_fd_sc_hd__or3_2
X_9699_ _9709_/CLK _9699_/D _4995_/X VGND VPWR _9699_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_21_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_44 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_334 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_83 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_218 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_43 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_94 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_87 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_543 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_384 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_192 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5380_ _9459_/Q _5376_/A _8930_/A1 _5376_/Y VGND VPWR _9459_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_172_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_356 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7050_ _7050_/A VGND VPWR _7059_/A VGND VPWR sky130_fd_sc_hd__buf_8
XFILLER_101_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6001_ _6001_/A VGND VPWR _6001_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_140_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_19 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7952_ _7952_/A VGND VPWR _8437_/B VGND VPWR sky130_fd_sc_hd__clkbuf_4
X_6903_ _6903_/A VGND VPWR _6903_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7883_ _8397_/A VGND VPWR _7886_/B VGND VPWR sky130_fd_sc_hd__inv_2
X_9622_ _9674_/CLK _9622_/D _9633_/SET_B VGND VPWR _9622_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_23_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_535 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6834_ _9733_/Q VGND VPWR _6834_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_50_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6765_ _6760_/Y _5306_/B _6761_/Y _5240_/B _6764_/X VGND VPWR _6783_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9553_ _9639_/CLK _9553_/D _9757_/SET_B VGND VPWR _9553_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_5716_ _9249_/Q VGND VPWR _5725_/B VGND VPWR sky130_fd_sc_hd__inv_2
X_8504_ _8501_/X _8504_/B _8504_/C VGND VPWR _8504_/X VGND VPWR sky130_fd_sc_hd__and3b_1
X_9484_ _9777_/CLK _9484_/D _9633_/SET_B VGND VPWR _9484_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_136_415 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_607 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6696_ _6694_/Y _5267_/B _6695_/Y _5442_/B VGND VPWR _6696_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_8435_ _8636_/B _8435_/B VGND VPWR _8436_/B VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_136_448 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_49 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5647_ _5647_/A _5651_/A _5751_/C VGND VPWR _5647_/X VGND VPWR sky130_fd_sc_hd__or3_2
XFILLER_123_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5578_ _9324_/Q _5574_/A _8925_/A1 _5574_/Y VGND VPWR _9324_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8366_ _8685_/B _8493_/B VGND VPWR _8675_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_144_470 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4529_ _9767_/Q _4526_/A _8844_/X _4526_/Y VGND VPWR _9767_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7317_ _6826_/Y _7079_/B _6928_/Y _7059_/A VGND VPWR _7317_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_8297_ _8651_/A _8606_/B VGND VPWR _8673_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_7248_ _6175_/Y _7048_/B _6215_/Y _7077_/A _7247_/X VGND VPWR _7255_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_172_48 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7179_ _8757_/A _7077_/C _6491_/Y _7077_/D _7178_/X VGND VPWR _7179_/X VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_105_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA_114 input85/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_103 input37/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_125 input86/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_121_52 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_147 _7698_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_158 _4814_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_136 input91/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_81_490 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_169 _6819_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_81_45 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_554 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_462 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_8 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_443 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xinput9 mask_rev_in[14] VGND VPWR input9/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_64_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_232 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_120 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4880_ _4877_/Y _5496_/B _4879_/Y _4517_/A VGND VPWR _4880_/X VGND VPWR sky130_fd_sc_hd__o22a_2
XFILLER_32_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_354 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_359 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6550_ _9539_/Q VGND VPWR _6550_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_5501_ _9377_/Q _5498_/A _8844_/X _5498_/Y VGND VPWR _9377_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_6481_ _6479_/Y _5916_/B _6480_/Y _5564_/B VGND VPWR _6481_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_10_19 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8220_ _8566_/B _8214_/Y _8217_/Y _8110_/C _8219_/Y VGND VPWR _8224_/C VGND VPWR
+ sky130_fd_sc_hd__o32a_2
X_5432_ _5432_/A VGND VPWR _5433_/A VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_105_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_418 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5363_ _9470_/Q _5357_/A _8841_/X _5357_/Y VGND VPWR _9470_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8151_ _8552_/A _8640_/B VGND VPWR _8674_/A VGND VPWR sky130_fd_sc_hd__nor2_1
Xoutput302 _9046_/Q VGND VPWR pwr_ctrl_out[2] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput324 _9760_/Q VGND VPWR sram_ro_clk VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput335 _9029_/Q VGND VPWR wb_dat_o[17] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput313 _7021_/X VGND VPWR spimemio_flash_io1_di VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_113_131 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7102_ _4833_/Y _7079_/B _4726_/Y _7059_/A VGND VPWR _7102_/X VGND VPWR sky130_fd_sc_hd__o22a_1
Xoutput357 _9012_/Q VGND VPWR wb_dat_o[8] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput346 _9039_/Q VGND VPWR wb_dat_o[27] VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_87_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5294_ _9518_/Q _5292_/A _5964_/B1 _5292_/Y VGND VPWR _9518_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8082_ _8082_/A _8186_/A VGND VPWR _8083_/C VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_101_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_7033_ _7033_/A VGND VPWR _7040_/B VGND VPWR sky130_fd_sc_hd__buf_8
XFILLER_142_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8984_ _9585_/Q _7699_/A VGND VPWR mgmt_gpio_out[7] VGND VPWR sky130_fd_sc_hd__ebufn_8
X_7935_ _8376_/A _7935_/B VGND VPWR _7936_/B VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_82_276 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7866_ _7866_/A VGND VPWR _8319_/A VGND VPWR sky130_fd_sc_hd__buf_2
X_9605_ _9617_/CLK _9605_/D _9295_/SET_B VGND VPWR _9605_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6817_ _6817_/A VGND VPWR _6817_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_23_387 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_9536_ _9768_/CLK _9536_/D _4628_/A VGND VPWR _9536_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_7797_ _7797_/A VGND VPWR _8188_/B VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_149_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_7 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6748_ _9288_/Q VGND VPWR _6748_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_183_307 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_551 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9467_ _9514_/CLK _9467_/D _4628_/A VGND VPWR _9467_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6679_ _6679_/A VGND VPWR _6679_/Y VGND VPWR sky130_fd_sc_hd__inv_4
X_8418_ _8686_/A VGND VPWR _8418_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9398_ _9758_/CLK _9398_/D _7011_/B VGND VPWR _9398_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_151_204 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8349_ _8640_/A _8349_/B VGND VPWR _8352_/B VGND VPWR sky130_fd_sc_hd__or2_2
XFILLER_4_5 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_67 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_243 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_82 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_60 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_112 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_60 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_212 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_571 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_70 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_112 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_75 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_435 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5981_ _9090_/Q _5981_/B _9091_/Q VGND VPWR _5981_/X VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_17_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_4932_ _4928_/Y _5458_/B _4930_/Y _5328_/B VGND VPWR _4932_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_7720_ _9087_/Q _7719_/B _7721_/A VGND VPWR _7720_/X VGND VPWR sky130_fd_sc_hd__o21a_1
XFILLER_177_101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7651_ _6743_/Y _7430_/X _6725_/Y _7432_/X _7650_/X VGND VPWR _7651_/X VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_4863_ _4855_/Y _5317_/B _4857_/Y _4491_/B _4862_/X VGND VPWR _4864_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_6602_ _6587_/Y _5480_/B _6590_/X _6596_/X _6601_/X VGND VPWR _6628_/C VGND VPWR
+ sky130_fd_sc_hd__o2111a_1
XANTENNA_14 _7309_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_4794_ _4911_/A _4929_/A VGND VPWR _5240_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_7582_ _6183_/Y _7441_/X _6195_/Y _7443_/X _7581_/X VGND VPWR _7589_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XANTENNA_36 _4804_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_25 _5259_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_47 _4922_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_6533_ _9657_/Q VGND VPWR _6533_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9321_ _9352_/CLK _9321_/D _9646_/SET_B VGND VPWR _9321_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XANTENNA_58 _6256_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_69 _6706_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_6464_ _9658_/Q VGND VPWR _6464_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9252_ _9278_/CLK _9252_/D _9633_/SET_B VGND VPWR _9252_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_8203_ _8203_/A VGND VPWR _8476_/B VGND VPWR sky130_fd_sc_hd__inv_2
X_5415_ _9436_/Q _5414_/A _8843_/X _5414_/Y VGND VPWR _9436_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_161_568 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6395_ _6390_/Y _5355_/B _6391_/Y _5374_/B _6394_/X VGND VPWR _6408_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9183_ _9613_/CLK _9183_/D _9646_/SET_B VGND VPWR _9183_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_5346_ _5346_/A VGND VPWR _5346_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_114_440 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_8134_ _8137_/B _8640_/B VGND VPWR _8642_/A VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_99_184 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_495 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5277_ _9528_/Q _5269_/A _8839_/X _5269_/Y VGND VPWR _9528_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8065_ _8065_/A _8703_/C VGND VPWR _8067_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_7016_ _7016_/A VGND VPWR _7017_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_55_232 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8967_ _7749_/X _8967_/A1 _8975_/S VGND VPWR _8967_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_7918_ _8515_/B _8254_/B VGND VPWR _8492_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_102_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_8898_ _9617_/Q _8846_/X _8930_/S VGND VPWR _8898_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_7849_ _8379_/D _8379_/B _8394_/C _8195_/A VGND VPWR _7850_/A VGND VPWR sky130_fd_sc_hd__or4_1
XFILLER_178_47 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9519_ _9771_/CLK _9519_/D _4628_/A VGND VPWR _9519_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_109_256 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_576 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_2_1_0_mgmt_gpio_in[4] clkbuf_2_1_0_mgmt_gpio_in[4]/A VGND VPWR _9709_/CLK
+ VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_30_622 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_156 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput12 mask_rev_in[17] VGND VPWR _6794_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput34 mask_rev_in[8] VGND VPWR input34/X VGND VPWR sky130_fd_sc_hd__buf_2
Xinput45 mgmt_gpio_in[18] VGND VPWR input45/X VGND VPWR sky130_fd_sc_hd__buf_2
Xinput23 mask_rev_in[27] VGND VPWR _6624_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput56 mgmt_gpio_in[28] VGND VPWR input56/X VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
Xinput78 spi_csb VGND VPWR input78/X VGND VPWR sky130_fd_sc_hd__buf_6
Xinput67 mgmt_gpio_in[3] VGND VPWR _4629_/C VGND VPWR sky130_fd_sc_hd__buf_12
Xinput89 spimemio_flash_io2_do VGND VPWR input89/X VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_6_350 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5200_ _9579_/Q _5193_/Y _8903_/X _5193_/A VGND VPWR _9579_/D VGND VPWR sky130_fd_sc_hd__o22a_1
X_6180_ _6178_/Y _5679_/B _6179_/Y _5660_/B VGND VPWR _6187_/B VGND VPWR sky130_fd_sc_hd__o22a_1
X_5131_ _9048_/Q _4951_/B _9708_/Q _9626_/Q _4951_/Y VGND VPWR _9626_/D VGND VPWR
+ sky130_fd_sc_hd__a32o_1
X_5062_ _5062_/A _5062_/B _5062_/C _5062_/D VGND VPWR _5063_/A VGND VPWR sky130_fd_sc_hd__or4_1
X_8821_ _9057_/Q _9078_/Q _9787_/Q VGND VPWR _8821_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_25_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8752_ _8752_/A VGND VPWR _8752_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_80_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5964_ _9104_/Q _5962_/A _5964_/B1 _5962_/Y VGND VPWR _9104_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7703_ _7703_/A VGND VPWR _7704_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_178_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5895_ _8959_/X VGND VPWR _5895_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_4915_ _6086_/B _4931_/B VGND VPWR _5420_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_8683_ _8683_/A _8683_/B VGND VPWR _8683_/X VGND VPWR sky130_fd_sc_hd__or2_1
X_4846_ _9528_/Q VGND VPWR _4846_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7634_ _6929_/Y _7425_/X _7631_/X _7633_/X VGND VPWR _7644_/C VGND VPWR sky130_fd_sc_hd__o211a_1
XFILLER_32_17 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7565_ _6277_/Y _7455_/X _6314_/Y _7457_/X VGND VPWR _7565_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4777_ _4773_/Y _5045_/B _4775_/Y _5916_/B VGND VPWR _4777_/X VGND VPWR sky130_fd_sc_hd__o22a_2
X_9304_ _9440_/CLK _9304_/D _9685_/SET_B VGND VPWR _9304_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6516_ _9104_/Q VGND VPWR _6516_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
XFILLER_134_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7496_ _6920_/Y _7461_/X _6832_/Y _7463_/X _7495_/X VGND VPWR _7499_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_161_332 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6447_ _6444_/Y _4832_/X _6445_/Y _5100_/B _6446_/Y VGND VPWR _6447_/X VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9235_ _9508_/CLK _9235_/D _9528_/SET_B VGND VPWR _9235_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_9166_ _9203_/CLK _9166_/D _9633_/SET_B VGND VPWR _9166_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6378_ _9285_/Q VGND VPWR _7392_/A VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_102_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8117_ _8117_/A _8117_/B VGND VPWR _8393_/A VGND VPWR sky130_fd_sc_hd__nand2_2
X_5329_ _5329_/A VGND VPWR _5330_/A VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_0_548 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_454 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9097_ _9501_/CLK _9097_/D _9647_/SET_B VGND VPWR _9097_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_8048_ _8554_/A _8389_/A _8047_/X VGND VPWR _8048_/Y VGND VPWR sky130_fd_sc_hd__o21ai_2
XFILLER_57_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_498 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_35 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_340 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_10 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_192 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_408 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_110 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_7 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_596 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_224 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_566 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4700_ _4931_/A _4843_/B VGND VPWR _5897_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_5680_ _5680_/A VGND VPWR _5681_/A VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_15_493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_90 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4631_ _6050_/A VGND VPWR _4994_/A VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_8_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_502 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7350_ _6652_/Y _7126_/X _6762_/Y _7128_/X VGND VPWR _7350_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4562_ _4562_/A VGND VPWR _9756_/D VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_6301_ _9223_/Q VGND VPWR _6301_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_4493_ _4493_/A VGND VPWR _4493_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7281_ _6127_/Y _7059_/D _6091_/Y _7116_/X _7280_/X VGND VPWR _7286_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_131_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9020_ _9027_/CLK _9020_/D VGND VPWR _9020_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_6232_ _9673_/Q VGND VPWR _6232_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_6163_ _9318_/Q VGND VPWR _6163_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_111_262 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5114_ _9638_/Q _5112_/A _8845_/X _5112_/Y VGND VPWR _9638_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_6094_ _6092_/Y _4577_/B _6093_/Y _4907_/X VGND VPWR _6094_/X VGND VPWR sky130_fd_sc_hd__o22a_2
X_5045_ _5960_/A _5045_/B VGND VPWR _5046_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_53_522 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_9784_ _9785_/CLK _9784_/D _9779_/SET_B VGND VPWR _9784_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_8804_ _8804_/A VGND VPWR _8804_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_6996_ _7075_/A _7094_/B VGND VPWR _6996_/Y VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_43_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5947_ _9115_/Q _5943_/A _8930_/A1 _5943_/Y VGND VPWR _9115_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8735_ _8735_/A _8735_/B _8735_/C _8735_/D VGND VPWR _8735_/X VGND VPWR sky130_fd_sc_hd__or4_1
XFILLER_33_290 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8666_ _8666_/A _8666_/B _8666_/C _8666_/D VGND VPWR _8735_/D VGND VPWR sky130_fd_sc_hd__or4_2
XFILLER_178_284 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7617_ _4848_/Y _7445_/X _4918_/Y _7447_/X VGND VPWR _7617_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_5878_ _9155_/Q _5874_/A _8925_/A1 _5874_/Y VGND VPWR _9155_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_193_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4829_ _4821_/Y _4822_/X _4823_/Y _5100_/B _4828_/X VGND VPWR _4830_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_8597_ _8597_/A _8597_/B _8597_/C _8597_/D VGND VPWR _8657_/D VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_175_26 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7548_ _6353_/Y _7451_/X _6415_/Y _7453_/X _7547_/X VGND VPWR _7553_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_4_128 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_438 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7479_ _4668_/Y _7471_/X _7121_/A _7473_/X _7478_/X VGND VPWR _7480_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_107_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_9218_ _9379_/CLK _9218_/D _9646_/SET_B VGND VPWR _9218_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_134_376 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_64 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9149_ _9280_/CLK _9149_/D _9757_/SET_B VGND VPWR _9149_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
Xinput202 wb_we_i VGND VPWR _7734_/A VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_102_262 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_102 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_74 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_40 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_252 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_230 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_274 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_263 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_435 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_296 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_82 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_608 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_324 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xhold1 hold1/A VGND VPWR hold1/X VGND VPWR sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_47_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_544 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6850_ _9787_/Q _6251_/Y _6849_/Y _6086_/X VGND VPWR _6850_/X VGND VPWR sky130_fd_sc_hd__o2bb2a_2
X_6781_ _6779_/Y _5290_/B _6780_/Y _5328_/B VGND VPWR _6781_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_5801_ _9210_/Q _5799_/A _8845_/X _5799_/Y VGND VPWR _9210_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8520_ _8472_/Y _8517_/Y _8518_/X _8444_/B VGND VPWR _8612_/B VGND VPWR sky130_fd_sc_hd__a31o_1
X_5732_ _9249_/Q _5731_/Y _5724_/Y VGND VPWR _9249_/D VGND VPWR sky130_fd_sc_hd__o21ba_1
Xclkbuf_1_1_1_mgmt_gpio_in[4] clkbuf_1_1_1_mgmt_gpio_in[4]/A VGND VPWR clkbuf_2_3_0_mgmt_gpio_in[4]/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_2
X_5663_ _9276_/Q _5662_/A _8846_/X _5662_/Y VGND VPWR _9276_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8451_ _8451_/A _8683_/A VGND VPWR _8453_/C VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_135_107 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7402_ _9254_/Q VGND VPWR _7413_/A VGND VPWR sky130_fd_sc_hd__inv_2
X_5594_ _5671_/A _5594_/B VGND VPWR _5595_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_8382_ _8705_/A _8382_/B VGND VPWR _8384_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_4614_ _4614_/A VGND VPWR _4615_/A VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_116_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4545_ _9067_/Q VGND VPWR _8812_/A VGND VPWR sky130_fd_sc_hd__inv_2
X_7333_ _6645_/Y _7077_/C _6756_/Y _7077_/D _7332_/X VGND VPWR _7333_/X VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_190_279 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_398 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4476_ _4787_/A _4891_/A _5259_/A VGND VPWR _4477_/S VGND VPWR sky130_fd_sc_hd__or3_1
X_7264_ _7264_/A _7264_/B _7264_/C _7264_/D VGND VPWR _7265_/C VGND VPWR sky130_fd_sc_hd__and4_1
X_9003_ _9596_/Q _8783_/A VGND VPWR mgmt_gpio_out[26] VGND VPWR sky130_fd_sc_hd__ebufn_8
XFILLER_89_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6215_ _9694_/Q VGND VPWR _6215_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7195_ _8793_/A _5728_/X _7705_/A _7040_/A _7194_/X VGND VPWR _7198_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_6146_ _6146_/A VGND VPWR _6974_/B VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_85_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_38 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6077_ _6072_/Y _5393_/B _6073_/Y _5317_/B _6076_/X VGND VPWR _6096_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_38_382 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5028_ _9686_/Q _5026_/A _8842_/X _5026_/Y VGND VPWR _9686_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_72_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_7 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6979_ _6326_/Y _6976_/A _9017_/Q _6976_/Y VGND VPWR _9017_/D VGND VPWR sky130_fd_sc_hd__o22a_1
X_9767_ _9769_/CLK _9767_/D _9757_/SET_B VGND VPWR _9767_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_9_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9698_ _9709_/CLK _9698_/D _5000_/X VGND VPWR _9698_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_8718_ _8347_/X _8717_/X _8223_/B _8312_/D VGND VPWR _8719_/B VGND VPWR sky130_fd_sc_hd__o211ai_1
XFILLER_166_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8649_ _8722_/A _8681_/B _8720_/B VGND VPWR _8649_/Y VGND VPWR sky130_fd_sc_hd__nor3_1
XFILLER_186_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_310 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_78 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_346 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_455 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_555 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_132 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_368 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6000_ _6040_/A VGND VPWR _6001_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_79_260 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_7951_ _8525_/A _8538_/B _8538_/C _8084_/A VGND VPWR _7952_/A VGND VPWR sky130_fd_sc_hd__or4_1
X_7882_ _8394_/D _8097_/B VGND VPWR _8397_/A VGND VPWR sky130_fd_sc_hd__or2_4
X_6902_ _9684_/Q VGND VPWR _6902_/Y VGND VPWR sky130_fd_sc_hd__inv_4
XFILLER_23_514 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9621_ _9674_/CLK _9621_/D _9633_/SET_B VGND VPWR _9621_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6833_ _9642_/Q VGND VPWR _6833_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_50_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6764_ _6762_/Y _5251_/B _6763_/Y _5393_/B VGND VPWR _6764_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_9552_ _9639_/CLK _9552_/D _9633_/SET_B VGND VPWR _9552_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_50_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5715_ _9250_/Q VGND VPWR _6994_/A VGND VPWR sky130_fd_sc_hd__inv_2
X_8503_ _8341_/A _8239_/B _8238_/A _8498_/B _7910_/X VGND VPWR _8504_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9483_ _9483_/CLK _9483_/D _9685_/SET_B VGND VPWR _9483_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6695_ _9413_/Q VGND VPWR _6695_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_148_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5646_ _9278_/Q VGND VPWR _5751_/C VGND VPWR sky130_fd_sc_hd__inv_2
X_8434_ _8434_/A _8636_/C VGND VPWR _8435_/B VGND VPWR sky130_fd_sc_hd__nor2_1
X_5577_ _9325_/Q _5574_/A _8844_/X _5574_/Y VGND VPWR _9325_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8365_ _8551_/A _8378_/B _8250_/A VGND VPWR _8577_/C VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_104_302 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4528_ _9768_/Q _4526_/A _8845_/X _4526_/Y VGND VPWR _9768_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7316_ _6866_/Y _7095_/X _6935_/Y _7068_/D _7315_/X VGND VPWR _7321_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_8296_ _8296_/A _8296_/B VGND VPWR _8296_/Y VGND VPWR sky130_fd_sc_hd__nand2_1
X_7247_ _6232_/Y _7040_/C _6224_/Y _7059_/C VGND VPWR _7247_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4459_ _4459_/A VGND VPWR _6111_/A VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_7178_ _8773_/A _7086_/X _8771_/A _7088_/X VGND VPWR _7178_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_58_411 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6129_ _9674_/Q VGND VPWR _6129_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_73_403 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_115 input85/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_104 _6505_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_121_42 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_374 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_148 _7698_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_126 input86/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_137 input91/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_41_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA_159 _4814_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_81_68 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_94 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_230 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_414 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5500_ _9378_/Q _5498_/A _8845_/X _5498_/Y VGND VPWR _9378_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_185_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6480_ _9331_/Q VGND VPWR _6480_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_145_257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5431_ _5545_/A _5431_/B VGND VPWR _5432_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_114_622 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5362_ _9471_/Q _5357_/A _8842_/X _5357_/Y VGND VPWR _9471_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8150_ _8150_/A _8685_/B VGND VPWR _8152_/A VGND VPWR sky130_fd_sc_hd__or2_1
Xoutput325 _9761_/Q VGND VPWR sram_ro_csb VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput303 _9047_/Q VGND VPWR pwr_ctrl_out[3] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput314 _8817_/X VGND VPWR spimemio_flash_io2_di VGND VPWR sky130_fd_sc_hd__buf_2
X_7101_ _4897_/Y _7095_/X _4779_/Y _7068_/D _7100_/X VGND VPWR _7108_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_8081_ _8188_/B _8640_/B VGND VPWR _8186_/A VGND VPWR sky130_fd_sc_hd__or2_1
Xoutput358 _9013_/Q VGND VPWR wb_dat_o[9] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput336 _9030_/Q VGND VPWR wb_dat_o[18] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput347 _9040_/Q VGND VPWR wb_dat_o[28] VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_59_208 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_143 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5293_ _9519_/Q _5292_/A _5963_/B1 _5292_/Y VGND VPWR _9519_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7032_ _7073_/C _7109_/B VGND VPWR _7033_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_87_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_116 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8983_ _8983_/A _7701_/A VGND VPWR mgmt_gpio_out[6] VGND VPWR sky130_fd_sc_hd__ebufn_8
XFILLER_70_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_7934_ _8282_/C _7836_/C _7831_/Y _7933_/X VGND VPWR _7935_/B VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_23_300 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_480 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7865_ _7959_/A _8528_/A _8525_/A _8189_/A VGND VPWR _7866_/A VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_50_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6816_ _6811_/Y _4613_/B _6812_/Y _4504_/B _6815_/X VGND VPWR _6829_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9604_ _9617_/CLK _9604_/D _9295_/SET_B VGND VPWR _9604_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_7796_ _8084_/A _8085_/A VGND VPWR _7797_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_6747_ _6742_/Y _5110_/B _6743_/Y _5916_/B _6746_/X VGND VPWR _6759_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_2
X_9535_ _9535_/CLK _9535_/D _9528_/SET_B VGND VPWR _9535_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_164_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_511 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6678_ _6673_/Y _5968_/B _6674_/Y _5864_/B _6677_/X VGND VPWR _6690_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9466_ _9514_/CLK _9466_/D _4628_/A VGND VPWR _9466_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_5629_ _9288_/Q _5623_/A _8955_/A1 _5623_/Y VGND VPWR _9288_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_9397_ _9509_/CLK _9397_/D _9528_/SET_B VGND VPWR _9397_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_8417_ _8667_/B _8577_/A VGND VPWR _8686_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_151_216 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8348_ _8378_/B _8347_/X _8216_/X VGND VPWR _8349_/B VGND VPWR sky130_fd_sc_hd__o21a_1
XFILLER_104_110 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8279_ _8279_/A _8378_/B _8279_/C VGND VPWR _8280_/C VGND VPWR sky130_fd_sc_hd__or3_1
XFILLER_116_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_79 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_572 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_12 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_83 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_50 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_94 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_124 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_566 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_583 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_544 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_282 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_270 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5980_ _5980_/A VGND VPWR _5980_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_4931_ _4931_/A _4931_/B VGND VPWR _5328_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_32_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7650_ _6779_/Y _7434_/X _6780_/Y _7436_/X VGND VPWR _7650_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4862_ _4858_/Y _5374_/B _4860_/Y _4861_/X VGND VPWR _4862_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_177_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6601_ _6597_/Y _5232_/B _8785_/A _5240_/B _6600_/X VGND VPWR _6601_/X VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9320_ _9613_/CLK _9320_/D _9646_/SET_B VGND VPWR _9320_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_7581_ _6225_/Y _7445_/X _6164_/Y _7447_/X VGND VPWR _7581_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4793_ _9546_/Q VGND VPWR _4793_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
XANTENNA_15 _7331_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_48 _4935_/D VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_37 _4833_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_26 _4481_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_20_347 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_358 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6532_ _9154_/Q VGND VPWR _7699_/A VGND VPWR sky130_fd_sc_hd__clkinv_4
XANTENNA_59 _6271_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_137_19 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9251_ _9278_/CLK _9251_/D _9633_/SET_B VGND VPWR _9251_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_6463_ _9671_/Q VGND VPWR _6463_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_173_374 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5414_ _5414_/A VGND VPWR _5414_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_8202_ _8202_/A _8213_/A VGND VPWR _8721_/A VGND VPWR sky130_fd_sc_hd__nor2_4
X_9182_ _9652_/CLK _9182_/D _9646_/SET_B VGND VPWR _9182_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_126_290 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8133_ _8133_/A VGND VPWR _8358_/A VGND VPWR sky130_fd_sc_hd__inv_2
X_6394_ _6392_/Y _6081_/B _6393_/Y _5602_/B VGND VPWR _6394_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_87_303 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5345_ _5345_/A VGND VPWR _5346_/A VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_101_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5276_ _9529_/Q _5269_/A _8930_/A1 _5269_/Y VGND VPWR _9529_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8064_ _8518_/A _8064_/B _8064_/C VGND VPWR _8703_/C VGND VPWR sky130_fd_sc_hd__and3_1
X_7015_ _9586_/Q _7015_/B VGND VPWR _7016_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_55_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_244 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_8966_ _7747_/X _8966_/A1 _8975_/S VGND VPWR _8966_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_55_299 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7917_ _8734_/A _7917_/B _8317_/A _8597_/A VGND VPWR _7917_/Y VGND VPWR sky130_fd_sc_hd__nor4_1
XFILLER_169_603 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8897_ _8896_/X _9149_/Q _9054_/Q VGND VPWR _8897_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_11_303 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7848_ _7848_/A _8077_/A VGND VPWR _7929_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_23_174 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_59 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7779_ _7832_/A _7837_/B _5934_/X VGND VPWR _8218_/B VGND VPWR sky130_fd_sc_hd__o21ai_2
X_9518_ _9545_/CLK _9518_/D _4628_/A VGND VPWR _9518_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_149_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9449_ _9785_/CLK _9449_/D _9779_/SET_B VGND VPWR _9449_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_137_599 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_62 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_130 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_450 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xinput13 mask_rev_in[18] VGND VPWR _6766_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_128_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput35 mask_rev_in[9] VGND VPWR _6849_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput24 mask_rev_in[28] VGND VPWR _6411_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput46 mgmt_gpio_in[19] VGND VPWR _6521_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput57 mgmt_gpio_in[29] VGND VPWR input57/X VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
Xinput79 spi_enabled VGND VPWR _8833_/S VGND VPWR sky130_fd_sc_hd__buf_6
Xinput68 mgmt_gpio_in[5] VGND VPWR _8801_/A VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_170_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5130_ _5130_/A VGND VPWR _5130_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_151_591 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5061_ _8812_/A _5058_/X _8811_/A _5060_/X VGND VPWR _5062_/C VGND VPWR sky130_fd_sc_hd__o22ai_1
XFILLER_37_200 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8820_ _9217_/Q _9069_/Q _9787_/Q VGND VPWR _8820_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_92_372 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5963_ _9105_/Q _5962_/A _5963_/B1 _5962_/Y VGND VPWR _9105_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8751_ _8751_/A VGND VPWR _8752_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xclkbuf_opt_4_0_csclk clkbuf_2_1_0_csclk/X VGND VPWR clkbuf_opt_4_0_csclk/X VGND VPWR
+ sky130_fd_sc_hd__clkbuf_16
X_4914_ _9424_/Q VGND VPWR _4914_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_7702_ _7702_/A VGND VPWR _7702_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_8682_ _8720_/B _8722_/A _8722_/B _8723_/A VGND VPWR _8682_/X VGND VPWR sky130_fd_sc_hd__or4_4
X_5894_ _5894_/A1 _8875_/X _8924_/X _9139_/Q VGND VPWR _9139_/D VGND VPWR sky130_fd_sc_hd__o22a_2
XFILLER_178_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_4845_ _4840_/Y _4841_/X _4842_/Y _5968_/B _4844_/X VGND VPWR _4864_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_7633_ _6922_/Y _7430_/X _6805_/Y _7432_/X _7632_/X VGND VPWR _7633_/X VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_193_425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4776_ _4925_/A _4843_/B VGND VPWR _5916_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_7564_ _6308_/Y _7441_/X _6256_/Y _7443_/X _7563_/X VGND VPWR _7571_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9303_ _9440_/CLK _9303_/D _9685_/SET_B VGND VPWR _9303_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6515_ _9272_/Q VGND VPWR _8759_/A VGND VPWR sky130_fd_sc_hd__inv_4
X_7495_ _6879_/Y _7465_/X _6825_/Y _7467_/X VGND VPWR _7495_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_106_9 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6446_ input56/X _6322_/Y _8817_/A _4680_/Y VGND VPWR _6446_/Y VGND VPWR sky130_fd_sc_hd__a22oi_4
X_9234_ _9371_/CLK _9234_/D _9295_/SET_B VGND VPWR _9234_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_106_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6377_ _9273_/Q VGND VPWR _6377_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9165_ _9203_/CLK _9165_/D _9633_/SET_B VGND VPWR _9165_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_0_527 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_9096_ _9501_/CLK _9096_/D _9647_/SET_B VGND VPWR _9096_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_8116_ _8116_/A _8116_/B VGND VPWR _8117_/B VGND VPWR sky130_fd_sc_hd__or2_2
X_5328_ _5671_/A _5328_/B VGND VPWR _5329_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_102_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_8047_ _8047_/A _8467_/A VGND VPWR _8047_/X VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_87_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5259_ _5259_/A _5259_/B VGND VPWR _5260_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_68_391 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_266 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_534 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_47 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_8949_ _9713_/Q _6629_/Y _8957_/S VGND VPWR _8949_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_73_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_494 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_436 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_488 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_352 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_22 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_122 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_103 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_531 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_211 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_578 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4630_ _6052_/B _7022_/B VGND VPWR _6050_/A VGND VPWR sky130_fd_sc_hd__nor2_8
XFILLER_116_514 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6300_ _6296_/Y _5621_/B _6297_/Y _5013_/B _6299_/X VGND VPWR _6307_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_4561_ _5967_/B1 _9756_/Q _4561_/S VGND VPWR _4562_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_128_374 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7280_ _6109_/Y _7118_/X _6068_/Y _7048_/C VGND VPWR _7280_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4492_ _4492_/A VGND VPWR _4493_/A VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_170_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6231_ _9638_/Q VGND VPWR _6231_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_170_130 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6162_ _6157_/Y _5089_/B _6158_/X _6161_/X VGND VPWR _6174_/B VGND VPWR sky130_fd_sc_hd__o211a_1
X_5113_ _9639_/Q _5112_/A _8846_/X _5112_/Y VGND VPWR _9639_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_6093_ _6093_/A VGND VPWR _6093_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_111_274 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5044_ _8969_/X _4551_/B _9675_/Q _5062_/D VGND VPWR _9675_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_72_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_8803_ _8803_/A _8833_/S VGND VPWR _8804_/A VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_25_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6995_ _9248_/Q _7056_/B _7125_/A VGND VPWR _7094_/B VGND VPWR sky130_fd_sc_hd__or3_1
X_9783_ _9785_/CLK _9783_/D _9779_/SET_B VGND VPWR _9783_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_53_534 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5946_ _9116_/Q _5943_/A _5965_/B1 _5943_/Y VGND VPWR _9116_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8734_ _8734_/A _8734_/B _8734_/C _8734_/D VGND VPWR _8735_/B VGND VPWR sky130_fd_sc_hd__or4_1
XFILLER_80_353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_606 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5877_ _9156_/Q _5874_/A _8844_/X _5874_/Y VGND VPWR _9156_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8665_ _8665_/A _8665_/B _7877_/X VGND VPWR _8666_/B VGND VPWR sky130_fd_sc_hd__or3b_1
XFILLER_139_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4828_ _8807_/A _5227_/B _4827_/Y _6251_/A VGND VPWR _4828_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_7616_ _4765_/Y _7425_/X _7613_/X _7615_/X VGND VPWR _7626_/C VGND VPWR sky130_fd_sc_hd__o211a_1
XFILLER_178_296 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8596_ _8077_/A _8239_/B _8236_/A _8304_/Y _8504_/B VGND VPWR _8727_/A VGND VPWR
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_193_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7547_ _6398_/Y _7455_/X _6439_/Y _7457_/X VGND VPWR _7547_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4759_ _9294_/Q VGND VPWR _7121_/A VGND VPWR sky130_fd_sc_hd__clkinv_4
XFILLER_175_38 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_300 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7478_ _4814_/Y _7475_/X _4726_/Y _7477_/X VGND VPWR _7478_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_9217_ _9280_/CLK _9217_/D _9757_/SET_B VGND VPWR _9217_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6429_ _9777_/Q VGND VPWR _6429_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
XFILLER_134_388 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_76 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9148_ _9280_/CLK _9148_/D _9757_/SET_B VGND VPWR _9148_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_0_357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_486 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9079_ _9790_/CLK _9079_/D _9757_/SET_B VGND VPWR _9079_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_56_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_242 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_231 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_220 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_286 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_275 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_264 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_403 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_442 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_94 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_428 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_311 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_355 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_163 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_539 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_420 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_580 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_550 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold2 hold2/A VGND VPWR hold2/X VGND VPWR sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_39_328 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_350 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_556 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_342 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5800_ _9211_/Q _5799_/A _8846_/X _5799_/Y VGND VPWR _9211_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_6780_ _9491_/Q VGND VPWR _6780_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_22_217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5731_ _9055_/Q _7041_/A _5713_/Y VGND VPWR _5731_/Y VGND VPWR sky130_fd_sc_hd__a21oi_1
X_5662_ _5662_/A VGND VPWR _5662_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_8450_ _8450_/A VGND VPWR _8683_/A VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_30_283 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5593_ _9312_/Q _5585_/A _8839_/X _5585_/Y VGND VPWR _9312_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7401_ _9252_/Q _7401_/B VGND VPWR _7466_/A VGND VPWR sky130_fd_sc_hd__or2_4
X_4613_ _5259_/A _4613_/B VGND VPWR _4614_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_8381_ _8722_/A _8381_/B VGND VPWR _8382_/B VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_163_428 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4544_ _9066_/Q VGND VPWR _8810_/A VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_163_439 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7332_ _6723_/Y _7086_/X _6695_/Y _7088_/X VGND VPWR _7332_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_190_247 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_355 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7263_ _6164_/Y _7124_/X _6163_/Y _7068_/B _7262_/X VGND VPWR _7264_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_171_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9002_ _9595_/Q _8781_/A VGND VPWR mgmt_gpio_out[25] VGND VPWR sky130_fd_sc_hd__ebufn_8
X_4475_ _6052_/A VGND VPWR _5259_/A VGND VPWR sky130_fd_sc_hd__buf_12
X_6214_ _9746_/Q VGND VPWR _6214_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_143_196 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_7194_ _8761_/A _7392_/B VGND VPWR _7194_/X VGND VPWR sky130_fd_sc_hd__or2_1
X_6145_ _6071_/Y _6145_/B _6145_/C _6145_/D VGND VPWR _6145_/Y VGND VPWR sky130_fd_sc_hd__nand4b_4
X_6076_ _6074_/Y _5420_/B _6075_/Y _4861_/X VGND VPWR _6076_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_57_103 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5027_ _9687_/Q _5026_/A _8925_/A1 _5026_/Y VGND VPWR _9687_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_38_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9766_ _9769_/CLK _9766_/D _9757_/SET_B VGND VPWR _9766_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_8717_ _8640_/A _8164_/A _8640_/A _8640_/B VGND VPWR _8717_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_6978_ _6237_/Y _6976_/A _9018_/Q _6976_/Y VGND VPWR _9018_/D VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_179_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9697_ _9709_/CLK _9697_/D _5004_/X VGND VPWR _9697_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_5929_ _7781_/A _7781_/B VGND VPWR _7837_/C VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_166_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8648_ _8566_/B _8214_/Y _8340_/C VGND VPWR _8681_/B VGND VPWR sky130_fd_sc_hd__o21a_1
X_8579_ _8708_/B _8579_/B _8579_/C VGND VPWR _8716_/A VGND VPWR sky130_fd_sc_hd__or3_2
XFILLER_119_31 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_322 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_491 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_358 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_187 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_103 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_61 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_534 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_71 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_531 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_415 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7950_ _8394_/D _8515_/B _8660_/C VGND VPWR _8187_/A VGND VPWR sky130_fd_sc_hd__or3_1
XFILLER_39_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7881_ _7881_/A VGND VPWR _8566_/A VGND VPWR sky130_fd_sc_hd__inv_2
X_6901_ _6901_/A _6901_/B _6901_/C _6901_/D VGND VPWR _6945_/A VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_35_364 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9620_ _9620_/CLK _9620_/D _9633_/SET_B VGND VPWR _9620_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6832_ _9521_/Q VGND VPWR _6832_/Y VGND VPWR sky130_fd_sc_hd__inv_6
XFILLER_50_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6763_ _9444_/Q VGND VPWR _6763_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9551_ _9639_/CLK _9551_/D _9757_/SET_B VGND VPWR _9551_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_50_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6694_ _9530_/Q VGND VPWR _6694_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_5714_ _7401_/B _9055_/Q _9251_/Q _5713_/Y VGND VPWR _9251_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8502_ _8230_/A _8498_/B _7877_/X _8233_/A VGND VPWR _8504_/B VGND VPWR sky130_fd_sc_hd__o211a_1
X_9482_ _9483_/CLK _9482_/D _9685_/SET_B VGND VPWR _9482_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_5645_ _6997_/A _5643_/Y _5724_/B _9054_/Q _8819_/X VGND VPWR _5651_/A VGND VPWR
+ sky130_fd_sc_hd__a32o_2
X_8433_ _8514_/A _8433_/B VGND VPWR _8636_/C VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_40_18 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_480 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_214 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5576_ _9326_/Q _5574_/A _8845_/X _5574_/Y VGND VPWR _9326_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8364_ _8364_/A _8730_/C _8575_/C _8364_/D VGND VPWR _8368_/A VGND VPWR sky130_fd_sc_hd__or4_1
XFILLER_116_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7315_ _6843_/Y _7097_/X _6845_/Y _7099_/X VGND VPWR _7315_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4527_ _9769_/Q _4526_/A _8846_/X _4526_/Y VGND VPWR _9769_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8295_ _8295_/A _8295_/B VGND VPWR _8296_/B VGND VPWR sky130_fd_sc_hd__and2_1
X_4458_ _4661_/C _8938_/X _4665_/C VGND VPWR _4459_/A VGND VPWR sky130_fd_sc_hd__or3_1
X_7246_ _6160_/Y _7082_/X _6195_/Y _7084_/X _7245_/X VGND VPWR _7265_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_77_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7177_ _7177_/A _7177_/B _7177_/C VGND VPWR _7177_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
XFILLER_100_520 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6128_ _9158_/Q VGND VPWR _6128_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_105_66 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_106 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6059_ _9100_/Q VGND VPWR _6059_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_58_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_139 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_105 _4629_/C VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_116 input85/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_138 _8955_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_149 _5960_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_127 input86/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_26_386 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_98 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_9749_ _9777_/CLK _9749_/D _9757_/SET_B VGND VPWR _9749_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_154_247 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_130 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_95 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_570 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_106 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_364 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_378 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5430_ _9424_/Q _5422_/A _8839_/X _5422_/Y VGND VPWR _9424_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_145_269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5361_ _9472_/Q _5357_/A _8925_/A1 _5357_/Y VGND VPWR _9472_/D VGND VPWR sky130_fd_sc_hd__a22o_1
Xoutput304 _4808_/A VGND VPWR reset VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput326 _9119_/Q VGND VPWR wb_ack_o VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput315 _8818_/X VGND VPWR spimemio_flash_io3_di VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_99_323 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5292_ _5292_/A VGND VPWR _5292_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7100_ _4926_/Y _7097_/X _4910_/Y _7099_/X VGND VPWR _7100_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_8080_ _8080_/A VGND VPWR _8640_/B VGND VPWR sky130_fd_sc_hd__buf_8
Xoutput337 _9031_/Q VGND VPWR wb_dat_o[19] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput348 _9041_/Q VGND VPWR wb_dat_o[29] VGND VPWR sky130_fd_sc_hd__buf_2
X_7031_ _7127_/A _7111_/C VGND VPWR _7109_/B VGND VPWR sky130_fd_sc_hd__or2_1
X_8982_ _9583_/Q _8745_/A VGND VPWR mgmt_gpio_out[5] VGND VPWR sky130_fd_sc_hd__ebufn_8
XFILLER_82_212 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_128 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7933_ _8662_/A _7933_/B VGND VPWR _7933_/X VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_55_437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_18 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_312 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7864_ _7864_/A VGND VPWR _7864_/X VGND VPWR sky130_fd_sc_hd__buf_6
XFILLER_168_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6815_ _6813_/Y _4870_/X _6814_/Y _4623_/B VGND VPWR _6815_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_7795_ _8538_/C _8516_/B VGND VPWR _8085_/A VGND VPWR sky130_fd_sc_hd__or2_2
X_9603_ _9617_/CLK _9603_/D _9295_/SET_B VGND VPWR _9603_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_50_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6746_ _6744_/Y _4841_/X _6745_/Y _5100_/B VGND VPWR _6746_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_9534_ _9534_/CLK _9534_/D _9647_/SET_B VGND VPWR _9534_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_51_28 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9465_ _9514_/CLK _9465_/D _4628_/A VGND VPWR _9465_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6677_ _6675_/Y _4613_/B _6676_/Y _4868_/X VGND VPWR _6677_/X VGND VPWR sky130_fd_sc_hd__o22a_2
XFILLER_164_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8416_ _8416_/A VGND VPWR _8667_/B VGND VPWR sky130_fd_sc_hd__inv_2
X_5628_ _9289_/Q _5623_/A _8842_/X _5623_/Y VGND VPWR _9289_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_9396_ _9509_/CLK _9396_/D _9528_/SET_B VGND VPWR _9396_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_164_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5559_ _9337_/Q _5558_/A _8843_/X _5558_/Y VGND VPWR _9337_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8347_ _8377_/B _8350_/C VGND VPWR _8347_/X VGND VPWR sky130_fd_sc_hd__or2_2
XFILLER_183_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_122 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_8278_ _8345_/A _8583_/C _8345_/B VGND VPWR _8279_/A VGND VPWR sky130_fd_sc_hd__or3b_1
XFILLER_116_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7229_ _6264_/Y _7079_/B _6316_/Y _7059_/A VGND VPWR _7229_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_76_25 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_231 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_584 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_372 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_24 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_40 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_1_0_wb_clk_i clkbuf_3_1_0_wb_clk_i/A VGND VPWR _9681_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_54_492 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_73 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_334 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_136 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_95 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_84 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_556 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_450 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_304 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_407 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_4930_ _9489_/Q VGND VPWR _4930_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_178_604 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4861_ _6111_/A _4925_/A VGND VPWR _4861_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_32_131 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6600_ _9069_/Q _6251_/Y _6599_/Y _4602_/B VGND VPWR _6600_/X VGND VPWR sky130_fd_sc_hd__o2bb2a_1
XFILLER_32_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4792_ _9748_/Q VGND VPWR _4792_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7580_ _6218_/Y _7425_/X _7577_/X _7579_/X VGND VPWR _7590_/C VGND VPWR sky130_fd_sc_hd__o211a_1
XANTENNA_16 _7353_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_38 _4835_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_27 _4481_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_158_372 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6531_ _6531_/A VGND VPWR _6531_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
XANTENNA_49 _6096_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_9250_ _9278_/CLK _9250_/D _9633_/SET_B VGND VPWR _9250_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6462_ _9692_/Q VGND VPWR _6462_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_8201_ _8377_/C VGND VPWR _8340_/C VGND VPWR sky130_fd_sc_hd__inv_2
X_6393_ _9306_/Q VGND VPWR _6393_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9181_ _9613_/CLK _9181_/D _9646_/SET_B VGND VPWR _9181_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_5413_ _5413_/A VGND VPWR _5414_/A VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_161_548 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_386 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8132_ _8164_/A _8137_/B VGND VPWR _8133_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_5344_ _5545_/A _5344_/B VGND VPWR _5345_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_99_164 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5275_ _9530_/Q _5269_/A _8841_/X _5269_/Y VGND VPWR _9530_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8063_ _8077_/A VGND VPWR _8518_/A VGND VPWR sky130_fd_sc_hd__clkinv_4
X_7014_ _7014_/A VGND VPWR _7014_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_8965_ _7745_/X _8965_/A1 _8975_/S VGND VPWR _8965_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_15_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_470 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7916_ _8077_/A _8254_/B VGND VPWR _8597_/A VGND VPWR sky130_fd_sc_hd__nor2_1
X_8896_ _7397_/Y _9631_/Q _8959_/S VGND VPWR _8896_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_7847_ _7847_/A VGND VPWR _8077_/A VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_11_315 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7778_ _7756_/B _7777_/Y _7837_/B _7777_/A VGND VPWR _7897_/A VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_137_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9517_ _9545_/CLK _9517_/D _4628_/A VGND VPWR _9517_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6729_ _9465_/Q VGND VPWR _6729_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_164_320 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_139 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_9448_ _9785_/CLK _9448_/D _9779_/SET_B VGND VPWR _9448_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_152_504 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_386 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9379_ _9379_/CLK _9379_/D _9779_/SET_B VGND VPWR _9379_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_87_13 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_318 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_74 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_94 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_60 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput36 mgmt_gpio_in[0] VGND VPWR _8805_/A VGND VPWR sky130_fd_sc_hd__buf_8
Xinput14 mask_rev_in[19] VGND VPWR _6570_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput25 mask_rev_in[29] VGND VPWR _6245_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_128_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput58 mgmt_gpio_in[2] VGND VPWR _4949_/A VGND VPWR sky130_fd_sc_hd__buf_12
Xinput69 mgmt_gpio_in[6] VGND VPWR input69/X VGND VPWR sky130_fd_sc_hd__buf_2
Xinput47 mgmt_gpio_in[1] VGND VPWR input47/X VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_6_374 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5060_ _5060_/A VGND VPWR _5060_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_37_212 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5962_ _5962_/A VGND VPWR _5962_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_8750_ _8750_/A VGND VPWR _8750_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_4913_ _4906_/Y _4907_/X _4908_/Y _4577_/B _4912_/X VGND VPWR _4934_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_2
X_7701_ _7701_/A VGND VPWR _7702_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_18_492 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_8681_ _8681_/A _8681_/B _8681_/C VGND VPWR _8723_/A VGND VPWR sky130_fd_sc_hd__or3_1
X_5893_ _5893_/A1 _8877_/X _8924_/X _9140_/Q VGND VPWR _9140_/D VGND VPWR sky130_fd_sc_hd__o22a_2
X_7632_ _6874_/Y _7434_/X _6843_/Y _7436_/X VGND VPWR _7632_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4844_ _4919_/A _6158_/A VGND VPWR _4844_/X VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_148_19 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_7563_ _6239_/Y _7445_/X _6269_/Y _7447_/X VGND VPWR _7563_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4775_ _9120_/Q VGND VPWR _4775_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_165_139 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9302_ _9440_/CLK _9302_/D _9685_/SET_B VGND VPWR _9302_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6514_ _9193_/Q VGND VPWR _8749_/A VGND VPWR sky130_fd_sc_hd__clkinv_4
XFILLER_119_578 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7494_ _6933_/Y _7451_/X _6853_/Y _7453_/X _7493_/X VGND VPWR _7499_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9233_ _9508_/CLK _9233_/D _9647_/SET_B VGND VPWR _9233_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6445_ _9645_/Q VGND VPWR _6445_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_164_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6376_ _6371_/Y _5679_/B _6372_/Y _5776_/B _6375_/X VGND VPWR _6376_/X VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9164_ _9203_/CLK _9164_/D _9633_/SET_B VGND VPWR _9164_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_8115_ _8401_/A VGND VPWR _8115_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_5327_ _9494_/Q _5319_/A _8839_/X _5319_/Y VGND VPWR _9494_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_9095_ _9508_/CLK _9095_/D _9295_/SET_B VGND VPWR _9095_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_8046_ _8624_/B _8554_/A VGND VPWR _8467_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_5258_ _9541_/Q _5253_/A _5967_/B1 _5253_/Y VGND VPWR _9541_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_75_307 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5189_ _6040_/A VGND VPWR _5190_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_73_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8948_ hold1/X _6237_/Y _8957_/S VGND VPWR _8948_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_188_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_546 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8879_ _8878_/X _9140_/Q _9054_/Q VGND VPWR _8879_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_11_123 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_331 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_448 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_138 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_364 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_63 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_74 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_334 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_322 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_231 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_134 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_340 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_220 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_415 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_331 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_498 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4560_ _4560_/A VGND VPWR _9757_/D VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_190_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_386 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_526 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4491_ _5960_/A _4491_/B VGND VPWR _4492_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_6230_ _9099_/Q VGND VPWR _6230_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_170_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6161_ _6159_/Y _5382_/B _6160_/Y _5317_/B VGND VPWR _6161_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_170_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5112_ _5112_/A VGND VPWR _5112_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_6092_ _9747_/Q VGND VPWR _6092_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_84_104 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_487 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5043_ _8970_/X _4551_/B _9676_/Q _5062_/D VGND VPWR _9676_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_38_576 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_8802_ _8802_/A VGND VPWR _8802_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_25_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6994_ _6994_/A _9249_/Q VGND VPWR _7075_/A VGND VPWR sky130_fd_sc_hd__or2_4
X_9782_ _9785_/CLK _9782_/D _9779_/SET_B VGND VPWR _9782_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_80_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_259 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8733_ _8733_/A VGND VPWR _8733_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_5945_ _9117_/Q _5943_/A _5964_/B1 _5943_/Y VGND VPWR _9117_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_5876_ _9157_/Q _5874_/A _8845_/X _5874_/Y VGND VPWR _9157_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8664_ _8664_/A VGND VPWR _8664_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_7615_ _4775_/Y _7430_/X _4836_/Y _7432_/X _7614_/X VGND VPWR _7615_/X VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_4827_ _9203_/Q VGND VPWR _4827_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_8595_ _8595_/A _8595_/B _8595_/C _7902_/X VGND VPWR _8659_/C VGND VPWR sky130_fd_sc_hd__or4b_1
XFILLER_5_609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7546_ _6368_/Y _7441_/X _6390_/Y _7443_/X _7545_/X VGND VPWR _7553_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_4758_ _4749_/Y _5602_/B _4751_/Y _5545_/B _4757_/X VGND VPWR _4790_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_4689_ _6086_/B _4843_/B VGND VPWR _5949_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_7477_ _7477_/A VGND VPWR _7477_/X VGND VPWR sky130_fd_sc_hd__buf_6
X_6428_ _9420_/Q VGND VPWR _6428_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_134_356 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9216_ _9655_/CLK _9216_/D _9779_/SET_B VGND VPWR _9216_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_9147_ _9280_/CLK _9147_/D _9757_/SET_B VGND VPWR _9147_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6359_ _6359_/A1 _6165_/A _6356_/Y _5621_/B _6358_/X VGND VPWR _6359_/X VGND VPWR
+ sky130_fd_sc_hd__o221a_2
XFILLER_130_562 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_9078_ _9790_/CLK _9078_/D _9757_/SET_B VGND VPWR _9078_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_8029_ _8624_/B _8550_/A VGND VPWR _8029_/X VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_88_498 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_30 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_192 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_210 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_243 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_232 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_276 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_254 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_415 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_454 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_106 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_298 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_287 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_487 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_175 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_432 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_435 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_70 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_354 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5730_ _5730_/A VGND VPWR _9250_/D VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_15_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7400_ _7400_/A VGND VPWR _7400_/X VGND VPWR sky130_fd_sc_hd__buf_6
X_5661_ _5661_/A VGND VPWR _5662_/A VGND VPWR sky130_fd_sc_hd__clkbuf_4
X_5592_ _9313_/Q _5585_/A _8930_/A1 _5585_/Y VGND VPWR _9313_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8380_ _8380_/A _8380_/B _8720_/C _8585_/A VGND VPWR _8381_/B VGND VPWR sky130_fd_sc_hd__or4_1
X_4612_ _6111_/A _6158_/B VGND VPWR _4613_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_4543_ _9064_/Q VGND VPWR _8811_/A VGND VPWR sky130_fd_sc_hd__inv_2
X_7331_ _7331_/A _7331_/B _7331_/C VGND VPWR _7331_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
X_7262_ _6188_/Y _7126_/X _6189_/Y _7128_/X VGND VPWR _7262_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_104_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4474_ _4729_/A _4729_/B _4669_/A _4729_/D VGND VPWR _4891_/A VGND VPWR sky130_fd_sc_hd__or4_4
X_9001_ _9594_/Q _8779_/A VGND VPWR mgmt_gpio_out[24] VGND VPWR sky130_fd_sc_hd__ebufn_8
X_6213_ _8823_/X VGND VPWR _6213_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_7193_ _7703_/A _7059_/D _8767_/A _7116_/X _7192_/X VGND VPWR _7198_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_6144_ _6144_/A _6144_/B _6144_/C _6144_/D VGND VPWR _6145_/D VGND VPWR sky130_fd_sc_hd__and4_1
X_6075_ _6075_/A VGND VPWR _6075_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
XFILLER_85_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5026_ _5026_/A VGND VPWR _5026_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_26_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9765_ _9768_/CLK _9765_/D _4628_/A VGND VPWR _9765_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_6977_ _6145_/Y _6976_/A _9019_/Q _6976_/Y VGND VPWR _9019_/D VGND VPWR sky130_fd_sc_hd__o22a_1
X_5928_ _7774_/C _7774_/D _5928_/C VGND VPWR _5936_/C VGND VPWR sky130_fd_sc_hd__or3_1
X_8716_ _8716_/A _8716_/B _8716_/C _8716_/D VGND VPWR _8729_/A VGND VPWR sky130_fd_sc_hd__or4_1
XFILLER_110_67 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_415 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_404 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_9696_ _8837_/A1 _9696_/D _5010_/X VGND VPWR _9696_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_186_16 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8647_ _8647_/A _8716_/C _8678_/C _8721_/C VGND VPWR _8647_/Y VGND VPWR sky130_fd_sc_hd__nor4_1
X_5859_ _5849_/X _8855_/X _8924_/X _9167_/Q VGND VPWR _9167_/D VGND VPWR sky130_fd_sc_hd__o22a_2
XFILLER_166_245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8578_ _8578_/A _8578_/B _8578_/C VGND VPWR _8645_/D VGND VPWR sky130_fd_sc_hd__or3_1
XFILLER_147_470 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_43 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_610 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7529_ _8765_/A _7455_/X _6517_/Y _7457_/X VGND VPWR _7529_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_79_14 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_115 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_75 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_392 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_73 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_384 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_94 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_543 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_9 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_495 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_240 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_178 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_287 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6900_ _6895_/Y _5572_/B _6896_/Y _5897_/B _6899_/X VGND VPWR _6901_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_7880_ _8394_/D _8272_/A VGND VPWR _7881_/A VGND VPWR sky130_fd_sc_hd__or2_2
X_6831_ _6831_/A VGND VPWR _6831_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_35_376 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9550_ _9655_/CLK _9550_/D _9633_/SET_B VGND VPWR _9550_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_50_357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8501_ _8594_/A _8695_/C _8501_/C _8501_/D VGND VPWR _8501_/X VGND VPWR sky130_fd_sc_hd__or4_2
X_6762_ _9543_/Q VGND VPWR _6762_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_9481_ _9527_/CLK _9481_/D _9685_/SET_B VGND VPWR _9481_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_5713_ _5713_/A VGND VPWR _5713_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_6693_ _9340_/Q VGND VPWR _6693_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_176_576 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8432_ _8562_/A _8672_/C _8432_/C VGND VPWR _8434_/A VGND VPWR sky130_fd_sc_hd__or3_1
X_5644_ _9055_/Q VGND VPWR _5724_/B VGND VPWR sky130_fd_sc_hd__clkinv_4
XFILLER_148_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8363_ _8627_/B _8490_/B VGND VPWR _8364_/D VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_129_492 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_19 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_131 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5575_ _9327_/Q _5574_/A _8846_/X _5574_/Y VGND VPWR _9327_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7314_ _6883_/Y _7048_/B _6800_/Y _7077_/A _7313_/X VGND VPWR _7321_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_4526_ _4526_/A VGND VPWR _4526_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_8294_ _8294_/A _8650_/C VGND VPWR _8295_/B VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_171_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_186 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4457_ _4456_/Y _8942_/X _8941_/X VGND VPWR _4665_/C VGND VPWR sky130_fd_sc_hd__a21o_1
X_7245_ _6178_/Y _7077_/C _6151_/Y _7077_/D _7244_/X VGND VPWR _7245_/X VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_172_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7176_ _7176_/A _7176_/B _7176_/C _7176_/D VGND VPWR _7177_/C VGND VPWR sky130_fd_sc_hd__and4_1
X_6127_ _9113_/Q VGND VPWR _6127_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_105_78 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6058_ _9044_/Q _6054_/A _8916_/A1 _6054_/Y VGND VPWR _9044_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_73_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_7 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA_106 input77/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_5009_ _6040_/A VGND VPWR _5010_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA_117 input85/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_128 input86/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_139 _6485_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_53_162 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_9748_ _9755_/CLK _9748_/D _9757_/SET_B VGND VPWR _9748_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_9679_ _9681_/CLK _9679_/D _6146_/A VGND VPWR _9679_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_182_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_142 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_258 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_431 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_178 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_542 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_70 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5360_ _9473_/Q _5357_/A _8844_/X _5357_/Y VGND VPWR _9473_/D VGND VPWR sky130_fd_sc_hd__a22o_1
Xoutput316 _9762_/Q VGND VPWR sram_ro_addr[0] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput305 _8802_/X VGND VPWR ser_rx VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_160_229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_484 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xoutput327 _9020_/Q VGND VPWR wb_dat_o[0] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput338 _9021_/Q VGND VPWR wb_dat_o[1] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput349 _9022_/Q VGND VPWR wb_dat_o[2] VGND VPWR sky130_fd_sc_hd__buf_2
X_5291_ _5291_/A VGND VPWR _5292_/A VGND VPWR sky130_fd_sc_hd__clkbuf_2
X_7030_ _7030_/A VGND VPWR _7040_/A VGND VPWR sky130_fd_sc_hd__buf_8
XFILLER_95_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8981_ _9582_/Q _7703_/A VGND VPWR mgmt_gpio_out[4] VGND VPWR sky130_fd_sc_hd__ebufn_8
XFILLER_55_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_224 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7932_ _8394_/B _8298_/A _7931_/X VGND VPWR _7933_/B VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_51_600 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_7863_ _8496_/A _8305_/A VGND VPWR _7864_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_23_324 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6814_ _9720_/Q VGND VPWR _6814_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7794_ _7823_/A _7823_/B _8538_/B VGND VPWR _8516_/B VGND VPWR sky130_fd_sc_hd__o21ai_2
X_9602_ _9617_/CLK _9602_/D _9295_/SET_B VGND VPWR _9602_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_50_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9533_ _9535_/CLK _9533_/D _9528_/SET_B VGND VPWR _9533_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6745_ _9643_/Q VGND VPWR _6745_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
X_9464_ _9514_/CLK _9464_/D _4628_/A VGND VPWR _9464_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_8415_ _8551_/A _8401_/B _8412_/X _8414_/Y VGND VPWR _8415_/X VGND VPWR sky130_fd_sc_hd__o211a_1
X_6676_ _6676_/A VGND VPWR _6676_/Y VGND VPWR sky130_fd_sc_hd__inv_4
XFILLER_191_332 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5627_ _9290_/Q _5623_/A _8925_/A1 _5623_/Y VGND VPWR _9290_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_9395_ _9509_/CLK _9395_/D _9528_/SET_B VGND VPWR _9395_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_5558_ _5558_/A VGND VPWR _5558_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_8346_ _8346_/A _8346_/B _8196_/X VGND VPWR _8350_/C VGND VPWR sky130_fd_sc_hd__or3b_1
X_4509_ _9775_/Q _4506_/A _5965_/B1 _4506_/Y VGND VPWR _9775_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8277_ _8525_/A _8189_/A _8213_/A _8583_/A _8189_/Y VGND VPWR _8345_/B VGND VPWR
+ sky130_fd_sc_hd__o32a_1
XFILLER_132_443 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7228_ _6290_/Y _7095_/X _6308_/Y _7068_/D _7227_/X VGND VPWR _7233_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_5489_ _5489_/A VGND VPWR _5490_/A VGND VPWR sky130_fd_sc_hd__clkbuf_2
X_7159_ _6667_/Y _7040_/C _6754_/Y _7059_/C VGND VPWR _7159_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_58_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_608 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_384 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_30 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_346 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_96 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_362 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_462 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_50 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_210 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_338 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_224 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_555 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_246 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_611 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4860_ _4860_/A VGND VPWR _4860_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_178_616 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4791_ _4791_/A _4791_/B _4791_/C _4791_/D VGND VPWR _4936_/B VGND VPWR sky130_fd_sc_hd__and4_1
X_6530_ _6528_/Y _5897_/B _6529_/Y _5024_/B VGND VPWR _6530_/X VGND VPWR sky130_fd_sc_hd__o22a_2
XANTENNA_17 _7375_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_39 _4842_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_28 _4481_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_6461_ _9342_/Q VGND VPWR _6461_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_173_310 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_384 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_343 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6392_ _9394_/Q VGND VPWR _6392_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9180_ _9613_/CLK _9180_/D _9646_/SET_B VGND VPWR _9180_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_8200_ _8218_/A _8200_/B _8200_/C VGND VPWR _8377_/C VGND VPWR sky130_fd_sc_hd__or3_2
X_5412_ _5671_/A _5412_/B VGND VPWR _5413_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_5343_ _9484_/Q _5338_/A _5967_/B1 _5338_/Y VGND VPWR _9484_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8131_ _8131_/A _8676_/A _8357_/A _8573_/A VGND VPWR _8136_/A VGND VPWR sky130_fd_sc_hd__or4_1
XFILLER_99_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_176 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5274_ _9531_/Q _5269_/A _8929_/A1 _5269_/Y VGND VPWR _9531_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8062_ _8062_/A _8062_/B VGND VPWR _8065_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_101_126 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7013_ _7013_/A VGND VPWR _7014_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_95_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_202 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8964_ _7743_/X _8964_/A1 _8975_/S VGND VPWR _8964_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_102_13 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8895_ _8894_/X _9148_/Q _9054_/Q VGND VPWR _8895_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_7915_ _8226_/C _8319_/A VGND VPWR _8254_/B VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_70_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_7846_ _8394_/A _8394_/B _8394_/C _8195_/A VGND VPWR _7847_/A VGND VPWR sky130_fd_sc_hd__or4_1
XFILLER_184_608 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7777_ _7777_/A VGND VPWR _7777_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_4989_ _9091_/Q _9090_/Q _9092_/Q VGND VPWR _4989_/X VGND VPWR sky130_fd_sc_hd__o21a_1
XFILLER_11_327 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6728_ _6723_/Y _5404_/B _6724_/Y _5496_/B _6727_/X VGND VPWR _6741_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9516_ _9771_/CLK _9516_/D _4628_/A VGND VPWR _9516_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_176_192 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6659_ _4921_/A _6158_/A _6658_/Y _4481_/B _6158_/X VGND VPWR _6659_/X VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9447_ _9791_/CLK _9447_/D _9633_/SET_B VGND VPWR _9447_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_9378_ _9378_/CLK _9378_/D _9646_/SET_B VGND VPWR _9378_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_8329_ _8662_/A _8600_/A _8329_/C VGND VPWR _8331_/A VGND VPWR sky130_fd_sc_hd__or3_1
XFILLER_117_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_402 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_36 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_500 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_382 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_471 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_460 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_50 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_360 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_72 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput37 mgmt_gpio_in[10] VGND VPWR input37/X VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
Xinput15 mask_rev_in[1] VGND VPWR _6813_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput26 mask_rev_in[2] VGND VPWR _6706_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_143_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_568 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput48 mgmt_gpio_in[20] VGND VPWR _6450_/A VGND VPWR sky130_fd_sc_hd__clkbuf_2
Xinput59 mgmt_gpio_in[30] VGND VPWR _6193_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_182_162 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_6 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_500 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_566 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5961_ _5961_/A VGND VPWR _5962_/A VGND VPWR sky130_fd_sc_hd__clkbuf_2
X_4912_ _6158_/A _4925_/A _4909_/Y _4910_/Y _5278_/B VGND VPWR _4912_/X VGND VPWR
+ sky130_fd_sc_hd__o32a_1
X_8680_ _8716_/D _8731_/D _8680_/C _8720_/A VGND VPWR _8680_/Y VGND VPWR sky130_fd_sc_hd__nor4_2
X_7700_ _7700_/A VGND VPWR _7700_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_7631_ _6856_/Y _7427_/X _6938_/Y _5699_/X VGND VPWR _7631_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_5892_ _5892_/A1 _8879_/X _8924_/X _9141_/Q VGND VPWR _9141_/D VGND VPWR sky130_fd_sc_hd__o22a_2
XFILLER_33_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4843_ _4929_/A _4843_/B VGND VPWR _5968_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_33_496 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7562_ _6315_/Y _7425_/X _7559_/X _7561_/X VGND VPWR _7572_/C VGND VPWR sky130_fd_sc_hd__o211a_1
X_4774_ _6158_/B _4843_/B VGND VPWR _5045_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_165_129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_168 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7493_ _6793_/Y _7455_/X _6908_/Y _7457_/X VGND VPWR _7493_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_6513_ _6508_/Y _5556_/B _8763_/A _5572_/B _6512_/X VGND VPWR _6526_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9301_ _9788_/CLK _9301_/D _9295_/SET_B VGND VPWR _9301_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_146_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6444_ _6444_/A VGND VPWR _6444_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9232_ _9508_/CLK _9232_/D _9528_/SET_B VGND VPWR _9232_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6375_ _6373_/Y _5789_/B _6374_/Y _5768_/B VGND VPWR _6375_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_9163_ _9532_/CLK _9163_/D _9647_/SET_B VGND VPWR _9163_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_8114_ _8164_/A VGND VPWR _8114_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_5326_ _9495_/Q _5319_/A _8930_/A1 _5319_/Y VGND VPWR _9495_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_9094_ _9501_/CLK _9094_/D _9647_/SET_B VGND VPWR _9094_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_87_102 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5257_ _9542_/Q _5253_/A _5966_/B1 _5253_/Y VGND VPWR _9542_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8045_ _8045_/A _8615_/B VGND VPWR _8047_/A VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_180_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5188_ _9587_/Q _5939_/A _5108_/X _4551_/X VGND VPWR _9587_/D VGND VPWR sky130_fd_sc_hd__a211o_1
XFILLER_56_500 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_544 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_38 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8947_ _9715_/Q _6326_/Y _8957_/S VGND VPWR _8947_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_73_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_49 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8878_ _7199_/Y _9635_/Q _8959_/S VGND VPWR _8878_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_11_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_7829_ _7829_/A VGND VPWR _8376_/A VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_11_102 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_135 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_75 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_471 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_64 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_376 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_102 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_243 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_202 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_430 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_82 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_343 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4490_ _4911_/A _4805_/A VGND VPWR _4491_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_170_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_379 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6160_ _9500_/Q VGND VPWR _6160_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_69_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5111_ _5111_/A VGND VPWR _5112_/A VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_69_146 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6091_ _9379_/Q VGND VPWR _6091_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_85_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_116 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5042_ _8971_/X _4551_/B _9677_/Q _5062_/D VGND VPWR _9677_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_38_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_352 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_599 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8801_ _8801_/A _8801_/B VGND VPWR _8802_/A VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_25_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_547 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6993_ _9054_/Q _8819_/X _9054_/Q _6997_/C _9055_/Q VGND VPWR _9054_/D VGND VPWR
+ sky130_fd_sc_hd__a221o_2
X_9781_ _9785_/CLK _9781_/D _9779_/SET_B VGND VPWR _9781_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_51_csclk _9329_/CLK VGND VPWR _9768_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_18_290 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8732_ _8732_/A VGND VPWR _8732_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_5944_ _9118_/Q _5943_/A _5963_/B1 _5943_/Y VGND VPWR _9118_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_80_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_400 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5875_ _9158_/Q _5874_/A _8846_/X _5874_/Y VGND VPWR _9158_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8663_ _8696_/C _8727_/C _8663_/C _8721_/A VGND VPWR _8664_/A VGND VPWR sky130_fd_sc_hd__or4_1
X_7614_ _4800_/Y _7434_/X _4930_/Y _7436_/X VGND VPWR _7614_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_8594_ _8594_/A _8594_/B _7896_/X VGND VPWR _8595_/A VGND VPWR sky130_fd_sc_hd__or3b_1
X_4826_ _6111_/A _4927_/A VGND VPWR _5227_/B VGND VPWR sky130_fd_sc_hd__or2_1
X_7545_ _6357_/Y _7445_/X _6328_/Y _7447_/X VGND VPWR _7545_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_21_499 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_354 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4757_ _4787_/A _4891_/A _4753_/Y _4754_/Y _6135_/A VGND VPWR _4757_/X VGND VPWR
+ sky130_fd_sc_hd__o32a_1
XFILLER_111_9 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7476_ _7476_/A _9251_/Q _7476_/C _9255_/Q VGND VPWR _7477_/A VGND VPWR sky130_fd_sc_hd__or4_1
X_4688_ _4729_/A _8944_/X _8934_/X _4729_/D VGND VPWR _6086_/B VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_108_12 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9215_ _9758_/CLK _9215_/D _9779_/SET_B VGND VPWR _9215_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6427_ _9498_/Q VGND VPWR _6427_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_161_143 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6358_ _9772_/Q _6251_/Y _6357_/Y _5420_/B VGND VPWR _6358_/X VGND VPWR sky130_fd_sc_hd__o2bb2a_2
X_9146_ _9280_/CLK _9146_/D _9757_/SET_B VGND VPWR _9146_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_102_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_315 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5309_ _9509_/Q _5308_/A _8846_/X _5308_/Y VGND VPWR _9509_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_9077_ _9687_/CLK _9077_/D _9685_/SET_B VGND VPWR _9077_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6289_ _9753_/Q VGND VPWR _6289_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_102_287 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8028_ _8521_/A _8550_/A VGND VPWR _8410_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_124_88 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_160 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_42 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_19_csclk clkbuf_2_3_0_csclk/X VGND VPWR _9509_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XPHY_200 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_222 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_211 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_411 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_266 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_255 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_244 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_299 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_288 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_235 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_466 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_499 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_110 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_316 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_187 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_444 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_606 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_447 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_7 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_108 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_536 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_92 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5660_ _6052_/A _5660_/B VGND VPWR _5661_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_4611_ _8934_/X _8932_/X _4729_/A _8944_/X VGND VPWR _6158_/B VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_175_268 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5591_ _9314_/Q _5585_/A _8841_/X _5585_/Y VGND VPWR _9314_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7330_ _7330_/A _7330_/B _7330_/C _7330_/D VGND VPWR _7331_/C VGND VPWR sky130_fd_sc_hd__and4_1
X_4542_ _9065_/Q VGND VPWR _7731_/A VGND VPWR sky130_fd_sc_hd__clkinv_2
X_7261_ _6200_/Y _5728_/X _6230_/Y _7040_/A _7260_/X VGND VPWR _7264_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_4473_ _8932_/X VGND VPWR _4729_/D VGND VPWR sky130_fd_sc_hd__clkinv_2
X_9000_ _9568_/Q _8777_/A VGND VPWR mgmt_gpio_out[23] VGND VPWR sky130_fd_sc_hd__ebufn_8
X_6212_ _9157_/Q VGND VPWR _6212_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
XFILLER_131_327 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7192_ _8779_/A _7118_/X _8799_/A _7048_/C VGND VPWR _7192_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_6143_ _7282_/A _5610_/B _6139_/Y _5679_/B _6142_/X VGND VPWR _6144_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_6074_ _9431_/Q VGND VPWR _6074_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
XFILLER_85_469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5025_ _5025_/A VGND VPWR _5026_/A VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_38_341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_491 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_374 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_18 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_9764_ _9770_/CLK _9764_/D _7011_/B VGND VPWR _9764_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_6976_ _6976_/A VGND VPWR _6976_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_26_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_8715_ _8715_/A _8715_/B _8715_/C VGND VPWR _8716_/B VGND VPWR sky130_fd_sc_hd__or3_1
X_5927_ _7771_/A _7771_/B _7771_/C _7771_/D VGND VPWR _5928_/C VGND VPWR sky130_fd_sc_hd__or4_1
X_9695_ _9695_/CLK _9695_/D _9779_/SET_B VGND VPWR _9695_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_139_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_427 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5858_ _5849_/X _8857_/X _8924_/X _9168_/Q VGND VPWR _9168_/D VGND VPWR sky130_fd_sc_hd__o22a_2
X_8646_ _8646_/A _8646_/B VGND VPWR _8678_/C VGND VPWR sky130_fd_sc_hd__or2_1
X_8577_ _8577_/A _8577_/B _8577_/C VGND VPWR _8675_/C VGND VPWR sky130_fd_sc_hd__or3_1
X_5789_ _5960_/A _5789_/B VGND VPWR _5790_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_4809_ _9541_/Q VGND VPWR _4809_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_5_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7528_ _8755_/A _7441_/X _8791_/A _7443_/X _7527_/X VGND VPWR _7535_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_147_482 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_132 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_66 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7459_ _4740_/Y _7451_/X _4916_/Y _7453_/X _7458_/X VGND VPWR _7480_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_107_368 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_9129_ _9129_/CLK _9129_/D _9779_/SET_B VGND VPWR _9129_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_76_414 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_330 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_127 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_344 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_130 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_580 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_555 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_94 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_89 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_60 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_296 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_299 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_355 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6830_ _6830_/A _6830_/B _6830_/C _6830_/D VGND VPWR _6946_/A VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_35_344 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_388 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_152 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6761_ _9548_/Q VGND VPWR _6761_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_8500_ _8695_/A _8659_/A _8594_/B _7892_/X VGND VPWR _8501_/D VGND VPWR sky130_fd_sc_hd__or4b_1
X_5712_ _5724_/B _5704_/Y _5710_/Y _9252_/Q _5713_/A VGND VPWR _9252_/D VGND VPWR
+ sky130_fd_sc_hd__o32a_1
XFILLER_188_360 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6692_ _9780_/Q VGND VPWR _6692_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9480_ _9527_/CLK _9480_/D _9685_/SET_B VGND VPWR _9480_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_5643_ _9056_/Q VGND VPWR _5643_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_8431_ _8431_/A _8431_/B VGND VPWR _8432_/C VGND VPWR sky130_fd_sc_hd__or2_1
X_5574_ _5574_/A VGND VPWR _5574_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_8362_ _8362_/A _8362_/B VGND VPWR _8575_/C VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_191_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_7313_ _6940_/Y _7040_/C _6922_/Y _7059_/C VGND VPWR _7313_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4525_ _4525_/A VGND VPWR _4526_/A VGND VPWR sky130_fd_sc_hd__clkbuf_4
X_8293_ _8377_/C _8204_/A _9067_/Q VGND VPWR _8650_/C VGND VPWR sky130_fd_sc_hd__o21ai_2
XFILLER_131_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_327 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4456_ _9587_/Q VGND VPWR _4456_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_171_271 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7244_ _6159_/Y _7086_/X _6225_/Y _7088_/X VGND VPWR _7244_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_7175_ _6767_/Y _7124_/X _6738_/Y _7068_/B _7174_/X VGND VPWR _7176_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_6126_ _9225_/Q VGND VPWR _6126_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_85_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_244 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6057_ _9045_/Q _6054_/A _8930_/A1 _6054_/Y VGND VPWR _9045_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XANTENNA_107 input77/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_5008_ _5008_/A VGND VPWR _9697_/D VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA_118 input86/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_129 input86/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_41_314 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_196 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9747_ _9777_/CLK _9747_/D _9757_/SET_B VGND VPWR _9747_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6959_ _6946_/Y _6952_/A _9029_/Q _6952_/Y VGND VPWR _9029_/D VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_14_32 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9678_ _9681_/CLK _9678_/D _6146_/A VGND VPWR _9678_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_8629_ _8710_/A _8629_/B _8686_/D _8628_/X VGND VPWR _8633_/A VGND VPWR sky130_fd_sc_hd__or4b_2
XFILLER_139_268 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_154 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_443 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_130 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_380 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_544 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_82 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xoutput317 _9763_/Q VGND VPWR sram_ro_addr[1] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput306 _8819_/X VGND VPWR serial_clock VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_5290_ _5671_/A _5290_/B VGND VPWR _5291_/A VGND VPWR sky130_fd_sc_hd__or2_1
Xoutput328 _9014_/Q VGND VPWR wb_dat_o[10] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput339 _9032_/Q VGND VPWR wb_dat_o[20] VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_141_455 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_292 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_308 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8980_ _9581_/Q _7705_/A VGND VPWR mgmt_gpio_out[3] VGND VPWR sky130_fd_sc_hd__ebufn_8
XFILLER_48_480 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7931_ _7931_/A _7931_/B VGND VPWR _7931_/X VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_70_409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_612 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7862_ _8260_/A VGND VPWR _7862_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9601_ _9601_/CLK _9601_/D _9295_/SET_B VGND VPWR _9601_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_90_291 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6813_ _6813_/A VGND VPWR _6813_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7793_ _8189_/A _7791_/B _7792_/B VGND VPWR _8538_/B VGND VPWR sky130_fd_sc_hd__a21o_2
X_6744_ _6744_/A VGND VPWR _6744_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9532_ _9532_/CLK _9532_/D _9647_/SET_B VGND VPWR _9532_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_167_19 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_380 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6675_ _9723_/Q VGND VPWR _6675_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9463_ _9514_/CLK _9463_/D _4628_/A VGND VPWR _9463_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_164_503 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_8414_ _8627_/C VGND VPWR _8414_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_5626_ _9291_/Q _5623_/A _8844_/X _5623_/Y VGND VPWR _9291_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_9394_ _9483_/CLK _9394_/D _9528_/SET_B VGND VPWR _9394_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_8345_ _8345_/A _8345_/B VGND VPWR _8377_/B VGND VPWR sky130_fd_sc_hd__or2_1
X_5557_ _5557_/A VGND VPWR _5558_/A VGND VPWR sky130_fd_sc_hd__clkbuf_2
X_4508_ _9776_/Q _4506_/A _5964_/B1 _4506_/Y VGND VPWR _9776_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8276_ _8660_/A _8660_/B _8496_/A VGND VPWR _8280_/B VGND VPWR sky130_fd_sc_hd__or3_2
X_5488_ _5671_/A _5488_/B VGND VPWR _5489_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_116_23 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_135 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_455 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7227_ _6240_/Y _7097_/X _6271_/Y _7099_/X VGND VPWR _7227_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_132_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7158_ _6717_/Y _7082_/X _6704_/Y _7084_/X _7157_/X VGND VPWR _7177_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_6109_ _9535_/Q VGND VPWR _6109_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7089_ _4916_/Y _7086_/X _4914_/Y _7088_/X VGND VPWR _7089_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_86_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_428 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_396 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_31 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_37 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_612 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_64 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_308 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_358 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_374 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_528 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_399 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_263 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_499 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_266 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_152 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4790_ _4790_/A _4790_/B _4790_/C _4790_/D VGND VPWR _4791_/D VGND VPWR sky130_fd_sc_hd__and4_1
XANTENNA_18 _7397_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_29 _5178_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_6460_ _8808_/B _6134_/A _6456_/Y _5949_/B _6459_/X VGND VPWR _6473_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_6391_ _9462_/Q VGND VPWR _6391_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_5411_ _9437_/Q _5406_/A _5967_/B1 _5406_/Y VGND VPWR _9437_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_161_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_208 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5342_ _9485_/Q _5338_/A _5966_/B1 _5338_/Y VGND VPWR _9485_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8130_ _8213_/A _8130_/B VGND VPWR _8573_/A VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_99_133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8061_ _8061_/A _8064_/B _8061_/C VGND VPWR _8062_/B VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_114_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5273_ _9532_/Q _5269_/A _8843_/X _5269_/Y VGND VPWR _9532_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7012_ _9626_/Q input86/X VGND VPWR _7013_/A VGND VPWR sky130_fd_sc_hd__or2b_1
XFILLER_68_553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_214 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_8963_ _7741_/X _8963_/A1 _8975_/S VGND VPWR _8963_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_102_25 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7914_ _8521_/B _8246_/B VGND VPWR _8317_/A VGND VPWR sky130_fd_sc_hd__nor2_1
X_8894_ _7375_/Y _9630_/Q _8959_/S VGND VPWR _8894_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_7845_ _7845_/A VGND VPWR _8305_/A VGND VPWR sky130_fd_sc_hd__buf_8
XFILLER_62_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7776_ _8189_/A _7791_/B _7966_/A _7966_/C VGND VPWR _7777_/A VGND VPWR sky130_fd_sc_hd__or4_1
X_4988_ _9700_/Q _9699_/Q VGND VPWR _5992_/B VGND VPWR sky130_fd_sc_hd__nor2_1
X_9515_ _9545_/CLK _9515_/D _4628_/A VGND VPWR _9515_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6727_ _6725_/Y _5232_/B _6726_/Y _4822_/X VGND VPWR _6727_/X VGND VPWR sky130_fd_sc_hd__o22a_2
XFILLER_127_7 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_160 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9446_ _9791_/CLK _9446_/D _9779_/SET_B VGND VPWR _9446_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6658_ _9788_/Q VGND VPWR _6658_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
X_5609_ _9302_/Q _5604_/A _5967_/B1 _5604_/Y VGND VPWR _9302_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_9377_ _9378_/CLK _9377_/D _9646_/SET_B VGND VPWR _9377_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_191_163 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_528 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6589_ _9466_/Q VGND VPWR _6589_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_8328_ _7848_/A _8300_/B _8327_/Y VGND VPWR _8329_/C VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_117_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_8259_ _8259_/A _8367_/B VGND VPWR _8261_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_87_48 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_414 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_512 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_87 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_483 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_414 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_188 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xinput16 mask_rev_in[20] VGND VPWR _6385_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput27 mask_rev_in[30] VGND VPWR _6207_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput38 mgmt_gpio_in[11] VGND VPWR _6505_/A VGND VPWR sky130_fd_sc_hd__buf_6
Xinput49 mgmt_gpio_in[21] VGND VPWR input49/X VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_143_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_580 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_526 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5960_ _5960_/A _5960_/B VGND VPWR _5961_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_65_578 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_91 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_548 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4911_ _4911_/A _6086_/B VGND VPWR _5278_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_5891_ _5891_/A1 _8881_/X _8924_/X _9142_/Q VGND VPWR _9142_/D VGND VPWR sky130_fd_sc_hd__o22a_2
X_7630_ _6932_/Y _7415_/X _6800_/Y _7417_/X _7629_/X VGND VPWR _7644_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_4842_ _9093_/Q VGND VPWR _4842_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
XFILLER_20_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4773_ _9667_/Q VGND VPWR _4773_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7561_ _6304_/Y _7430_/X _6263_/Y _7432_/X _7560_/X VGND VPWR _7561_/X VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_6512_ _6510_/Y _5671_/B _8753_/A _5776_/B VGND VPWR _6512_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_7492_ _6939_/Y _7441_/X _6787_/Y _7443_/X _7491_/X VGND VPWR _7499_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9300_ _9788_/CLK _9300_/D _9295_/SET_B VGND VPWR _9300_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_9231_ _9508_/CLK _9231_/D _9528_/SET_B VGND VPWR _9231_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6443_ _6438_/Y _4841_/X _6439_/Y _5089_/B _6442_/X VGND VPWR _6443_/X VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_173_196 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6374_ _9230_/Q VGND VPWR _6374_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9162_ _9358_/CLK _9162_/D _9685_/SET_B VGND VPWR _9162_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_5325_ _9496_/Q _5319_/A _8841_/X _5319_/Y VGND VPWR _9496_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_9093_ _9501_/CLK _9093_/D _9647_/SET_B VGND VPWR _9093_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_8113_ _8401_/A _8378_/B VGND VPWR _8354_/A VGND VPWR sky130_fd_sc_hd__nor2_1
X_5256_ _9543_/Q _5253_/A _5965_/B1 _5253_/Y VGND VPWR _9543_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8044_ _8521_/A _8554_/A VGND VPWR _8615_/B VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_102_469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_9 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_350 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5187_ _9059_/Q VGND VPWR _5939_/A VGND VPWR sky130_fd_sc_hd__inv_2
X_8946_ _8945_/X _9676_/Q _9587_/Q VGND VPWR _8946_/X VGND VPWR sky130_fd_sc_hd__mux2_4
XFILLER_56_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_8877_ _8876_/X _9139_/Q _9054_/Q VGND VPWR _8877_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_464 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7828_ _8097_/B _8660_/B _8660_/C VGND VPWR _7829_/A VGND VPWR sky130_fd_sc_hd__or3_1
X_7759_ _8525_/A _7894_/B _7903_/C _8528_/A VGND VPWR _8394_/D VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_11_147 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_620 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_9429_ _9508_/CLK _9429_/D _9295_/SET_B VGND VPWR _9429_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_137_388 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_358 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_230 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_512 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_236 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_375 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_442 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_288 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6090_ _9405_/Q VGND VPWR _6090_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_5110_ _5545_/A _5110_/B VGND VPWR _5111_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_5041_ _8972_/X _4551_/B _9678_/Q _5062_/D VGND VPWR _9678_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_69_158 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_128 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_364 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9780_ _9785_/CLK _9780_/D _9779_/SET_B VGND VPWR _9780_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
Xclkbuf_0_wb_clk_i wb_clk_i VGND VPWR clkbuf_0_wb_clk_i/X VGND VPWR sky130_fd_sc_hd__clkbuf_16
X_8800_ _8800_/A VGND VPWR _8800_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_25_217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8731_ _8731_/A _8731_/B _8731_/C _8731_/D VGND VPWR _8731_/X VGND VPWR sky130_fd_sc_hd__or4_1
X_6992_ _5643_/Y _5753_/B _9053_/Q _6991_/Y VGND VPWR _9053_/D VGND VPWR sky130_fd_sc_hd__a2bb2o_1
XFILLER_80_334 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5943_ _5943_/A VGND VPWR _5943_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_178_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5874_ _5874_/A VGND VPWR _5874_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_8662_ _8662_/A _8662_/B _8662_/C _8661_/X VGND VPWR _8663_/C VGND VPWR sky130_fd_sc_hd__or4b_2
X_4825_ _9559_/Q VGND VPWR _8807_/A VGND VPWR sky130_fd_sc_hd__inv_2
X_8593_ _7836_/B _8591_/Y _8641_/A _8501_/C VGND VPWR _8695_/D VGND VPWR sky130_fd_sc_hd__a211o_1
X_7613_ _4858_/Y _7427_/X _4718_/Y _5699_/X VGND VPWR _7613_/X VGND VPWR sky130_fd_sc_hd__o22a_2
XFILLER_193_236 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_7544_ _6456_/Y _7425_/X _7541_/X _7543_/X VGND VPWR _7554_/C VGND VPWR sky130_fd_sc_hd__o211a_1
X_4756_ _4756_/A VGND VPWR _6135_/A VGND VPWR sky130_fd_sc_hd__buf_8
XFILLER_162_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_366 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7475_ _7475_/A VGND VPWR _7475_/X VGND VPWR sky130_fd_sc_hd__buf_8
X_4687_ _9106_/Q VGND VPWR _4687_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_108_24 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_9214_ _9655_/CLK _9214_/D _9779_/SET_B VGND VPWR _9214_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6426_ _6421_/Y _5496_/B _6422_/Y _5393_/B _6425_/X VGND VPWR _6433_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_6357_ _9428_/Q VGND VPWR _6357_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9145_ _9203_/CLK _9145_/D _9633_/SET_B VGND VPWR _9145_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_161_199 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_520 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5308_ _5308_/A VGND VPWR _5308_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_130_542 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6288_ _9209_/Q VGND VPWR _6288_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9076_ _9687_/CLK _9076_/D _9685_/SET_B VGND VPWR _9076_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_48_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5239_ _9554_/Q _5234_/A _5967_/B1 _5234_/Y VGND VPWR _9554_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8027_ _8389_/A _8137_/B _8097_/B _8137_/B _8026_/X VGND VPWR _8027_/X VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_84_38 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_556 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_55 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8929_ _9613_/Q _8929_/A1 _8930_/S VGND VPWR _8929_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XPHY_234 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_223 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_212 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_267 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_256 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_278 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_247 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_40 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_459 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_4610_ _9726_/Q _4604_/A _5967_/B1 _4604_/Y VGND VPWR _9726_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_5590_ _9315_/Q _5585_/A _8929_/A1 _5585_/Y VGND VPWR _9315_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_30_275 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_206 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4541_ _4541_/A VGND VPWR _9760_/D VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_190_239 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_100 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7260_ _7260_/A _7392_/B VGND VPWR _7260_/X VGND VPWR sky130_fd_sc_hd__or2_1
X_4472_ _8934_/X VGND VPWR _4669_/A VGND VPWR sky130_fd_sc_hd__clkinv_2
X_7191_ _8747_/A _7040_/D _8765_/A _7110_/X _7190_/X VGND VPWR _7198_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_6211_ _6211_/A _6211_/B _6211_/C _6211_/D VGND VPWR _6237_/C VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_143_188 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6142_ _6140_/Y _5818_/B _6141_/Y _5572_/B VGND VPWR _6142_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_6073_ _9501_/Q VGND VPWR _6073_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_57_139 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5024_ _5259_/A _5024_/B VGND VPWR _5025_/A VGND VPWR sky130_fd_sc_hd__or2_2
XFILLER_38_353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9763_ _9770_/CLK _9763_/D _7011_/B VGND VPWR _9763_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_6975_ _6975_/A VGND VPWR _6976_/A VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_80_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5926_ _7770_/A _7770_/B _7768_/A _7768_/B VGND VPWR _5936_/B VGND VPWR sky130_fd_sc_hd__or4_1
X_8714_ _8714_/A _8714_/B _8714_/C _8714_/D VGND VPWR _8739_/A VGND VPWR sky130_fd_sc_hd__or4_1
X_9694_ _9695_/CLK _9694_/D _9779_/SET_B VGND VPWR _9694_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_8645_ _8645_/A _8645_/B _8645_/C _8645_/D VGND VPWR _8716_/C VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_80_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_439 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5857_ _5849_/X _8859_/X _8924_/X _9169_/Q VGND VPWR _9169_/D VGND VPWR sky130_fd_sc_hd__o22a_2
X_4808_ _4808_/A VGND VPWR _4808_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_186_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_8576_ _8576_/A _8642_/D _8730_/D _8576_/D VGND VPWR _8580_/A VGND VPWR sky130_fd_sc_hd__or4_1
X_5788_ _9277_/Q _9056_/Q _5787_/Y _9217_/Q _5755_/A VGND VPWR _9217_/D VGND VPWR
+ sky130_fd_sc_hd__a32o_1
X_7527_ _8771_/A _7445_/X _8769_/A _7447_/X VGND VPWR _7527_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4739_ _4739_/A VGND VPWR _6134_/A VGND VPWR sky130_fd_sc_hd__buf_6
X_7458_ _4804_/Y _7455_/X _4769_/Y _7457_/X VGND VPWR _7458_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_6409_ _9415_/Q VGND VPWR _6409_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_7389_ _6434_/Y _7040_/D _6363_/Y _7110_/X _7388_/X VGND VPWR _7396_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_103_520 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_9128_ _9379_/CLK _9128_/D _9779_/SET_B VGND VPWR _9128_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_9059_ _4450_/A1 _9059_/D _6146_/A VGND VPWR _9059_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_88_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_356 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_142 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_164 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_592 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_518 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_50_csclk _9329_/CLK VGND VPWR _9770_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_69_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_72 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_106 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_164 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6760_ _9504_/Q VGND VPWR _6760_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
XFILLER_62_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5711_ _9053_/Q _9055_/Q VGND VPWR _5713_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_6691_ _6691_/A _6691_/B _6691_/C _6691_/D VGND VPWR _6785_/B VGND VPWR sky130_fd_sc_hd__and4_1
X_5642_ _9054_/Q VGND VPWR _6997_/A VGND VPWR sky130_fd_sc_hd__inv_2
X_8430_ _8430_/A _8560_/B VGND VPWR _8431_/B VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_176_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8361_ _8361_/A _8361_/B VGND VPWR _8730_/C VGND VPWR sky130_fd_sc_hd__or2_1
X_5573_ _5573_/A VGND VPWR _5574_/A VGND VPWR sky130_fd_sc_hd__clkbuf_4
X_7312_ _6848_/Y _7082_/X _6824_/Y _7084_/X _7311_/X VGND VPWR _7331_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_4524_ _5960_/A _4524_/B VGND VPWR _4525_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_8292_ _8514_/A _8292_/B VGND VPWR _8294_/A VGND VPWR sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_18_csclk clkbuf_2_3_0_csclk/X VGND VPWR _9483_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_104_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_4455_ _8936_/X VGND VPWR _4661_/C VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_131_103 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7243_ _7243_/A _7243_/B _7243_/C VGND VPWR _7243_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
XFILLER_104_339 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7174_ _6650_/Y _7126_/X _6692_/Y _7128_/X VGND VPWR _7174_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_131_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_14 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6125_ _6120_/Y _5013_/B _6121_/Y _5797_/B _6124_/X VGND VPWR _6144_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_100_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_256 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6056_ _9046_/Q _6054_/A _8955_/A1 _6054_/Y VGND VPWR _9046_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_5007_ _4949_/A _9697_/Q _5007_/S VGND VPWR _5008_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_119 input86/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_108 input77/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_121_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9746_ _9777_/CLK _9746_/D _9757_/SET_B VGND VPWR _9746_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_157_7 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6958_ _6785_/Y _6952_/A _9030_/Q _6952_/Y VGND VPWR _9030_/D VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_41_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_359 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_44 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5909_ _9131_/Q _5907_/A _8845_/X _5907_/Y VGND VPWR _9131_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_9677_ _9681_/CLK _9677_/D _6146_/A VGND VPWR _9677_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6889_ _9152_/Q VGND VPWR _6889_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_139_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_534 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8628_ _8130_/B _8554_/B _8454_/B _8133_/A _8408_/Y VGND VPWR _8628_/X VGND VPWR
+ sky130_fd_sc_hd__o2111a_1
XFILLER_108_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_8559_ _8559_/A _8709_/A _8631_/B _8688_/B VGND VPWR _8563_/A VGND VPWR sky130_fd_sc_hd__or4_1
XFILLER_5_216 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_431 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_400 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_466 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_75 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_40 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_136 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_158 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_331 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_392 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_94 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput307 _8822_/X VGND VPWR serial_data_1 VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput318 _9764_/Q VGND VPWR sram_ro_addr[2] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput329 _9015_/Q VGND VPWR wb_dat_o[11] VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_99_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_467 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7930_ _7848_/A _8305_/A _7929_/Y VGND VPWR _7931_/B VGND VPWR sky130_fd_sc_hd__o21ba_1
XFILLER_48_492 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7861_ _8305_/A VGND VPWR _8299_/B VGND VPWR sky130_fd_sc_hd__inv_2
X_9600_ _9601_/CLK _9600_/D _9295_/SET_B VGND VPWR _9600_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6812_ _9774_/Q VGND VPWR _6812_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
XFILLER_23_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7792_ _8525_/A _7792_/B VGND VPWR _7823_/B VGND VPWR sky130_fd_sc_hd__nor2_1
X_9531_ _9535_/CLK _9531_/D _9528_/SET_B VGND VPWR _9531_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_6743_ _9122_/Q VGND VPWR _6743_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_176_342 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6674_ _9161_/Q VGND VPWR _6674_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9462_ _9532_/CLK _9462_/D _9647_/SET_B VGND VPWR _9462_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_5625_ _9292_/Q _5623_/A _8845_/X _5623_/Y VGND VPWR _9292_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8413_ _8614_/B _8575_/A VGND VPWR _8627_/C VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_176_397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9393_ _9509_/CLK _9393_/D _9528_/SET_B VGND VPWR _9393_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_191_367 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_8344_ _8279_/A _8378_/B _8640_/A _8279_/C _8311_/B VGND VPWR _8352_/A VGND VPWR
+ sky130_fd_sc_hd__o32a_2
X_5556_ _5671_/A _5556_/B VGND VPWR _5557_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_132_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5487_ _9385_/Q _5482_/A _5967_/B1 _5482_/Y VGND VPWR _9385_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_4507_ _9777_/Q _4506_/A _5963_/B1 _4506_/Y VGND VPWR _9777_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8275_ _8275_/A _8693_/B VGND VPWR _8275_/X VGND VPWR sky130_fd_sc_hd__or2_2
X_7226_ _6298_/Y _7048_/B _6297_/Y _7077_/A _7225_/X VGND VPWR _7233_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_132_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_467 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_510 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7157_ _6664_/Y _7077_/C _6693_/Y _7077_/D _7156_/X VGND VPWR _7157_/X VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_76_17 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6108_ _6103_/Y _5431_/B _6104_/Y _6027_/B _6107_/X VGND VPWR _6119_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_7088_ _7088_/A VGND VPWR _7088_/X VGND VPWR sky130_fd_sc_hd__buf_8
XFILLER_132_34 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_270 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_98 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_9729_ _9774_/CLK _9729_/D _9757_/SET_B VGND VPWR _9729_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_41_189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_386 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_275 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_19 _7500_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_146_537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5410_ _9438_/Q _5406_/A _5966_/B1 _5406_/Y VGND VPWR _9438_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_6390_ _9472_/Q VGND VPWR _6390_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
XFILLER_161_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5341_ _9486_/Q _5338_/A _5965_/B1 _5338_/Y VGND VPWR _9486_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8060_ _8060_/A VGND VPWR _8061_/C VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_99_145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5272_ _9533_/Q _5269_/A _8844_/X _5269_/Y VGND VPWR _9533_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7011_ _9586_/Q _7011_/B VGND VPWR _7011_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_141_275 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_106 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_139 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_8962_ _7739_/X _8962_/A1 _8975_/S VGND VPWR _8962_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_7913_ _8077_/A _8246_/B _7864_/X _8316_/A _7912_/X VGND VPWR _7917_/B VGND VPWR
+ sky130_fd_sc_hd__o221ai_1
X_8893_ _8892_/X _9147_/Q _9054_/Q VGND VPWR _8893_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_7844_ _8394_/A _8379_/B _8394_/C _8195_/A VGND VPWR _7845_/A VGND VPWR sky130_fd_sc_hd__or4_1
XFILLER_24_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_443 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_19 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7775_ _8193_/A _7775_/B _7775_/C _7775_/D VGND VPWR _7966_/C VGND VPWR sky130_fd_sc_hd__or4_1
X_9514_ _9514_/CLK _9514_/D _4628_/A VGND VPWR _9514_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6726_ _6726_/A VGND VPWR _6726_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_4987_ _4987_/A VGND VPWR _4987_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_6657_ _9434_/Q VGND VPWR _6657_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9445_ _9791_/CLK _9445_/D _9633_/SET_B VGND VPWR _9445_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_164_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5608_ _9303_/Q _5604_/A _5966_/B1 _5604_/Y VGND VPWR _9303_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_9376_ _9379_/CLK _9376_/D _9779_/SET_B VGND VPWR _9376_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6588_ _9505_/Q VGND VPWR _8777_/A VGND VPWR sky130_fd_sc_hd__inv_6
XFILLER_105_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_570 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5539_ _9351_/Q _5536_/A _8844_/X _5536_/Y VGND VPWR _9351_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8327_ _8327_/A _8599_/C _8506_/C _8693_/C VGND VPWR _8327_/Y VGND VPWR sky130_fd_sc_hd__nor4_2
XFILLER_127_89 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_264 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_8258_ _8510_/A _8262_/B VGND VPWR _8367_/B VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_59_521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7209_ _6372_/Y _7068_/A _6402_/Y _7105_/X VGND VPWR _7209_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_8189_ _8189_/A _8213_/A VGND VPWR _8189_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_143_44 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_524 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_426 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xinput17 mask_rev_in[21] VGND VPWR _6262_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput28 mask_rev_in[31] VGND VPWR _6106_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput39 mgmt_gpio_in[12] VGND VPWR _6455_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_143_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_451 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_387 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5890_ _5890_/A1 _8883_/X _8924_/X _9143_/Q VGND VPWR _9143_/D VGND VPWR sky130_fd_sc_hd__o22a_2
X_4910_ _9520_/Q VGND VPWR _4910_/Y VGND VPWR sky130_fd_sc_hd__inv_4
XFILLER_45_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4841_ _6111_/A _4900_/B VGND VPWR _4841_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_33_432 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_115 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_7560_ _6275_/Y _7434_/X _6240_/Y _7436_/X VGND VPWR _7560_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4772_ _4787_/A _6086_/B VGND VPWR _5583_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_7491_ _6855_/Y _7445_/X _6871_/Y _7447_/X VGND VPWR _7491_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_6511_ _9221_/Q VGND VPWR _8753_/A VGND VPWR sky130_fd_sc_hd__inv_6
XFILLER_9_160 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6442_ _6440_/Y _5526_/B _6441_/Y _5897_/B VGND VPWR _6442_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_9230_ _9440_/CLK _9230_/D _9685_/SET_B VGND VPWR _9230_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_173_164 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_9161_ _9532_/CLK _9161_/D _9528_/SET_B VGND VPWR _9161_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_161_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8112_ _8640_/B VGND VPWR _8390_/B VGND VPWR sky130_fd_sc_hd__inv_4
Xclkbuf_3_0_0_wb_clk_i clkbuf_3_1_0_wb_clk_i/A VGND VPWR _9203_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_2
X_6373_ _9216_/Q VGND VPWR _6373_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_114_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_231 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5324_ _9497_/Q _5319_/A _8929_/A1 _5319_/Y VGND VPWR _9497_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_9092_ _8837_/A1 _9092_/D _5980_/X VGND VPWR _9092_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_114_275 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5255_ _9544_/Q _5253_/A _5964_/B1 _5253_/Y VGND VPWR _9544_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8043_ _8097_/B _8552_/A _8042_/X VGND VPWR _8045_/A VGND VPWR sky130_fd_sc_hd__o21ai_1
X_5186_ _9588_/Q _5180_/A _8916_/A1 _5180_/Y VGND VPWR _9588_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_113_36 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_14 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8945_ _9083_/Q _9082_/Q _9051_/Q VGND VPWR _8945_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8876_ _7177_/Y _9634_/Q _8959_/S VGND VPWR _8876_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_83_398 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7827_ _8175_/A VGND VPWR _8476_/A VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_51_251 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7758_ _8660_/C VGND VPWR _8282_/C VGND VPWR sky130_fd_sc_hd__clkinv_2
X_7689_ _6409_/Y _7445_/X _6404_/Y _7447_/X VGND VPWR _7689_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_6709_ _6704_/Y _5355_/B _6705_/Y _5336_/B _6708_/X VGND VPWR _6716_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_11_159 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_120 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9428_ _9508_/CLK _9428_/D _9647_/SET_B VGND VPWR _9428_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_152_304 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_570 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_99 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9359_ _9493_/CLK _9359_/D _4628_/A VGND VPWR _9359_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_105_242 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_524 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_384 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_270 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_410 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_62 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_152 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_356 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_130 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_175 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_584 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_402 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5040_ _8973_/X _4551_/B _9679_/Q _5062_/D VGND VPWR _9679_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_26_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6991_ _9791_/Q VGND VPWR _6991_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_38_568 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_162 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_376 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8730_ _8730_/A _8730_/B _8730_/C _8730_/D VGND VPWR _8731_/B VGND VPWR sky130_fd_sc_hd__or4_2
X_5942_ _5942_/A VGND VPWR _5943_/A VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_21_413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_262 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8661_ _8660_/C _8341_/A _8660_/B _8660_/X _8556_/Y VGND VPWR _8661_/X VGND VPWR
+ sky130_fd_sc_hd__o311a_1
X_5873_ _5873_/A VGND VPWR _5874_/A VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_178_245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8592_ _8592_/A VGND VPWR _8641_/A VGND VPWR sky130_fd_sc_hd__inv_2
X_4824_ _6111_/A _4891_/A VGND VPWR _5100_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_7612_ _4712_/Y _7415_/X _4784_/Y _7417_/X _7611_/X VGND VPWR _7626_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_138_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7543_ _6337_/Y _7430_/X _6402_/Y _7432_/X _7542_/X VGND VPWR _7543_/X VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_4755_ _4787_/A _4931_/A VGND VPWR _4756_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_174_451 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7474_ _7476_/A _9251_/Q _7474_/C _7474_/D VGND VPWR _7475_/A VGND VPWR sky130_fd_sc_hd__or4_1
X_4686_ _4921_/A _4780_/B VGND VPWR _5810_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_9213_ _9758_/CLK _9213_/D _9779_/SET_B VGND VPWR _9213_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_146_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6425_ _6423_/Y _5450_/B _6424_/Y _5518_/B VGND VPWR _6425_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_6356_ _9290_/Q VGND VPWR _6356_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9144_ _9278_/CLK _9144_/D _9633_/SET_B VGND VPWR _9144_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_161_189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9075_ _9358_/CLK _9075_/D _9685_/SET_B VGND VPWR _9075_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_5307_ _5307_/A VGND VPWR _5308_/A VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_68_18 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6287_ _9343_/Q VGND VPWR _6287_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_130_554 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_8026_ _8097_/B _8130_/B _8023_/X _8407_/A _8454_/B VGND VPWR _8026_/X VGND VPWR
+ sky130_fd_sc_hd__o2111a_1
X_5238_ _9555_/Q _5234_/A _5966_/B1 _5234_/Y VGND VPWR _9555_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_5169_ _5169_/A VGND VPWR _5169_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_56_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8928_ _9615_/Q _8844_/X _8930_/S VGND VPWR _8928_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XPHY_224 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_202 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_8859_ _8858_/X _9168_/Q _9054_/Q VGND VPWR _8859_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_268 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_246 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_235 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_43 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_279 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_31 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_326 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_454 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_40 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_118 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_96 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_516 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_324 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_210 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_131 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4540_ _5966_/B1 _9760_/Q _4540_/S VGND VPWR _4541_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_128_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_4471_ _4471_/A VGND VPWR _4787_/A VGND VPWR sky130_fd_sc_hd__buf_8
XFILLER_171_443 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_134 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7190_ _8763_/A _7112_/X _7699_/A _7077_/B VGND VPWR _7190_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_6210_ _6205_/Y _5507_/B _6206_/Y _6086_/X _6209_/X VGND VPWR _6211_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_2
XFILLER_131_307 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6141_ _9327_/Q VGND VPWR _6141_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_85_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6072_ _9449_/Q VGND VPWR _6072_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_5023_ _9688_/Q _5015_/A _8916_/A1 _5015_/Y VGND VPWR _9688_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_81_611 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_471 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_9762_ _9770_/CLK _9762_/D _7011_/B VGND VPWR _9762_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_6974_ _6974_/A _6974_/B VGND VPWR _6975_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_8713_ _8713_/A _8713_/B _8713_/C _8713_/D VGND VPWR _8714_/B VGND VPWR sky130_fd_sc_hd__or4_1
X_5925_ _7768_/C _7768_/D _5925_/C input148/X VGND VPWR _5936_/A VGND VPWR sky130_fd_sc_hd__or4b_1
X_9693_ _9695_/CLK _9693_/D _9779_/SET_B VGND VPWR _9693_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_21_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_37 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_8644_ _8677_/D _8719_/C _8731_/A _8675_/D VGND VPWR _8647_/A VGND VPWR sky130_fd_sc_hd__or4_4
X_5856_ _5849_/X _8861_/X _8924_/X _9170_/Q VGND VPWR _9170_/D VGND VPWR sky130_fd_sc_hd__o22a_2
X_4807_ _4807_/A VGND VPWR _4808_/A VGND VPWR sky130_fd_sc_hd__buf_2
X_5787_ _5787_/A VGND VPWR _5787_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_8575_ _8575_/A _8575_/B _8575_/C VGND VPWR _8576_/D VGND VPWR sky130_fd_sc_hd__or3_1
X_7526_ _7703_/A _7425_/X _7523_/X _7525_/X VGND VPWR _7536_/C VGND VPWR sky130_fd_sc_hd__o211a_1
X_4738_ _4787_/A _4927_/A VGND VPWR _4739_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_21_298 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4669_ _4669_/A _4729_/D _8946_/X _8944_/X VGND VPWR _4927_/A VGND VPWR sky130_fd_sc_hd__or4_4
X_7457_ _7457_/A VGND VPWR _7457_/X VGND VPWR sky130_fd_sc_hd__buf_8
XFILLER_119_79 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6408_ _6408_/A _6408_/B _6408_/C _6408_/D VGND VPWR _6474_/A VGND VPWR sky130_fd_sc_hd__and4_1
X_7388_ _6361_/Y _7112_/X _6441_/Y _7077_/B VGND VPWR _7388_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_9127_ _9379_/CLK _9127_/D _9646_/SET_B VGND VPWR _9127_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_103_543 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6339_ _6334_/Y _5968_/B _6335_/Y _5488_/B _6338_/X VGND VPWR _6352_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9058_ _9058_/CLK _9058_/D _6041_/X VGND VPWR _9058_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_76_438 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_32 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8009_ _8009_/A _8060_/A VGND VPWR _8009_/X VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_151_66 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_276 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_362 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_140 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_600 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_176 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5710_ _7472_/A VGND VPWR _5710_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_176_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6690_ _6690_/A _6690_/B _6690_/C _6690_/D VGND VPWR _6691_/D VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_31_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5641_ _9277_/Q VGND VPWR _5647_/A VGND VPWR sky130_fd_sc_hd__inv_2
X_8360_ _8360_/A _8573_/C _8642_/C _8574_/C VGND VPWR _8364_/A VGND VPWR sky130_fd_sc_hd__or4_1
X_5572_ _6052_/A _5572_/B VGND VPWR _5573_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_144_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8291_ _8672_/C _8650_/B _8291_/C VGND VPWR _8292_/B VGND VPWR sky130_fd_sc_hd__or3_1
X_4523_ _6111_/A _6111_/B VGND VPWR _4524_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_7311_ _6927_/Y _7077_/C _6904_/Y _7077_/D _7310_/X VGND VPWR _7311_/X VGND VPWR
+ sky130_fd_sc_hd__o221a_1
Xclkbuf_1_0_1_csclk clkbuf_1_0_1_csclk/A VGND VPWR clkbuf_2_1_0_csclk/A VGND VPWR
+ sky130_fd_sc_hd__clkbuf_2
X_7242_ _7242_/A _7242_/B _7242_/C _7242_/D VGND VPWR _7243_/C VGND VPWR sky130_fd_sc_hd__and4_1
X_4454_ _6052_/A VGND VPWR _5960_/A VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_131_126 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7173_ _6763_/Y _5728_/X _6673_/Y _7040_/A _7172_/X VGND VPWR _7176_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_6124_ _6122_/Y _5757_/B _6123_/Y _5905_/B VGND VPWR _6124_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_6055_ _9047_/Q _6054_/A _8929_/A1 _6054_/Y VGND VPWR _9047_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_100_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_268 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5006_ _5006_/A VGND VPWR _5007_/S VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_93_290 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA_109 input77/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_121_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_463 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9745_ _9777_/CLK _9745_/D _9757_/SET_B VGND VPWR _9745_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6957_ _6629_/Y _6952_/A _9031_/Q _6952_/Y VGND VPWR _9031_/D VGND VPWR sky130_fd_sc_hd__o22a_1
X_5908_ _9132_/Q _5907_/A _8846_/X _5907_/Y VGND VPWR _9132_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_6888_ _6883_/Y _5829_/B _6884_/Y _5583_/B _6887_/X VGND VPWR _6901_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9676_ _9681_/CLK _9676_/D _6146_/A VGND VPWR _9676_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_139_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_78 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5839_ _5839_/A VGND VPWR _5839_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_8627_ _8627_/A _8627_/B _8627_/C _8627_/D VGND VPWR _8686_/D VGND VPWR sky130_fd_sc_hd__or4_2
X_8558_ _8558_/A VGND VPWR _8688_/B VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_147_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7509_ _6710_/Y _7445_/X _6767_/Y _7447_/X VGND VPWR _7509_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_135_443 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_8489_ _8720_/A _8713_/A _8703_/A VGND VPWR _8603_/A VGND VPWR sky130_fd_sc_hd__or3_1
XFILLER_1_478 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_52 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_379 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_360 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_95 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput308 _8823_/X VGND VPWR serial_data_2 VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput319 _9765_/Q VGND VPWR sram_ro_addr[3] VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_141_479 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_159 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_235 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_7860_ _8515_/B _8262_/B VGND VPWR _8667_/A VGND VPWR sky130_fd_sc_hd__nor2_1
X_6811_ _9722_/Q VGND VPWR _6811_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_50_102 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_7791_ _8189_/A _7791_/B VGND VPWR _7792_/B VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_23_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6742_ _9634_/Q VGND VPWR _6742_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9530_ _9532_/CLK _9530_/D _9647_/SET_B VGND VPWR _9530_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_9461_ _9789_/CLK _9461_/D _9647_/SET_B VGND VPWR _9461_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6673_ _9095_/Q VGND VPWR _6673_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_176_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_354 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5624_ _9293_/Q _5623_/A _8846_/X _5623_/Y VGND VPWR _9293_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8412_ _8550_/A _8401_/B _8409_/X _8411_/Y VGND VPWR _8412_/X VGND VPWR sky130_fd_sc_hd__o211a_1
X_9392_ _9483_/CLK _9392_/D _9528_/SET_B VGND VPWR _9392_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_31_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_8343_ _7886_/B _8003_/Y _8110_/C VGND VPWR _8343_/Y VGND VPWR sky130_fd_sc_hd__o21ai_2
XFILLER_117_443 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5555_ _9338_/Q _5547_/A _8839_/X _5547_/Y VGND VPWR _9338_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_191_379 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4506_ _4506_/A VGND VPWR _4506_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_5486_ _9386_/Q _5482_/A _5966_/B1 _5482_/Y VGND VPWR _9386_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8274_ _8510_/A _8660_/B _8496_/A VGND VPWR _8693_/B VGND VPWR sky130_fd_sc_hd__nor3_1
X_7225_ _6282_/Y _7040_/C _6304_/Y _7059_/C VGND VPWR _7225_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_7156_ _6713_/Y _7086_/X _6710_/Y _7088_/X VGND VPWR _7156_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_76_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6107_ _6105_/Y _5110_/B _6106_/Y _4822_/X VGND VPWR _6107_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_86_522 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7087_ _7127_/C _7087_/B VGND VPWR _7088_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_6038_ _9069_/Q _4466_/A _8929_/A1 _4466_/Y VGND VPWR _9069_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_132_46 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_22 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_260 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_7989_ _8098_/A _8386_/B VGND VPWR _8050_/B VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_81_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_88 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_9728_ _9769_/CLK _9728_/D _7011_/B VGND VPWR _9728_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_167_332 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_99 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_9659_ _4450_/A1 _9659_/D _6146_/A VGND VPWR _9659_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_10_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_37 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_216 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_622 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_17_csclk clkbuf_2_3_0_csclk/X VGND VPWR _9508_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_60_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_364 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5340_ _9487_/Q _5338_/A _5964_/B1 _5338_/Y VGND VPWR _9487_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_99_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5271_ _9534_/Q _5269_/A _8845_/X _5269_/Y VGND VPWR _9534_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_99_157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_608 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7010_ _9626_/Q _7011_/B VGND VPWR _7010_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_68_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8961_ _7737_/X _8961_/A1 _8975_/S VGND VPWR _8961_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_7912_ _8238_/A _7864_/X _7909_/X _7910_/X _8454_/A VGND VPWR _7912_/X VGND VPWR
+ sky130_fd_sc_hd__o2111a_1
XFILLER_48_290 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_8892_ _7353_/Y _9629_/Q _8959_/S VGND VPWR _8892_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_63_260 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7843_ _8515_/B _7848_/A VGND VPWR _7931_/A VGND VPWR sky130_fd_sc_hd__or2_2
XFILLER_23_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_455 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7774_ _7959_/A _8583_/A _7774_/C _7774_/D VGND VPWR _7775_/D VGND VPWR sky130_fd_sc_hd__nand4bb_1
X_4986_ _4994_/A VGND VPWR _4987_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_149_310 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9513_ _9514_/CLK _9513_/D _4628_/A VGND VPWR _9513_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6725_ _9556_/Q VGND VPWR _6725_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_6656_ _9764_/Q VGND VPWR _6656_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9444_ _9785_/CLK _9444_/D _9779_/SET_B VGND VPWR _9444_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6587_ _9388_/Q VGND VPWR _6587_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_5607_ _9304_/Q _5604_/A _5965_/B1 _5604_/Y VGND VPWR _9304_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_9375_ _9379_/CLK _9375_/D _9779_/SET_B VGND VPWR _9375_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_11_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5538_ _9352_/Q _5536_/A _8845_/X _5536_/Y VGND VPWR _9352_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8326_ _8468_/A _8715_/B VGND VPWR _8693_/C VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_145_582 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_8257_ _8257_/A _8674_/B VGND VPWR _8259_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_7208_ _6356_/Y _7059_/B _6392_/Y _7068_/C _7207_/X VGND VPWR _7211_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_5469_ _5545_/A _6081_/B VGND VPWR _5470_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_132_276 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_511 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_8188_ _8305_/A _8188_/B VGND VPWR _8606_/B VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_59_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7139_ _6854_/Y _7097_/X _6832_/Y _7099_/X VGND VPWR _7139_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_100_162 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_430 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_75 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xinput18 mask_rev_in[22] VGND VPWR _6208_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_155_324 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput29 mask_rev_in[3] VGND VPWR _6618_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_155_368 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_319 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_298 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_514 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_219 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_444 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4840_ _4840_/A VGND VPWR _4840_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_21_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4771_ _9312_/Q VGND VPWR _4771_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_6510_ _9267_/Q VGND VPWR _6510_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_146_302 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7490_ _6919_/Y _7425_/X _7487_/X _7489_/X VGND VPWR _7500_/C VGND VPWR sky130_fd_sc_hd__o211a_1
XFILLER_146_324 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6441_ _9137_/Q VGND VPWR _6441_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_173_154 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_9160_ _9358_/CLK _9160_/D _9528_/SET_B VGND VPWR _9160_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6372_ _9222_/Q VGND VPWR _6372_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_161_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5323_ _9498_/Q _5319_/A _8925_/A1 _5319_/Y VGND VPWR _9498_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8111_ _8378_/B VGND VPWR _8544_/B VGND VPWR sky130_fd_sc_hd__clkinv_4
XFILLER_114_243 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9091_ _8837_/A1 _9091_/D _5984_/X VGND VPWR _9091_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_142_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5254_ _9545_/Q _5253_/A _5963_/B1 _5253_/Y VGND VPWR _9545_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8042_ _8389_/A _8552_/A _8041_/Y VGND VPWR _8042_/X VGND VPWR sky130_fd_sc_hd__o21a_1
X_5185_ _9589_/Q _5180_/A _8840_/X _5180_/Y VGND VPWR _9589_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_110_460 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_374 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_344 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_558 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_48 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_8944_ _8943_/X _9675_/Q _9587_/Q VGND VPWR _8944_/X VGND VPWR sky130_fd_sc_hd__mux2_4
XFILLER_83_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8875_ _8874_/X _9138_/Q _9054_/Q VGND VPWR _8875_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_7826_ _8515_/A _8272_/A VGND VPWR _8175_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_24_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_438 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7757_ _7757_/A VGND VPWR _8660_/C VGND VPWR sky130_fd_sc_hd__buf_4
X_4969_ _4969_/A VGND VPWR _4969_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_6708_ _6706_/Y _4870_/X _6707_/Y _5602_/B VGND VPWR _6708_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_7688_ _6458_/Y _7425_/X _7685_/X _7687_/X VGND VPWR _7698_/C VGND VPWR sky130_fd_sc_hd__o211a_1
X_9427_ _9527_/CLK _9427_/D _9528_/SET_B VGND VPWR _9427_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6639_ _9220_/Q VGND VPWR _6639_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_138_56 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_49 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_582 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_9358_ _9358_/CLK _9358_/D _9685_/SET_B VGND VPWR _9358_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_105_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_8309_ _7864_/X _8498_/A _8341_/B _8498_/B VGND VPWR _8309_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_9289_ _9596_/CLK _9289_/D _9528_/SET_B VGND VPWR _9289_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_3_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_254 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_30 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_466 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_74 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_187 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_360 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_202 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_414 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6990_ _9709_/Q _6023_/Y _4953_/Y _9049_/Q VGND VPWR _9049_/D VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_65_388 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5941_ _5960_/A _5941_/B VGND VPWR _5942_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_92_174 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8660_ _8660_/A _8660_/B _8660_/C VGND VPWR _8660_/X VGND VPWR sky130_fd_sc_hd__or3_1
X_5872_ _6052_/A _5872_/B VGND VPWR _5873_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_4823_ _9641_/Q VGND VPWR _4823_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7611_ _4677_/Y _7419_/X _4809_/Y _7421_/X VGND VPWR _7611_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_8591_ _8510_/A _8498_/A _7879_/B _8397_/A VGND VPWR _8591_/Y VGND VPWR sky130_fd_sc_hd__o211ai_1
XFILLER_21_425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4754_ _4754_/A VGND VPWR _4754_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7542_ _6346_/Y _7434_/X _6329_/Y _7436_/X VGND VPWR _7542_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_146_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7473_ _7473_/A VGND VPWR _7473_/X VGND VPWR sky130_fd_sc_hd__buf_8
XFILLER_174_463 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4685_ _9198_/Q VGND VPWR _4685_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9212_ _9655_/CLK _9212_/D _9779_/SET_B VGND VPWR _9212_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_161_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6424_ _9363_/Q VGND VPWR _6424_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_6355_ _6354_/Y _5121_/B _4844_/X _6158_/X VGND VPWR _6355_/X VGND VPWR sky130_fd_sc_hd__o211a_1
X_9143_ _9203_/CLK _9143_/D _9633_/SET_B VGND VPWR _9143_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6286_ _6281_/Y _6165_/A _6282_/Y _5045_/B _6285_/X VGND VPWR _6307_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9074_ _9687_/CLK _9074_/D _9685_/SET_B VGND VPWR _9074_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_5306_ _5545_/A _5306_/B VGND VPWR _5307_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_0_329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5237_ _9556_/Q _5234_/A _5965_/B1 _5234_/Y VGND VPWR _9556_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8025_ _8624_/B _8137_/B VGND VPWR _8454_/B VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_68_182 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5168_ _5168_/A VGND VPWR _5169_/A VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_44_506 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5099_ _9646_/Q _5091_/A _8916_/A1 _5091_/Y VGND VPWR _9646_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_56_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8927_ _9616_/Q _8845_/X _8930_/S VGND VPWR _8927_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_71_347 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_68 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_214 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_203 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_8858_ _7572_/Y _9637_/Q _8978_/S VGND VPWR _8858_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XPHY_258 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_247 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_236 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_7809_ _7903_/C _8528_/A _8525_/A _8189_/A VGND VPWR _7878_/A VGND VPWR sky130_fd_sc_hd__or4_1
X_8789_ _8789_/A VGND VPWR _8790_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XPHY_269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_132 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_52 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_528 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_580 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_222 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_463 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4470_ _8936_/X _4665_/B _4801_/C VGND VPWR _4471_/A VGND VPWR sky130_fd_sc_hd__or3_1
XFILLER_143_146 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6140_ _9197_/Q VGND VPWR _6140_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_97_211 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6071_ _6071_/A _6071_/B VGND VPWR _6071_/Y VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_66_620 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5022_ _9689_/Q _5015_/A _8930_/A1 _5015_/Y VGND VPWR _9689_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_65_130 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6973_ _9061_/Q VGND VPWR _6974_/A VGND VPWR sky130_fd_sc_hd__inv_2
X_9761_ _9770_/CLK _9761_/D _7011_/B VGND VPWR _9761_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
XFILLER_53_325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5924_ _9065_/D VGND VPWR _6147_/B VGND VPWR sky130_fd_sc_hd__inv_2
X_8712_ _8738_/A _8712_/B VGND VPWR _8712_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
X_9692_ _9695_/CLK _9692_/D _9779_/SET_B VGND VPWR _9692_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_8643_ _7987_/Y _8390_/B _8317_/B _8364_/D _8576_/D VGND VPWR _8675_/D VGND VPWR
+ sky130_fd_sc_hd__a2111o_2
X_5855_ _5849_/X _8863_/X _8924_/X _9171_/Q VGND VPWR _9171_/D VGND VPWR sky130_fd_sc_hd__o22a_2
X_4806_ _9770_/Q _9708_/Q _9626_/Q VGND VPWR _4807_/A VGND VPWR sky130_fd_sc_hd__or3_1
XFILLER_119_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_8574_ _8574_/A _8574_/B _8574_/C VGND VPWR _8730_/D VGND VPWR sky130_fd_sc_hd__or3_1
X_5786_ _9218_/Q _5778_/A _8916_/A1 _5778_/Y VGND VPWR _9218_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7525_ _7701_/A _7430_/X _8785_/A _7432_/X _7524_/X VGND VPWR _7525_/X VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_4737_ _4737_/A VGND VPWR _4737_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_4668_ _9151_/Q VGND VPWR _4668_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7456_ _7456_/A _7466_/A _9255_/Q VGND VPWR _7457_/A VGND VPWR sky130_fd_sc_hd__or3_1
XFILLER_162_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6407_ _6402_/Y _5240_/B _6403_/Y _4491_/B _6406_/X VGND VPWR _6408_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_4599_ _9733_/Q _4592_/A _5966_/B1 _4592_/Y VGND VPWR _9733_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_9126_ _9129_/CLK _9126_/D _9779_/SET_B VGND VPWR _9126_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_7387_ _7387_/A _7387_/B _7387_/C _7387_/D VGND VPWR _7397_/B VGND VPWR sky130_fd_sc_hd__and4_1
X_6338_ _6336_/Y _4893_/X _6337_/Y _5905_/B VGND VPWR _6338_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_103_555 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9057_ _9280_/CLK _9057_/D _9757_/SET_B VGND VPWR _9057_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6269_ _9403_/Q VGND VPWR _6269_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
X_8008_ _8218_/A _8218_/B _8008_/C VGND VPWR _8060_/A VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_69_491 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_3_0_csclk clkbuf_2_3_0_csclk/A VGND VPWR clkbuf_2_3_0_csclk/X VGND VPWR
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_56_130 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_99 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_308 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_78 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_575 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_496 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_91 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_374 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_119 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_288 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_7 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_612 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5640_ _9279_/Q VGND VPWR _5649_/B VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_31_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5571_ _9328_/Q _5566_/A _5967_/B1 _5566_/Y VGND VPWR _9328_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_184_580 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7310_ _6873_/Y _7086_/X _6867_/Y _7088_/X VGND VPWR _7310_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4522_ _8946_/X _4729_/B _8934_/X _4729_/D VGND VPWR _6111_/B VGND VPWR sky130_fd_sc_hd__or4_4
X_8290_ _8606_/B _8290_/B VGND VPWR _8291_/C VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_156_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7241_ _6269_/Y _7124_/X _6311_/Y _7068_/B _7240_/X VGND VPWR _7242_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_4453_ _5133_/A VGND VPWR _6052_/A VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_7_270 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_138 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7172_ _7172_/A _7392_/B VGND VPWR _7172_/X VGND VPWR sky130_fd_sc_hd__or2_1
X_6123_ _9132_/Q VGND VPWR _6123_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_6054_ _6054_/A VGND VPWR _6054_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_105_38 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5005_ _9091_/Q _6022_/C _9092_/Q _6022_/B VGND VPWR _5006_/A VGND VPWR sky130_fd_sc_hd__or4_1
XFILLER_54_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_155 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_475 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6956_ _6475_/Y _6952_/A _9032_/Q _6952_/Y VGND VPWR _9032_/D VGND VPWR sky130_fd_sc_hd__o22a_2
X_9744_ _9777_/CLK _9744_/D _9757_/SET_B VGND VPWR _9744_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_5907_ _5907_/A VGND VPWR _5907_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_22_542 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_374 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_514 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6887_ _6885_/Y _5564_/B _6886_/Y _6052_/C VGND VPWR _6887_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_9675_ _9681_/CLK _9675_/D _6146_/A VGND VPWR _9675_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_14_68 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8626_ _8401_/A _8624_/X _8117_/A _8625_/Y VGND VPWR _8629_/B VGND VPWR sky130_fd_sc_hd__o22ai_2
X_5838_ _5838_/A VGND VPWR _5839_/A VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_139_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_8557_ _8386_/A _7971_/A _8389_/A _7829_/A _8556_/Y VGND VPWR _8558_/A VGND VPWR
+ sky130_fd_sc_hd__o311a_1
X_5769_ _5769_/A VGND VPWR _5770_/A VGND VPWR sky130_fd_sc_hd__clkbuf_2
X_7508_ _6775_/Y _7425_/X _7505_/X _7507_/X VGND VPWR _7518_/C VGND VPWR sky130_fd_sc_hd__o211a_1
XFILLER_147_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8488_ _8488_/A VGND VPWR _8488_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_7439_ _4687_/Y _7425_/X _7428_/X _7438_/X VGND VPWR _7481_/C VGND VPWR sky130_fd_sc_hd__o211a_1
XFILLER_135_499 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_116 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_531 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_436 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9109_ _9379_/CLK _9109_/D _9779_/SET_B VGND VPWR _9109_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_29_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_92 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_568 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xoutput309 _8820_/X VGND VPWR serial_load VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_96_71 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_160 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6810_ _6805_/Y _5232_/B _6806_/Y _4841_/X _6809_/X VGND VPWR _6829_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_7790_ _8528_/B _7900_/A VGND VPWR _8538_/C VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_50_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6741_ _6741_/A _6741_/B _6741_/C _6741_/D VGND VPWR _6784_/B VGND VPWR sky130_fd_sc_hd__and4_1
X_9460_ _9532_/CLK _9460_/D _9647_/SET_B VGND VPWR _9460_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6672_ _6667_/Y _5045_/B _6668_/Y _5488_/B _6671_/X VGND VPWR _6690_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_5623_ _5623_/A VGND VPWR _5623_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9391_ _9483_/CLK _9391_/D _9528_/SET_B VGND VPWR _9391_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_8411_ _8734_/B _8574_/A VGND VPWR _8411_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_117_411 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8342_ _8114_/Y _8115_/Y _8594_/B VGND VPWR _8356_/A VGND VPWR sky130_fd_sc_hd__a21o_1
XFILLER_129_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5554_ _9339_/Q _5547_/A _8930_/A1 _5547_/Y VGND VPWR _9339_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_105_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5485_ _9387_/Q _5482_/A _5965_/B1 _5482_/Y VGND VPWR _9387_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8273_ _8273_/A _8715_/B VGND VPWR _8275_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_4505_ _4505_/A VGND VPWR _4506_/A VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_116_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7224_ _6244_/Y _7082_/X _6256_/Y _7084_/X _7223_/X VGND VPWR _7243_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_7155_ _7155_/A _7155_/B _7155_/C VGND VPWR _7155_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
X_6106_ _6106_/A VGND VPWR _6106_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_58_247 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_171 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7086_ _7086_/A VGND VPWR _7086_/X VGND VPWR sky130_fd_sc_hd__buf_8
XFILLER_86_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6037_ _9070_/Q _6029_/A _8839_/X _6029_/Y VGND VPWR _9070_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_132_58 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_12 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_7 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_250 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_23 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7988_ _7988_/A _8091_/B VGND VPWR _8386_/B VGND VPWR sky130_fd_sc_hd__or2b_2
XPHY_89 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_9727_ _9769_/CLK _9727_/D _7011_/B VGND VPWR _9727_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6939_ _9232_/Q VGND VPWR _6939_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_25_89 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9658_ _9779_/CLK _9658_/D _9779_/SET_B VGND VPWR _9658_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_8609_ _8609_/A VGND VPWR _8666_/C VGND VPWR sky130_fd_sc_hd__inv_2
X_9589_ _9617_/CLK _9589_/D _9295_/SET_B VGND VPWR _9589_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_10_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_0_csclk _8847_/X VGND VPWR clkbuf_0_csclk/X VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_123_436 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_210 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_274 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_49 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_0_0_csclk clkbuf_0_csclk/X VGND VPWR clkbuf_1_0_1_csclk/A VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_66_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_376 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_6 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_230 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5270_ _9535_/Q _5269_/A _8846_/X _5269_/Y VGND VPWR _9535_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_141_266 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_331 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8960_ _7735_/X _5060_/X _8960_/S VGND VPWR _8960_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_7911_ _8521_/B _8239_/B VGND VPWR _8454_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_8891_ _8890_/X _9146_/Q _9054_/Q VGND VPWR _8891_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_7842_ _8660_/B _8496_/A VGND VPWR _7848_/A VGND VPWR sky130_fd_sc_hd__or2_2
XFILLER_23_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4985_ _9701_/Q _4966_/A _4949_/A _4966_/Y VGND VPWR _9701_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7773_ _8525_/A VGND VPWR _8583_/A VGND VPWR sky130_fd_sc_hd__inv_6
XFILLER_51_467 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9512_ _9514_/CLK _9512_/D _4628_/A VGND VPWR _9512_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6724_ _9374_/Q VGND VPWR _6724_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_9443_ _9791_/CLK _9443_/D _9779_/SET_B VGND VPWR _9443_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_192_612 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6655_ _6650_/Y _6027_/B _6651_/Y _4602_/B _6654_/X VGND VPWR _6691_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_5606_ _9305_/Q _5604_/A _5964_/B1 _5604_/Y VGND VPWR _9305_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_6586_ _6586_/A _6586_/B _6586_/C VGND VPWR _6628_/B VGND VPWR sky130_fd_sc_hd__and3_1
X_9374_ _9379_/CLK _9374_/D _9646_/SET_B VGND VPWR _9374_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_8325_ _8325_/A VGND VPWR _8468_/A VGND VPWR sky130_fd_sc_hd__inv_2
X_5537_ _9353_/Q _5536_/A _8846_/X _5536_/Y VGND VPWR _9353_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_117_274 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8256_ _8260_/A _8264_/B VGND VPWR _8674_/B VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_11_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5468_ _9398_/Q _5460_/A _5967_/B1 _5460_/Y VGND VPWR _9398_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7207_ _6428_/Y _7079_/B _6377_/Y _7059_/A VGND VPWR _7207_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_59_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_8187_ _8187_/A VGND VPWR _8650_/B VGND VPWR sky130_fd_sc_hd__inv_2
X_5399_ _9446_/Q _5395_/A _5963_/B1 _5395_/Y VGND VPWR _9446_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_59_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7138_ _6933_/Y _7048_/B _6921_/Y _7077_/A _7137_/X VGND VPWR _7145_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_100_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7069_ _7073_/C _7085_/B VGND VPWR _7070_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_100_174 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_442 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xinput19 mask_rev_in[23] VGND VPWR _6093_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_136_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_42 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_288 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_526 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_50 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4770_ _4805_/A _4843_/B VGND VPWR _5089_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_158_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6440_ _9358_/Q VGND VPWR _6440_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_127_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_358 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6371_ _9260_/Q VGND VPWR _6371_/Y VGND VPWR sky130_fd_sc_hd__inv_4
X_5322_ _9499_/Q _5319_/A _8844_/X _5319_/Y VGND VPWR _9499_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8110_ _8625_/A _8282_/B _8110_/C VGND VPWR _8708_/B VGND VPWR sky130_fd_sc_hd__and3_2
X_9090_ _9709_/CLK _9090_/D _5988_/X VGND VPWR _9090_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_5253_ _5253_/A VGND VPWR _5253_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_8041_ _8041_/A _8685_/A VGND VPWR _8041_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_87_128 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5184_ _9590_/Q _5180_/A _8841_/X _5180_/Y VGND VPWR _9590_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_83_301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_356 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8943_ _9082_/Q _4949_/A _9051_/Q VGND VPWR _8943_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_83_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_8874_ _7155_/Y _9633_/Q _8959_/S VGND VPWR _8874_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_7825_ _7825_/A VGND VPWR _8515_/A VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_184_409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7756_ _7832_/A _7756_/B _7837_/C VGND VPWR _7757_/A VGND VPWR sky130_fd_sc_hd__or3_1
X_4968_ _4994_/A VGND VPWR _4969_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_137_303 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6707_ _9304_/Q VGND VPWR _6707_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7687_ _6331_/Y _7430_/X _6412_/Y _7432_/X _7686_/X VGND VPWR _7687_/X VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_4899_ _9437_/Q VGND VPWR _4899_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_9426_ _9527_/CLK _9426_/D _9528_/SET_B VGND VPWR _9426_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6638_ _9228_/Q VGND VPWR _6638_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_138_46 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_155 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9357_ _9358_/CLK _9357_/D _9685_/SET_B VGND VPWR _9357_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6569_ _9735_/Q VGND VPWR _6569_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_8308_ _7836_/A _8299_/A _7836_/B _7879_/Y VGND VPWR _8497_/A VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_133_531 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9288_ _9483_/CLK _9288_/D _9528_/SET_B VGND VPWR _9288_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_16_csclk clkbuf_2_3_0_csclk/X VGND VPWR _9344_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_154_23 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_266 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8239_ _8341_/A _8239_/B VGND VPWR _8361_/B VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_59_320 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_42 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_31 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_478 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_472 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_604 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_199 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_176 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_372 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_426 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_214 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_504 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5940_ _9059_/Q _7731_/A _9119_/Q _5938_/Y _5939_/X VGND VPWR _9119_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_92_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5871_ _9159_/Q _5866_/A _8839_/X _5866_/Y VGND VPWR _9159_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7610_ _4920_/Y _7400_/X _4731_/A _7405_/X _7609_/X VGND VPWR _7626_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_33_275 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4822_ _6158_/A _4929_/A VGND VPWR _4822_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_8590_ _8605_/B _8543_/Y _8564_/X _8589_/X VGND VPWR _8590_/Y VGND VPWR sky130_fd_sc_hd__o211ai_1
XFILLER_147_612 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_303 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4753_ _9789_/Q VGND VPWR _4753_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7541_ _6422_/Y _7427_/X _6360_/Y _5699_/X VGND VPWR _7541_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_7472_ _7472_/A _7476_/C _9255_/Q VGND VPWR _7473_/A VGND VPWR sky130_fd_sc_hd__or3_1
X_4684_ _4675_/Y _5507_/B _4677_/Y _5080_/B _4683_/X VGND VPWR _4705_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9211_ _9613_/CLK _9211_/D _9646_/SET_B VGND VPWR _9211_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6423_ _9410_/Q VGND VPWR _6423_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_146_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_103 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6354_ _9631_/Q VGND VPWR _6354_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9142_ _9278_/CLK _9142_/D _9757_/SET_B VGND VPWR _9142_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_5305_ _9510_/Q _5300_/A _5967_/B1 _5300_/Y VGND VPWR _9510_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_6285_ _7238_/A _5610_/B _6284_/Y _5837_/B VGND VPWR _6285_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_9073_ _9687_/CLK _9073_/D _9685_/SET_B VGND VPWR _9073_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_88_437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5236_ _9557_/Q _5234_/A _5964_/B1 _5234_/Y VGND VPWR _9557_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8024_ _8521_/A _8137_/B VGND VPWR _8407_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_88_459 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5167_ _5545_/A _6322_/A VGND VPWR _5168_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_5098_ _9647_/Q _5091_/A _8930_/A1 _5091_/Y VGND VPWR _9647_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_56_334 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_518 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8926_ _9605_/Q _8842_/X _8926_/S VGND VPWR _8926_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_17_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_215 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_204 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_359 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8857_ _8856_/X _9167_/Q _9054_/Q VGND VPWR _8857_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XPHY_259 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_248 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_226 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_23 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8788_ _8788_/A VGND VPWR _8788_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_7808_ _8660_/C _8119_/A VGND VPWR _8587_/A VGND VPWR sky130_fd_sc_hd__nor2_2
X_7739_ _9068_/Q _7739_/A2 _9067_/Q _7739_/B2 _7738_/X VGND VPWR _7739_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_137_144 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9409_ _9493_/CLK _9409_/D _4628_/A VGND VPWR _9409_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_4_603 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_467 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_99 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_512 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_356 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_131 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_80 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_7 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_234 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_71 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_158 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_180 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_267 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_556 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6070_ _6065_/Y _5837_/B _6066_/Y _5660_/B _6069_/X VGND VPWR _6071_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_66_610 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5021_ _9690_/Q _5015_/A _8955_/A1 _5015_/Y VGND VPWR _9690_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_93_440 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_142 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_9760_ _9770_/CLK _9760_/D _7011_/B VGND VPWR _9760_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_53_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6972_ _4936_/Y _6964_/A _9020_/Q _6964_/Y VGND VPWR _9020_/D VGND VPWR sky130_fd_sc_hd__o22a_1
X_8711_ _8117_/A _8624_/X _8117_/B _8625_/Y _8710_/Y VGND VPWR _8712_/B VGND VPWR
+ sky130_fd_sc_hd__o221ai_4
X_5923_ _9120_/Q _5918_/A _5967_/B1 _5918_/Y VGND VPWR _9120_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_9691_ _9695_/CLK _9691_/D _9779_/SET_B VGND VPWR _9691_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_34_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5854_ _5849_/X _8865_/X _8924_/X _9172_/Q VGND VPWR _9172_/D VGND VPWR sky130_fd_sc_hd__o22a_2
X_8642_ _8642_/A _8642_/B _8642_/C _8642_/D VGND VPWR _8731_/A VGND VPWR sky130_fd_sc_hd__or4_2
X_8573_ _8573_/A _8573_/B _8573_/C VGND VPWR _8642_/D VGND VPWR sky130_fd_sc_hd__or3_1
X_4805_ _4805_/A _4931_/B VGND VPWR _5534_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_7524_ _8779_/A _7434_/X _8777_/A _7436_/X VGND VPWR _7524_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_5785_ _9219_/Q _5778_/A _8930_/A1 _5778_/Y VGND VPWR _9219_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_9_91 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4736_ _4732_/Y _5621_/B _4734_/Y _5797_/B VGND VPWR _4736_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_162_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4667_ _4898_/A _4843_/B VGND VPWR _5905_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_7455_ _7455_/A VGND VPWR _7455_/X VGND VPWR sky130_fd_sc_hd__buf_8
XFILLER_162_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6406_ _6404_/Y _5480_/B _6405_/Y _4577_/B VGND VPWR _6406_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_7386_ _6369_/Y _7048_/D _6445_/Y _7040_/B _7385_/X VGND VPWR _7387_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_115_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4598_ _9734_/Q _4592_/A _5965_/B1 _4592_/Y VGND VPWR _9734_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_9125_ _9379_/CLK _9125_/D _9646_/SET_B VGND VPWR _9125_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6337_ _9129_/Q VGND VPWR _6337_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_88_223 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_9056_ _9203_/CLK _9056_/D _9633_/SET_B VGND VPWR _9056_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_6268_ _9767_/Q VGND VPWR _6268_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_28_12 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6199_ _9552_/Q VGND VPWR _6199_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_8007_ _8003_/Y _8566_/B _8064_/C VGND VPWR _8016_/A VGND VPWR sky130_fd_sc_hd__o21a_1
X_5219_ _9568_/Q _5218_/Y _8917_/X _5218_/A VGND VPWR _9568_/D VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_29_312 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8909_ _7730_/Y _9699_/Q _9048_/Q VGND VPWR _8909_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_40_565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_238 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_98 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_350 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_320 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_212 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_386 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_164 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_326 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_443 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_134 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_206 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_548 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5570_ _9329_/Q _5566_/A _5966_/B1 _5566_/Y VGND VPWR _9329_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_144_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4521_ _4521_/A VGND VPWR _9770_/D VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_171_220 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7240_ _6291_/Y _7126_/X _6241_/Y _7128_/X VGND VPWR _7240_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4452_ _8939_/X VGND VPWR _5133_/A VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_144_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7171_ _6775_/Y _7059_/D _6724_/Y _7116_/X _7170_/X VGND VPWR _7176_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_124_180 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6122_ _9238_/Q VGND VPWR _6122_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_6053_ _6053_/A VGND VPWR _6054_/A VGND VPWR sky130_fd_sc_hd__clkbuf_2
X_5004_ _5004_/A VGND VPWR _5004_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_38_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9743_ _9777_/CLK _9743_/D _9757_/SET_B VGND VPWR _9743_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6955_ _6326_/Y _6952_/A _9033_/Q _6952_/Y VGND VPWR _9033_/D VGND VPWR sky130_fd_sc_hd__o22a_1
X_9674_ _9674_/CLK _9674_/D _9633_/SET_B VGND VPWR _9674_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_5906_ _5906_/A VGND VPWR _5907_/A VGND VPWR sky130_fd_sc_hd__clkbuf_4
X_6886_ _9045_/Q VGND VPWR _6886_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_8625_ _8625_/A _8625_/B VGND VPWR _8625_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_167_526 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5837_ _6052_/A _5837_/B VGND VPWR _5838_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_8556_ _8601_/D VGND VPWR _8556_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_5768_ _5960_/A _5768_/B VGND VPWR _5769_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_4719_ _4903_/B _4780_/B VGND VPWR _5594_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_7507_ _6754_/Y _7430_/X _6761_/Y _7432_/X _7506_/X VGND VPWR _7507_/X VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_8487_ _8487_/A _8486_/X VGND VPWR _8488_/A VGND VPWR sky130_fd_sc_hd__or2b_1
X_7438_ _4664_/Y _7430_/X _4793_/Y _7432_/X _7437_/X VGND VPWR _7438_/X VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_5699_ _5699_/A VGND VPWR _5699_/X VGND VPWR sky130_fd_sc_hd__buf_8
XFILLER_162_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_456 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_584 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_79 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_128 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_426 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7369_ _6516_/Y _7059_/D _6555_/Y _7116_/X _7368_/X VGND VPWR _7374_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_89_543 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_9108_ _9379_/CLK _9108_/D _9779_/SET_B VGND VPWR _9108_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_130_150 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9039_ _9039_/CLK _9039_/D VGND VPWR _9039_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_183_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_89 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_42 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_75 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_106 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_491 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_410 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6740_ _6735_/Y _5278_/B _6736_/Y _5344_/B _6739_/X VGND VPWR _6741_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_50_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6671_ _6669_/Y _4832_/X _6670_/Y _4590_/B VGND VPWR _6671_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_8410_ _8410_/A VGND VPWR _8734_/B VGND VPWR sky130_fd_sc_hd__inv_2
X_9390_ _9483_/CLK _9390_/D _9528_/SET_B VGND VPWR _9390_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_5622_ _5622_/A VGND VPWR _5623_/A VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_136_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5553_ _9340_/Q _5547_/A _8841_/X _5547_/Y VGND VPWR _9340_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8341_ _8341_/A _8341_/B _8496_/A VGND VPWR _8594_/B VGND VPWR sky130_fd_sc_hd__nor3_1
XFILLER_117_423 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4504_ _5259_/A _4504_/B VGND VPWR _4505_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_144_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_456 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5484_ _9388_/Q _5482_/A _5964_/B1 _5482_/Y VGND VPWR _9388_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8272_ _8272_/A _8660_/B _8496_/A VGND VPWR _8715_/B VGND VPWR sky130_fd_sc_hd__nor3_1
X_7223_ _6309_/Y _7077_/C _6287_/Y _7077_/D _7222_/X VGND VPWR _7223_/X VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_7154_ _7154_/A _7154_/B _7154_/C _7154_/D VGND VPWR _7155_/C VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_100_301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6105_ _9639_/Q VGND VPWR _6105_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_112_183 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7085_ _7127_/C _7085_/B VGND VPWR _7086_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_100_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6036_ _9071_/Q _6029_/A _8840_/X _6029_/Y VGND VPWR _9071_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_54_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_13 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_35 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7987_ _8551_/A VGND VPWR _7987_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XPHY_79 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_9726_ _9769_/CLK _9726_/D _7011_/B VGND VPWR _9726_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_6938_ _9308_/Q VGND VPWR _6938_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_6869_ _6867_/Y _5442_/B _6868_/Y _5251_/B VGND VPWR _6869_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_9657_ _9779_/CLK _9657_/D _9779_/SET_B VGND VPWR _9657_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_22_384 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_8608_ _8496_/A _8515_/B _8305_/B _8019_/C _8447_/X VGND VPWR _8609_/A VGND VPWR
+ sky130_fd_sc_hd__o311a_1
X_9588_ _9601_/CLK _9588_/D _9295_/SET_B VGND VPWR _9588_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_8539_ _8539_/A _8721_/C _8538_/X VGND VPWR _8705_/D VGND VPWR sky130_fd_sc_hd__or3b_2
XFILLER_182_326 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_359 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_546 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_590 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_123 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_92 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_96 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_388 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_6 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_242 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_8890_ _7331_/Y _9628_/Q _8959_/S VGND VPWR _8890_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_7910_ _8515_/B _8239_/B VGND VPWR _7910_/X VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_36_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7841_ _7841_/A VGND VPWR _8515_/B VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_102_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7772_ _7903_/C VGND VPWR _7959_/A VGND VPWR sky130_fd_sc_hd__inv_2
X_4984_ _4984_/A VGND VPWR _4984_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_6723_ _9439_/Q VGND VPWR _6723_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9511_ _9514_/CLK _9511_/D _4628_/A VGND VPWR _9511_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_176_131 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6654_ _6652_/Y _4504_/B _6653_/Y _5178_/B VGND VPWR _6654_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_9442_ _9791_/CLK _9442_/D _9633_/SET_B VGND VPWR _9442_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_164_304 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5605_ _9306_/Q _5604_/A _8843_/X _5604_/Y VGND VPWR _9306_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_191_134 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9373_ _9379_/CLK _9373_/D _9779_/SET_B VGND VPWR _9373_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6585_ _8745_/A _5013_/B _6581_/Y _5789_/B _6584_/X VGND VPWR _6586_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_5536_ _5536_/A VGND VPWR _5536_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_8324_ _8324_/A _8498_/B VGND VPWR _8506_/C VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_127_26 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_426 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5467_ _9399_/Q _5460_/A _5966_/B1 _5460_/Y VGND VPWR _9399_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8255_ _8255_/A _8493_/B VGND VPWR _8257_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_7206_ _6396_/Y _7095_/X _6368_/Y _7068_/D _7205_/X VGND VPWR _7211_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_5398_ _9447_/Q _5395_/A _8844_/X _5395_/Y VGND VPWR _9447_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8186_ _8186_/A VGND VPWR _8672_/C VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_98_192 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_492 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7137_ _6910_/Y _7040_/C _6799_/Y _7059_/C VGND VPWR _7137_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_59_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_131 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7068_ _7068_/A _7068_/B _7068_/C _7068_/D VGND VPWR _7078_/C VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_86_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_186 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6019_ _6019_/A VGND VPWR _9081_/D VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_100_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_498 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_148 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_9709_ _9709_/CLK _9709_/D _4948_/X VGND VPWR _9709_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_146_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_192 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_123 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_99 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_54 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_92 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_302 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_196 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6370_ _6368_/Y _5757_/B _6369_/Y _5810_/B VGND VPWR _6370_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_127_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5321_ _9500_/Q _5319_/A _8845_/X _5319_/Y VGND VPWR _9500_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8040_ _8624_/B _8552_/A VGND VPWR _8685_/A VGND VPWR sky130_fd_sc_hd__nor2_1
X_5252_ _5252_/A VGND VPWR _5253_/A VGND VPWR sky130_fd_sc_hd__clkbuf_2
X_5183_ _9591_/Q _5180_/A _8842_/X _5180_/Y VGND VPWR _9591_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_3_60 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_484 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_8942_ _9089_/Q _9088_/Q _9051_/Q VGND VPWR _8942_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_36_262 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8873_ _8872_/X _9175_/Q _9054_/Q VGND VPWR _8873_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_7824_ _8538_/C _7899_/A _8084_/A VGND VPWR _7825_/A VGND VPWR sky130_fd_sc_hd__or3_1
XFILLER_24_446 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_243 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7755_ _8660_/A VGND VPWR _8299_/A VGND VPWR sky130_fd_sc_hd__inv_2
X_4967_ _9707_/Q _4966_/A _9706_/Q _4966_/Y VGND VPWR _9707_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7686_ _6330_/Y _7434_/X _6347_/Y _7436_/X VGND VPWR _7686_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4898_ _4898_/A _4931_/B VGND VPWR _5344_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_6706_ _6706_/A VGND VPWR _6706_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
XFILLER_137_315 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6637_ _9206_/Q VGND VPWR _6637_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_192_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9425_ _9527_/CLK _9425_/D _9647_/SET_B VGND VPWR _9425_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_9356_ _9358_/CLK _9356_/D _9685_/SET_B VGND VPWR _9356_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6568_ _9497_/Q VGND VPWR _8789_/A VGND VPWR sky130_fd_sc_hd__clkinv_8
XFILLER_164_167 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_8307_ _8305_/B _8264_/B _8441_/A VGND VPWR _8310_/B VGND VPWR sky130_fd_sc_hd__o21ai_1
X_5519_ _5519_/A VGND VPWR _5520_/A VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_105_212 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_543 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6499_ _6497_/Y _5742_/B _6498_/Y _5810_/B VGND VPWR _6499_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_9287_ _9483_/CLK _9287_/D _9528_/SET_B VGND VPWR _9287_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_8238_ _8238_/A _8260_/B VGND VPWR _8574_/B VGND VPWR sky130_fd_sc_hd__nor2_1
X_8169_ _8169_/A VGND VPWR _8373_/A VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_59_332 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_484 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_50 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_262 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_43 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_287 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_440 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_612 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_80 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_318 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_188 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_384 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_438 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5870_ _9160_/Q _5866_/A _5966_/B1 _5866_/Y VGND VPWR _9160_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_4821_ _4821_/A VGND VPWR _4821_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_61_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_602 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4752_ _4787_/A _4929_/A VGND VPWR _5545_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_7540_ _6372_/Y _7415_/X _6462_/Y _7417_/X _7539_/X VGND VPWR _7554_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_119_315 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4683_ input61/X _4680_/Y _4681_/Y _6052_/C VGND VPWR _4683_/X VGND VPWR sky130_fd_sc_hd__o2bb2a_1
X_7471_ _7471_/A VGND VPWR _7471_/X VGND VPWR sky130_fd_sc_hd__buf_8
X_9210_ _9652_/CLK _9210_/D _9647_/SET_B VGND VPWR _9210_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6422_ _9446_/Q VGND VPWR _6422_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_134_329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_9141_ _9278_/CLK _9141_/D _9757_/SET_B VGND VPWR _9141_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6353_ _9194_/Q VGND VPWR _6353_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_161_159 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_351 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6284_ _9182_/Q VGND VPWR _6284_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_5304_ _9511_/Q _5300_/A _5966_/B1 _5300_/Y VGND VPWR _9511_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_9072_ _9358_/CLK _9072_/D _9685_/SET_B VGND VPWR _9072_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_88_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5235_ _9558_/Q _5234_/A _5963_/B1 _5234_/Y VGND VPWR _9558_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8023_ _8389_/A _8130_/B _8020_/X _8403_/A _8450_/A VGND VPWR _8023_/X VGND VPWR
+ sky130_fd_sc_hd__o2111a_1
X_5166_ _9602_/Q _5158_/A _8916_/A1 _5158_/Y VGND VPWR _9602_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_5097_ _9648_/Q _5091_/A _8955_/A1 _5091_/Y VGND VPWR _9648_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_71_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8925_ _9606_/Q _8925_/A1 _8926_/S VGND VPWR _8925_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_17_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_216 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_8856_ _7554_/Y _9636_/Q _8978_/S VGND VPWR _8856_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XPHY_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_238 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_227 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5999_ _9088_/Q _5995_/A _8913_/X _5995_/Y VGND VPWR _9088_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7807_ _8394_/D _8521_/A VGND VPWR _8119_/A VGND VPWR sky130_fd_sc_hd__or2_2
X_8787_ _8787_/A VGND VPWR _8788_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_33_35 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_7738_ _9066_/Q _7738_/B VGND VPWR _7738_/X VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_177_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_460 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_218 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9408_ _9493_/CLK _9408_/D _4628_/A VGND VPWR _9408_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_7669_ _6479_/Y _7430_/X _6597_/Y _7432_/X _7668_/X VGND VPWR _7669_/X VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_137_156 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9339_ _9508_/CLK _9339_/D _9647_/SET_B VGND VPWR _9339_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_3_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xoutput290 _9756_/Q VGND VPWR pll_trim[24] VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_75_611 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_184 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_64 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_360 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_63 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_50 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_192 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5020_ _9691_/Q _5015_/A _8929_/A1 _5015_/Y VGND VPWR _9691_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_78_471 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_579 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_154 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_102 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_8710_ _8710_/A VGND VPWR _8710_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_6971_ _6946_/Y _6964_/A _9021_/Q _6964_/Y VGND VPWR _9021_/D VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_179_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5922_ _9121_/Q _5918_/A _8930_/A1 _5918_/Y VGND VPWR _9121_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_9690_ _9695_/CLK _9690_/D _9779_/SET_B VGND VPWR _9690_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_34_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_179 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8641_ _8641_/A _8641_/B _8641_/C _8343_/Y VGND VPWR _8719_/C VGND VPWR sky130_fd_sc_hd__or4b_2
X_5853_ _5849_/X _8867_/X _8924_/X _9173_/Q VGND VPWR _9173_/D VGND VPWR sky130_fd_sc_hd__o22a_2
Xclkbuf_leaf_15_csclk clkbuf_2_3_0_csclk/X VGND VPWR _9501_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_61_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5784_ _9220_/Q _5778_/A _8955_/A1 _5778_/Y VGND VPWR _9220_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8572_ _8641_/B _8719_/A _8572_/C _8677_/C VGND VPWR _8576_/A VGND VPWR sky130_fd_sc_hd__or4_1
X_4804_ _9346_/Q VGND VPWR _4804_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
X_7523_ _8793_/A _7427_/X _8763_/A _5699_/X VGND VPWR _7523_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4735_ _6158_/B _4780_/B VGND VPWR _5797_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_162_413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7454_ _7456_/A _7466_/A _7474_/D VGND VPWR _7455_/A VGND VPWR sky130_fd_sc_hd__or3_1
X_4666_ _4666_/A VGND VPWR _4843_/B VGND VPWR sky130_fd_sc_hd__buf_8
X_6405_ _9744_/Q VGND VPWR _6405_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7385_ _6373_/Y _7068_/A _6412_/Y _7105_/X VGND VPWR _7385_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4597_ _9735_/Q _4592_/A _5964_/B1 _4592_/Y VGND VPWR _9735_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_1_607 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6336_ _6336_/A VGND VPWR _6336_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_162_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9124_ _9655_/CLK _9124_/D _7011_/B VGND VPWR _9124_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_115_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9055_ _9203_/CLK _9055_/D _9633_/SET_B VGND VPWR _9055_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_95_19 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_490 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6267_ _6262_/Y _4907_/X _6263_/Y _5240_/B _6266_/X VGND VPWR _6280_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_57_611 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5218_ _5218_/A VGND VPWR _5218_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_130_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6198_ _6193_/Y _6322_/A _6194_/Y _5837_/B _6197_/X VGND VPWR _6211_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_8006_ _8525_/C VGND VPWR _8064_/C VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_151_14 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_346 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_590 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5149_ _9616_/Q _5147_/A _8845_/X _5147_/Y VGND VPWR _9616_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_151_36 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_316 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8908_ _7726_/Y _4949_/A _9048_/Q VGND VPWR _8908_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_52_360 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_8839_ _4949_/A _9659_/Q _9587_/Q VGND VPWR _8839_/X VGND VPWR sky130_fd_sc_hd__mux2_8
XFILLER_185_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_246 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_88 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_210 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_17 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_243 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_332 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_600 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_176 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_390 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_218 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4520_ _5967_/B1 _9770_/Q _4520_/S VGND VPWR _4521_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_4451_ _9575_/Q _4901_/A _9081_/Q VGND VPWR _8990_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_7170_ _6694_/Y _7118_/X _6686_/Y _7048_/C VGND VPWR _7170_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_98_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6121_ _9211_/Q VGND VPWR _6121_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_124_192 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6052_ _6052_/A _6052_/B _6052_/C VGND VPWR _6053_/A VGND VPWR sky130_fd_sc_hd__or3_2
XFILLER_85_216 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5003_ _6040_/A VGND VPWR _5004_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_53_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_17 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_9742_ _9777_/CLK _9742_/D _9757_/SET_B VGND VPWR _9742_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6954_ _6237_/Y _6952_/A _9034_/Q _6952_/Y VGND VPWR _9034_/D VGND VPWR sky130_fd_sc_hd__o22a_1
X_9673_ _9674_/CLK _9673_/D _9633_/SET_B VGND VPWR _9673_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_5905_ _6052_/A _5905_/B VGND VPWR _5906_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_6885_ _9329_/Q VGND VPWR _6885_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_8624_ _8632_/A _8624_/B VGND VPWR _8624_/X VGND VPWR sky130_fd_sc_hd__and2_1
X_5836_ _9185_/Q _5831_/A _5967_/B1 _5831_/Y VGND VPWR _9185_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_5767_ _9231_/Q _5759_/A _8839_/X _5759_/Y VGND VPWR _9231_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8555_ _8119_/A _8397_/B _8168_/A _8401_/B _8169_/A VGND VPWR _8631_/B VGND VPWR
+ sky130_fd_sc_hd__o221ai_1
X_4718_ _9307_/Q VGND VPWR _4718_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7506_ _6694_/Y _7434_/X _6760_/Y _7436_/X VGND VPWR _7506_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_5698_ _7456_/A _7462_/A _7474_/D VGND VPWR _5699_/A VGND VPWR sky130_fd_sc_hd__or3_1
X_8486_ _8514_/B _8485_/X VGND VPWR _8486_/X VGND VPWR sky130_fd_sc_hd__or2b_1
XFILLER_162_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7437_ _4846_/Y _7434_/X _4926_/Y _7436_/X VGND VPWR _7437_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4649_ _9714_/Q _4636_/A _8949_/X _4636_/Y VGND VPWR _9714_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_135_468 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_416 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7368_ _6606_/Y _7118_/X _6503_/Y _7048_/C VGND VPWR _7368_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_89_555 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_23 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9107_ _9378_/CLK _9107_/D _9646_/SET_B VGND VPWR _9107_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6319_ _6314_/Y _5089_/B _6315_/Y _5949_/B _6318_/X VGND VPWR _6325_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_7299_ _7299_/A _7299_/B _7299_/C _7299_/D VGND VPWR _7309_/B VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_130_162 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9038_ _9664_/CLK _9038_/D VGND VPWR _9038_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_29_154 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_208 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_11 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_544 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_87 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_446 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_470 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_216 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_463 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_430 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_422 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_527 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6670_ _9734_/Q VGND VPWR _6670_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_5621_ _6052_/A _5621_/B VGND VPWR _5622_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_5552_ _9341_/Q _5547_/A _8929_/A1 _5547_/Y VGND VPWR _9341_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8340_ _8079_/C _8340_/B _8340_/C _8394_/A VGND VPWR _8722_/A VGND VPWR sky130_fd_sc_hd__and4b_1
X_4503_ _4911_/A _4921_/A VGND VPWR _4504_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_8271_ _8271_/A _8506_/B VGND VPWR _8273_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_117_468 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5483_ _9389_/Q _5482_/A _5963_/B1 _5482_/Y VGND VPWR _9389_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_144_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7222_ _6274_/Y _7086_/X _6239_/Y _7088_/X VGND VPWR _7222_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_7153_ _6871_/Y _7124_/X _6884_/Y _7068_/B _7152_/X VGND VPWR _7154_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_7084_ _7084_/A VGND VPWR _7084_/X VGND VPWR sky130_fd_sc_hd__buf_8
X_6104_ _9077_/Q VGND VPWR _6104_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
X_6035_ _9072_/Q _6029_/A _8841_/X _6029_/Y VGND VPWR _9072_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_100_357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_47 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_9725_ _9769_/CLK _9725_/D _9757_/SET_B VGND VPWR _9725_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_7986_ _7986_/A VGND VPWR _8551_/A VGND VPWR sky130_fd_sc_hd__buf_2
XPHY_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_47 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6937_ _6932_/Y _5789_/B _6933_/Y _5818_/B _6936_/X VGND VPWR _6944_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_6868_ _9542_/Q VGND VPWR _6868_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9656_ _9779_/CLK _9656_/D _9779_/SET_B VGND VPWR _9656_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_9587_ _4450_/A1 _9587_/D _6146_/A VGND VPWR _9587_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_8607_ _8607_/A _8607_/B _8607_/C _7910_/X VGND VPWR _8735_/A VGND VPWR sky130_fd_sc_hd__or4b_2
X_5819_ _5819_/A VGND VPWR _5820_/A VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_155_519 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6799_ _9126_/Q VGND VPWR _6799_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_8538_ _8583_/A _8538_/B _8538_/C _8538_/D VGND VPWR _8538_/X VGND VPWR sky130_fd_sc_hd__or4_1
XFILLER_157_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_254 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8469_ _7848_/A _8305_/A _8097_/B _8554_/A VGND VPWR _8698_/A VGND VPWR sky130_fd_sc_hd__o22ai_1
XFILLER_150_235 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_374 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_154 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_327 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_344 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xinput190 wb_dat_i[4] VGND VPWR _8965_/A1 VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_7840_ _8379_/D _8394_/B _8394_/C _8195_/A VGND VPWR _7841_/A VGND VPWR sky130_fd_sc_hd__or4_1
XFILLER_36_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7771_ _7771_/A _7771_/B _7771_/C _7771_/D VGND VPWR _7775_/C VGND VPWR sky130_fd_sc_hd__nand4_1
X_4983_ _4994_/A VGND VPWR _4984_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_6722_ _6717_/Y _5317_/B _6718_/Y _5518_/B _6721_/X VGND VPWR _6741_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9510_ _9514_/CLK _9510_/D _4628_/A VGND VPWR _9510_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6653_ _8803_/A VGND VPWR _6653_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9441_ _9514_/CLK _9441_/D _9685_/SET_B VGND VPWR _9441_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_149_379 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5604_ _5604_/A VGND VPWR _5604_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_191_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9372_ _9379_/CLK _9372_/D _9779_/SET_B VGND VPWR _9372_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6584_ _6582_/Y _5621_/B _6583_/Y _5526_/B VGND VPWR _6584_/X VGND VPWR sky130_fd_sc_hd__o22a_2
XFILLER_11_49 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8323_ _8463_/A _8645_/B VGND VPWR _8599_/C VGND VPWR sky130_fd_sc_hd__or2_1
X_5535_ _5535_/A VGND VPWR _5536_/A VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_145_596 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5466_ _9400_/Q _5460_/A _5965_/B1 _5460_/Y VGND VPWR _9400_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8254_ _8341_/A _8254_/B VGND VPWR _8493_/B VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_105_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_438 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7205_ _6329_/Y _7097_/X _6349_/Y _7099_/X VGND VPWR _7205_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_8185_ _8185_/A VGND VPWR _8514_/A VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_160_577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5397_ _9448_/Q _5395_/A _8845_/X _5395_/Y VGND VPWR _9448_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_101_611 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7136_ _6825_/Y _7082_/X _6787_/Y _7084_/X _7135_/X VGND VPWR _7155_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_86_344 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7067_ _7067_/A VGND VPWR _7068_/D VGND VPWR sky130_fd_sc_hd__clkbuf_16
X_6018_ _8916_/A1 _9081_/Q _6018_/S VGND VPWR _6019_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_15_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7969_ _7969_/A _8120_/B VGND VPWR _7970_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_9708_ _9709_/CLK _9708_/D _4957_/X VGND VPWR _9708_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_9639_ _9639_/CLK _9639_/D _9633_/SET_B VGND VPWR _9639_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_167_154 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_135 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_276 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_66 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_600 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_308 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5320_ _9501_/Q _5319_/A _8846_/X _5319_/Y VGND VPWR _9501_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_142_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5251_ _5259_/A _5251_/B VGND VPWR _5252_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_87_119 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5182_ _9592_/Q _5180_/A _8925_/A1 _5180_/Y VGND VPWR _9592_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_3_72 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6999__13 _6997_/X VGND VPWR _7000_/B2 VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_95_163 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_8941_ _8940_/X _9681_/Q _9587_/Q VGND VPWR _8941_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_83_325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_8872_ _7698_/Y _9631_/Q _8978_/S VGND VPWR _8872_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_51_211 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_274 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_414 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7823_ _7823_/A _7823_/B _8538_/B VGND VPWR _7899_/A VGND VPWR sky130_fd_sc_hd__or3b_1
X_7754_ _8379_/D _8394_/B _7838_/B VGND VPWR _8660_/A VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_51_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_4966_ _4966_/A VGND VPWR _4966_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_6705_ _9486_/Q VGND VPWR _6705_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
XFILLER_22_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7685_ _6391_/Y _7427_/X _6361_/Y _5699_/X VGND VPWR _7685_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4897_ _9476_/Q VGND VPWR _4897_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
X_9424_ _9535_/CLK _9424_/D _9528_/SET_B VGND VPWR _9424_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6636_ _7172_/A _5610_/B _6632_/Y _5594_/B _6635_/X VGND VPWR _6649_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_6567_ _6567_/A _6567_/B _6567_/C _6567_/D VGND VPWR _6628_/A VGND VPWR sky130_fd_sc_hd__and4_1
X_9355_ _9358_/CLK _9355_/D _9685_/SET_B VGND VPWR _9355_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_192_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8306_ _8521_/B _7885_/B _8447_/B _8215_/X _8397_/A VGND VPWR _8306_/X VGND VPWR
+ sky130_fd_sc_hd__o2111a_1
X_5518_ _5671_/A _5518_/B VGND VPWR _5519_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_145_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_9286_ _9483_/CLK _9286_/D _9528_/SET_B VGND VPWR _9286_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6498_ _9201_/Q VGND VPWR _6498_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_133_555 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5449_ _9411_/Q _5444_/A _5967_/B1 _5444_/Y VGND VPWR _9411_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8237_ _8237_/A _8358_/B _8642_/B _8359_/B VGND VPWR _8241_/A VGND VPWR sky130_fd_sc_hd__or4_1
X_8168_ _8168_/A _8378_/B VGND VPWR _8169_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_86_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_344 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_12 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7119_ _4846_/Y _7118_/X _4675_/Y _7048_/C VGND VPWR _7119_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_8099_ _8195_/A _8099_/B VGND VPWR _8100_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_47_89 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_84 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_406 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_102 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_599 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_238 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_80 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4820_ _4813_/Y _4537_/B _4814_/Y _6027_/B _4819_/X VGND VPWR _4830_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_159_441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4751_ _9338_/Q VGND VPWR _4751_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_159_474 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_260 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7470_ _7472_/A _7470_/B _9255_/Q VGND VPWR _7471_/A VGND VPWR sky130_fd_sc_hd__or3_1
X_4682_ _4787_/A _4876_/B VGND VPWR _6052_/C VGND VPWR sky130_fd_sc_hd__or2_4
X_6421_ _9376_/Q VGND VPWR _6421_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_174_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9140_ _9278_/CLK _9140_/D _9757_/SET_B VGND VPWR _9140_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_161_127 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6352_ _6352_/A _6352_/B _6352_/C _6352_/D VGND VPWR _6475_/A VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_154_190 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5303_ _9512_/Q _5300_/A _5965_/B1 _5300_/Y VGND VPWR _9512_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_9071_ _9358_/CLK _9071_/D _9685_/SET_B VGND VPWR _9071_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6283_ _9299_/Q VGND VPWR _7238_/A VGND VPWR sky130_fd_sc_hd__clkinv_2
X_5234_ _5234_/A VGND VPWR _5234_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_8022_ _8624_/B _8130_/B VGND VPWR _8450_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_5165_ _9603_/Q _5158_/A _8840_/X _5158_/Y VGND VPWR _9603_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_68_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_100 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5096_ _9649_/Q _5091_/A _8929_/A1 _5091_/Y VGND VPWR _9649_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_37_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8924_ _9055_/Q _8819_/X _9054_/Q VGND VPWR _8924_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_83_199 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8855_ _8854_/X _9166_/Q _9054_/Q VGND VPWR _8855_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XPHY_206 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_7806_ _7806_/A VGND VPWR _8521_/A VGND VPWR sky130_fd_sc_hd__buf_8
XPHY_239 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_228 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5998_ _5998_/A VGND VPWR _5998_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_8786_ _8786_/A VGND VPWR _8786_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_7737_ _9068_/Q _7737_/A2 _9067_/Q _7737_/B2 _7736_/X VGND VPWR _7737_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_4949_ _4949_/A VGND VPWR _4949_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_130_7 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_102 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7668_ _6606_/Y _7434_/X _6604_/Y _7436_/X VGND VPWR _7668_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_20_472 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6619_ _6617_/Y _5121_/B _6618_/Y _4870_/X VGND VPWR _6619_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_9407_ _9493_/CLK _9407_/D _4628_/A VGND VPWR _9407_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_153_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7599_ _6074_/Y _7445_/X _6090_/Y _7447_/X VGND VPWR _7599_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_106_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9338_ _9535_/CLK _9338_/D _9528_/SET_B VGND VPWR _9338_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_3_126 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_79 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9269_ _9535_/CLK _9269_/D _9528_/SET_B VGND VPWR _9269_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_160_160 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xoutput280 _9747_/Q VGND VPWR pll_trim[15] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput291 _9757_/Q VGND VPWR pll_trim[25] VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_87_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_196 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_76 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_247 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_75 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_40 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_90 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_5 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_494 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6970_ _6785_/Y _6964_/A _9022_/Q _6964_/Y VGND VPWR _9022_/D VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_19_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5921_ _9122_/Q _5918_/A _5965_/B1 _5918_/Y VGND VPWR _9122_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_179_536 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8640_ _8640_/A _8640_/B _8640_/C VGND VPWR _8641_/C VGND VPWR sky130_fd_sc_hd__nor3_1
X_5852_ _5849_/X _8869_/X _8924_/X _9174_/Q VGND VPWR _9174_/D VGND VPWR sky130_fd_sc_hd__o22a_2
XFILLER_21_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8571_ _8571_/A _8571_/B _8571_/C VGND VPWR _8677_/C VGND VPWR sky130_fd_sc_hd__or3_1
X_5783_ _9221_/Q _5778_/A _8929_/A1 _5778_/Y VGND VPWR _9221_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_4803_ _4903_/B _4931_/B VGND VPWR _5290_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_9_71 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4734_ _9204_/Q VGND VPWR _4734_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7522_ _8753_/A _7415_/X _8745_/A _7417_/X _7521_/X VGND VPWR _7536_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_119_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4665_ _8936_/X _4665_/B _4665_/C VGND VPWR _4666_/A VGND VPWR sky130_fd_sc_hd__or3_1
X_7453_ _7453_/A VGND VPWR _7453_/X VGND VPWR sky130_fd_sc_hd__buf_8
X_4596_ _9736_/Q _4592_/A _5963_/B1 _4592_/Y VGND VPWR _9736_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7384_ _6393_/Y _7059_/B _6423_/Y _7068_/C _7383_/X VGND VPWR _7387_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_6404_ _9389_/Q VGND VPWR _6404_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_6335_ _9384_/Q VGND VPWR _6335_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9123_ _9655_/CLK _9123_/D _9779_/SET_B VGND VPWR _9123_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_115_385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_9054_ _9278_/CLK _9054_/D _9633_/SET_B VGND VPWR _9054_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_88_236 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8005_ _8005_/A VGND VPWR _8566_/B VGND VPWR sky130_fd_sc_hd__inv_2
X_6266_ _6264_/Y _5431_/B _6265_/Y _4602_/B VGND VPWR _6266_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_57_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6197_ _6195_/Y _5355_/B _6196_/Y _5344_/B VGND VPWR _6197_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_5217_ _6135_/A _6322_/A _5259_/A _8976_/X VGND VPWR _5218_/A VGND VPWR sky130_fd_sc_hd__a211o_4
X_5148_ _9617_/Q _5147_/A _8846_/X _5147_/Y VGND VPWR _9617_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_151_26 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_48 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5079_ _5079_/A VGND VPWR _9659_/D VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_29_358 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8907_ _7725_/X _9088_/Q _9051_/Q VGND VPWR _8907_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_71_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8838_ input85/X _4949_/A _9626_/Q VGND VPWR _8838_/X VGND VPWR sky130_fd_sc_hd__mux2_2
X_8769_ _8769_/A VGND VPWR _8770_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_40_512 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_523 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_466 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_222 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_612 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_464 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_188 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_422 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_291 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4450_ _9576_/Q _4450_/A1 _9788_/Q VGND VPWR _8991_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_6120_ _9695_/Q VGND VPWR _6120_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_152_480 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_206 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6051_ _6051_/A VGND VPWR _6051_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_112_399 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5002_ _5002_/A VGND VPWR _9698_/D VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_38_133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9741_ _9777_/CLK _9741_/D _9757_/SET_B VGND VPWR _9741_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6953_ _6145_/Y _6952_/A _9035_/Q _6952_/Y VGND VPWR _9035_/D VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_53_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5904_ _9133_/Q _5899_/A _8839_/X _5899_/Y VGND VPWR _9133_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_9672_ _9695_/CLK _9672_/D _9779_/SET_B VGND VPWR _9672_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6884_ _9313_/Q VGND VPWR _6884_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_179_344 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5835_ _9186_/Q _5831_/A _5966_/B1 _5831_/Y VGND VPWR _9186_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8623_ _8098_/A _8622_/X _8547_/X VGND VPWR _8710_/A VGND VPWR sky130_fd_sc_hd__o21ai_2
XFILLER_139_219 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_567 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5766_ _9232_/Q _5759_/A _8840_/X _5759_/Y VGND VPWR _9232_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8554_ _8554_/A _8554_/B VGND VPWR _8709_/A VGND VPWR sky130_fd_sc_hd__nor2_1
X_5697_ _9255_/Q VGND VPWR _7474_/D VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_175_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7505_ _6763_/Y _7427_/X _6661_/Y _5699_/X VGND VPWR _7505_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4717_ _4876_/B _4843_/B VGND VPWR _5837_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_8485_ _8485_/A _8514_/C VGND VPWR _8485_/X VGND VPWR sky130_fd_sc_hd__or2_1
X_7436_ _7436_/A VGND VPWR _7436_/X VGND VPWR sky130_fd_sc_hd__buf_6
X_4648_ _4648_/A VGND VPWR _4648_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_162_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9106_ _9379_/CLK _9106_/D _9646_/SET_B VGND VPWR _9106_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_7367_ _6486_/Y _7040_/D _6508_/Y _7110_/X _7366_/X VGND VPWR _7374_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_4579_ _4579_/A VGND VPWR _4579_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_115_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6318_ _6316_/Y _5660_/B _6317_/Y _6134_/A VGND VPWR _6318_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_7298_ _4685_/Y _7048_/D _4823_/Y _7040_/B _7297_/X VGND VPWR _7299_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_1_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_355 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_206 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_35 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6249_ _6249_/A VGND VPWR _6249_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9037_ _9664_/CLK _9037_/D VGND VPWR _9037_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_72_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_434 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_62 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_556 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_550 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_542 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_458 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_428 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_575 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_119 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_439 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_14_csclk clkbuf_2_2_0_csclk/X VGND VPWR _9534_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_96_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_29_csclk clkbuf_2_3_0_csclk/X VGND VPWR _9653_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_63_456 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_174 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_539 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5620_ _9294_/Q _5612_/A _8916_/A1 _5612_/Y VGND VPWR _9294_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_157_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5551_ _9342_/Q _5547_/A _8925_/A1 _5547_/Y VGND VPWR _9342_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8270_ _8341_/A _8270_/B VGND VPWR _8506_/B VGND VPWR sky130_fd_sc_hd__nor2_1
X_4502_ _8934_/X _8932_/X _8946_/X _4729_/B VGND VPWR _4921_/A VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_105_609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5482_ _5482_/A VGND VPWR _5482_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7221_ _7221_/A _7221_/B _7221_/C VGND VPWR _7221_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
XFILLER_144_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7152_ _6823_/Y _7126_/X _6844_/Y _7128_/X VGND VPWR _7152_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_112_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7083_ _7098_/C _7125_/A _7127_/C VGND VPWR _7084_/A VGND VPWR sky130_fd_sc_hd__or3_1
X_6103_ _9423_/Q VGND VPWR _6103_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
X_6034_ _9073_/Q _6029_/A _8842_/X _6029_/Y VGND VPWR _9073_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_94_581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_412 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_7985_ _7997_/B _7992_/B VGND VPWR _7986_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_14_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_37 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6936_ _7326_/A _5632_/B _6935_/Y _5768_/B VGND VPWR _6936_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_9724_ _9769_/CLK _9724_/D _9757_/SET_B VGND VPWR _9724_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XPHY_59 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_139 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_303 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9655_ _9655_/CLK _9655_/D _9779_/SET_B VGND VPWR _9655_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6867_ _9412_/Q VGND VPWR _6867_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_41_14 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_9586_ _8837_/A1 _9586_/D _5190_/X VGND VPWR _9586_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_6798_ _6793_/Y _5534_/B _6794_/Y _4907_/X _6797_/X VGND VPWR _6830_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_5818_ _6052_/A _5818_/B VGND VPWR _5819_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_8606_ _8672_/B _8606_/B VGND VPWR _8705_/B VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_148_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5749_ _9240_/Q _5744_/A _8839_/X _5744_/Y VGND VPWR _9240_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8537_ _7836_/A _8299_/B _8061_/C _8536_/Y _8474_/B VGND VPWR _8617_/B VGND VPWR
+ sky130_fd_sc_hd__a311o_1
XFILLER_6_519 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8468_ _8468_/A _8630_/A VGND VPWR _8470_/B VGND VPWR sky130_fd_sc_hd__or2_1
X_8399_ _8213_/A _8117_/B _8395_/X _8398_/Y VGND VPWR _8399_/X VGND VPWR sky130_fd_sc_hd__o211a_1
X_7419_ _7419_/A VGND VPWR _7419_/X VGND VPWR sky130_fd_sc_hd__buf_6
XFILLER_150_247 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_246 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_472 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_386 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_507 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_518 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_55 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_423 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_61 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_6 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_428 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_480 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_356 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput180 wb_dat_i[24] VGND VPWR _7737_/A2 VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput191 wb_dat_i[5] VGND VPWR _8966_/A1 VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_91_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_540 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4982_ _9702_/Q _4966_/A _9701_/Q _4966_/Y VGND VPWR _9702_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7770_ _7770_/A _7770_/B VGND VPWR _7775_/B VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_189_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6721_ _6719_/Y _5450_/B _6720_/Y _5431_/B VGND VPWR _6721_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_189_494 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9440_ _9440_/CLK _9440_/D _4628_/A VGND VPWR _9440_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6652_ _9775_/Q VGND VPWR _6652_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
XFILLER_149_369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9371_ _9371_/CLK _9371_/D _9295_/SET_B VGND VPWR _9371_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_5603_ _5603_/A VGND VPWR _5604_/A VGND VPWR sky130_fd_sc_hd__clkbuf_2
X_8322_ _7862_/Y _8302_/Y _8318_/X _8493_/C _8657_/A VGND VPWR _8327_/A VGND VPWR
+ sky130_fd_sc_hd__a2111o_2
X_6583_ _9357_/Q VGND VPWR _6583_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
X_5534_ _5545_/A _5534_/B VGND VPWR _5535_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_5465_ _9401_/Q _5460_/A _5964_/B1 _5460_/Y VGND VPWR _9401_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8253_ _8253_/A _8577_/B VGND VPWR _8255_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_160_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7204_ _6353_/Y _7048_/B _6462_/Y _7077_/A _7203_/X VGND VPWR _7211_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_8184_ _8184_/A _8636_/B VGND VPWR _8295_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_5396_ _9449_/Q _5395_/A _8846_/X _5395_/Y VGND VPWR _9449_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7135_ _6891_/Y _7077_/C _6916_/Y _7077_/D _7134_/X VGND VPWR _7135_/X VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_86_323 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7066_ _9246_/Q _9245_/Q _7098_/C _7073_/C VGND VPWR _7067_/A VGND VPWR sky130_fd_sc_hd__or4_1
XFILLER_86_356 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6017_ _9082_/Q _5995_/A _8902_/X _5995_/Y VGND VPWR _9082_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_54_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7968_ _7968_/A _8218_/A VGND VPWR _8120_/B VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_52_13 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7899_ _7899_/A _8525_/C VGND VPWR _8472_/A VGND VPWR sky130_fd_sc_hd__or2_2
X_9707_ _4446_/A1 _9707_/D _4963_/X VGND VPWR _9707_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6919_ _9107_/Q VGND VPWR _6919_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_9638_ _9639_/CLK _9638_/D _9633_/SET_B VGND VPWR _9638_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_183_604 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_9569_ _8837_/A1 _9569_/D _5213_/X VGND VPWR _9569_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_10_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_191 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_75 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_612 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_492 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5250_ _9546_/Q _5242_/A _5967_/B1 _5242_/Y VGND VPWR _9546_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_5_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_40 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5181_ _9593_/Q _5180_/A _8844_/X _5180_/Y VGND VPWR _9593_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8940_ _9088_/Q _9087_/Q _9051_/Q VGND VPWR _8940_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_3_84 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_231 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8871_ _8870_/X _9174_/Q _9054_/Q VGND VPWR _8871_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_36_286 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7822_ _8202_/A _8272_/A VGND VPWR _8703_/A VGND VPWR sky130_fd_sc_hd__nor2_4
X_7753_ _8394_/C _7839_/A VGND VPWR _7838_/B VGND VPWR sky130_fd_sc_hd__or2_2
X_4965_ _4965_/A VGND VPWR _4966_/A VGND VPWR sky130_fd_sc_hd__buf_8
X_6704_ _9470_/Q VGND VPWR _6704_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_177_431 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7684_ _6373_/Y _7415_/X _6416_/Y _7417_/X _7683_/X VGND VPWR _7698_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_4896_ _4896_/A _4896_/B _4896_/C _4896_/D VGND VPWR _4935_/C VGND VPWR sky130_fd_sc_hd__and4_1
X_9423_ _9684_/CLK _9423_/D _9685_/SET_B VGND VPWR _9423_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6635_ _6633_/Y _5660_/B _6634_/Y _5671_/B VGND VPWR _6635_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_164_136 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_520 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6566_ _6561_/Y _4832_/X _8791_/A _5355_/B _6565_/X VGND VPWR _6567_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9354_ _9354_/CLK _9354_/D _9685_/SET_B VGND VPWR _9354_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_152_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5517_ _9364_/Q _5509_/A _8839_/X _5509_/Y VGND VPWR _9364_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_9285_ _9687_/CLK _9285_/D _9528_/SET_B VGND VPWR _9285_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_8305_ _8305_/A _8305_/B VGND VPWR _8447_/B VGND VPWR sky130_fd_sc_hd__or2_1
X_8236_ _8236_/A VGND VPWR _8359_/B VGND VPWR sky130_fd_sc_hd__inv_2
X_6497_ _9243_/Q VGND VPWR _6497_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_5448_ _9412_/Q _5444_/A _5966_/B1 _5444_/Y VGND VPWR _9412_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_87_610 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5379_ _9460_/Q _5376_/A _8841_/X _5376_/Y VGND VPWR _9460_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8167_ _8167_/A _8715_/A VGND VPWR _8172_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_99_492 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8098_ _8098_/A _8098_/B VGND VPWR _8688_/A VGND VPWR sky130_fd_sc_hd__nor2_1
X_7118_ _7118_/A VGND VPWR _7118_/X VGND VPWR sky130_fd_sc_hd__buf_8
XFILLER_86_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_356 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_24 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7049_ _7098_/C _7125_/A _7073_/C VGND VPWR _7050_/A VGND VPWR sky130_fd_sc_hd__or3_1
XFILLER_74_326 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_30 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_96 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_383 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_164 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_315 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_80 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_264 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_212 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4750_ _4787_/A _4900_/B VGND VPWR _5602_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_186_272 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4681_ _9044_/Q VGND VPWR _4681_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
X_6420_ _6415_/Y _5382_/B _6416_/Y _5941_/B _6419_/X VGND VPWR _6433_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_115_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6351_ _6346_/Y _5267_/B _6347_/Y _5328_/B _6350_/X VGND VPWR _6352_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_127_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5302_ _9513_/Q _5300_/A _5964_/B1 _5300_/Y VGND VPWR _9513_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_9070_ _9687_/CLK _9070_/D _9685_/SET_B VGND VPWR _9070_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6282_ _9672_/Q VGND VPWR _6282_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_8021_ _8521_/A _8130_/B VGND VPWR _8403_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_5233_ _5233_/A VGND VPWR _5234_/A VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_124_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5164_ _9604_/Q _5158_/A _8841_/X _5158_/Y VGND VPWR _9604_/D VGND VPWR sky130_fd_sc_hd__a22o_1
Xclkbuf_opt_3_0_csclk clkbuf_2_1_0_csclk/X VGND VPWR clkbuf_opt_3_0_csclk/X VGND VPWR
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_68_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_462 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5095_ _9650_/Q _5091_/A _8925_/A1 _5091_/Y VGND VPWR _9650_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8923_ _9621_/Q _8929_/A1 _8955_/S VGND VPWR _8923_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_71_329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8854_ _7536_/Y _9635_/Q _8978_/S VGND VPWR _8854_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XPHY_207 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_7805_ _7839_/A _8632_/A VGND VPWR _7806_/A VGND VPWR sky130_fd_sc_hd__or2_1
XPHY_229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_218 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5997_ _6040_/A VGND VPWR _5998_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_8785_ _8785_/A VGND VPWR _8786_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_7736_ _9066_/Q _7736_/B VGND VPWR _7736_/X VGND VPWR sky130_fd_sc_hd__and2_1
X_4948_ _4948_/A VGND VPWR _4948_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_177_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4879_ _9771_/Q VGND VPWR _4879_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7667_ _6543_/Y _7427_/X _6484_/Y _5699_/X VGND VPWR _7667_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_123_7 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6618_ _6618_/A VGND VPWR _6618_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9406_ _9493_/CLK _9406_/D _4628_/A VGND VPWR _9406_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_192_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7598_ _6127_/Y _7425_/X _7595_/X _7597_/X VGND VPWR _7608_/C VGND VPWR sky130_fd_sc_hd__o211a_1
XFILLER_152_128 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_383 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6549_ _9776_/Q VGND VPWR _6549_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9337_ _9532_/CLK _9337_/D _9528_/SET_B VGND VPWR _9337_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_106_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9268_ _9354_/CLK _9268_/D _9685_/SET_B VGND VPWR _9268_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_160_172 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8219_ _8279_/C _8311_/B VGND VPWR _8219_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
X_9199_ _9789_/CLK _9199_/D _4628_/A VGND VPWR _9199_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
Xoutput270 _9719_/Q VGND VPWR pll_ena VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput292 _9734_/Q VGND VPWR pll_trim[2] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput281 _9748_/Q VGND VPWR pll_trim[16] VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_181_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_484 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_495 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_191 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_540 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5920_ _9123_/Q _5918_/A _5964_/B1 _5918_/Y VGND VPWR _9123_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_0_74 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_548 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5851_ _5849_/X _8871_/X _8924_/X _9175_/Q VGND VPWR _9175_/D VGND VPWR sky130_fd_sc_hd__o22a_2
XFILLER_21_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5782_ _9222_/Q _5778_/A _8925_/A1 _5778_/Y VGND VPWR _9222_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8570_ _8213_/A _8117_/A _8341_/B _8260_/B _8352_/B VGND VPWR _8572_/C VGND VPWR
+ sky130_fd_sc_hd__o221ai_4
X_4802_ _4802_/A VGND VPWR _4931_/B VGND VPWR sky130_fd_sc_hd__buf_6
XFILLER_166_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_103 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7521_ _8743_/A _7419_/X _8781_/A _7421_/X VGND VPWR _7521_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4733_ _4787_/A _4917_/A VGND VPWR _5621_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_9_83 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7452_ _7466_/A _7470_/B _7474_/D VGND VPWR _7453_/A VGND VPWR sky130_fd_sc_hd__or3_1
XFILLER_119_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6403_ _9782_/Q VGND VPWR _6403_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_4664_ _9125_/Q VGND VPWR _4664_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_134_106 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4595_ _9737_/Q _4592_/A _8844_/X _4592_/Y VGND VPWR _9737_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7383_ _6417_/Y _7079_/B _6379_/Y _7059_/A VGND VPWR _7383_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_6334_ _9097_/Q VGND VPWR _6334_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9122_ _9785_/CLK _9122_/D _7011_/B VGND VPWR _9122_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_130_301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6265_ _9731_/Q VGND VPWR _6265_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9053_ _9278_/CLK _9053_/D _9633_/SET_B VGND VPWR _9053_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_88_248 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5216_ _9569_/Q _5214_/Y _5985_/B _5215_/Y VGND VPWR _9569_/D VGND VPWR sky130_fd_sc_hd__o22a_1
X_8004_ _8394_/D _8164_/A VGND VPWR _8005_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_6196_ _9482_/Q VGND VPWR _6196_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_130_356 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5147_ _5147_/A VGND VPWR _5147_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_96_292 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5078_ _8961_/X _9659_/Q _5078_/S VGND VPWR _5079_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_84_465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8906_ _9614_/Q _8925_/A1 _8930_/S VGND VPWR _8906_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_44_47 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8837_ input83/X _8837_/A1 _9586_/Q VGND VPWR _8837_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_8768_ _8768_/A VGND VPWR _8768_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_178_570 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7719_ _9087_/Q _7719_/B VGND VPWR _7721_/A VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_40_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8699_ _8699_/A _8699_/B _8699_/C _8699_/D VGND VPWR _8732_/A VGND VPWR sky130_fd_sc_hd__or4_1
XFILLER_69_11 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_248 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_70 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_456 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_492 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6050_ _6050_/A VGND VPWR _6051_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_112_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5001_ _8908_/X _9698_/Q _5001_/S VGND VPWR _5002_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_38_189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_9740_ _9777_/CLK _9740_/D _9757_/SET_B VGND VPWR _9740_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6952_ _6952_/A VGND VPWR _6952_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_6883_ _9186_/Q VGND VPWR _6883_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_5903_ _9134_/Q _5899_/A _5966_/B1 _5899_/Y VGND VPWR _9134_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_9671_ _9674_/CLK _9671_/D _9633_/SET_B VGND VPWR _9671_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_5834_ _9187_/Q _5831_/A _5965_/B1 _5831_/Y VGND VPWR _9187_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8622_ _7971_/A _8116_/B _8624_/B _8397_/A _8395_/B VGND VPWR _8622_/X VGND VPWR
+ sky130_fd_sc_hd__o311a_1
XFILLER_61_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5765_ _9233_/Q _5759_/A _8841_/X _5759_/Y VGND VPWR _9233_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8553_ _8553_/A _8627_/D _8686_/C _8630_/D VGND VPWR _8559_/A VGND VPWR sky130_fd_sc_hd__or4_2
XFILLER_22_579 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5696_ _5724_/B _7462_/A _7456_/A VGND VPWR _5696_/Y VGND VPWR sky130_fd_sc_hd__nor3_1
X_8484_ _8188_/B _8389_/A _8086_/B VGND VPWR _8514_/C VGND VPWR sky130_fd_sc_hd__o21ai_1
X_7504_ _6639_/Y _7415_/X _6681_/Y _7417_/X _7503_/X VGND VPWR _7518_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_4716_ _9177_/Q VGND VPWR _4716_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_7435_ _7472_/A _7470_/B _7474_/D VGND VPWR _7436_/A VGND VPWR sky130_fd_sc_hd__or3_1
X_4647_ _4994_/A VGND VPWR _4648_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_30_38 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7366_ _6484_/Y _7112_/X _6528_/Y _7077_/B VGND VPWR _7366_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_162_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_9 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6317_ _6317_/A VGND VPWR _6317_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9105_ _9777_/CLK _9105_/D _7011_/B VGND VPWR _9105_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_4578_ _4578_/A VGND VPWR _4579_/A VGND VPWR sky130_fd_sc_hd__clkbuf_4
X_7297_ _4712_/Y _7068_/A _4836_/Y _7105_/X VGND VPWR _7297_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_9036_ _9664_/CLK _9036_/D VGND VPWR _9036_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_6248_ _6243_/Y _4577_/B _6244_/Y _5317_/B _6247_/X VGND VPWR _6248_/X VGND VPWR
+ sky130_fd_sc_hd__o221a_2
XFILLER_39_47 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_218 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_378 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6179_ _9275_/Q VGND VPWR _6179_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_130_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_12 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_398 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_554 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_532 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_587 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_468 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_120 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_186 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5550_ _9343_/Q _5547_/A _8844_/X _5547_/Y VGND VPWR _9343_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_157_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4501_ _9778_/Q _4493_/A _5967_/B1 _4493_/Y VGND VPWR _9778_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_5481_ _5481_/A VGND VPWR _5482_/A VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_6_40 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7220_ _7220_/A _7220_/B _7220_/C _7220_/D VGND VPWR _7221_/C VGND VPWR sky130_fd_sc_hd__and4_1
XANTENNA_0 user_clock VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_125_481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_610 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7151_ _6818_/Y _5728_/X _6913_/Y _7040_/A _7150_/X VGND VPWR _7154_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_98_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6102_ _6097_/Y _4832_/X _6098_/Y _5534_/B _6101_/X VGND VPWR _6119_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_2
X_7082_ _7082_/A VGND VPWR _7082_/X VGND VPWR sky130_fd_sc_hd__buf_8
XFILLER_140_462 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6033_ _9074_/Q _6029_/A _8843_/X _6029_/Y VGND VPWR _9074_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_112_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7984_ _8525_/A _8091_/B _8098_/A VGND VPWR _7997_/B VGND VPWR sky130_fd_sc_hd__or3_2
XPHY_38 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6935_ _9227_/Q VGND VPWR _6935_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9723_ _9769_/CLK _9723_/D _9757_/SET_B VGND VPWR _9723_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XPHY_49 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_9654_ _9779_/CLK _9654_/D _9779_/SET_B VGND VPWR _9654_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6866_ _9464_/Q VGND VPWR _6866_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_167_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_315 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_186 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5817_ _9198_/Q _5812_/A _8839_/X _5812_/Y VGND VPWR _9198_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_9585_ _9674_/CLK _9585_/D _9633_/SET_B VGND VPWR _9585_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_6797_ _6795_/Y _4537_/B _6796_/Y _4564_/B VGND VPWR _6797_/X VGND VPWR sky130_fd_sc_hd__o22a_2
X_8605_ _8605_/A _8605_/B VGND VPWR _8707_/B VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_22_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_376 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8536_ _8536_/A VGND VPWR _8536_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_5748_ _9241_/Q _5744_/A _8930_/A1 _5744_/Y VGND VPWR _9241_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_148_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8467_ _8467_/A VGND VPWR _8630_/A VGND VPWR sky130_fd_sc_hd__inv_2
X_5679_ _6052_/A _5679_/B VGND VPWR _5680_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_123_407 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7418_ _7476_/A _9251_/Q _7456_/A _9255_/Q VGND VPWR _7419_/A VGND VPWR sky130_fd_sc_hd__or4_1
X_8398_ _8396_/Y _8397_/Y _8121_/Y VGND VPWR _8398_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
X_7349_ _6712_/Y _5728_/X _6685_/Y _7040_/A _7348_/X VGND VPWR _7352_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_173_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9019_ _9039_/CLK _9019_/D VGND VPWR _9019_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_106_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_402 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_55 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_88 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_314 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_492 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_598 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_379 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput170 wb_dat_i[15] VGND VPWR _7751_/B2 VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput181 wb_dat_i[25] VGND VPWR _7739_/A2 VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput192 wb_dat_i[6] VGND VPWR _8967_/A1 VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_91_552 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_298 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4981_ _4981_/A VGND VPWR _4981_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_51_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6720_ _9418_/Q VGND VPWR _6720_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_149_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6651_ _9728_/Q VGND VPWR _6651_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_6582_ _9289_/Q VGND VPWR _6582_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9370_ _9371_/CLK _9370_/D _9295_/SET_B VGND VPWR _9370_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_5602_ _5671_/A _5602_/B VGND VPWR _5603_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_31_173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5533_ _9354_/Q _5528_/A _8839_/X _5528_/Y VGND VPWR _9354_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8321_ _8461_/A _8674_/B VGND VPWR _8657_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_5464_ _9402_/Q _5460_/A _5963_/B1 _5460_/Y VGND VPWR _9402_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8252_ _8319_/A _8260_/B VGND VPWR _8577_/B VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_132_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5395_ _5395_/A VGND VPWR _5395_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7203_ _6463_/Y _7040_/C _6337_/Y _7059_/C VGND VPWR _7203_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_8183_ _8096_/A _8386_/A _8097_/B _9066_/Q VGND VPWR _8636_/B VGND VPWR sky130_fd_sc_hd__o31ai_4
XFILLER_160_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7134_ _6853_/Y _7086_/X _6855_/Y _7088_/X VGND VPWR _7134_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_7065_ _7065_/A VGND VPWR _7068_/C VGND VPWR sky130_fd_sc_hd__buf_8
X_6016_ _6016_/A VGND VPWR _6016_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_36_37 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_210 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_608 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_7967_ _7756_/B _8102_/B _7756_/B _8102_/B VGND VPWR _7968_/A VGND VPWR sky130_fd_sc_hd__o2bb2a_1
XFILLER_54_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_7 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7898_ _8008_/C _7898_/B VGND VPWR _8525_/C VGND VPWR sky130_fd_sc_hd__or2_4
X_6918_ _6913_/Y _5968_/B _6914_/Y _5621_/B _6917_/X VGND VPWR _6925_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9706_ _4446_/A1 _9706_/D _4969_/X VGND VPWR _9706_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_52_25 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6849_ _6849_/A VGND VPWR _6849_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9637_ _9791_/CLK _9637_/D _9633_/SET_B VGND VPWR _9637_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_13_csclk clkbuf_2_2_0_csclk/X VGND VPWR _9532_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_22_173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9568_ _9617_/CLK _9568_/D _9295_/SET_B VGND VPWR _9568_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_8519_ _8516_/Y _8517_/Y _8518_/X _8453_/C VGND VPWR _8607_/A VGND VPWR sky130_fd_sc_hd__a31o_1
X_9499_ _9501_/CLK _9499_/D _9647_/SET_B VGND VPWR _9499_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_28_csclk clkbuf_opt_6_0_csclk/X VGND VPWR _9378_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_123_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_338 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_184 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_80 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_622 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5180_ _5180_/A VGND VPWR _5180_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_3_52 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_508 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_198 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_176 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8870_ _7680_/Y _9630_/Q _8978_/S VGND VPWR _8870_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_7821_ _8394_/A _8394_/B _7838_/B VGND VPWR _8272_/A VGND VPWR sky130_fd_sc_hd__or3_4
X_7752_ _8379_/B VGND VPWR _8394_/B VGND VPWR sky130_fd_sc_hd__inv_2
X_4964_ _9048_/Q _4964_/B _9051_/Q VGND VPWR _4965_/A VGND VPWR sky130_fd_sc_hd__or3_1
XFILLER_36_298 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6703_ _6698_/Y _6251_/A _6699_/Y _4577_/B _6702_/X VGND VPWR _6716_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_4
XFILLER_177_443 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_123 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7683_ _6464_/Y _7419_/X _6341_/Y _7421_/X VGND VPWR _7683_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4895_ _4887_/Y _4590_/B _4888_/Y _5298_/B _4894_/X VGND VPWR _4896_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9422_ _9684_/CLK _9422_/D _9685_/SET_B VGND VPWR _9422_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6634_ _9266_/Q VGND VPWR _6634_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_6565_ _8783_/A _6027_/B _6564_/Y _4861_/X VGND VPWR _6565_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_9353_ _9378_/CLK _9353_/D _9646_/SET_B VGND VPWR _9353_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_5516_ _9365_/Q _5509_/A _8930_/A1 _5509_/Y VGND VPWR _9365_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8304_ _8451_/A _8642_/B VGND VPWR _8304_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
X_9284_ _9358_/CLK _9284_/D _9528_/SET_B VGND VPWR _9284_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6496_ _9128_/Q VGND VPWR _7701_/A VGND VPWR sky130_fd_sc_hd__clkinv_4
XFILLER_160_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_384 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5447_ _9413_/Q _5444_/A _5965_/B1 _5444_/Y VGND VPWR _9413_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8235_ _8510_/A _8239_/B VGND VPWR _8236_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_160_387 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_207 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5378_ _9461_/Q _5376_/A _8842_/X _5376_/Y VGND VPWR _9461_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8166_ _8168_/A _8640_/B VGND VPWR _8715_/A VGND VPWR sky130_fd_sc_hd__nor2_1
X_7117_ _9246_/Q _9245_/Q _7127_/B _7127_/C VGND VPWR _7118_/A VGND VPWR sky130_fd_sc_hd__or4_1
X_8097_ _8170_/A _8097_/B VGND VPWR _8098_/B VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_59_368 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_36 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7048_ _7392_/B _7048_/B _7048_/C _7048_/D VGND VPWR _7078_/A VGND VPWR sky130_fd_sc_hd__and4_1
X_8999_ _9567_/Q _8775_/A VGND VPWR mgmt_gpio_out[22] VGND VPWR sky130_fd_sc_hd__ebufn_8
XFILLER_70_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_118 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_61 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_98 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_292 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_327 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_91 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4680_ _5178_/B VGND VPWR _4680_/Y VGND VPWR sky130_fd_sc_hd__inv_4
XFILLER_146_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_284 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6350_ _6348_/Y _5404_/B _6349_/Y _5278_/B VGND VPWR _6350_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_154_170 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5301_ _9514_/Q _5300_/A _5963_/B1 _5300_/Y VGND VPWR _9514_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_115_535 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6281_ _8801_/A VGND VPWR _6281_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_69_611 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_8020_ _8401_/A _8389_/A _8097_/B _8401_/A _8019_/X VGND VPWR _8020_/X VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_5232_ _5259_/A _5232_/B VGND VPWR _5233_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_124_19 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5163_ _9605_/Q _5158_/A _8842_/X _5158_/Y VGND VPWR _9605_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_96_441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5094_ _9651_/Q _5091_/A _8844_/X _5091_/Y VGND VPWR _9651_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_56_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8922_ _9604_/Q _8841_/X _8926_/S VGND VPWR _8922_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_64_360 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_8853_ _8852_/X _9165_/Q _9054_/Q VGND VPWR _8853_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_7804_ _8379_/C _8394_/A _8379_/B VGND VPWR _8632_/A VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_24_213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_566 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_219 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_208 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5996_ _9089_/Q _5995_/A _8907_/X _5995_/Y VGND VPWR _9089_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8784_ _8784_/A VGND VPWR _8784_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_7735_ _9067_/Q _5058_/X _7733_/X _7734_/X VGND VPWR _7735_/X VGND VPWR sky130_fd_sc_hd__a211o_1
X_4947_ _4994_/A VGND VPWR _4948_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_4878_ _6158_/B _4931_/B VGND VPWR _5496_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_7666_ _6581_/Y _7415_/X _6539_/Y _7417_/X _7665_/X VGND VPWR _7680_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_177_273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6617_ _9630_/Q VGND VPWR _6617_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9405_ _9758_/CLK _9405_/D _7011_/B VGND VPWR _9405_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_192_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7597_ _6123_/Y _7430_/X _6083_/Y _7432_/X _7596_/X VGND VPWR _7597_/X VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9336_ _9532_/CLK _9336_/D _9647_/SET_B VGND VPWR _9336_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_118_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6548_ _6543_/Y _5374_/B _6544_/Y _5110_/B _6547_/X VGND VPWR _6567_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_6479_ _9123_/Q VGND VPWR _6479_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_106_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9267_ _9354_/CLK _9267_/D _9685_/SET_B VGND VPWR _9267_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_106_568 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8218_ _8218_/A _8218_/B _8218_/C VGND VPWR _8279_/C VGND VPWR sky130_fd_sc_hd__or3_2
X_9198_ _9440_/CLK _9198_/D _4628_/A VGND VPWR _9198_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
Xoutput271 _9726_/Q VGND VPWR pll_sel[0] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput260 _9729_/Q VGND VPWR pll90_sel[0] VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_160_184 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_538 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8149_ _8164_/A _8552_/A VGND VPWR _8685_/B VGND VPWR sky130_fd_sc_hd__nor2_1
Xoutput293 _9735_/Q VGND VPWR pll_trim[3] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput282 _9749_/Q VGND VPWR pll_trim[17] VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_87_496 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_40 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_232 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_463 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_316 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_596 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5850_ _9176_/Q _8924_/X _8873_/X _5849_/X VGND VPWR _9176_/D VGND VPWR sky130_fd_sc_hd__o22a_2
X_4801_ _8936_/X _8938_/X _4801_/C VGND VPWR _4802_/A VGND VPWR sky130_fd_sc_hd__or3_1
X_5781_ _9223_/Q _5778_/A _8844_/X _5778_/Y VGND VPWR _9223_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_9_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4732_ _9286_/Q VGND VPWR _4732_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7520_ _8775_/A _7408_/X _7705_/A _7410_/X _7519_/X VGND VPWR _7536_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_174_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_284 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4663_ _4891_/A _4780_/B VGND VPWR _5556_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_7451_ _7451_/A VGND VPWR _7451_/X VGND VPWR sky130_fd_sc_hd__buf_8
XFILLER_147_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_19 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6402_ _9550_/Q VGND VPWR _6402_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_4594_ _9738_/Q _4592_/A _8845_/X _4592_/Y VGND VPWR _9738_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7382_ _6399_/Y _7095_/X _6374_/Y _7068_/D _7381_/X VGND VPWR _7387_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_6333_ _6328_/Y _5458_/B _6329_/Y _5306_/B _6332_/X VGND VPWR _6352_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9121_ _9655_/CLK _9121_/D _9779_/SET_B VGND VPWR _9121_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_9052_ _9709_/CLK _9052_/D _6043_/X VGND VPWR _9052_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6264_ _9421_/Q VGND VPWR _6264_/Y VGND VPWR sky130_fd_sc_hd__inv_6
XFILLER_142_184 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8003_ _8009_/A VGND VPWR _8003_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_5215_ _9048_/Q _7008_/A VGND VPWR _5215_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
X_6195_ _9474_/Q VGND VPWR _6195_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_5146_ _5146_/A VGND VPWR _5147_/A VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_28_49 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5077_ _5077_/A VGND VPWR _9660_/D VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_84_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_8905_ _9612_/Q _8955_/A1 _8930_/S VGND VPWR _8905_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_37_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_59 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8836_ input84/X _4629_/C _9626_/Q VGND VPWR _8836_/X VGND VPWR sky130_fd_sc_hd__mux2_2
X_5979_ _6040_/A VGND VPWR _5980_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_8767_ _8767_/A VGND VPWR _8768_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_8_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7718_ _7718_/A VGND VPWR _7719_/B VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_178_582 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8698_ _8698_/A _8708_/A _7931_/A VGND VPWR _8699_/B VGND VPWR sky130_fd_sc_hd__or3b_1
X_7649_ _6712_/Y _7427_/X _6632_/Y _5699_/X VGND VPWR _7649_/X VGND VPWR sky130_fd_sc_hd__o22a_2
XFILLER_153_427 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_52 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_23 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9319_ _9344_/CLK _9319_/D _9295_/SET_B VGND VPWR _9319_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_106_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_582 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_33 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_66 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_360 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_499 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_190 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_160 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_468 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_596 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_107 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_460 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_151 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_508 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5000_ _5000_/A VGND VPWR _5000_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_22_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_390 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_488 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6951_ _6951_/A VGND VPWR _6952_/A VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_34_330 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5902_ _9135_/Q _5899_/A _8841_/X _5899_/Y VGND VPWR _9135_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_6882_ _6879_/Y _5797_/B _7150_/A _5610_/B _6881_/Y VGND VPWR _6901_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9670_ _9674_/CLK _9670_/D _9633_/SET_B VGND VPWR _9670_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_34_385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_8621_ _8713_/D VGND VPWR _8621_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_5833_ _9188_/Q _5831_/A _5964_/B1 _5831_/Y VGND VPWR _9188_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_61_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8552_ _8552_/A _8554_/B VGND VPWR _8630_/D VGND VPWR sky130_fd_sc_hd__nor2_1
X_7503_ _6667_/Y _7419_/X _6692_/Y _7421_/X VGND VPWR _7503_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_5764_ _9234_/Q _5759_/A _8929_/A1 _5759_/Y VGND VPWR _9234_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_5695_ _9254_/Q _9253_/Q VGND VPWR _7456_/A VGND VPWR sky130_fd_sc_hd__or2_4
X_4715_ _4706_/Y _5671_/B _4708_/Y _5776_/B _4714_/X VGND VPWR _4791_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_8483_ _8483_/A _8605_/A VGND VPWR _8485_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_30_580 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_118 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4646_ _9715_/Q _4636_/A _8950_/X _4636_/Y VGND VPWR _9715_/D VGND VPWR sky130_fd_sc_hd__a22o_2
X_7434_ _7434_/A VGND VPWR _7434_/X VGND VPWR sky130_fd_sc_hd__buf_6
XFILLER_190_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_7365_ _7365_/A _7365_/B _7365_/C _7365_/D VGND VPWR _7375_/B VGND VPWR sky130_fd_sc_hd__and4_1
X_4577_ _5960_/A _4577_/B VGND VPWR _4578_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_190_577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_9104_ _9775_/CLK _9104_/D _7011_/B VGND VPWR _9104_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6316_ _9274_/Q VGND VPWR _6316_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_143_493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_471 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7296_ _4749_/Y _7059_/B _4890_/Y _7068_/C _7295_/X VGND VPWR _7299_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_2
X_6247_ _6245_/Y _4822_/X _6246_/Y _5393_/B VGND VPWR _6247_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_9035_ _9039_/CLK _9035_/D VGND VPWR _9035_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_6178_ _9262_/Q VGND VPWR _6178_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_57_444 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5129_ _6040_/A VGND VPWR _5130_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_55_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8819_ _9239_/Q _9772_/Q _9787_/Q VGND VPWR _8819_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_9_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_24 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_256 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_599 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_484 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_71 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_436 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_127 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_132 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_380 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_327 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4500_ _9779_/Q _4493_/A _8930_/A1 _4493_/Y VGND VPWR _9779_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_5480_ _5671_/A _5480_/B VGND VPWR _5481_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_172_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_52 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_1 wb_clk_i VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_7150_ _7150_/A _7392_/B VGND VPWR _7150_/X VGND VPWR sky130_fd_sc_hd__or2_1
X_6101_ _6099_/Y _4893_/X _6100_/Y _4841_/X VGND VPWR _6101_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_7081_ _7098_/C _7127_/A _7127_/C VGND VPWR _7082_/A VGND VPWR sky130_fd_sc_hd__or3_1
XFILLER_112_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6032_ _9075_/Q _6029_/A _8844_/X _6029_/Y VGND VPWR _9075_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_79_580 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_19 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_499 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7983_ _8097_/B VGND VPWR _8544_/A VGND VPWR sky130_fd_sc_hd__clkinv_4
XPHY_28 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_190 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_9722_ _9769_/CLK _9722_/D _7011_/B VGND VPWR _9722_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_6934_ _9282_/Q VGND VPWR _7326_/A VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_41_108 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_9653_ _9653_/CLK _9653_/D _9646_/SET_B VGND VPWR _9653_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6865_ _9477_/Q VGND VPWR _6865_/Y VGND VPWR sky130_fd_sc_hd__inv_4
X_8604_ _8604_/A VGND VPWR _8604_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_6796_ _9749_/Q VGND VPWR _6796_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_5816_ _9199_/Q _5812_/A _5966_/B1 _5812_/Y VGND VPWR _9199_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_9584_ _9674_/CLK _9584_/D _9633_/SET_B VGND VPWR _9584_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_10_528 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5747_ _9242_/Q _5744_/A _8841_/X _5744_/Y VGND VPWR _9242_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8535_ _8535_/A _8668_/C _8615_/D _8699_/A VGND VPWR _8541_/A VGND VPWR sky130_fd_sc_hd__or4_2
XFILLER_148_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_49 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8466_ _8466_/A _8615_/C VGND VPWR _8470_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_163_544 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5678_ _9264_/Q _5673_/A _8839_/X _5673_/Y VGND VPWR _9264_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7417_ _7417_/A VGND VPWR _7417_/X VGND VPWR sky130_fd_sc_hd__buf_6
XFILLER_123_419 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_8397_ _8397_/A _8397_/B VGND VPWR _8397_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
X_4629_ _9789_/Q _9096_/Q _4629_/C VGND VPWR _7022_/B VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_104_622 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_26 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7348_ _7348_/A _7392_/B VGND VPWR _7348_/X VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_131_430 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7279_ _6065_/Y _7040_/D _6098_/Y _7110_/X _7278_/X VGND VPWR _7286_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_103_143 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9018_ _9039_/CLK _9018_/D VGND VPWR _9018_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_66_68 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_252 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_274 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_74 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_23 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_67 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_174 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_360 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_574 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_408 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xinput160 wb_adr_i[7] VGND VPWR _8528_/A VGND VPWR sky130_fd_sc_hd__buf_6
Xinput171 wb_dat_i[16] VGND VPWR _7736_/B VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput193 wb_dat_i[7] VGND VPWR _8968_/A1 VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput182 wb_dat_i[26] VGND VPWR _7741_/A2 VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_36_458 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4980_ _4994_/A VGND VPWR _4981_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_6650_ _9072_/Q VGND VPWR _6650_/Y VGND VPWR sky130_fd_sc_hd__inv_4
XFILLER_149_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6581_ _9215_/Q VGND VPWR _6581_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_5601_ _9307_/Q _5596_/A _8839_/X _5596_/Y VGND VPWR _9307_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_176_168 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_8320_ _8320_/A VGND VPWR _8461_/A VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_157_360 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5532_ _9355_/Q _5528_/A _5966_/B1 _5528_/Y VGND VPWR _9355_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_5463_ _9403_/Q _5460_/A _8844_/X _5460_/Y VGND VPWR _9403_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8251_ _8251_/A _8597_/B VGND VPWR _8253_/A VGND VPWR sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_9_csclk clkbuf_2_2_0_csclk/X VGND VPWR _9687_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_99_620 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8182_ _8433_/B _8182_/B VGND VPWR _8184_/A VGND VPWR sky130_fd_sc_hd__nor2_1
X_7202_ _6427_/Y _7082_/X _6390_/Y _7084_/X _7201_/X VGND VPWR _7221_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_2
X_5394_ _5394_/A VGND VPWR _5395_/A VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_132_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_7133_ _7133_/A VGND VPWR _7133_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_113_463 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7064_ _7075_/A _7109_/B VGND VPWR _7065_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_67_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6015_ _6040_/A VGND VPWR _6016_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_82_520 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_594 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_222 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_564 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_428 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7966_ _7966_/A _7966_/B _7966_/C VGND VPWR _8102_/B VGND VPWR sky130_fd_sc_hd__or3_1
X_9705_ _4446_/A1 _9705_/D _4972_/X VGND VPWR _9705_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_7897_ _7897_/A VGND VPWR _8008_/C VGND VPWR sky130_fd_sc_hd__inv_2
X_6917_ _6915_/Y _5507_/B _6916_/Y _5545_/B VGND VPWR _6917_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_167_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_9636_ _9639_/CLK _9636_/D _9633_/SET_B VGND VPWR _9636_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6848_ _9511_/Q VGND VPWR _6848_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_168_48 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9567_ _9617_/CLK _9567_/D _9295_/SET_B VGND VPWR _9567_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_183_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6779_ _9517_/Q VGND VPWR _6779_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_8518_ _8518_/A _8518_/B VGND VPWR _8518_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_9498_ _9534_/CLK _9498_/D _9647_/SET_B VGND VPWR _9498_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_8449_ _8449_/A _8449_/B VGND VPWR _8453_/B VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_123_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_216 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_463 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_174 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_73 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_210 input83/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_45_299 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_371 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_6 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_290 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_271 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_188 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7820_ _8660_/B VGND VPWR _8282_/B VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_91_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7751_ _9068_/Q _7751_/A2 _9067_/Q _7751_/B2 _7750_/X VGND VPWR _7751_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_4963_ _4963_/A VGND VPWR _4963_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_7682_ _6424_/Y _7400_/X _6362_/Y _7405_/X _7681_/X VGND VPWR _7698_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_6702_ _6700_/Y _5480_/B _6701_/Y _5564_/B VGND VPWR _6702_/X VGND VPWR sky130_fd_sc_hd__o22a_2
XFILLER_51_269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_455 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_4894_ _4890_/Y _5450_/B _4892_/Y _4893_/X VGND VPWR _4894_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_9421_ _9684_/CLK _9421_/D _9528_/SET_B VGND VPWR _9421_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_6633_ _9271_/Q VGND VPWR _6633_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_22_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_403 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_436 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6564_ _6564_/A VGND VPWR _6564_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9352_ _9352_/CLK _9352_/D _9646_/SET_B VGND VPWR _9352_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6495_ _9284_/Q VGND VPWR _7370_/A VGND VPWR sky130_fd_sc_hd__inv_2
X_8303_ _8303_/A VGND VPWR _8451_/A VGND VPWR sky130_fd_sc_hd__inv_2
X_5515_ _9366_/Q _5509_/A _8955_/A1 _5509_/Y VGND VPWR _9366_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_9283_ _9687_/CLK _9283_/D _9528_/SET_B VGND VPWR _9283_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_5446_ _9414_/Q _5444_/A _5964_/B1 _5444_/Y VGND VPWR _9414_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8234_ _8238_/A _8264_/B VGND VPWR _8642_/B VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_160_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_219 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5377_ _9462_/Q _5376_/A _8843_/X _5376_/Y VGND VPWR _9462_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8165_ _8165_/A _8708_/D VGND VPWR _8167_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_160_399 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8096_ _8096_/A _8096_/B VGND VPWR _8170_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_7116_ _7116_/A VGND VPWR _7116_/X VGND VPWR sky130_fd_sc_hd__buf_8
X_7047_ _7047_/A VGND VPWR _7048_/D VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_47_48 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_8998_ _9566_/Q _8773_/A VGND VPWR mgmt_gpio_out[21] VGND VPWR sky130_fd_sc_hd__ebufn_8
XFILLER_70_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7949_ _8188_/B _8378_/B VGND VPWR _8185_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_187_208 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_567 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_319 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_9619_ _9674_/CLK _9619_/D _9633_/SET_B VGND VPWR _9619_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_183_425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_73 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_536 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_77 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_260 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_580 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_61 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_512 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_296 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5300_ _5300_/A VGND VPWR _5300_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_5_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_547 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6280_ _6280_/A _6280_/B _6280_/C _6280_/D VGND VPWR _6326_/B VGND VPWR sky130_fd_sc_hd__and4_2
XFILLER_142_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5231_ _5231_/A VGND VPWR _9559_/D VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_123_580 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5162_ _9606_/Q _5158_/A _8925_/A1 _5158_/Y VGND VPWR _9606_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_110_241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5093_ _9652_/Q _5091_/A _8845_/X _5091_/Y VGND VPWR _9652_/D VGND VPWR sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_12_csclk clkbuf_2_2_0_csclk/X VGND VPWR _9535_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_56_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_8921_ _9607_/Q _8844_/X _8926_/S VGND VPWR _8921_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_83_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_18 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_19 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_8852_ _7518_/Y _9634_/Q _8978_/S VGND VPWR _8852_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_27_csclk clkbuf_2_3_0_csclk/X VGND VPWR _9352_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_83_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7803_ _8188_/B _8624_/B VGND VPWR _8562_/A VGND VPWR sky130_fd_sc_hd__nor2_1
X_8783_ _8783_/A VGND VPWR _8784_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XPHY_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5995_ _5995_/A VGND VPWR _5995_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7734_ _7734_/A _7734_/B _9068_/Q VGND VPWR _7734_/X VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_52_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4946_ _9710_/Q _9696_/Q _9050_/Q _5993_/B VGND VPWR _9710_/D VGND VPWR sky130_fd_sc_hd__o211a_1
X_4877_ _9372_/Q VGND VPWR _4877_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7665_ _6533_/Y _7419_/X _6609_/Y _7421_/X VGND VPWR _7665_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_192_211 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7596_ _6109_/Y _7434_/X _6110_/Y _7436_/X VGND VPWR _7596_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_9404_ _9758_/CLK _9404_/D _7011_/B VGND VPWR _9404_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_6616_ _9445_/Q VGND VPWR _8793_/A VGND VPWR sky130_fd_sc_hd__clkinv_8
XFILLER_153_609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_9335_ _9535_/CLK _9335_/D _9528_/SET_B VGND VPWR _9335_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6547_ _6545_/Y _4613_/B _6546_/Y _4577_/B VGND VPWR _6547_/X VGND VPWR sky130_fd_sc_hd__o22a_2
XFILLER_3_107 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_9266_ _9354_/CLK _9266_/D _9685_/SET_B VGND VPWR _9266_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6478_ _9259_/Q VGND VPWR _8757_/A VGND VPWR sky130_fd_sc_hd__inv_6
XFILLER_160_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5429_ _9425_/Q _5422_/A _8930_/A1 _5422_/Y VGND VPWR _9425_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8217_ _8341_/A _8341_/B _8009_/A _8215_/X _8216_/X VGND VPWR _8217_/Y VGND VPWR
+ sky130_fd_sc_hd__o2111ai_1
X_9197_ _9653_/CLK _9197_/D _9646_/SET_B VGND VPWR _9197_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
Xoutput261 _9730_/Q VGND VPWR pll90_sel[1] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput250 _8837_/X VGND VPWR pad_flash_clk VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_8148_ _8148_/A _8577_/A VGND VPWR _8150_/A VGND VPWR sky130_fd_sc_hd__or2_1
Xoutput272 _9727_/Q VGND VPWR pll_sel[1] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput294 _9736_/Q VGND VPWR pll_trim[4] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput283 _9750_/Q VGND VPWR pll_trim[18] VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_181_48 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_8079_ _8379_/D _8394_/B _8079_/C VGND VPWR _8080_/A VGND VPWR sky130_fd_sc_hd__or3_1
XFILLER_114_64 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_564 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_52 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_23 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_50 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_244 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_72 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_1_wb_clk_i clkbuf_1_1_1_wb_clk_i/A VGND VPWR clkbuf_2_3_0_wb_clk_i/A VGND
+ VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_48_80 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_91 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_6 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_372 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4800_ _9515_/Q VGND VPWR _4800_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_34_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5780_ _9224_/Q _5778_/A _8845_/X _5778_/Y VGND VPWR _9224_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_187_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4731_ _4731_/A _5742_/B VGND VPWR _4731_/X VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_147_425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_296 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7450_ _7474_/C _7466_/A _9255_/Q VGND VPWR _7451_/A VGND VPWR sky130_fd_sc_hd__or3_1
X_4662_ _4662_/A VGND VPWR _4780_/B VGND VPWR sky130_fd_sc_hd__buf_8
XFILLER_174_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6401_ _6396_/Y _5344_/B _6397_/Y _5298_/B _6400_/X VGND VPWR _6408_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_174_288 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7381_ _6347_/Y _7097_/X _6340_/Y _7099_/X VGND VPWR _7381_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4593_ _9739_/Q _4592_/A _8846_/X _4592_/Y VGND VPWR _9739_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_9120_ _9655_/CLK _9120_/D _7011_/B VGND VPWR _9120_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_127_182 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6332_ _6330_/Y _5290_/B _6331_/Y _5916_/B VGND VPWR _6332_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_135_19 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9051_ _8837_/A1 _9051_/D _6045_/X VGND VPWR _9051_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_6263_ _9551_/Q VGND VPWR _6263_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
XFILLER_88_217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5214_ _5214_/A _5985_/B VGND VPWR _5214_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
X_8002_ _8394_/D _8077_/A VGND VPWR _8009_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_6194_ _9183_/Q VGND VPWR _6194_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_111_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5145_ _6134_/A _5156_/B VGND VPWR _5146_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_5076_ _8962_/X _9660_/Q _5078_/S VGND VPWR _5077_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_8904_ _9624_/Q _8845_/X _8955_/S VGND VPWR _8904_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_44_16 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_8835_ _6582_/Y input92/X _8835_/S VGND VPWR _8835_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_5978_ _9093_/Q _5970_/A _8839_/X _5970_/Y VGND VPWR _9093_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8766_ _8766_/A VGND VPWR _8766_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_100_33 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7717_ _9086_/Q _7716_/B _7718_/A VGND VPWR _7717_/X VGND VPWR sky130_fd_sc_hd__o21a_1
X_4929_ _4929_/A _4931_/B VGND VPWR _5458_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_8697_ _8697_/A VGND VPWR _8697_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_7648_ _6640_/Y _7415_/X _6772_/Y _7417_/X _7647_/X VGND VPWR _7662_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_100_99 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_288 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7579_ _6224_/Y _7430_/X _6199_/Y _7432_/X _7578_/X VGND VPWR _7579_/X VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_118_182 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_171 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_439 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9318_ _9508_/CLK _9318_/D _9295_/SET_B VGND VPWR _9318_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_161_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_35 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9249_ _9278_/CLK _9249_/D _9633_/SET_B VGND VPWR _9249_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_106_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_79 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_78 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_523 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_320 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_542 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_210 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_119 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_247 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6950_ _6974_/B _6950_/B VGND VPWR _6951_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_5901_ _9136_/Q _5899_/A _8842_/X _5899_/Y VGND VPWR _9136_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_46_180 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_342 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6881_ input47/X _8955_/S input53/X _6322_/Y VGND VPWR _6881_/Y VGND VPWR sky130_fd_sc_hd__a22oi_1
XFILLER_61_161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5832_ _9189_/Q _5831_/A _5963_/B1 _5831_/Y VGND VPWR _9189_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8620_ _8706_/A _8705_/B _8703_/B _8620_/D VGND VPWR _8620_/Y VGND VPWR sky130_fd_sc_hd__nor4_1
X_5763_ _9235_/Q _5759_/A _8925_/A1 _5759_/Y VGND VPWR _9235_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8551_ _8551_/A _8554_/B VGND VPWR _8686_/C VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_14_19 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_211 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4714_ _7304_/A _5632_/B _4712_/Y _5789_/B VGND VPWR _4714_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_7502_ _6724_/Y _7400_/X _6664_/Y _7405_/X _7501_/X VGND VPWR _7518_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_108_609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_8482_ _8562_/A _8650_/B VGND VPWR _8605_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_5694_ _5694_/A VGND VPWR _7462_/A VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_147_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7433_ _7462_/A _7474_/C _7474_/D VGND VPWR _7434_/A VGND VPWR sky130_fd_sc_hd__or3_1
X_4645_ _4645_/A VGND VPWR _4645_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_30_18 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4576_ _6158_/A _4876_/B VGND VPWR _4577_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_7364_ _6498_/Y _7048_/D _6551_/Y _7040_/B _7363_/X VGND VPWR _7365_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_190_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9103_ _9777_/CLK _9103_/D _9633_/SET_B VGND VPWR _9103_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6315_ _9111_/Q VGND VPWR _6315_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_143_483 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7295_ _4902_/Y _7079_/B _4706_/Y _7059_/A VGND VPWR _7295_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_9034_ _9664_/CLK _9034_/D VGND VPWR _9034_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_130_144 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6246_ _9447_/Q VGND VPWR _6246_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_6177_ _6175_/Y _5818_/B _6176_/Y _5572_/B VGND VPWR _6187_/A VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_29_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5128_ _9627_/Q _5123_/A _5967_/B1 _5123_/Y VGND VPWR _9627_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_84_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_478 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_106 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5059_ _7734_/A _5059_/B VGND VPWR _5060_/A VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_111_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8818_ _8818_/A VGND VPWR _8818_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_158_509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_36 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8749_ _8749_/A VGND VPWR _8750_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_138_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_268 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_463 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_267 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_150 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_386 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_370 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_350 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_2 _8977_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_6_64 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6100_ _6100_/A VGND VPWR _6100_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_152_280 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7080_ _7080_/A VGND VPWR _8959_/S VGND VPWR sky130_fd_sc_hd__buf_6
XFILLER_140_486 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6031_ _9076_/Q _6029_/A _8845_/X _6029_/Y VGND VPWR _9076_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_66_220 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7982_ _7982_/A VGND VPWR _8552_/A VGND VPWR sky130_fd_sc_hd__clkbuf_4
XPHY_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6933_ _9191_/Q VGND VPWR _6933_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9721_ _9769_/CLK _9721_/D _9757_/SET_B VGND VPWR _9721_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_22_301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6864_ _6859_/Y _5496_/B _6860_/Y _5240_/B _6863_/X VGND VPWR _6877_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9652_ _9652_/CLK _9652_/D _9647_/SET_B VGND VPWR _9652_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_179_133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5815_ _9200_/Q _5812_/A _8841_/X _5812_/Y VGND VPWR _9200_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8603_ _8603_/A _8603_/B _8603_/C _8603_/D VGND VPWR _8604_/A VGND VPWR sky130_fd_sc_hd__or4_1
X_6795_ _9760_/Q VGND VPWR _6795_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9583_ _9674_/CLK _9583_/D _9633_/SET_B VGND VPWR _9583_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_5746_ _9243_/Q _5744_/A _8842_/X _5744_/Y VGND VPWR _9243_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8534_ _8471_/Y _8523_/Y _8518_/X _8470_/B VGND VPWR _8699_/A VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_175_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_17 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5677_ _9265_/Q _5673_/A _5966_/B1 _5673_/Y VGND VPWR _9265_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8465_ _8305_/A _8270_/B _8097_/B _8552_/A VGND VPWR _8615_/C VGND VPWR sky130_fd_sc_hd__o22ai_1
XFILLER_135_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_4628_ _4628_/A VGND VPWR _6052_/B VGND VPWR sky130_fd_sc_hd__inv_2
X_7416_ _7466_/A _7470_/B _9255_/Q VGND VPWR _7417_/A VGND VPWR sky130_fd_sc_hd__or3_1
XFILLER_163_556 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_8396_ _8396_/A VGND VPWR _8396_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_89_301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7347_ _6731_/Y _7059_/D _6718_/Y _7116_/X _7346_/X VGND VPWR _7352_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_4559_ _5966_/B1 _9757_/Q _4561_/S VGND VPWR _4560_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_173_38 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_442 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7278_ _6141_/Y _7112_/X _6128_/Y _7077_/B VGND VPWR _7278_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_103_155 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_9017_ _9664_/CLK _9017_/D VGND VPWR _9017_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_6229_ _6224_/Y _5905_/B _6225_/Y _5420_/B _6228_/X VGND VPWR _6236_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_66_47 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_20 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_415 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_407 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_79 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_492 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_103 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_186 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_586 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_331 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_94 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_220 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xinput161 wb_adr_i[8] VGND VPWR _7774_/D VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput150 wb_adr_i[27] VGND VPWR _5930_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput172 wb_dat_i[17] VGND VPWR _7738_/B VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput194 wb_dat_i[8] VGND VPWR _7737_/B2 VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput183 wb_dat_i[27] VGND VPWR _7743_/A2 VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_189_442 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5600_ _9308_/Q _5596_/A _8930_/A1 _5596_/Y VGND VPWR _9308_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_6580_ _9691_/Q VGND VPWR _8745_/A VGND VPWR sky130_fd_sc_hd__clkinv_4
XFILLER_164_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5531_ _9356_/Q _5528_/A _8841_/X _5528_/Y VGND VPWR _9356_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8250_ _8250_/A VGND VPWR _8597_/B VGND VPWR sky130_fd_sc_hd__inv_2
X_5462_ _9404_/Q _5460_/A _8845_/X _5460_/Y VGND VPWR _9404_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7201_ _6371_/Y _7077_/C _6461_/Y _7077_/D _7200_/X VGND VPWR _7201_/X VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_132_217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_8181_ _8651_/A _8562_/A _8636_/A _8180_/Y VGND VPWR _8182_/B VGND VPWR sky130_fd_sc_hd__or4b_1
X_5393_ _5545_/A _5393_/B VGND VPWR _5394_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_7132_ _7132_/A _7132_/B _7132_/C VGND VPWR _7133_/A VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_98_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_475 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7063_ _7063_/A VGND VPWR _7068_/B VGND VPWR sky130_fd_sc_hd__buf_8
XFILLER_143_19 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_294 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6014_ _9083_/Q _5995_/A _8900_/X _5995_/Y VGND VPWR _9083_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_39_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_234 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7965_ _8583_/A _8091_/B VGND VPWR _7971_/A VGND VPWR sky130_fd_sc_hd__or2_2
X_9704_ _4446_/A1 _9704_/D _4975_/X VGND VPWR _9704_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_35_470 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6916_ _9339_/Q VGND VPWR _6916_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7896_ _7896_/A _8341_/B VGND VPWR _7896_/X VGND VPWR sky130_fd_sc_hd__or2_1
X_9635_ _9791_/CLK _9635_/D _9633_/SET_B VGND VPWR _9635_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6847_ _6847_/A VGND VPWR _6847_/Y VGND VPWR sky130_fd_sc_hd__inv_4
XFILLER_50_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_7 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6778_ _6778_/A VGND VPWR _6778_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9566_ _9617_/CLK _9566_/D _9295_/SET_B VGND VPWR _9566_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_22_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_348 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8517_ _8517_/A VGND VPWR _8517_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_155_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5729_ _6994_/A _5692_/Y _5724_/Y _5724_/B _5728_/X VGND VPWR _5730_/A VGND VPWR
+ sky130_fd_sc_hd__o32a_1
X_9497_ _9501_/CLK _9497_/D _9647_/SET_B VGND VPWR _9497_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_163_331 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_342 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8448_ _8612_/A _8448_/B _8448_/C _8447_/X VGND VPWR _8449_/B VGND VPWR sky130_fd_sc_hd__or4b_1
XFILLER_136_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8379_ _8202_/A _8379_/B _8379_/C _8379_/D VGND VPWR _8585_/A VGND VPWR sky130_fd_sc_hd__and4b_1
XFILLER_117_31 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_24 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_186 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_404 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_200 input83/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_73_565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_211 input83/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_45_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_180 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_10 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_283 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_540 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_223 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7750_ _9066_/Q _7750_/B VGND VPWR _7750_/X VGND VPWR sky130_fd_sc_hd__and2_1
X_4962_ _4994_/A VGND VPWR _4963_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_32_451 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6701_ _9330_/Q VGND VPWR _6701_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7681_ _6399_/Y _7408_/X _6418_/Y _7410_/X VGND VPWR _7681_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4893_ _6111_/A _4917_/A VGND VPWR _4893_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_9420_ _9684_/CLK _9420_/D _9685_/SET_B VGND VPWR _9420_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6632_ _9309_/Q VGND VPWR _6632_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_149_147 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6563_ _9073_/Q VGND VPWR _8783_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_118_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9351_ _9613_/CLK _9351_/D _9646_/SET_B VGND VPWR _9351_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_8302_ _8498_/B VGND VPWR _8302_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_5514_ _9367_/Q _5509_/A _8929_/A1 _5509_/Y VGND VPWR _9367_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_6494_ _8797_/A _6081_/B _7705_/A _5968_/B _6493_/X VGND VPWR _6501_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_2
X_9282_ _9687_/CLK _9282_/D _9685_/SET_B VGND VPWR _9282_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_118_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8233_ _8233_/A VGND VPWR _8358_/B VGND VPWR sky130_fd_sc_hd__inv_2
X_5445_ _9415_/Q _5444_/A _5963_/B1 _5444_/Y VGND VPWR _9415_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_160_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8164_ _8164_/A _8168_/A VGND VPWR _8708_/D VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_154_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5376_ _5376_/A VGND VPWR _5376_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7115_ _7127_/C _7115_/B VGND VPWR _7116_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_113_272 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8095_ _8521_/A _8437_/B VGND VPWR _8560_/A VGND VPWR sky130_fd_sc_hd__nor2_1
X_7046_ _7125_/A _7127_/B _7073_/C VGND VPWR _7047_/A VGND VPWR sky130_fd_sc_hd__or3_1
X_6039__1 _9709_/CLK VGND VPWR _9058_/CLK VGND VPWR sky130_fd_sc_hd__inv_4
XFILLER_86_178 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8997_ _9565_/Q _8771_/A VGND VPWR mgmt_gpio_out[20] VGND VPWR sky130_fd_sc_hd__ebufn_8
XFILLER_55_598 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7948_ _7948_/A VGND VPWR _8378_/B VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_70_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_579 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7879_ _7879_/A _7879_/B VGND VPWR _7879_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
X_9618_ _9674_/CLK _9618_/D _9633_/SET_B VGND VPWR _9618_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_7_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_9549_ _9639_/CLK _9549_/D _9757_/SET_B VGND VPWR _9549_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_170_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_183 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_89 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_272 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_115 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_95 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_362 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_8_csclk clkbuf_2_2_0_csclk/X VGND VPWR _9358_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_18_278 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_220 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5230_ _5967_/B1 _9559_/Q _5230_/S VGND VPWR _5231_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_102_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5161_ _9607_/Q _5158_/A _8844_/X _5158_/Y VGND VPWR _9607_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_5092_ _9653_/Q _5091_/A _8846_/X _5091_/Y VGND VPWR _9653_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_110_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_264 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8920_ _9622_/Q _8925_/A1 _8955_/S VGND VPWR _8920_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_83_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_148 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8851_ _8850_/X _9164_/Q _9054_/Q VGND VPWR _8851_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_91_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5994_ _9051_/Q _5993_/X _6022_/B VGND VPWR _5995_/A VGND VPWR sky130_fd_sc_hd__o21ai_4
X_5848__4 _8924_/X VGND VPWR _5896_/B1 VGND VPWR sky130_fd_sc_hd__inv_4
X_7802_ _7802_/A VGND VPWR _8624_/B VGND VPWR sky130_fd_sc_hd__buf_6
X_8782_ _8782_/A VGND VPWR _8782_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_52_524 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7733_ _7733_/A _7734_/A _9066_/Q VGND VPWR _7733_/X VGND VPWR sky130_fd_sc_hd__and3_1
X_4945_ _7008_/A VGND VPWR _5993_/B VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_20_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4876_ _6111_/A _4876_/B VGND VPWR _5110_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_7664_ _6555_/Y _7400_/X _6497_/Y _7405_/X _7663_/X VGND VPWR _7680_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_2
XFILLER_20_410 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_223 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7595_ _6072_/Y _7427_/X _6141_/Y _5699_/X VGND VPWR _7595_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_9403_ _9758_/CLK _9403_/D _7011_/B VGND VPWR _9403_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6615_ _9487_/Q VGND VPWR _6615_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
X_6546_ _9743_/Q VGND VPWR _6546_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9334_ _9532_/CLK _9334_/D _9647_/SET_B VGND VPWR _9334_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_192_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9265_ _9789_/CLK _9265_/D _9685_/SET_B VGND VPWR _9265_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6477_ _9229_/Q VGND VPWR _6477_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_5428_ _9426_/Q _5422_/A _8841_/X _5422_/Y VGND VPWR _9426_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8216_ _8510_/A _8341_/B VGND VPWR _8216_/X VGND VPWR sky130_fd_sc_hd__or2_2
X_9196_ _9653_/CLK _9196_/D _9646_/SET_B VGND VPWR _9196_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
Xoutput251 _7011_/Y VGND VPWR pad_flash_clk_oeb VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput262 _9731_/Q VGND VPWR pll90_sel[2] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput240 _8746_/X VGND VPWR mgmt_gpio_oeb[5] VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_99_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5359_ _9474_/Q _5357_/A _8845_/X _5357_/Y VGND VPWR _9474_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8147_ _8213_/A _8551_/A VGND VPWR _8577_/A VGND VPWR sky130_fd_sc_hd__nor2_1
Xoutput273 _9728_/Q VGND VPWR pll_sel[2] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput295 _9737_/Q VGND VPWR pll_trim[5] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput284 _9751_/Q VGND VPWR pll_trim[19] VGND VPWR sky130_fd_sc_hd__buf_2
X_8078_ _8078_/A _8672_/B VGND VPWR _8082_/A VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_101_275 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_264 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7029_ _7073_/C _7123_/B VGND VPWR _7030_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_74_104 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_14 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_76 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_256 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_22 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_11 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_418 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_84 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_470 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_218 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_66 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_384 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_376 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4730_ _4900_/B _4780_/B VGND VPWR _5742_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_159_275 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4661_ _4665_/B _4665_/C _4661_/C VGND VPWR _4662_/A VGND VPWR sky130_fd_sc_hd__or3_1
XFILLER_80_90 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6400_ _6398_/Y _5534_/B _6399_/Y _5366_/B VGND VPWR _6400_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_7380_ _6467_/Y _7048_/B _6416_/Y _7077_/A _7379_/X VGND VPWR _7387_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_4592_ _4592_/A VGND VPWR _4592_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_6331_ _9124_/Q VGND VPWR _6331_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_155_481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_323 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9050_ _8837_/A1 _9050_/D _6047_/X VGND VPWR _9050_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_6262_ _6262_/A VGND VPWR _6262_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_142_175 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6193_ _6193_/A VGND VPWR _6193_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_8001_ _8097_/B _8117_/A VGND VPWR _8612_/A VGND VPWR sky130_fd_sc_hd__nor2_1
X_5213_ _5213_/A VGND VPWR _5213_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_69_443 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5144_ _9618_/Q _5136_/A _8916_/A1 _5136_/Y VGND VPWR _9618_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_5075_ _5075_/A VGND VPWR _9661_/D VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_8903_ _9619_/Q _8930_/A1 _8955_/S VGND VPWR _8903_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_71_118 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8834_ _6485_/Y input90/X _8835_/S VGND VPWR _8834_/X VGND VPWR sky130_fd_sc_hd__mux2_2
XFILLER_64_192 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_387 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5977_ _9094_/Q _5970_/A _8930_/A1 _5970_/Y VGND VPWR _9094_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8765_ _8765_/A VGND VPWR _8766_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_4928_ _9398_/Q VGND VPWR _4928_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_8696_ _8696_/A _8696_/B _8696_/C _8727_/D VGND VPWR _8697_/A VGND VPWR sky130_fd_sc_hd__or4_1
X_7716_ _9086_/Q _7716_/B VGND VPWR _7718_/A VGND VPWR sky130_fd_sc_hd__nand2_1
X_7647_ _6732_/Y _7419_/X _6762_/Y _7421_/X VGND VPWR _7647_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_121_7 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_4859_ _4931_/A _4911_/A VGND VPWR _5374_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_193_565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_7578_ _6171_/Y _7434_/X _6169_/Y _7436_/X VGND VPWR _7578_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_9317_ _9501_/CLK _9317_/D _9647_/SET_B VGND VPWR _9317_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6529_ _9686_/Q VGND VPWR _6529_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
XFILLER_133_131 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_47 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_9248_ _9278_/CLK _9248_/D _9779_/SET_B VGND VPWR _9248_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_192_48 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9179_ _9652_/CLK _9179_/D _9646_/SET_B VGND VPWR _9179_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_87_251 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_402 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_332 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_74 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_11_csclk clkbuf_2_2_0_csclk/X VGND VPWR _9527_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_171_259 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_26_csclk clkbuf_2_3_0_csclk/X VGND VPWR _9613_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_140_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_90 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5900_ _9137_/Q _5899_/A _8843_/X _5899_/Y VGND VPWR _9137_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_81_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6880_ _9295_/Q VGND VPWR _7150_/A VGND VPWR sky130_fd_sc_hd__inv_2
X_5831_ _5831_/A VGND VPWR _5831_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_5762_ _9236_/Q _5759_/A _8844_/X _5759_/Y VGND VPWR _9236_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8550_ _8550_/A _8554_/B VGND VPWR _8627_/D VGND VPWR sky130_fd_sc_hd__nor2_1
X_7501_ _6736_/Y _7408_/X _6673_/Y _7410_/X VGND VPWR _7501_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4713_ _4919_/A _4780_/B VGND VPWR _5789_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_5693_ _9252_/Q _9251_/Q VGND VPWR _5694_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_8481_ _8481_/A _8706_/A VGND VPWR _8483_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_7432_ _7432_/A VGND VPWR _7432_/X VGND VPWR sky130_fd_sc_hd__buf_6
X_4644_ _4994_/A VGND VPWR _4645_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_7363_ _6581_/Y _7068_/A _6597_/Y _7105_/X VGND VPWR _7363_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4575_ _4669_/A _4729_/D _4729_/A _8944_/X VGND VPWR _4876_/B VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_89_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6314_ _9651_/Q VGND VPWR _6314_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7294_ _4924_/Y _7095_/X _4722_/Y _7068_/D _7293_/X VGND VPWR _7299_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9102_ _9775_/CLK _9102_/D _7011_/B VGND VPWR _9102_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_9033_ _9664_/CLK _9033_/D VGND VPWR _9033_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_6245_ _6245_/A VGND VPWR _6245_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_103_326 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6176_ _9326_/Q VGND VPWR _6176_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_5127_ _9628_/Q _5123_/A _5966_/B1 _5123_/Y VGND VPWR _9628_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_5058_ _7734_/A _5058_/B VGND VPWR _5058_/X VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_84_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_118 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_298 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_471 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_33 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8817_ _8817_/A VGND VPWR _8817_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_80_493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8748_ _8748_/A VGND VPWR _8748_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_71_48 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_8679_ _8721_/A _8720_/C _8721_/C _8723_/C VGND VPWR _8680_/C VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_138_245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_131 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_442 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_232 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_276 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_279 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_2_0_mgmt_gpio_in[4] clkbuf_2_3_0_mgmt_gpio_in[4]/A VGND VPWR _9089_/CLK
+ VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_43_162 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_360 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_368 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_382 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_371 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_582 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_542 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_3 _8930_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_172_568 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_76 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_80 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_292 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6030_ _9077_/Q _6029_/A _8846_/X _6029_/Y VGND VPWR _9077_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_140_498 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_232 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7981_ _7995_/B _7992_/B VGND VPWR _7982_/A VGND VPWR sky130_fd_sc_hd__or2_1
XPHY_19 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6932_ _9213_/Q VGND VPWR _6932_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9720_ _9770_/CLK _9720_/D _7011_/B VGND VPWR _9720_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6863_ _6861_/Y _4577_/B _8808_/A _5227_/B VGND VPWR _6863_/X VGND VPWR sky130_fd_sc_hd__o22a_2
X_9651_ _9653_/CLK _9651_/D _9646_/SET_B VGND VPWR _9651_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_179_145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5814_ _9201_/Q _5812_/A _5964_/B1 _5812_/Y VGND VPWR _9201_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8602_ _8202_/A _8341_/A _8660_/C _7881_/A _8334_/X VGND VPWR _8603_/D VGND VPWR
+ sky130_fd_sc_hd__o221ai_1
X_6794_ _6794_/A VGND VPWR _6794_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9582_ _9674_/CLK _9582_/D _9633_/SET_B VGND VPWR _9582_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_5745_ _9244_/Q _5744_/A _8843_/X _5744_/Y VGND VPWR _9244_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8533_ _8516_/Y _8528_/Y _8518_/X _8464_/D VGND VPWR _8615_/D VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_157_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5676_ _9266_/Q _5673_/A _8841_/X _5673_/Y VGND VPWR _9266_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8464_ _8464_/A _8464_/B _8668_/A _8464_/D VGND VPWR _8466_/A VGND VPWR sky130_fd_sc_hd__or4_1
X_7415_ _7415_/A VGND VPWR _7415_/X VGND VPWR sky130_fd_sc_hd__buf_6
X_4627_ _4627_/A VGND VPWR _9719_/D VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_190_354 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_8395_ _8496_/A _8395_/B VGND VPWR _8395_/X VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_190_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7346_ _6779_/Y _7118_/X _6668_/Y _7048_/C VGND VPWR _7346_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4558_ _5259_/A _4558_/B VGND VPWR _4561_/S VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_103_123 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4489_ _8934_/X _8932_/X _8946_/X _8944_/X VGND VPWR _4805_/A VGND VPWR sky130_fd_sc_hd__or4_4
X_7277_ _7277_/A _7277_/B _7277_/C _7277_/D VGND VPWR _7287_/B VGND VPWR sky130_fd_sc_hd__and4_1
X_9016_ _9039_/CLK _9016_/D VGND VPWR _9016_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_6228_ _6226_/Y _4524_/B _6227_/Y _4832_/X VGND VPWR _6228_/X VGND VPWR sky130_fd_sc_hd__o22a_2
X_6159_ _9456_/Q VGND VPWR _6159_/Y VGND VPWR sky130_fd_sc_hd__inv_2
Xrepeater370 _7011_/B VGND VPWR _9779_/SET_B VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_82_14 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_460 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_534 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_272 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_294 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xinput162 wb_adr_i[9] VGND VPWR _7774_/C VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput140 wb_adr_i[18] VGND VPWR _7768_/D VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput151 wb_adr_i[28] VGND VPWR _5930_/B VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput195 wb_dat_i[9] VGND VPWR _7739_/B2 VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput173 wb_dat_i[18] VGND VPWR _7740_/B VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput184 wb_dat_i[28] VGND VPWR _7745_/A2 VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_76_574 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_611 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_190 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_148 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_390 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5530_ _9357_/Q _5528_/A _8842_/X _5528_/Y VGND VPWR _9357_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_5461_ _9405_/Q _5460_/A _8846_/X _5460_/Y VGND VPWR _9405_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_172_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7200_ _6415_/Y _7086_/X _6357_/Y _7088_/X VGND VPWR _7200_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_172_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_516 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5392_ _9450_/Q _5384_/A _8916_/A1 _5384_/Y VGND VPWR _9450_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8180_ _8544_/A _8092_/Y _8179_/X VGND VPWR _8180_/Y VGND VPWR sky130_fd_sc_hd__a21oi_1
XFILLER_125_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7131_ _7131_/A _7131_/B _7131_/C _7131_/D VGND VPWR _7132_/C VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_86_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_7062_ _7075_/A _7087_/B VGND VPWR _7063_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_6013_ _6013_/A VGND VPWR _6013_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_67_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_18 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7964_ _8189_/A _8099_/B _7966_/B VGND VPWR _8091_/B VGND VPWR sky130_fd_sc_hd__a21bo_2
XFILLER_36_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_246 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_9703_ _4446_/A1 _9703_/D _4978_/X VGND VPWR _9703_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6915_ _9365_/Q VGND VPWR _6915_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_35_493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7895_ _7895_/A VGND VPWR _8341_/B VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_50_441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6846_ _6844_/Y _4491_/B _6845_/Y _5259_/B VGND VPWR _6846_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_9634_ _9655_/CLK _9634_/D _9633_/SET_B VGND VPWR _9634_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_9565_ _9617_/CLK _9565_/D _9295_/SET_B VGND VPWR _9565_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_6777_ _6772_/Y _5941_/B _6773_/Y _5089_/B _6776_/X VGND VPWR _6783_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_8516_ _8525_/C _8516_/B VGND VPWR _8516_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
X_5728_ _5728_/A VGND VPWR _5728_/X VGND VPWR sky130_fd_sc_hd__buf_8
XFILLER_6_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9496_ _9532_/CLK _9496_/D _9647_/SET_B VGND VPWR _9496_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_108_248 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5659_ _5647_/A _5651_/A _9277_/Q _5659_/B2 _5651_/X VGND VPWR _9277_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_2
X_8447_ _8496_/A _8447_/B VGND VPWR _8447_/X VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_163_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8378_ _8565_/A _8378_/B VGND VPWR _8720_/C VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_117_43 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7329_ _6872_/Y _7124_/X _6885_/Y _7068_/B _7328_/X VGND VPWR _7330_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_131_251 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_36 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_198 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_416 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA_201 input83/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_212 _6135_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_26_460 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_103 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_72 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_192 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_207 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_338 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_295 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_552 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_246 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4961_ _9092_/Q _9048_/Q _4949_/A _4958_/Y _4960_/X VGND VPWR _9708_/D VGND VPWR
+ sky130_fd_sc_hd__a41o_1
X_4892_ _4892_/A VGND VPWR _4892_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_6700_ _9387_/Q VGND VPWR _6700_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7680_ _7680_/A _7680_/B _7680_/C _7680_/D VGND VPWR _7680_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
XFILLER_32_463 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6631_ _9296_/Q VGND VPWR _7172_/A VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_149_159 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9350_ _9352_/CLK _9350_/D _9646_/SET_B VGND VPWR _9350_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6562_ _9471_/Q VGND VPWR _8791_/A VGND VPWR sky130_fd_sc_hd__inv_12
X_8301_ _8301_/A VGND VPWR _8498_/B VGND VPWR sky130_fd_sc_hd__buf_6
X_5513_ _9368_/Q _5509_/A _8925_/A1 _5509_/Y VGND VPWR _9368_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_6493_ _6491_/Y _5545_/B _8751_/A _5797_/B VGND VPWR _6493_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_9281_ _9687_/CLK _9281_/D _9528_/SET_B VGND VPWR _9281_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_133_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5444_ _5444_/A VGND VPWR _5444_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_8232_ _8341_/A _8232_/B VGND VPWR _8233_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_8163_ _8708_/B _8163_/B VGND VPWR _8165_/A VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_160_357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7114_ _4716_/Y _7040_/D _4804_/Y _7110_/X _7113_/X VGND VPWR _7131_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_5375_ _5375_/A VGND VPWR _5376_/A VGND VPWR sky130_fd_sc_hd__clkbuf_2
X_8094_ _8094_/A VGND VPWR _8720_/A VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_101_435 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7045_ _7045_/A VGND VPWR _7048_/C VGND VPWR sky130_fd_sc_hd__buf_8
XFILLER_170_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_522 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8996_ _9564_/Q _8769_/A VGND VPWR mgmt_gpio_out[19] VGND VPWR sky130_fd_sc_hd__ebufn_8
XFILLER_82_374 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7947_ _8379_/D _8379_/B _8079_/C VGND VPWR _7948_/A VGND VPWR sky130_fd_sc_hd__or3_1
XFILLER_35_290 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7878_ _7878_/A _8341_/A VGND VPWR _7879_/B VGND VPWR sky130_fd_sc_hd__or2_2
X_6829_ _6829_/A _6829_/B _6829_/C _6829_/D VGND VPWR _6830_/D VGND VPWR sky130_fd_sc_hd__and4_1
X_9617_ _9617_/CLK _9617_/D _9295_/SET_B VGND VPWR _9617_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_23_496 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_106 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_524 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9548_ _9639_/CLK _9548_/D _9633_/SET_B VGND VPWR _9548_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_183_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_170 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9479_ _9684_/CLK _9479_/D _9685_/SET_B VGND VPWR _9479_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_12_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_324 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_195 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_284 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_511 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_374 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_427 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_107 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_302 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_508 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5160_ _9608_/Q _5158_/A _8845_/X _5158_/Y VGND VPWR _9608_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_68_135 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5091_ _5091_/A VGND VPWR _5091_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_96_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_276 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_8850_ _7500_/Y _9633_/Q _8978_/S VGND VPWR _8850_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_227 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5993_ _9050_/Q _5993_/B _7008_/B VGND VPWR _5993_/X VGND VPWR sky130_fd_sc_hd__and3_1
X_7801_ _8394_/B _8093_/A VGND VPWR _7802_/A VGND VPWR sky130_fd_sc_hd__or2_1
X_5848__5 _8924_/X VGND VPWR _5894_/A1 VGND VPWR sky130_fd_sc_hd__inv_4
X_8781_ _8781_/A VGND VPWR _8782_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_64_374 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4944_ _4944_/A VGND VPWR _7008_/A VGND VPWR sky130_fd_sc_hd__clkbuf_4
X_7732_ _7732_/A VGND VPWR _8960_/S VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_149_19 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4875_ _9632_/Q VGND VPWR _4875_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7663_ _6589_/Y _7408_/X _6529_/Y _7410_/X VGND VPWR _7663_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_9402_ _9758_/CLK _9402_/D _7011_/B VGND VPWR _9402_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6614_ _6609_/Y _5251_/B _8765_/A _5534_/B _6613_/X VGND VPWR _6627_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_7594_ _6126_/Y _7415_/X _6120_/Y _7417_/X _7593_/X VGND VPWR _7608_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_165_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_246 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_235 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6545_ _9724_/Q VGND VPWR _6545_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9333_ _9535_/CLK _9333_/D _9528_/SET_B VGND VPWR _9333_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_118_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_9264_ _9354_/CLK _9264_/D _9685_/SET_B VGND VPWR _9264_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_133_324 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_162 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6476_ _6149_/A _6475_/Y _9040_/Q _6149_/Y VGND VPWR _9040_/D VGND VPWR sky130_fd_sc_hd__o22a_2
X_8215_ _8660_/A _8498_/A VGND VPWR _8215_/X VGND VPWR sky130_fd_sc_hd__or2_2
XFILLER_160_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5427_ _9427_/Q _5422_/A _8929_/A1 _5422_/Y VGND VPWR _9427_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_9195_ _9653_/CLK _9195_/D _9646_/SET_B VGND VPWR _9195_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
Xoutput252 _8836_/X VGND VPWR pad_flash_csb VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput241 _7702_/X VGND VPWR mgmt_gpio_oeb[6] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput230 _8792_/X VGND VPWR mgmt_gpio_oeb[30] VGND VPWR sky130_fd_sc_hd__buf_2
X_5358_ _9475_/Q _5357_/A _8846_/X _5357_/Y VGND VPWR _9475_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8146_ _7987_/Y _8544_/B _8145_/X VGND VPWR _8148_/A VGND VPWR sky130_fd_sc_hd__a21o_1
Xoutput274 _9732_/Q VGND VPWR pll_trim[0] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput285 _9733_/Q VGND VPWR pll_trim[1] VGND VPWR sky130_fd_sc_hd__buf_2
Xoutput263 _9758_/Q VGND VPWR pll_bypass VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_59_102 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8077_ _8077_/A _8437_/B VGND VPWR _8672_/B VGND VPWR sky130_fd_sc_hd__nor2_1
Xoutput296 _9738_/Q VGND VPWR pll_trim[6] VGND VPWR sky130_fd_sc_hd__buf_2
X_7028_ _7104_/A _7111_/C VGND VPWR _7123_/B VGND VPWR sky130_fd_sc_hd__or2_1
X_5289_ _6052_/A VGND VPWR _5671_/A VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_75_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_599 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_8979_ _9580_/Q _8743_/A VGND VPWR mgmt_gpio_out[2] VGND VPWR sky130_fd_sc_hd__ebufn_8
XFILLER_15_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_608 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_416 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_202 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_268 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_376 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_131 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_9 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_455 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_50 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_396 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xnet299_2 _4446_/A1 VGND VPWR _7022_/A VGND VPWR sky130_fd_sc_hd__inv_4
XFILLER_61_388 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_232 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4660_ _9333_/Q VGND VPWR _4660_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_147_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4591_ _4591_/A VGND VPWR _4592_/A VGND VPWR sky130_fd_sc_hd__buf_2
X_6330_ _9519_/Q VGND VPWR _6330_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_142_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_6261_ _6256_/Y _5355_/B _6257_/Y _4870_/X _6260_/X VGND VPWR _6280_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_130_327 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6192_ _6188_/Y _6027_/B _6189_/Y _4491_/B _6191_/X VGND VPWR _6211_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_8000_ _8000_/A VGND VPWR _8117_/A VGND VPWR sky130_fd_sc_hd__buf_6
X_5212_ _6040_/A VGND VPWR _5213_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_5143_ _9619_/Q _5136_/A _8930_/A1 _5136_/Y VGND VPWR _9619_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_57_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5074_ _8963_/X _9661_/Q _5078_/S VGND VPWR _5075_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_37_330 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8902_ _7708_/Y _4949_/A _9051_/Q VGND VPWR _8902_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_8833_ _6491_/Y input82/X _8833_/S VGND VPWR _8833_/X VGND VPWR sky130_fd_sc_hd__mux2_4
XFILLER_44_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5976_ _9095_/Q _5970_/A _8841_/X _5970_/Y VGND VPWR _9095_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8764_ _8764_/A VGND VPWR _8764_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_178_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8695_ _8695_/A _8695_/B _8695_/C _8695_/D VGND VPWR _8727_/D VGND VPWR sky130_fd_sc_hd__or4_1
X_7715_ _7716_/B _7715_/B VGND VPWR _7715_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
X_4927_ _4927_/A _4931_/B VGND VPWR _5306_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_52_399 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_79 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4858_ _9458_/Q VGND VPWR _4858_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7646_ _6718_/Y _7400_/X _6645_/Y _7405_/X _7645_/X VGND VPWR _7662_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_2
X_7577_ _6200_/Y _7427_/X _6176_/Y _5699_/X VGND VPWR _7577_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_4789_ _4779_/Y _5757_/B _4781_/Y _6322_/A _4788_/X VGND VPWR _4790_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9316_ _9534_/CLK _9316_/D _9647_/SET_B VGND VPWR _9316_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6528_ _9136_/Q VGND VPWR _6528_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_6459_ _6457_/Y _5837_/B _6458_/Y _5960_/B VGND VPWR _6459_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_9247_ _9278_/CLK _9247_/D _9779_/SET_B VGND VPWR _9247_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_7_csclk clkbuf_2_2_0_csclk/X VGND VPWR _9354_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_161_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9178_ _9613_/CLK _9178_/D _9646_/SET_B VGND VPWR _9178_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_121_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_8129_ _8130_/B _8378_/B VGND VPWR _8357_/A VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_87_263 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_235 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_162 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_440 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_620 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5830_ _5830_/A VGND VPWR _5831_/A VGND VPWR sky130_fd_sc_hd__clkbuf_2
X_5761_ _9237_/Q _5759_/A _8845_/X _5759_/Y VGND VPWR _9237_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_4712_ _9212_/Q VGND VPWR _4712_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_8480_ _8515_/B _8437_/B _8521_/B _8437_/B VGND VPWR _8706_/A VGND VPWR sky130_fd_sc_hd__o22ai_4
X_7500_ _7500_/A _7500_/B _7500_/C _7500_/D VGND VPWR _7500_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
XFILLER_175_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5692_ _5692_/A VGND VPWR _5692_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_7431_ _7474_/C _7472_/A _7474_/D VGND VPWR _7432_/A VGND VPWR sky130_fd_sc_hd__or3_1
XFILLER_175_577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_4643_ hold1/A _4636_/A _8947_/X _4636_/Y VGND VPWR _9716_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_128_460 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4574_ _9748_/Q _4566_/A _5967_/B1 _4566_/Y VGND VPWR _9748_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7362_ _6522_/Y _7059_/B _6557_/Y _7068_/C _7361_/X VGND VPWR _7365_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_143_441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7293_ _4930_/Y _7097_/X _4883_/Y _7099_/X VGND VPWR _7293_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_6313_ _6308_/Y _5757_/B _6309_/Y _5679_/B _6312_/X VGND VPWR _6325_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_9101_ _9777_/CLK _9101_/D _7011_/B VGND VPWR _9101_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_9032_ _9039_/CLK _9032_/D VGND VPWR _9032_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_6244_ _9499_/Q VGND VPWR _6244_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
XFILLER_89_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_102 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_550 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6175_ _9196_/Q VGND VPWR _6175_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_29_105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5126_ _9629_/Q _5123_/A _5965_/B1 _5123_/Y VGND VPWR _9629_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_111_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_222 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5057_ _7734_/A _7734_/B _8813_/A VGND VPWR _5062_/B VGND VPWR sky130_fd_sc_hd__a21oi_1
XFILLER_176_9 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_28 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_45 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_8816_ _8816_/A VGND VPWR _8816_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_5959_ _9106_/Q _5951_/A _8916_/A1 _5951_/Y VGND VPWR _9106_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8747_ _8747_/A VGND VPWR _8748_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_185_319 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_8678_ _8678_/A _8678_/B _8678_/C VGND VPWR _8723_/C VGND VPWR sky130_fd_sc_hd__or3_2
X_7629_ _6940_/Y _7419_/X _6868_/Y _7421_/X VGND VPWR _7629_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_4_248 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_64 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_498 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_171 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_472 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_350 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_383 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_372 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_268 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_11 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA_4 _7155_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_140_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_102 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_244 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7980_ _8528_/A _7994_/A VGND VPWR _7992_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_6931_ _6926_/Y _5660_/B _6927_/Y _5742_/B _6930_/X VGND VPWR _6944_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_81_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_9650_ _9653_/CLK _9650_/D _9646_/SET_B VGND VPWR _9650_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6862_ _9560_/Q VGND VPWR _8808_/A VGND VPWR sky130_fd_sc_hd__clkinv_2
X_5813_ _9202_/Q _5812_/A _8843_/X _5812_/Y VGND VPWR _9202_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8601_ _8601_/A _8696_/A _8662_/C _8601_/D VGND VPWR _8603_/B VGND VPWR sky130_fd_sc_hd__or4_1
X_9581_ _9620_/CLK _9581_/D _9633_/SET_B VGND VPWR _9581_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_8532_ _8528_/Y _8525_/Y _8518_/X _8464_/B VGND VPWR _8668_/C VGND VPWR sky130_fd_sc_hd__a31o_1
X_6793_ _9347_/Q VGND VPWR _6793_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
X_5744_ _5744_/A VGND VPWR _5744_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_5675_ _9267_/Q _5673_/A _8842_/X _5673_/Y VGND VPWR _9267_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_8463_ _8463_/A _8685_/A VGND VPWR _8464_/D VGND VPWR sky130_fd_sc_hd__or2_1
XFILLER_135_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7414_ _7474_/C _7472_/A _9255_/Q VGND VPWR _7415_/A VGND VPWR sky130_fd_sc_hd__or3_1
X_8394_ _8394_/A _8394_/B _8394_/C _8394_/D VGND VPWR _8395_/B VGND VPWR sky130_fd_sc_hd__or4_2
X_4626_ _5967_/B1 _9719_/Q _4626_/S VGND VPWR _4627_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_163_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7345_ _6674_/Y _7040_/D _6662_/Y _7110_/X _7344_/X VGND VPWR _7352_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_190_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_219 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4557_ _6111_/A _4805_/A VGND VPWR _4558_/B VGND VPWR sky130_fd_sc_hd__or2_2
XFILLER_171_580 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_7276_ _6121_/Y _7048_/D _6062_/Y _7040_/B _7275_/X VGND VPWR _7277_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_4488_ _4488_/A VGND VPWR _4911_/A VGND VPWR sky130_fd_sc_hd__buf_6
X_6227_ _6227_/A VGND VPWR _6227_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_9015_ _9039_/CLK _9015_/D VGND VPWR _9015_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_97_380 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6158_ _6158_/A _6158_/B VGND VPWR _6158_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_111_190 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5109_ _9640_/Q _5108_/X _7731_/A _5062_/D VGND VPWR _9640_/D VGND VPWR sky130_fd_sc_hd__o211a_2
Xclkbuf_leaf_10_csclk clkbuf_2_2_0_csclk/X VGND VPWR _9684_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_181_7 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6089_ _6083_/Y _5240_/B _6084_/Y _4590_/B _6088_/X VGND VPWR _6096_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_2
Xrepeater371 _9647_/SET_B VGND VPWR _9295_/SET_B VGND VPWR sky130_fd_sc_hd__buf_12
Xrepeater360 _8843_/X VGND VPWR _8925_/A1 VGND VPWR sky130_fd_sc_hd__buf_12
Xclkbuf_leaf_25_csclk clkbuf_2_3_0_csclk/X VGND VPWR _9652_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_41_612 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_9779_ _9779_/CLK _9779_/D _9779_/SET_B VGND VPWR _9779_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_31_52 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_430 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_546 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_290 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput163 wb_cyc_i VGND VPWR input163/X VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
Xinput141 wb_adr_i[19] VGND VPWR _7768_/C VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput152 wb_adr_i[29] VGND VPWR input152/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput130 usr2_vdd_pwrgood VGND VPWR _4867_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_36_406 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xinput196 wb_rstn_i VGND VPWR _6146_/A VGND VPWR sky130_fd_sc_hd__buf_12
Xinput174 wb_dat_i[19] VGND VPWR _7742_/B VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput185 wb_dat_i[29] VGND VPWR _7747_/A2 VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_16_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_400 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_494 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_191 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_180 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5460_ _5460_/A VGND VPWR _5460_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_8_395 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_528 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
X_5391_ _9451_/Q _5384_/A _8840_/X _5384_/Y VGND VPWR _9451_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_7130_ _4928_/Y _7124_/X _4771_/Y _7068_/B _7129_/X VGND VPWR _7131_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_7061_ _7061_/A VGND VPWR _7068_/A VGND VPWR sky130_fd_sc_hd__buf_8
XFILLER_101_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6012_ _6040_/A VGND VPWR _6013_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
.ends

.subckt caravel clock flash_clk flash_csb flash_io0 flash_io1 gpio mprj_io[0] mprj_io[10]
+ mprj_io[11] mprj_io[12] mprj_io[13] mprj_io[14] mprj_io[15] mprj_io[16] mprj_io[17]
+ mprj_io[18] mprj_io[19] mprj_io[1] mprj_io[20] mprj_io[21] mprj_io[22] mprj_io[23]
+ mprj_io[24] mprj_io[25] mprj_io[26] mprj_io[27] mprj_io[28] mprj_io[29] mprj_io[2]
+ mprj_io[30] mprj_io[31] mprj_io[32] mprj_io[33] mprj_io[34] mprj_io[35] mprj_io[36]
+ mprj_io[37] mprj_io[3] mprj_io[4] mprj_io[5] mprj_io[6] mprj_io[7] mprj_io[8] mprj_io[9]
+ resetb vccd vccd1 vccd2 vdda vdda1 vdda1_2 vdda2 vddio vddio_2 vssa vssa1 vssa1_2
+ vssa2 vssd vssd1 vssd2 vssio vssio_2
Xgpio_control_in_2\[0\] gpio_defaults_block_19/gpio_defaults[0] gpio_defaults_block_19/gpio_defaults[10]
+ gpio_defaults_block_19/gpio_defaults[11] gpio_defaults_block_19/gpio_defaults[12]
+ gpio_defaults_block_19/gpio_defaults[1] gpio_defaults_block_19/gpio_defaults[2]
+ gpio_defaults_block_19/gpio_defaults[3] gpio_defaults_block_19/gpio_defaults[4]
+ gpio_defaults_block_19/gpio_defaults[5] gpio_defaults_block_19/gpio_defaults[6]
+ gpio_defaults_block_19/gpio_defaults[7] gpio_defaults_block_19/gpio_defaults[8]
+ gpio_defaults_block_19/gpio_defaults[9] housekeeping/mgmt_gpio_in[19] gpio_control_in_2\[0\]/one
+ housekeeping/mgmt_gpio_in[19] gpio_control_in_2\[0\]/one padframe/mprj_io_analog_en[19]
+ padframe/mprj_io_analog_pol[19] padframe/mprj_io_analog_sel[19] padframe/mprj_io_dm[57]
+ padframe/mprj_io_dm[58] padframe/mprj_io_dm[59] padframe/mprj_io_holdover[19] padframe/mprj_io_ib_mode_sel[19]
+ padframe/mprj_io_in[19] padframe/mprj_io_inp_dis[19] padframe/mprj_io_out[19] padframe/mprj_io_oeb[19]
+ padframe/mprj_io_slow_sel[19] padframe/mprj_io_vtrip_sel[19] gpio_control_in_2\[0\]/resetn
+ gpio_control_in_2\[0\]/resetn_out gpio_control_in_2\[0\]/serial_clock gpio_control_in_2\[0\]/serial_clock_out
+ gpio_control_in_2\[0\]/serial_data_in gpio_control_in_2\[0\]/serial_data_out gpio_control_in_2\[0\]/serial_load
+ gpio_control_in_2\[0\]/serial_load_out mprj/io_in[19] mprj/io_oeb[19] mprj/io_out[19]
+ vccd1_core VSUBS gpio_control_in_2\[0\]/zero dw_304538_1027427# vccd_core vssd1_core
+ gpio_control_block
Xgpio_defaults_block_22 VSUBS gpio_defaults_block_22/gpio_defaults[0] gpio_defaults_block_22/gpio_defaults[10]
+ gpio_defaults_block_22/gpio_defaults[11] gpio_defaults_block_22/gpio_defaults[12]
+ gpio_defaults_block_22/gpio_defaults[1] gpio_defaults_block_22/gpio_defaults[2]
+ gpio_defaults_block_22/gpio_defaults[3] gpio_defaults_block_22/gpio_defaults[4]
+ gpio_defaults_block_22/gpio_defaults[5] gpio_defaults_block_22/gpio_defaults[6]
+ gpio_defaults_block_22/gpio_defaults[7] gpio_defaults_block_22/gpio_defaults[8]
+ gpio_defaults_block_22/gpio_defaults[9] vccd_core gpio_defaults_block
Xgpio_defaults_block_11 VSUBS gpio_defaults_block_11/gpio_defaults[0] gpio_defaults_block_11/gpio_defaults[10]
+ gpio_defaults_block_11/gpio_defaults[11] gpio_defaults_block_11/gpio_defaults[12]
+ gpio_defaults_block_11/gpio_defaults[1] gpio_defaults_block_11/gpio_defaults[2]
+ gpio_defaults_block_11/gpio_defaults[3] gpio_defaults_block_11/gpio_defaults[4]
+ gpio_defaults_block_11/gpio_defaults[5] gpio_defaults_block_11/gpio_defaults[6]
+ gpio_defaults_block_11/gpio_defaults[7] gpio_defaults_block_11/gpio_defaults[8]
+ gpio_defaults_block_11/gpio_defaults[9] vccd_core gpio_defaults_block
Xgpio_defaults_block_33 VSUBS gpio_defaults_block_33/gpio_defaults[0] gpio_defaults_block_33/gpio_defaults[10]
+ gpio_defaults_block_33/gpio_defaults[11] gpio_defaults_block_33/gpio_defaults[12]
+ gpio_defaults_block_33/gpio_defaults[1] gpio_defaults_block_33/gpio_defaults[2]
+ gpio_defaults_block_33/gpio_defaults[3] gpio_defaults_block_33/gpio_defaults[4]
+ gpio_defaults_block_33/gpio_defaults[5] gpio_defaults_block_33/gpio_defaults[6]
+ gpio_defaults_block_33/gpio_defaults[7] gpio_defaults_block_33/gpio_defaults[8]
+ gpio_defaults_block_33/gpio_defaults[9] vccd_core gpio_defaults_block
Xgpio_defaults_block_23 VSUBS gpio_defaults_block_23/gpio_defaults[0] gpio_defaults_block_23/gpio_defaults[10]
+ gpio_defaults_block_23/gpio_defaults[11] gpio_defaults_block_23/gpio_defaults[12]
+ gpio_defaults_block_23/gpio_defaults[1] gpio_defaults_block_23/gpio_defaults[2]
+ gpio_defaults_block_23/gpio_defaults[3] gpio_defaults_block_23/gpio_defaults[4]
+ gpio_defaults_block_23/gpio_defaults[5] gpio_defaults_block_23/gpio_defaults[6]
+ gpio_defaults_block_23/gpio_defaults[7] gpio_defaults_block_23/gpio_defaults[8]
+ gpio_defaults_block_23/gpio_defaults[9] vccd_core gpio_defaults_block
Xgpio_control_in_1\[6\] gpio_defaults_block_14/gpio_defaults[0] gpio_defaults_block_14/gpio_defaults[10]
+ gpio_defaults_block_14/gpio_defaults[11] gpio_defaults_block_14/gpio_defaults[12]
+ gpio_defaults_block_14/gpio_defaults[1] gpio_defaults_block_14/gpio_defaults[2]
+ gpio_defaults_block_14/gpio_defaults[3] gpio_defaults_block_14/gpio_defaults[4]
+ gpio_defaults_block_14/gpio_defaults[5] gpio_defaults_block_14/gpio_defaults[6]
+ gpio_defaults_block_14/gpio_defaults[7] gpio_defaults_block_14/gpio_defaults[8]
+ gpio_defaults_block_14/gpio_defaults[9] housekeeping/mgmt_gpio_in[14] gpio_control_in_1\[6\]/one
+ housekeeping/mgmt_gpio_in[14] gpio_control_in_1\[6\]/one padframe/mprj_io_analog_en[14]
+ padframe/mprj_io_analog_pol[14] padframe/mprj_io_analog_sel[14] padframe/mprj_io_dm[42]
+ padframe/mprj_io_dm[43] padframe/mprj_io_dm[44] padframe/mprj_io_holdover[14] padframe/mprj_io_ib_mode_sel[14]
+ padframe/mprj_io_in[14] padframe/mprj_io_inp_dis[14] padframe/mprj_io_out[14] padframe/mprj_io_oeb[14]
+ padframe/mprj_io_slow_sel[14] padframe/mprj_io_vtrip_sel[14] gpio_control_in_1\[6\]/resetn
+ gpio_control_in_1\[7\]/resetn gpio_control_in_1\[6\]/serial_clock gpio_control_in_1\[7\]/serial_clock
+ gpio_control_in_1\[6\]/serial_data_in gpio_control_in_1\[7\]/serial_data_in gpio_control_in_1\[6\]/serial_load
+ gpio_control_in_1\[7\]/serial_load mprj/io_in[14] mprj/io_oeb[14] mprj/io_out[14]
+ vccd1_core VSUBS gpio_control_in_1\[6\]/zero dw_707553_929138# vccd_core vssd1_core
+ gpio_control_block
Xgpio_defaults_block_12 VSUBS gpio_defaults_block_12/gpio_defaults[0] gpio_defaults_block_12/gpio_defaults[10]
+ gpio_defaults_block_12/gpio_defaults[11] gpio_defaults_block_12/gpio_defaults[12]
+ gpio_defaults_block_12/gpio_defaults[1] gpio_defaults_block_12/gpio_defaults[2]
+ gpio_defaults_block_12/gpio_defaults[3] gpio_defaults_block_12/gpio_defaults[4]
+ gpio_defaults_block_12/gpio_defaults[5] gpio_defaults_block_12/gpio_defaults[6]
+ gpio_defaults_block_12/gpio_defaults[7] gpio_defaults_block_12/gpio_defaults[8]
+ gpio_defaults_block_12/gpio_defaults[9] vccd_core gpio_defaults_block
Xgpio_defaults_defaults_block_34 VSUBS gpio_control_in_2\[15\]/gpio_defaults[0] gpio_control_in_2\[15\]/gpio_defaults[10]
+ gpio_control_in_2\[15\]/gpio_defaults[11] gpio_control_in_2\[15\]/gpio_defaults[12]
+ gpio_control_in_2\[15\]/gpio_defaults[1] gpio_control_in_2\[15\]/gpio_defaults[2]
+ gpio_control_in_2\[15\]/gpio_defaults[3] gpio_control_in_2\[15\]/gpio_defaults[4]
+ gpio_control_in_2\[15\]/gpio_defaults[5] gpio_control_in_2\[15\]/gpio_defaults[6]
+ gpio_control_in_2\[15\]/gpio_defaults[7] gpio_control_in_2\[15\]/gpio_defaults[8]
+ gpio_control_in_2\[15\]/gpio_defaults[9] vccd_core gpio_defaults_block
Xpll pll/clockp[0] pll/clockp[1] pll/dco pll/div[0] pll/div[1] pll/div[2] pll/div[3]
+ pll/div[4] pll/enable pll/ext_trim[0] pll/ext_trim[10] pll/ext_trim[11] pll/ext_trim[12]
+ pll/ext_trim[13] pll/ext_trim[14] pll/ext_trim[15] pll/ext_trim[16] pll/ext_trim[17]
+ pll/ext_trim[18] pll/ext_trim[19] pll/ext_trim[1] pll/ext_trim[20] pll/ext_trim[21]
+ pll/ext_trim[22] pll/ext_trim[23] pll/ext_trim[24] pll/ext_trim[25] pll/ext_trim[2]
+ pll/ext_trim[3] pll/ext_trim[4] pll/ext_trim[5] pll/ext_trim[6] pll/ext_trim[7]
+ pll/ext_trim[8] pll/ext_trim[9] pll/osc pll/resetb vccd_core VSUBS digital_pll
Xpadframe clock pll/osc por/por_l flash_clk padframe/flash_clk_core padframe/flash_clk_ieb_core
+ padframe/flash_clk_oeb_core flash_csb padframe/flash_csb_core padframe/flash_csb_ieb_core
+ padframe/flash_csb_oeb_core flash_io0 padframe/flash_io0_di_core padframe/flash_io0_do_core
+ padframe/flash_io0_oeb_core flash_io1 padframe/flash_io1_di_core padframe/flash_io1_do_core
+ padframe/flash_io1_oeb_core gpio soc/gpio_in_pad soc/gpio_inenb_pad soc/gpio_mode0_pad
+ soc/gpio_mode1_pad soc/gpio_out_pad soc/gpio_outenb_pad vccd vdda vddio vddio_2
+ vssa vssd vssio vssio_2 mprj_io[0] padframe/mprj_io_analog_en[0] padframe/mprj_io_analog_pol[0]
+ padframe/mprj_io_analog_sel[0] padframe/mprj_io_dm[0] padframe/mprj_io_dm[1] padframe/mprj_io_dm[2]
+ padframe/mprj_io_holdover[0] padframe/mprj_io_ib_mode_sel[0] padframe/mprj_io_inp_dis[0]
+ padframe/mprj_io_oeb[0] padframe/mprj_io_out[0] padframe/mprj_io_slow_sel[0] padframe/mprj_io_vtrip_sel[0]
+ padframe/mprj_io_in[0] mprj/analog_io[3] mprj_io[10] padframe/mprj_io_analog_en[10]
+ padframe/mprj_io_analog_pol[10] padframe/mprj_io_analog_sel[10] padframe/mprj_io_dm[30]
+ padframe/mprj_io_dm[31] padframe/mprj_io_dm[32] padframe/mprj_io_holdover[10] padframe/mprj_io_ib_mode_sel[10]
+ padframe/mprj_io_inp_dis[10] padframe/mprj_io_oeb[10] padframe/mprj_io_out[10] padframe/mprj_io_slow_sel[10]
+ padframe/mprj_io_vtrip_sel[10] padframe/mprj_io_in[10] mprj/analog_io[4] mprj_io[11]
+ padframe/mprj_io_analog_en[11] padframe/mprj_io_analog_pol[11] padframe/mprj_io_analog_sel[11]
+ padframe/mprj_io_dm[33] padframe/mprj_io_dm[34] padframe/mprj_io_dm[35] padframe/mprj_io_holdover[11]
+ padframe/mprj_io_ib_mode_sel[11] padframe/mprj_io_inp_dis[11] padframe/mprj_io_oeb[11]
+ padframe/mprj_io_out[11] padframe/mprj_io_slow_sel[11] padframe/mprj_io_vtrip_sel[11]
+ padframe/mprj_io_in[11] mprj/analog_io[5] mprj_io[12] padframe/mprj_io_analog_en[12]
+ padframe/mprj_io_analog_pol[12] padframe/mprj_io_analog_sel[12] padframe/mprj_io_dm[36]
+ padframe/mprj_io_dm[37] padframe/mprj_io_dm[38] padframe/mprj_io_holdover[12] padframe/mprj_io_ib_mode_sel[12]
+ padframe/mprj_io_inp_dis[12] padframe/mprj_io_oeb[12] padframe/mprj_io_out[12] padframe/mprj_io_slow_sel[12]
+ padframe/mprj_io_vtrip_sel[12] padframe/mprj_io_in[12] mprj/analog_io[6] mprj_io[13]
+ padframe/mprj_io_analog_en[13] padframe/mprj_io_analog_pol[13] padframe/mprj_io_analog_sel[13]
+ padframe/mprj_io_dm[39] padframe/mprj_io_dm[40] padframe/mprj_io_dm[41] padframe/mprj_io_holdover[13]
+ padframe/mprj_io_ib_mode_sel[13] padframe/mprj_io_inp_dis[13] padframe/mprj_io_oeb[13]
+ padframe/mprj_io_out[13] padframe/mprj_io_slow_sel[13] padframe/mprj_io_vtrip_sel[13]
+ padframe/mprj_io_in[13] mprj/analog_io[7] mprj_io[14] padframe/mprj_io_analog_en[14]
+ padframe/mprj_io_analog_pol[14] padframe/mprj_io_analog_sel[14] padframe/mprj_io_dm[42]
+ padframe/mprj_io_dm[43] padframe/mprj_io_dm[44] padframe/mprj_io_holdover[14] padframe/mprj_io_ib_mode_sel[14]
+ padframe/mprj_io_inp_dis[14] padframe/mprj_io_oeb[14] padframe/mprj_io_out[14] padframe/mprj_io_slow_sel[14]
+ padframe/mprj_io_vtrip_sel[14] padframe/mprj_io_in[14] mprj/analog_io[8] mprj_io[15]
+ padframe/mprj_io_analog_en[15] padframe/mprj_io_analog_pol[15] padframe/mprj_io_analog_sel[15]
+ padframe/mprj_io_dm[45] padframe/mprj_io_dm[46] padframe/mprj_io_dm[47] padframe/mprj_io_holdover[15]
+ padframe/mprj_io_ib_mode_sel[15] padframe/mprj_io_inp_dis[15] padframe/mprj_io_oeb[15]
+ padframe/mprj_io_out[15] padframe/mprj_io_slow_sel[15] padframe/mprj_io_vtrip_sel[15]
+ padframe/mprj_io_in[15] mprj/analog_io[9] mprj_io[16] padframe/mprj_io_analog_en[16]
+ padframe/mprj_io_analog_pol[16] padframe/mprj_io_analog_sel[16] padframe/mprj_io_dm[48]
+ padframe/mprj_io_dm[49] padframe/mprj_io_dm[50] padframe/mprj_io_holdover[16] padframe/mprj_io_ib_mode_sel[16]
+ padframe/mprj_io_inp_dis[16] padframe/mprj_io_oeb[16] padframe/mprj_io_out[16] padframe/mprj_io_slow_sel[16]
+ padframe/mprj_io_vtrip_sel[16] padframe/mprj_io_in[16] mprj/analog_io[10] mprj_io[17]
+ padframe/mprj_io_analog_en[17] padframe/mprj_io_analog_pol[17] padframe/mprj_io_analog_sel[17]
+ padframe/mprj_io_dm[51] padframe/mprj_io_dm[52] padframe/mprj_io_dm[53] padframe/mprj_io_holdover[17]
+ padframe/mprj_io_ib_mode_sel[17] padframe/mprj_io_inp_dis[17] padframe/mprj_io_oeb[17]
+ padframe/mprj_io_out[17] padframe/mprj_io_slow_sel[17] padframe/mprj_io_vtrip_sel[17]
+ padframe/mprj_io_in[17] mprj/analog_io[11] mprj_io[18] padframe/mprj_io_analog_en[18]
+ padframe/mprj_io_analog_pol[18] padframe/mprj_io_analog_sel[18] padframe/mprj_io_dm[54]
+ padframe/mprj_io_dm[55] padframe/mprj_io_dm[56] padframe/mprj_io_holdover[18] padframe/mprj_io_ib_mode_sel[18]
+ padframe/mprj_io_inp_dis[18] padframe/mprj_io_oeb[18] padframe/mprj_io_out[18] padframe/mprj_io_slow_sel[18]
+ padframe/mprj_io_vtrip_sel[18] padframe/mprj_io_in[18] mprj_io[1] padframe/mprj_io_analog_en[1]
+ padframe/mprj_io_analog_pol[1] padframe/mprj_io_analog_sel[1] padframe/mprj_io_dm[3]
+ padframe/mprj_io_dm[4] padframe/mprj_io_dm[5] padframe/mprj_io_holdover[1] padframe/mprj_io_ib_mode_sel[1]
+ padframe/mprj_io_inp_dis[1] padframe/mprj_io_oeb[1] padframe/mprj_io_out[1] padframe/mprj_io_slow_sel[1]
+ padframe/mprj_io_vtrip_sel[1] padframe/mprj_io_in[1] mprj_io[2] padframe/mprj_io_analog_en[2]
+ padframe/mprj_io_analog_pol[2] padframe/mprj_io_analog_sel[2] padframe/mprj_io_dm[6]
+ padframe/mprj_io_dm[7] padframe/mprj_io_dm[8] padframe/mprj_io_holdover[2] padframe/mprj_io_ib_mode_sel[2]
+ padframe/mprj_io_inp_dis[2] padframe/mprj_io_oeb[2] padframe/mprj_io_out[2] padframe/mprj_io_slow_sel[2]
+ padframe/mprj_io_vtrip_sel[2] padframe/mprj_io_in[2] mprj_io[3] padframe/mprj_io_analog_en[3]
+ padframe/mprj_io_analog_pol[3] padframe/mprj_io_analog_sel[3] padframe/mprj_io_dm[10]
+ padframe/mprj_io_dm[11] padframe/mprj_io_dm[9] padframe/mprj_io_holdover[3] padframe/mprj_io_ib_mode_sel[3]
+ padframe/mprj_io_inp_dis[3] padframe/mprj_io_oeb[3] padframe/mprj_io_out[3] padframe/mprj_io_slow_sel[3]
+ padframe/mprj_io_vtrip_sel[3] padframe/mprj_io_in[3] mprj_io[4] padframe/mprj_io_analog_en[4]
+ padframe/mprj_io_analog_pol[4] padframe/mprj_io_analog_sel[4] padframe/mprj_io_dm[12]
+ padframe/mprj_io_dm[13] padframe/mprj_io_dm[14] padframe/mprj_io_holdover[4] padframe/mprj_io_ib_mode_sel[4]
+ padframe/mprj_io_inp_dis[4] padframe/mprj_io_oeb[4] padframe/mprj_io_out[4] padframe/mprj_io_slow_sel[4]
+ padframe/mprj_io_vtrip_sel[4] padframe/mprj_io_in[4] mprj_io[5] padframe/mprj_io_analog_en[5]
+ padframe/mprj_io_analog_pol[5] padframe/mprj_io_analog_sel[5] padframe/mprj_io_dm[15]
+ padframe/mprj_io_dm[16] padframe/mprj_io_dm[17] padframe/mprj_io_holdover[5] padframe/mprj_io_ib_mode_sel[5]
+ padframe/mprj_io_inp_dis[5] padframe/mprj_io_oeb[5] padframe/mprj_io_out[5] padframe/mprj_io_slow_sel[5]
+ padframe/mprj_io_vtrip_sel[5] padframe/mprj_io_in[5] mprj_io[6] padframe/mprj_io_analog_en[6]
+ padframe/mprj_io_analog_pol[6] padframe/mprj_io_analog_sel[6] padframe/mprj_io_dm[18]
+ padframe/mprj_io_dm[19] padframe/mprj_io_dm[20] padframe/mprj_io_holdover[6] padframe/mprj_io_ib_mode_sel[6]
+ padframe/mprj_io_inp_dis[6] padframe/mprj_io_oeb[6] padframe/mprj_io_out[6] padframe/mprj_io_slow_sel[6]
+ padframe/mprj_io_vtrip_sel[6] padframe/mprj_io_in[6] mprj/analog_io[0] mprj_io[7]
+ padframe/mprj_io_analog_en[7] padframe/mprj_io_analog_pol[7] padframe/mprj_io_analog_sel[7]
+ padframe/mprj_io_dm[21] padframe/mprj_io_dm[22] padframe/mprj_io_dm[23] padframe/mprj_io_holdover[7]
+ padframe/mprj_io_ib_mode_sel[7] padframe/mprj_io_inp_dis[7] padframe/mprj_io_oeb[7]
+ padframe/mprj_io_out[7] padframe/mprj_io_slow_sel[7] padframe/mprj_io_vtrip_sel[7]
+ padframe/mprj_io_in[7] mprj/analog_io[1] mprj_io[8] padframe/mprj_io_analog_en[8]
+ padframe/mprj_io_analog_pol[8] padframe/mprj_io_analog_sel[8] padframe/mprj_io_dm[24]
+ padframe/mprj_io_dm[25] padframe/mprj_io_dm[26] padframe/mprj_io_holdover[8] padframe/mprj_io_ib_mode_sel[8]
+ padframe/mprj_io_inp_dis[8] padframe/mprj_io_oeb[8] padframe/mprj_io_out[8] padframe/mprj_io_slow_sel[8]
+ padframe/mprj_io_vtrip_sel[8] padframe/mprj_io_in[8] mprj/analog_io[2] mprj_io[9]
+ padframe/mprj_io_analog_en[9] padframe/mprj_io_analog_pol[9] padframe/mprj_io_analog_sel[9]
+ padframe/mprj_io_dm[27] padframe/mprj_io_dm[28] padframe/mprj_io_dm[29] padframe/mprj_io_holdover[9]
+ padframe/mprj_io_ib_mode_sel[9] padframe/mprj_io_inp_dis[9] padframe/mprj_io_oeb[9]
+ padframe/mprj_io_out[9] padframe/mprj_io_slow_sel[9] padframe/mprj_io_vtrip_sel[9]
+ padframe/mprj_io_in[9] mprj/analog_io[12] mprj_io[19] padframe/mprj_io_analog_en[19]
+ padframe/mprj_io_analog_pol[19] padframe/mprj_io_analog_sel[19] padframe/mprj_io_dm[57]
+ padframe/mprj_io_dm[58] padframe/mprj_io_dm[59] padframe/mprj_io_holdover[19] padframe/mprj_io_ib_mode_sel[19]
+ padframe/mprj_io_inp_dis[19] padframe/mprj_io_oeb[19] padframe/mprj_io_out[19] padframe/mprj_io_slow_sel[19]
+ padframe/mprj_io_vtrip_sel[19] padframe/mprj_io_in[19] mprj/analog_io[22] mprj_io[29]
+ padframe/mprj_io_analog_en[29] padframe/mprj_io_analog_pol[29] padframe/mprj_io_analog_sel[29]
+ padframe/mprj_io_dm[87] padframe/mprj_io_dm[88] padframe/mprj_io_dm[89] padframe/mprj_io_holdover[29]
+ padframe/mprj_io_ib_mode_sel[29] padframe/mprj_io_inp_dis[29] padframe/mprj_io_oeb[29]
+ padframe/mprj_io_out[29] padframe/mprj_io_slow_sel[29] padframe/mprj_io_vtrip_sel[29]
+ padframe/mprj_io_in[29] mprj/analog_io[23] mprj_io[30] padframe/mprj_io_analog_en[30]
+ padframe/mprj_io_analog_pol[30] padframe/mprj_io_analog_sel[30] padframe/mprj_io_dm[90]
+ padframe/mprj_io_dm[91] padframe/mprj_io_dm[92] padframe/mprj_io_holdover[30] padframe/mprj_io_ib_mode_sel[30]
+ padframe/mprj_io_inp_dis[30] padframe/mprj_io_oeb[30] padframe/mprj_io_out[30] padframe/mprj_io_slow_sel[30]
+ padframe/mprj_io_vtrip_sel[30] padframe/mprj_io_in[30] mprj/analog_io[24] mprj_io[31]
+ padframe/mprj_io_analog_en[31] padframe/mprj_io_analog_pol[31] padframe/mprj_io_analog_sel[31]
+ padframe/mprj_io_dm[93] padframe/mprj_io_dm[94] padframe/mprj_io_dm[95] padframe/mprj_io_holdover[31]
+ padframe/mprj_io_ib_mode_sel[31] padframe/mprj_io_inp_dis[31] padframe/mprj_io_oeb[31]
+ padframe/mprj_io_out[31] padframe/mprj_io_slow_sel[31] padframe/mprj_io_vtrip_sel[31]
+ padframe/mprj_io_in[31] mprj/analog_io[25] mprj_io[32] padframe/mprj_io_analog_en[32]
+ padframe/mprj_io_analog_pol[32] padframe/mprj_io_analog_sel[32] padframe/mprj_io_dm[96]
+ padframe/mprj_io_dm[97] padframe/mprj_io_dm[98] padframe/mprj_io_holdover[32] padframe/mprj_io_ib_mode_sel[32]
+ padframe/mprj_io_inp_dis[32] padframe/mprj_io_oeb[32] padframe/mprj_io_out[32] padframe/mprj_io_slow_sel[32]
+ padframe/mprj_io_vtrip_sel[32] padframe/mprj_io_in[32] mprj/analog_io[26] mprj_io[33]
+ padframe/mprj_io_analog_en[33] padframe/mprj_io_analog_pol[33] padframe/mprj_io_analog_sel[33]
+ padframe/mprj_io_dm[100] padframe/mprj_io_dm[101] padframe/mprj_io_dm[99] padframe/mprj_io_holdover[33]
+ padframe/mprj_io_ib_mode_sel[33] padframe/mprj_io_inp_dis[33] padframe/mprj_io_oeb[33]
+ padframe/mprj_io_out[33] padframe/mprj_io_slow_sel[33] padframe/mprj_io_vtrip_sel[33]
+ padframe/mprj_io_in[33] mprj/analog_io[27] mprj_io[34] padframe/mprj_io_analog_en[34]
+ padframe/mprj_io_analog_pol[34] padframe/mprj_io_analog_sel[34] padframe/mprj_io_dm[102]
+ padframe/mprj_io_dm[103] padframe/mprj_io_dm[104] padframe/mprj_io_holdover[34]
+ padframe/mprj_io_ib_mode_sel[34] padframe/mprj_io_inp_dis[34] padframe/mprj_io_oeb[34]
+ padframe/mprj_io_out[34] padframe/mprj_io_slow_sel[34] padframe/mprj_io_vtrip_sel[34]
+ padframe/mprj_io_in[34] mprj/analog_io[28] mprj_io[35] padframe/mprj_io_analog_en[35]
+ padframe/mprj_io_analog_pol[35] padframe/mprj_io_analog_sel[35] padframe/mprj_io_dm[105]
+ padframe/mprj_io_dm[106] padframe/mprj_io_dm[107] padframe/mprj_io_holdover[35]
+ padframe/mprj_io_ib_mode_sel[35] padframe/mprj_io_inp_dis[35] padframe/mprj_io_oeb[35]
+ padframe/mprj_io_out[35] padframe/mprj_io_slow_sel[35] padframe/mprj_io_vtrip_sel[35]
+ padframe/mprj_io_in[35] mprj_io[36] padframe/mprj_io_analog_en[36] padframe/mprj_io_analog_pol[36]
+ padframe/mprj_io_analog_sel[36] padframe/mprj_io_dm[108] padframe/mprj_io_dm[109]
+ padframe/mprj_io_dm[110] padframe/mprj_io_holdover[36] padframe/mprj_io_ib_mode_sel[36]
+ padframe/mprj_io_inp_dis[36] padframe/mprj_io_oeb[36] padframe/mprj_io_out[36] padframe/mprj_io_slow_sel[36]
+ padframe/mprj_io_vtrip_sel[36] padframe/mprj_io_in[36] mprj_io[37] padframe/mprj_io_analog_en[37]
+ padframe/mprj_io_analog_pol[37] padframe/mprj_io_analog_sel[37] padframe/mprj_io_dm[111]
+ padframe/mprj_io_dm[112] padframe/mprj_io_dm[113] padframe/mprj_io_holdover[37]
+ padframe/mprj_io_ib_mode_sel[37] padframe/mprj_io_inp_dis[37] padframe/mprj_io_oeb[37]
+ padframe/mprj_io_out[37] padframe/mprj_io_slow_sel[37] padframe/mprj_io_vtrip_sel[37]
+ padframe/mprj_io_in[37] mprj/analog_io[13] mprj_io[20] padframe/mprj_io_analog_en[20]
+ padframe/mprj_io_analog_pol[20] padframe/mprj_io_analog_sel[20] padframe/mprj_io_dm[60]
+ padframe/mprj_io_dm[61] padframe/mprj_io_dm[62] padframe/mprj_io_holdover[20] padframe/mprj_io_ib_mode_sel[20]
+ padframe/mprj_io_inp_dis[20] padframe/mprj_io_oeb[20] padframe/mprj_io_out[20] padframe/mprj_io_slow_sel[20]
+ padframe/mprj_io_vtrip_sel[20] padframe/mprj_io_in[20] mprj/analog_io[14] mprj_io[21]
+ padframe/mprj_io_analog_en[21] padframe/mprj_io_analog_pol[21] padframe/mprj_io_analog_sel[21]
+ padframe/mprj_io_dm[63] padframe/mprj_io_dm[64] padframe/mprj_io_dm[65] padframe/mprj_io_holdover[21]
+ padframe/mprj_io_ib_mode_sel[21] padframe/mprj_io_inp_dis[21] padframe/mprj_io_oeb[21]
+ padframe/mprj_io_out[21] padframe/mprj_io_slow_sel[21] padframe/mprj_io_vtrip_sel[21]
+ padframe/mprj_io_in[21] mprj/analog_io[15] mprj_io[22] padframe/mprj_io_analog_en[22]
+ padframe/mprj_io_analog_pol[22] padframe/mprj_io_analog_sel[22] padframe/mprj_io_dm[66]
+ padframe/mprj_io_dm[67] padframe/mprj_io_dm[68] padframe/mprj_io_holdover[22] padframe/mprj_io_ib_mode_sel[22]
+ padframe/mprj_io_inp_dis[22] padframe/mprj_io_oeb[22] padframe/mprj_io_out[22] padframe/mprj_io_slow_sel[22]
+ padframe/mprj_io_vtrip_sel[22] padframe/mprj_io_in[22] mprj/analog_io[16] mprj_io[23]
+ padframe/mprj_io_analog_en[23] padframe/mprj_io_analog_pol[23] padframe/mprj_io_analog_sel[23]
+ padframe/mprj_io_dm[69] padframe/mprj_io_dm[70] padframe/mprj_io_dm[71] padframe/mprj_io_holdover[23]
+ padframe/mprj_io_ib_mode_sel[23] padframe/mprj_io_inp_dis[23] padframe/mprj_io_oeb[23]
+ padframe/mprj_io_out[23] padframe/mprj_io_slow_sel[23] padframe/mprj_io_vtrip_sel[23]
+ padframe/mprj_io_in[23] mprj/analog_io[17] mprj_io[24] padframe/mprj_io_analog_en[24]
+ padframe/mprj_io_analog_pol[24] padframe/mprj_io_analog_sel[24] padframe/mprj_io_dm[72]
+ padframe/mprj_io_dm[73] padframe/mprj_io_dm[74] padframe/mprj_io_holdover[24] padframe/mprj_io_ib_mode_sel[24]
+ padframe/mprj_io_inp_dis[24] padframe/mprj_io_oeb[24] padframe/mprj_io_out[24] padframe/mprj_io_slow_sel[24]
+ padframe/mprj_io_vtrip_sel[24] padframe/mprj_io_in[24] mprj/analog_io[18] mprj_io[25]
+ padframe/mprj_io_analog_en[25] padframe/mprj_io_analog_pol[25] padframe/mprj_io_analog_sel[25]
+ padframe/mprj_io_dm[75] padframe/mprj_io_dm[76] padframe/mprj_io_dm[77] padframe/mprj_io_holdover[25]
+ padframe/mprj_io_ib_mode_sel[25] padframe/mprj_io_inp_dis[25] padframe/mprj_io_oeb[25]
+ padframe/mprj_io_out[25] padframe/mprj_io_slow_sel[25] padframe/mprj_io_vtrip_sel[25]
+ padframe/mprj_io_in[25] mprj/analog_io[19] mprj_io[26] padframe/mprj_io_analog_en[26]
+ padframe/mprj_io_analog_pol[26] padframe/mprj_io_analog_sel[26] padframe/mprj_io_dm[78]
+ padframe/mprj_io_dm[79] padframe/mprj_io_dm[80] padframe/mprj_io_holdover[26] padframe/mprj_io_ib_mode_sel[26]
+ padframe/mprj_io_inp_dis[26] padframe/mprj_io_oeb[26] padframe/mprj_io_out[26] padframe/mprj_io_slow_sel[26]
+ padframe/mprj_io_vtrip_sel[26] padframe/mprj_io_in[26] mprj/analog_io[20] mprj_io[27]
+ padframe/mprj_io_analog_en[27] padframe/mprj_io_analog_pol[27] padframe/mprj_io_analog_sel[27]
+ padframe/mprj_io_dm[81] padframe/mprj_io_dm[82] padframe/mprj_io_dm[83] padframe/mprj_io_holdover[27]
+ padframe/mprj_io_ib_mode_sel[27] padframe/mprj_io_inp_dis[27] padframe/mprj_io_oeb[27]
+ padframe/mprj_io_out[27] padframe/mprj_io_slow_sel[27] padframe/mprj_io_vtrip_sel[27]
+ padframe/mprj_io_in[27] mprj/analog_io[21] mprj_io[28] padframe/mprj_io_analog_en[28]
+ padframe/mprj_io_analog_pol[28] padframe/mprj_io_analog_sel[28] padframe/mprj_io_dm[84]
+ padframe/mprj_io_dm[85] padframe/mprj_io_dm[86] padframe/mprj_io_holdover[28] padframe/mprj_io_ib_mode_sel[28]
+ padframe/mprj_io_inp_dis[28] padframe/mprj_io_oeb[28] padframe/mprj_io_out[28] padframe/mprj_io_slow_sel[28]
+ padframe/mprj_io_vtrip_sel[28] padframe/mprj_io_in[28] por/porb_h resetb rstb_level/A
+ padframe/vdda padframe/vssa vccd1 vdda1 vdda1_2 vssa1 vssa1_2 vccd1_core vdda1_core
+ vssd1_core vssd1 vccd2 vdda2 vssa2 vccd2_core vdda2_core por/vdd3v3 vssd2_core vssd2
+ vssa2_core padframe/flash_io0_ieb_core por/vss3v3 vssa1_core padframe/flash_io1_ieb_core
+ vccd_core VSUBS chip_io
Xgpio_defaults_block_24 VSUBS gpio_defaults_block_24/gpio_defaults[0] gpio_defaults_block_24/gpio_defaults[10]
+ gpio_defaults_block_24/gpio_defaults[11] gpio_defaults_block_24/gpio_defaults[12]
+ gpio_defaults_block_24/gpio_defaults[1] gpio_defaults_block_24/gpio_defaults[2]
+ gpio_defaults_block_24/gpio_defaults[3] gpio_defaults_block_24/gpio_defaults[4]
+ gpio_defaults_block_24/gpio_defaults[5] gpio_defaults_block_24/gpio_defaults[6]
+ gpio_defaults_block_24/gpio_defaults[7] gpio_defaults_block_24/gpio_defaults[8]
+ gpio_defaults_block_24/gpio_defaults[9] vccd_core gpio_defaults_block
Xgpio_defaults_block_13 VSUBS gpio_defaults_block_13/gpio_defaults[0] gpio_defaults_block_13/gpio_defaults[10]
+ gpio_defaults_block_13/gpio_defaults[11] gpio_defaults_block_13/gpio_defaults[12]
+ gpio_defaults_block_13/gpio_defaults[1] gpio_defaults_block_13/gpio_defaults[2]
+ gpio_defaults_block_13/gpio_defaults[3] gpio_defaults_block_13/gpio_defaults[4]
+ gpio_defaults_block_13/gpio_defaults[5] gpio_defaults_block_13/gpio_defaults[6]
+ gpio_defaults_block_13/gpio_defaults[7] gpio_defaults_block_13/gpio_defaults[8]
+ gpio_defaults_block_13/gpio_defaults[9] vccd_core gpio_defaults_block
Xgpio_control_in_1a\[3\] gpio_defaults_block_5/gpio_defaults[0] gpio_defaults_block_5/gpio_defaults[10]
+ gpio_defaults_block_5/gpio_defaults[11] gpio_defaults_block_5/gpio_defaults[12]
+ gpio_defaults_block_5/gpio_defaults[1] gpio_defaults_block_5/gpio_defaults[2] gpio_defaults_block_5/gpio_defaults[3]
+ gpio_defaults_block_5/gpio_defaults[4] gpio_defaults_block_5/gpio_defaults[5] gpio_defaults_block_5/gpio_defaults[6]
+ gpio_defaults_block_5/gpio_defaults[7] gpio_defaults_block_5/gpio_defaults[8] gpio_defaults_block_5/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[5] gpio_control_in_1a\[3\]/one housekeeping/mgmt_gpio_in[5]
+ gpio_control_in_1a\[3\]/one padframe/mprj_io_analog_en[5] padframe/mprj_io_analog_pol[5]
+ padframe/mprj_io_analog_sel[5] padframe/mprj_io_dm[15] padframe/mprj_io_dm[16] padframe/mprj_io_dm[17]
+ padframe/mprj_io_holdover[5] padframe/mprj_io_ib_mode_sel[5] padframe/mprj_io_in[5]
+ padframe/mprj_io_inp_dis[5] padframe/mprj_io_out[5] padframe/mprj_io_oeb[5] padframe/mprj_io_slow_sel[5]
+ padframe/mprj_io_vtrip_sel[5] gpio_control_in_1a\[3\]/resetn gpio_control_in_1a\[4\]/resetn
+ gpio_control_in_1a\[3\]/serial_clock gpio_control_in_1a\[4\]/serial_clock gpio_control_in_1a\[3\]/serial_data_in
+ gpio_control_in_1a\[4\]/serial_data_in gpio_control_in_1a\[3\]/serial_load gpio_control_in_1a\[4\]/serial_load
+ mprj/io_in[5] mprj/io_oeb[5] mprj/io_out[5] vccd1_core VSUBS gpio_control_in_1a\[3\]/zero
+ dw_707553_347938# vccd_core vssd1_core gpio_control_block
Xgpio_control_in_2\[14\] gpio_defaults_block_33/gpio_defaults[0] gpio_defaults_block_33/gpio_defaults[10]
+ gpio_defaults_block_33/gpio_defaults[11] gpio_defaults_block_33/gpio_defaults[12]
+ gpio_defaults_block_33/gpio_defaults[1] gpio_defaults_block_33/gpio_defaults[2]
+ gpio_defaults_block_33/gpio_defaults[3] gpio_defaults_block_33/gpio_defaults[4]
+ gpio_defaults_block_33/gpio_defaults[5] gpio_defaults_block_33/gpio_defaults[6]
+ gpio_defaults_block_33/gpio_defaults[7] gpio_defaults_block_33/gpio_defaults[8]
+ gpio_defaults_block_33/gpio_defaults[9] housekeeping/mgmt_gpio_in[33] gpio_control_in_2\[14\]/one
+ housekeeping/mgmt_gpio_in[33] gpio_control_in_2\[14\]/one padframe/mprj_io_analog_en[33]
+ padframe/mprj_io_analog_pol[33] padframe/mprj_io_analog_sel[33] padframe/mprj_io_dm[99]
+ padframe/mprj_io_dm[100] padframe/mprj_io_dm[101] padframe/mprj_io_holdover[33]
+ padframe/mprj_io_ib_mode_sel[33] padframe/mprj_io_in[33] padframe/mprj_io_inp_dis[33]
+ padframe/mprj_io_out[33] padframe/mprj_io_oeb[33] padframe/mprj_io_slow_sel[33]
+ padframe/mprj_io_vtrip_sel[33] gpio_control_in_2\[14\]/resetn gpio_control_in_2\[13\]/resetn
+ gpio_control_in_2\[14\]/serial_clock gpio_control_in_2\[13\]/serial_clock gpio_control_in_2\[14\]/serial_data_in
+ gpio_control_in_2\[13\]/serial_data_in gpio_control_in_2\[14\]/serial_load gpio_control_in_2\[13\]/serial_load
+ mprj/io_in[33] mprj/io_oeb[33] mprj/io_out[33] vccd1_core VSUBS gpio_control_in_2\[14\]/zero
+ dw_8741_376938# vccd_core vssd1_core gpio_control_block
Xgpio_defaults_block_35 VSUBS gpio_defaults_block_35/gpio_defaults[0] gpio_defaults_block_35/gpio_defaults[10]
+ gpio_defaults_block_35/gpio_defaults[11] gpio_defaults_block_35/gpio_defaults[12]
+ gpio_defaults_block_35/gpio_defaults[1] gpio_defaults_block_35/gpio_defaults[2]
+ gpio_defaults_block_35/gpio_defaults[3] gpio_defaults_block_35/gpio_defaults[4]
+ gpio_defaults_block_35/gpio_defaults[5] gpio_defaults_block_35/gpio_defaults[6]
+ gpio_defaults_block_35/gpio_defaults[7] gpio_defaults_block_35/gpio_defaults[8]
+ gpio_defaults_block_35/gpio_defaults[9] vccd_core gpio_defaults_block
Xgpio_control_bidir_2\[0\] gpio_defaults_block_35/gpio_defaults[0] gpio_defaults_block_35/gpio_defaults[10]
+ gpio_defaults_block_35/gpio_defaults[11] gpio_defaults_block_35/gpio_defaults[12]
+ gpio_defaults_block_35/gpio_defaults[1] gpio_defaults_block_35/gpio_defaults[2]
+ gpio_defaults_block_35/gpio_defaults[3] gpio_defaults_block_35/gpio_defaults[4]
+ gpio_defaults_block_35/gpio_defaults[5] gpio_defaults_block_35/gpio_defaults[6]
+ gpio_defaults_block_35/gpio_defaults[7] gpio_defaults_block_35/gpio_defaults[8]
+ gpio_defaults_block_35/gpio_defaults[9] housekeeping/mgmt_gpio_in[35] housekeeping/mgmt_gpio_oeb[35]
+ housekeeping/mgmt_gpio_out[35] gpio_control_bidir_2\[0\]/one padframe/mprj_io_analog_en[35]
+ padframe/mprj_io_analog_pol[35] padframe/mprj_io_analog_sel[35] padframe/mprj_io_dm[105]
+ padframe/mprj_io_dm[106] padframe/mprj_io_dm[107] padframe/mprj_io_holdover[35]
+ padframe/mprj_io_ib_mode_sel[35] padframe/mprj_io_in[35] padframe/mprj_io_inp_dis[35]
+ padframe/mprj_io_out[35] padframe/mprj_io_oeb[35] padframe/mprj_io_slow_sel[35]
+ padframe/mprj_io_vtrip_sel[35] gpio_control_bidir_2\[0\]/resetn gpio_control_in_2\[15\]/resetn
+ gpio_control_bidir_2\[0\]/serial_clock gpio_control_in_2\[15\]/serial_clock gpio_control_bidir_2\[0\]/serial_data_in
+ gpio_control_in_2\[15\]/serial_data_in gpio_control_bidir_2\[0\]/serial_load gpio_control_in_2\[15\]/serial_load
+ mprj/io_in[35] mprj/io_oeb[35] mprj/io_out[35] vccd1_core VSUBS gpio_control_bidir_2\[0\]/zero
+ dw_8741_290538# vccd_core vssd1_core gpio_control_block
Xspare_logic_block_0 spare_logic_block_0/spare_xfq[0] spare_logic_block_0/spare_xfq[1]
+ spare_logic_block_0/spare_xfqn[0] spare_logic_block_0/spare_xfqn[1] spare_logic_block_0/spare_xi[0]
+ spare_logic_block_0/spare_xi[1] spare_logic_block_0/spare_xi[2] spare_logic_block_0/spare_xi[3]
+ spare_logic_block_0/spare_xib spare_logic_block_0/spare_xmx[0] spare_logic_block_0/spare_xmx[1]
+ spare_logic_block_0/spare_xna[0] spare_logic_block_0/spare_xna[1] spare_logic_block_0/spare_xno[0]
+ spare_logic_block_0/spare_xno[1] spare_logic_block_0/spare_xz[0] spare_logic_block_0/spare_xz[10]
+ spare_logic_block_0/spare_xz[11] spare_logic_block_0/spare_xz[12] spare_logic_block_0/spare_xz[13]
+ spare_logic_block_0/spare_xz[14] spare_logic_block_0/spare_xz[15] spare_logic_block_0/spare_xz[16]
+ spare_logic_block_0/spare_xz[17] spare_logic_block_0/spare_xz[18] spare_logic_block_0/spare_xz[19]
+ spare_logic_block_0/spare_xz[1] spare_logic_block_0/spare_xz[20] spare_logic_block_0/spare_xz[21]
+ spare_logic_block_0/spare_xz[22] spare_logic_block_0/spare_xz[23] spare_logic_block_0/spare_xz[24]
+ spare_logic_block_0/spare_xz[25] spare_logic_block_0/spare_xz[26] spare_logic_block_0/spare_xz[2]
+ spare_logic_block_0/spare_xz[3] spare_logic_block_0/spare_xz[4] spare_logic_block_0/spare_xz[5]
+ spare_logic_block_0/spare_xz[6] spare_logic_block_0/spare_xz[7] spare_logic_block_0/spare_xz[8]
+ spare_logic_block_0/spare_xz[9] VSUBS vccd_core spare_logic_block
Xsoc VSUBS vccd_core soc/core_clk soc/core_rstn soc/debug_in soc/debug_mode soc/debug_oeb
+ soc/debug_out soc/flash_clk soc/flash_csb soc/flash_io0_di soc/flash_io0_do soc/flash_io0_oeb
+ soc/flash_io1_di soc/flash_io1_do soc/flash_io1_oeb soc/flash_io2_di soc/flash_io2_do
+ soc/flash_io2_oeb soc/flash_io3_di soc/flash_io3_do soc/flash_io3_oeb soc/gpio_in_pad
+ soc/gpio_inenb_pad soc/gpio_mode0_pad soc/gpio_mode1_pad soc/gpio_out_pad soc/gpio_outenb_pad
+ soc/hk_ack_i soc/hk_cyc_o soc/hk_dat_i[0] soc/hk_dat_i[10] soc/hk_dat_i[11] soc/hk_dat_i[12]
+ soc/hk_dat_i[13] soc/hk_dat_i[14] soc/hk_dat_i[15] soc/hk_dat_i[16] soc/hk_dat_i[17]
+ soc/hk_dat_i[18] soc/hk_dat_i[19] soc/hk_dat_i[1] soc/hk_dat_i[20] soc/hk_dat_i[21]
+ soc/hk_dat_i[22] soc/hk_dat_i[23] soc/hk_dat_i[24] soc/hk_dat_i[25] soc/hk_dat_i[26]
+ soc/hk_dat_i[27] soc/hk_dat_i[28] soc/hk_dat_i[29] soc/hk_dat_i[2] soc/hk_dat_i[30]
+ soc/hk_dat_i[31] soc/hk_dat_i[3] soc/hk_dat_i[4] soc/hk_dat_i[5] soc/hk_dat_i[6]
+ soc/hk_dat_i[7] soc/hk_dat_i[8] soc/hk_dat_i[9] soc/hk_stb_o soc/irq[0] soc/irq[1]
+ soc/irq[2] soc/irq[3] soc/irq[4] soc/irq[5] soc/la_iena[0] soc/la_iena[100] soc/la_iena[101]
+ soc/la_iena[102] soc/la_iena[103] soc/la_iena[104] soc/la_iena[105] soc/la_iena[106]
+ soc/la_iena[107] soc/la_iena[108] soc/la_iena[109] soc/la_iena[10] soc/la_iena[110]
+ soc/la_iena[111] soc/la_iena[112] soc/la_iena[113] soc/la_iena[114] soc/la_iena[115]
+ soc/la_iena[116] soc/la_iena[117] soc/la_iena[118] soc/la_iena[119] soc/la_iena[11]
+ soc/la_iena[120] soc/la_iena[121] soc/la_iena[122] soc/la_iena[123] soc/la_iena[124]
+ soc/la_iena[125] soc/la_iena[126] soc/la_iena[127] soc/la_iena[12] soc/la_iena[13]
+ soc/la_iena[14] soc/la_iena[15] soc/la_iena[16] soc/la_iena[17] soc/la_iena[18]
+ soc/la_iena[19] soc/la_iena[1] soc/la_iena[20] soc/la_iena[21] soc/la_iena[22] soc/la_iena[23]
+ soc/la_iena[24] soc/la_iena[25] soc/la_iena[26] soc/la_iena[27] soc/la_iena[28]
+ soc/la_iena[29] soc/la_iena[2] soc/la_iena[30] soc/la_iena[31] soc/la_iena[32] soc/la_iena[33]
+ soc/la_iena[34] soc/la_iena[35] soc/la_iena[36] soc/la_iena[37] soc/la_iena[38]
+ soc/la_iena[39] soc/la_iena[3] soc/la_iena[40] soc/la_iena[41] soc/la_iena[42] soc/la_iena[43]
+ soc/la_iena[44] soc/la_iena[45] soc/la_iena[46] soc/la_iena[47] soc/la_iena[48]
+ soc/la_iena[49] soc/la_iena[4] soc/la_iena[50] soc/la_iena[51] soc/la_iena[52] soc/la_iena[53]
+ soc/la_iena[54] soc/la_iena[55] soc/la_iena[56] soc/la_iena[57] soc/la_iena[58]
+ soc/la_iena[59] soc/la_iena[5] soc/la_iena[60] soc/la_iena[61] soc/la_iena[62] soc/la_iena[63]
+ soc/la_iena[64] soc/la_iena[65] soc/la_iena[66] soc/la_iena[67] soc/la_iena[68]
+ soc/la_iena[69] soc/la_iena[6] soc/la_iena[70] soc/la_iena[71] soc/la_iena[72] soc/la_iena[73]
+ soc/la_iena[74] soc/la_iena[75] soc/la_iena[76] soc/la_iena[77] soc/la_iena[78]
+ soc/la_iena[79] soc/la_iena[7] soc/la_iena[80] soc/la_iena[81] soc/la_iena[82] soc/la_iena[83]
+ soc/la_iena[84] soc/la_iena[85] soc/la_iena[86] soc/la_iena[87] soc/la_iena[88]
+ soc/la_iena[89] soc/la_iena[8] soc/la_iena[90] soc/la_iena[91] soc/la_iena[92] soc/la_iena[93]
+ soc/la_iena[94] soc/la_iena[95] soc/la_iena[96] soc/la_iena[97] soc/la_iena[98]
+ soc/la_iena[99] soc/la_iena[9] soc/la_input[0] soc/la_input[100] soc/la_input[101]
+ soc/la_input[102] soc/la_input[103] soc/la_input[104] soc/la_input[105] soc/la_input[106]
+ soc/la_input[107] soc/la_input[108] soc/la_input[109] soc/la_input[10] soc/la_input[110]
+ soc/la_input[111] soc/la_input[112] soc/la_input[113] soc/la_input[114] soc/la_input[115]
+ soc/la_input[116] soc/la_input[117] soc/la_input[118] soc/la_input[119] soc/la_input[11]
+ soc/la_input[120] soc/la_input[121] soc/la_input[122] soc/la_input[123] soc/la_input[124]
+ soc/la_input[125] soc/la_input[126] soc/la_input[127] soc/la_input[12] soc/la_input[13]
+ soc/la_input[14] soc/la_input[15] soc/la_input[16] soc/la_input[17] soc/la_input[18]
+ soc/la_input[19] soc/la_input[1] soc/la_input[20] soc/la_input[21] soc/la_input[22]
+ soc/la_input[23] soc/la_input[24] soc/la_input[25] soc/la_input[26] soc/la_input[27]
+ soc/la_input[28] soc/la_input[29] soc/la_input[2] soc/la_input[30] soc/la_input[31]
+ soc/la_input[32] soc/la_input[33] soc/la_input[34] soc/la_input[35] soc/la_input[36]
+ soc/la_input[37] soc/la_input[38] soc/la_input[39] soc/la_input[3] soc/la_input[40]
+ soc/la_input[41] soc/la_input[42] soc/la_input[43] soc/la_input[44] soc/la_input[45]
+ soc/la_input[46] soc/la_input[47] soc/la_input[48] soc/la_input[49] soc/la_input[4]
+ soc/la_input[50] soc/la_input[51] soc/la_input[52] soc/la_input[53] soc/la_input[54]
+ soc/la_input[55] soc/la_input[56] soc/la_input[57] soc/la_input[58] soc/la_input[59]
+ soc/la_input[5] soc/la_input[60] soc/la_input[61] soc/la_input[62] soc/la_input[63]
+ soc/la_input[64] soc/la_input[65] soc/la_input[66] soc/la_input[67] soc/la_input[68]
+ soc/la_input[69] soc/la_input[6] soc/la_input[70] soc/la_input[71] soc/la_input[72]
+ soc/la_input[73] soc/la_input[74] soc/la_input[75] soc/la_input[76] soc/la_input[77]
+ soc/la_input[78] soc/la_input[79] soc/la_input[7] soc/la_input[80] soc/la_input[81]
+ soc/la_input[82] soc/la_input[83] soc/la_input[84] soc/la_input[85] soc/la_input[86]
+ soc/la_input[87] soc/la_input[88] soc/la_input[89] soc/la_input[8] soc/la_input[90]
+ soc/la_input[91] soc/la_input[92] soc/la_input[93] soc/la_input[94] soc/la_input[95]
+ soc/la_input[96] soc/la_input[97] soc/la_input[98] soc/la_input[99] soc/la_input[9]
+ soc/la_oenb[0] soc/la_oenb[100] soc/la_oenb[101] soc/la_oenb[102] soc/la_oenb[103]
+ soc/la_oenb[104] soc/la_oenb[105] soc/la_oenb[106] soc/la_oenb[107] soc/la_oenb[108]
+ soc/la_oenb[109] soc/la_oenb[10] soc/la_oenb[110] soc/la_oenb[111] soc/la_oenb[112]
+ soc/la_oenb[113] soc/la_oenb[114] soc/la_oenb[115] soc/la_oenb[116] soc/la_oenb[117]
+ soc/la_oenb[118] soc/la_oenb[119] soc/la_oenb[11] soc/la_oenb[120] soc/la_oenb[121]
+ soc/la_oenb[122] soc/la_oenb[123] soc/la_oenb[124] soc/la_oenb[125] soc/la_oenb[126]
+ soc/la_oenb[127] soc/la_oenb[12] soc/la_oenb[13] soc/la_oenb[14] soc/la_oenb[15]
+ soc/la_oenb[16] soc/la_oenb[17] soc/la_oenb[18] soc/la_oenb[19] soc/la_oenb[1] soc/la_oenb[20]
+ soc/la_oenb[21] soc/la_oenb[22] soc/la_oenb[23] soc/la_oenb[24] soc/la_oenb[25]
+ soc/la_oenb[26] soc/la_oenb[27] soc/la_oenb[28] soc/la_oenb[29] soc/la_oenb[2] soc/la_oenb[30]
+ soc/la_oenb[31] soc/la_oenb[32] soc/la_oenb[33] soc/la_oenb[34] soc/la_oenb[35]
+ soc/la_oenb[36] soc/la_oenb[37] soc/la_oenb[38] soc/la_oenb[39] soc/la_oenb[3] soc/la_oenb[40]
+ soc/la_oenb[41] soc/la_oenb[42] soc/la_oenb[43] soc/la_oenb[44] soc/la_oenb[45]
+ soc/la_oenb[46] soc/la_oenb[47] soc/la_oenb[48] soc/la_oenb[49] soc/la_oenb[4] soc/la_oenb[50]
+ soc/la_oenb[51] soc/la_oenb[52] soc/la_oenb[53] soc/la_oenb[54] soc/la_oenb[55]
+ soc/la_oenb[56] soc/la_oenb[57] soc/la_oenb[58] soc/la_oenb[59] soc/la_oenb[5] soc/la_oenb[60]
+ soc/la_oenb[61] soc/la_oenb[62] soc/la_oenb[63] soc/la_oenb[64] soc/la_oenb[65]
+ soc/la_oenb[66] soc/la_oenb[67] soc/la_oenb[68] soc/la_oenb[69] soc/la_oenb[6] soc/la_oenb[70]
+ soc/la_oenb[71] soc/la_oenb[72] soc/la_oenb[73] soc/la_oenb[74] soc/la_oenb[75]
+ soc/la_oenb[76] soc/la_oenb[77] soc/la_oenb[78] soc/la_oenb[79] soc/la_oenb[7] soc/la_oenb[80]
+ soc/la_oenb[81] soc/la_oenb[82] soc/la_oenb[83] soc/la_oenb[84] soc/la_oenb[85]
+ soc/la_oenb[86] soc/la_oenb[87] soc/la_oenb[88] soc/la_oenb[89] soc/la_oenb[8] soc/la_oenb[90]
+ soc/la_oenb[91] soc/la_oenb[92] soc/la_oenb[93] soc/la_oenb[94] soc/la_oenb[95]
+ soc/la_oenb[96] soc/la_oenb[97] soc/la_oenb[98] soc/la_oenb[99] soc/la_oenb[9] soc/la_output[0]
+ soc/la_output[100] soc/la_output[101] soc/la_output[102] soc/la_output[103] soc/la_output[104]
+ soc/la_output[105] soc/la_output[106] soc/la_output[107] soc/la_output[108] soc/la_output[109]
+ soc/la_output[10] soc/la_output[110] soc/la_output[111] soc/la_output[112] soc/la_output[113]
+ soc/la_output[114] soc/la_output[115] soc/la_output[116] soc/la_output[117] soc/la_output[118]
+ soc/la_output[119] soc/la_output[11] soc/la_output[120] soc/la_output[121] soc/la_output[122]
+ soc/la_output[123] soc/la_output[124] soc/la_output[125] soc/la_output[126] soc/la_output[127]
+ soc/la_output[12] soc/la_output[13] soc/la_output[14] soc/la_output[15] soc/la_output[16]
+ soc/la_output[17] soc/la_output[18] soc/la_output[19] soc/la_output[1] soc/la_output[20]
+ soc/la_output[21] soc/la_output[22] soc/la_output[23] soc/la_output[24] soc/la_output[25]
+ soc/la_output[26] soc/la_output[27] soc/la_output[28] soc/la_output[29] soc/la_output[2]
+ soc/la_output[30] soc/la_output[31] soc/la_output[32] soc/la_output[33] soc/la_output[34]
+ soc/la_output[35] soc/la_output[36] soc/la_output[37] soc/la_output[38] soc/la_output[39]
+ soc/la_output[3] soc/la_output[40] soc/la_output[41] soc/la_output[42] soc/la_output[43]
+ soc/la_output[44] soc/la_output[45] soc/la_output[46] soc/la_output[47] soc/la_output[48]
+ soc/la_output[49] soc/la_output[4] soc/la_output[50] soc/la_output[51] soc/la_output[52]
+ soc/la_output[53] soc/la_output[54] soc/la_output[55] soc/la_output[56] soc/la_output[57]
+ soc/la_output[58] soc/la_output[59] soc/la_output[5] soc/la_output[60] soc/la_output[61]
+ soc/la_output[62] soc/la_output[63] soc/la_output[64] soc/la_output[65] soc/la_output[66]
+ soc/la_output[67] soc/la_output[68] soc/la_output[69] soc/la_output[6] soc/la_output[70]
+ soc/la_output[71] soc/la_output[72] soc/la_output[73] soc/la_output[74] soc/la_output[75]
+ soc/la_output[76] soc/la_output[77] soc/la_output[78] soc/la_output[79] soc/la_output[7]
+ soc/la_output[80] soc/la_output[81] soc/la_output[82] soc/la_output[83] soc/la_output[84]
+ soc/la_output[85] soc/la_output[86] soc/la_output[87] soc/la_output[88] soc/la_output[89]
+ soc/la_output[8] soc/la_output[90] soc/la_output[91] soc/la_output[92] soc/la_output[93]
+ soc/la_output[94] soc/la_output[95] soc/la_output[96] soc/la_output[97] soc/la_output[98]
+ soc/la_output[99] soc/la_output[9] soc/mprj_ack_i soc/mprj_adr_o[0] soc/mprj_adr_o[10]
+ soc/mprj_adr_o[11] soc/mprj_adr_o[12] soc/mprj_adr_o[13] soc/mprj_adr_o[14] soc/mprj_adr_o[15]
+ soc/mprj_adr_o[16] soc/mprj_adr_o[17] soc/mprj_adr_o[18] soc/mprj_adr_o[19] soc/mprj_adr_o[1]
+ soc/mprj_adr_o[20] soc/mprj_adr_o[21] soc/mprj_adr_o[22] soc/mprj_adr_o[23] soc/mprj_adr_o[24]
+ soc/mprj_adr_o[25] soc/mprj_adr_o[26] soc/mprj_adr_o[27] soc/mprj_adr_o[28] soc/mprj_adr_o[29]
+ soc/mprj_adr_o[2] soc/mprj_adr_o[30] soc/mprj_adr_o[31] soc/mprj_adr_o[3] soc/mprj_adr_o[4]
+ soc/mprj_adr_o[5] soc/mprj_adr_o[6] soc/mprj_adr_o[7] soc/mprj_adr_o[8] soc/mprj_adr_o[9]
+ soc/mprj_cyc_o soc/mprj_dat_i[0] soc/mprj_dat_i[10] soc/mprj_dat_i[11] soc/mprj_dat_i[12]
+ soc/mprj_dat_i[13] soc/mprj_dat_i[14] soc/mprj_dat_i[15] soc/mprj_dat_i[16] soc/mprj_dat_i[17]
+ soc/mprj_dat_i[18] soc/mprj_dat_i[19] soc/mprj_dat_i[1] soc/mprj_dat_i[20] soc/mprj_dat_i[21]
+ soc/mprj_dat_i[22] soc/mprj_dat_i[23] soc/mprj_dat_i[24] soc/mprj_dat_i[25] soc/mprj_dat_i[26]
+ soc/mprj_dat_i[27] soc/mprj_dat_i[28] soc/mprj_dat_i[29] soc/mprj_dat_i[2] soc/mprj_dat_i[30]
+ soc/mprj_dat_i[31] soc/mprj_dat_i[3] soc/mprj_dat_i[4] soc/mprj_dat_i[5] soc/mprj_dat_i[6]
+ soc/mprj_dat_i[7] soc/mprj_dat_i[8] soc/mprj_dat_i[9] soc/mprj_dat_o[0] soc/mprj_dat_o[10]
+ soc/mprj_dat_o[11] soc/mprj_dat_o[12] soc/mprj_dat_o[13] soc/mprj_dat_o[14] soc/mprj_dat_o[15]
+ soc/mprj_dat_o[16] soc/mprj_dat_o[17] soc/mprj_dat_o[18] soc/mprj_dat_o[19] soc/mprj_dat_o[1]
+ soc/mprj_dat_o[20] soc/mprj_dat_o[21] soc/mprj_dat_o[22] soc/mprj_dat_o[23] soc/mprj_dat_o[24]
+ soc/mprj_dat_o[25] soc/mprj_dat_o[26] soc/mprj_dat_o[27] soc/mprj_dat_o[28] soc/mprj_dat_o[29]
+ soc/mprj_dat_o[2] soc/mprj_dat_o[30] soc/mprj_dat_o[31] soc/mprj_dat_o[3] soc/mprj_dat_o[4]
+ soc/mprj_dat_o[5] soc/mprj_dat_o[6] soc/mprj_dat_o[7] soc/mprj_dat_o[8] soc/mprj_dat_o[9]
+ soc/mprj_sel_o[0] soc/mprj_sel_o[1] soc/mprj_sel_o[2] soc/mprj_sel_o[3] soc/mprj_stb_o
+ soc/mprj_wb_iena soc/mprj_we_o soc/qspi_enabled soc/ser_rx soc/ser_tx soc/spi_csb
+ soc/spi_enabled soc/spi_sck soc/spi_sdi soc/spi_sdo soc/spi_sdoenb soc/sram_ro_addr[0]
+ soc/sram_ro_addr[1] soc/sram_ro_addr[2] soc/sram_ro_addr[3] soc/sram_ro_addr[4]
+ soc/sram_ro_addr[5] soc/sram_ro_addr[6] soc/sram_ro_addr[7] soc/sram_ro_clk soc/sram_ro_csb
+ soc/sram_ro_data[0] soc/sram_ro_data[10] soc/sram_ro_data[11] soc/sram_ro_data[12]
+ soc/sram_ro_data[13] soc/sram_ro_data[14] soc/sram_ro_data[15] soc/sram_ro_data[16]
+ soc/sram_ro_data[17] soc/sram_ro_data[18] soc/sram_ro_data[19] soc/sram_ro_data[1]
+ soc/sram_ro_data[20] soc/sram_ro_data[21] soc/sram_ro_data[22] soc/sram_ro_data[23]
+ soc/sram_ro_data[24] soc/sram_ro_data[25] soc/sram_ro_data[26] soc/sram_ro_data[27]
+ soc/sram_ro_data[28] soc/sram_ro_data[29] soc/sram_ro_data[2] soc/sram_ro_data[30]
+ soc/sram_ro_data[31] soc/sram_ro_data[3] soc/sram_ro_data[4] soc/sram_ro_data[5]
+ soc/sram_ro_data[6] soc/sram_ro_data[7] soc/sram_ro_data[8] soc/sram_ro_data[9]
+ soc/trap soc/uart_enabled soc/user_irq_ena[0] soc/user_irq_ena[1] soc/user_irq_ena[2]
+ mgmt_core_wrapper
Xgpio_defaults_block_14 VSUBS gpio_defaults_block_14/gpio_defaults[0] gpio_defaults_block_14/gpio_defaults[10]
+ gpio_defaults_block_14/gpio_defaults[11] gpio_defaults_block_14/gpio_defaults[12]
+ gpio_defaults_block_14/gpio_defaults[1] gpio_defaults_block_14/gpio_defaults[2]
+ gpio_defaults_block_14/gpio_defaults[3] gpio_defaults_block_14/gpio_defaults[4]
+ gpio_defaults_block_14/gpio_defaults[5] gpio_defaults_block_14/gpio_defaults[6]
+ gpio_defaults_block_14/gpio_defaults[7] gpio_defaults_block_14/gpio_defaults[8]
+ gpio_defaults_block_14/gpio_defaults[9] vccd_core gpio_defaults_block
Xgpio_defaults_block_25 VSUBS gpio_defaults_block_25/gpio_defaults[0] gpio_defaults_block_25/gpio_defaults[10]
+ gpio_defaults_block_25/gpio_defaults[11] gpio_defaults_block_25/gpio_defaults[12]
+ gpio_defaults_block_25/gpio_defaults[1] gpio_defaults_block_25/gpio_defaults[2]
+ gpio_defaults_block_25/gpio_defaults[3] gpio_defaults_block_25/gpio_defaults[4]
+ gpio_defaults_block_25/gpio_defaults[5] gpio_defaults_block_25/gpio_defaults[6]
+ gpio_defaults_block_25/gpio_defaults[7] gpio_defaults_block_25/gpio_defaults[8]
+ gpio_defaults_block_25/gpio_defaults[9] vccd_core gpio_defaults_block
Xgpio_control_in_2\[9\] gpio_defaults_block_28/gpio_defaults[0] gpio_defaults_block_28/gpio_defaults[10]
+ gpio_defaults_block_28/gpio_defaults[11] gpio_defaults_block_28/gpio_defaults[12]
+ gpio_defaults_block_28/gpio_defaults[1] gpio_defaults_block_28/gpio_defaults[2]
+ gpio_defaults_block_28/gpio_defaults[3] gpio_defaults_block_28/gpio_defaults[4]
+ gpio_defaults_block_28/gpio_defaults[5] gpio_defaults_block_28/gpio_defaults[6]
+ gpio_defaults_block_28/gpio_defaults[7] gpio_defaults_block_28/gpio_defaults[8]
+ gpio_defaults_block_28/gpio_defaults[9] housekeeping/mgmt_gpio_in[28] gpio_control_in_2\[9\]/one
+ housekeeping/mgmt_gpio_in[28] gpio_control_in_2\[9\]/one padframe/mprj_io_analog_en[28]
+ padframe/mprj_io_analog_pol[28] padframe/mprj_io_analog_sel[28] padframe/mprj_io_dm[84]
+ padframe/mprj_io_dm[85] padframe/mprj_io_dm[86] padframe/mprj_io_holdover[28] padframe/mprj_io_ib_mode_sel[28]
+ padframe/mprj_io_in[28] padframe/mprj_io_inp_dis[28] padframe/mprj_io_out[28] padframe/mprj_io_oeb[28]
+ padframe/mprj_io_slow_sel[28] padframe/mprj_io_vtrip_sel[28] gpio_control_in_2\[9\]/resetn
+ gpio_control_in_2\[8\]/resetn gpio_control_in_2\[9\]/serial_clock gpio_control_in_2\[8\]/serial_clock
+ gpio_control_in_2\[9\]/serial_data_in gpio_control_in_2\[8\]/serial_data_in gpio_control_in_2\[9\]/serial_load
+ gpio_control_in_2\[8\]/serial_load mprj/io_in[28] mprj/io_oeb[28] mprj/io_out[28]
+ vccd1_core VSUBS gpio_control_in_2\[9\]/zero dw_8741_677338# vccd_core vssd1_core
+ gpio_control_block
Xgpio_defaults_block_36 VSUBS gpio_defaults_block_36/gpio_defaults[0] gpio_defaults_block_36/gpio_defaults[10]
+ gpio_defaults_block_36/gpio_defaults[11] gpio_defaults_block_36/gpio_defaults[12]
+ gpio_defaults_block_36/gpio_defaults[1] gpio_defaults_block_36/gpio_defaults[2]
+ gpio_defaults_block_36/gpio_defaults[3] gpio_defaults_block_36/gpio_defaults[4]
+ gpio_defaults_block_36/gpio_defaults[5] gpio_defaults_block_36/gpio_defaults[6]
+ gpio_defaults_block_36/gpio_defaults[7] gpio_defaults_block_36/gpio_defaults[8]
+ gpio_defaults_block_36/gpio_defaults[9] vccd_core gpio_defaults_block
Xspare_logic_block_1 spare_logic_block_1/spare_xfq[0] spare_logic_block_1/spare_xfq[1]
+ spare_logic_block_1/spare_xfqn[0] spare_logic_block_1/spare_xfqn[1] spare_logic_block_1/spare_xi[0]
+ spare_logic_block_1/spare_xi[1] spare_logic_block_1/spare_xi[2] spare_logic_block_1/spare_xi[3]
+ spare_logic_block_1/spare_xib spare_logic_block_1/spare_xmx[0] spare_logic_block_1/spare_xmx[1]
+ spare_logic_block_1/spare_xna[0] spare_logic_block_1/spare_xna[1] spare_logic_block_1/spare_xno[0]
+ spare_logic_block_1/spare_xno[1] spare_logic_block_1/spare_xz[0] spare_logic_block_1/spare_xz[10]
+ spare_logic_block_1/spare_xz[11] spare_logic_block_1/spare_xz[12] spare_logic_block_1/spare_xz[13]
+ spare_logic_block_1/spare_xz[14] spare_logic_block_1/spare_xz[15] spare_logic_block_1/spare_xz[16]
+ spare_logic_block_1/spare_xz[17] spare_logic_block_1/spare_xz[18] spare_logic_block_1/spare_xz[19]
+ spare_logic_block_1/spare_xz[1] spare_logic_block_1/spare_xz[20] spare_logic_block_1/spare_xz[21]
+ spare_logic_block_1/spare_xz[22] spare_logic_block_1/spare_xz[23] spare_logic_block_1/spare_xz[24]
+ spare_logic_block_1/spare_xz[25] spare_logic_block_1/spare_xz[26] spare_logic_block_1/spare_xz[2]
+ spare_logic_block_1/spare_xz[3] spare_logic_block_1/spare_xz[4] spare_logic_block_1/spare_xz[5]
+ spare_logic_block_1/spare_xz[6] spare_logic_block_1/spare_xz[7] spare_logic_block_1/spare_xz[8]
+ spare_logic_block_1/spare_xz[9] VSUBS vccd_core spare_logic_block
Xgpio_defaults_block_15 VSUBS gpio_defaults_block_15/gpio_defaults[0] gpio_defaults_block_15/gpio_defaults[10]
+ gpio_defaults_block_15/gpio_defaults[11] gpio_defaults_block_15/gpio_defaults[12]
+ gpio_defaults_block_15/gpio_defaults[1] gpio_defaults_block_15/gpio_defaults[2]
+ gpio_defaults_block_15/gpio_defaults[3] gpio_defaults_block_15/gpio_defaults[4]
+ gpio_defaults_block_15/gpio_defaults[5] gpio_defaults_block_15/gpio_defaults[6]
+ gpio_defaults_block_15/gpio_defaults[7] gpio_defaults_block_15/gpio_defaults[8]
+ gpio_defaults_block_15/gpio_defaults[9] vccd_core gpio_defaults_block
Xgpio_control_in_1\[4\] gpio_defaults_block_12/gpio_defaults[0] gpio_defaults_block_12/gpio_defaults[10]
+ gpio_defaults_block_12/gpio_defaults[11] gpio_defaults_block_12/gpio_defaults[12]
+ gpio_defaults_block_12/gpio_defaults[1] gpio_defaults_block_12/gpio_defaults[2]
+ gpio_defaults_block_12/gpio_defaults[3] gpio_defaults_block_12/gpio_defaults[4]
+ gpio_defaults_block_12/gpio_defaults[5] gpio_defaults_block_12/gpio_defaults[6]
+ gpio_defaults_block_12/gpio_defaults[7] gpio_defaults_block_12/gpio_defaults[8]
+ gpio_defaults_block_12/gpio_defaults[9] housekeeping/mgmt_gpio_in[12] gpio_control_in_1\[4\]/one
+ housekeeping/mgmt_gpio_in[12] gpio_control_in_1\[4\]/one padframe/mprj_io_analog_en[12]
+ padframe/mprj_io_analog_pol[12] padframe/mprj_io_analog_sel[12] padframe/mprj_io_dm[36]
+ padframe/mprj_io_dm[37] padframe/mprj_io_dm[38] padframe/mprj_io_holdover[12] padframe/mprj_io_ib_mode_sel[12]
+ padframe/mprj_io_in[12] padframe/mprj_io_inp_dis[12] padframe/mprj_io_out[12] padframe/mprj_io_oeb[12]
+ padframe/mprj_io_slow_sel[12] padframe/mprj_io_vtrip_sel[12] gpio_control_in_1\[4\]/resetn
+ gpio_control_in_1\[5\]/resetn gpio_control_in_1\[4\]/serial_clock gpio_control_in_1\[5\]/serial_clock
+ gpio_control_in_1\[4\]/serial_data_in gpio_control_in_1\[5\]/serial_data_in gpio_control_in_1\[4\]/serial_load
+ gpio_control_in_1\[5\]/serial_load mprj/io_in[12] mprj/io_oeb[12] mprj/io_out[12]
+ vccd1_core VSUBS gpio_control_in_1\[4\]/zero dw_707553_705738# vccd_core vssd1_core
+ gpio_control_block
Xgpio_defaults_block_26 VSUBS gpio_defaults_block_26/gpio_defaults[0] gpio_defaults_block_26/gpio_defaults[10]
+ gpio_defaults_block_26/gpio_defaults[11] gpio_defaults_block_26/gpio_defaults[12]
+ gpio_defaults_block_26/gpio_defaults[1] gpio_defaults_block_26/gpio_defaults[2]
+ gpio_defaults_block_26/gpio_defaults[3] gpio_defaults_block_26/gpio_defaults[4]
+ gpio_defaults_block_26/gpio_defaults[5] gpio_defaults_block_26/gpio_defaults[6]
+ gpio_defaults_block_26/gpio_defaults[7] gpio_defaults_block_26/gpio_defaults[8]
+ gpio_defaults_block_26/gpio_defaults[9] vccd_core gpio_defaults_block
Xspare_logic_block_2 spare_logic_block_2/spare_xfq[0] spare_logic_block_2/spare_xfq[1]
+ spare_logic_block_2/spare_xfqn[0] spare_logic_block_2/spare_xfqn[1] spare_logic_block_2/spare_xi[0]
+ spare_logic_block_2/spare_xi[1] spare_logic_block_2/spare_xi[2] spare_logic_block_2/spare_xi[3]
+ spare_logic_block_2/spare_xib spare_logic_block_2/spare_xmx[0] spare_logic_block_2/spare_xmx[1]
+ spare_logic_block_2/spare_xna[0] spare_logic_block_2/spare_xna[1] spare_logic_block_2/spare_xno[0]
+ spare_logic_block_2/spare_xno[1] spare_logic_block_2/spare_xz[0] spare_logic_block_2/spare_xz[10]
+ spare_logic_block_2/spare_xz[11] spare_logic_block_2/spare_xz[12] spare_logic_block_2/spare_xz[13]
+ spare_logic_block_2/spare_xz[14] spare_logic_block_2/spare_xz[15] spare_logic_block_2/spare_xz[16]
+ spare_logic_block_2/spare_xz[17] spare_logic_block_2/spare_xz[18] spare_logic_block_2/spare_xz[19]
+ spare_logic_block_2/spare_xz[1] spare_logic_block_2/spare_xz[20] spare_logic_block_2/spare_xz[21]
+ spare_logic_block_2/spare_xz[22] spare_logic_block_2/spare_xz[23] spare_logic_block_2/spare_xz[24]
+ spare_logic_block_2/spare_xz[25] spare_logic_block_2/spare_xz[26] spare_logic_block_2/spare_xz[2]
+ spare_logic_block_2/spare_xz[3] spare_logic_block_2/spare_xz[4] spare_logic_block_2/spare_xz[5]
+ spare_logic_block_2/spare_xz[6] spare_logic_block_2/spare_xz[7] spare_logic_block_2/spare_xz[8]
+ spare_logic_block_2/spare_xz[9] VSUBS vccd_core spare_logic_block
Xgpio_defaults_block_37 VSUBS gpio_defaults_block_37/gpio_defaults[0] gpio_defaults_block_37/gpio_defaults[10]
+ gpio_defaults_block_37/gpio_defaults[11] gpio_defaults_block_37/gpio_defaults[12]
+ gpio_defaults_block_37/gpio_defaults[1] gpio_defaults_block_37/gpio_defaults[2]
+ gpio_defaults_block_37/gpio_defaults[3] gpio_defaults_block_37/gpio_defaults[4]
+ gpio_defaults_block_37/gpio_defaults[5] gpio_defaults_block_37/gpio_defaults[6]
+ gpio_defaults_block_37/gpio_defaults[7] gpio_defaults_block_37/gpio_defaults[8]
+ gpio_defaults_block_37/gpio_defaults[9] vccd_core gpio_defaults_block
Xpor vccd_core por/vdd3v3 por/vss3v3 por/porb_h por/por_l por/porb_l VSUBS simple_por
Xgpio_defaults_block_16 VSUBS gpio_defaults_block_16/gpio_defaults[0] gpio_defaults_block_16/gpio_defaults[10]
+ gpio_defaults_block_16/gpio_defaults[11] gpio_defaults_block_16/gpio_defaults[12]
+ gpio_defaults_block_16/gpio_defaults[1] gpio_defaults_block_16/gpio_defaults[2]
+ gpio_defaults_block_16/gpio_defaults[3] gpio_defaults_block_16/gpio_defaults[4]
+ gpio_defaults_block_16/gpio_defaults[5] gpio_defaults_block_16/gpio_defaults[6]
+ gpio_defaults_block_16/gpio_defaults[7] gpio_defaults_block_16/gpio_defaults[8]
+ gpio_defaults_block_16/gpio_defaults[9] vccd_core gpio_defaults_block
Xgpio_defaults_block_27 VSUBS gpio_defaults_block_27/gpio_defaults[0] gpio_defaults_block_27/gpio_defaults[10]
+ gpio_defaults_block_27/gpio_defaults[11] gpio_defaults_block_27/gpio_defaults[12]
+ gpio_defaults_block_27/gpio_defaults[1] gpio_defaults_block_27/gpio_defaults[2]
+ gpio_defaults_block_27/gpio_defaults[3] gpio_defaults_block_27/gpio_defaults[4]
+ gpio_defaults_block_27/gpio_defaults[5] gpio_defaults_block_27/gpio_defaults[6]
+ gpio_defaults_block_27/gpio_defaults[7] gpio_defaults_block_27/gpio_defaults[8]
+ gpio_defaults_block_27/gpio_defaults[9] vccd_core gpio_defaults_block
Xgpio_control_in_2\[12\] gpio_defaults_block_31/gpio_defaults[0] gpio_defaults_block_31/gpio_defaults[10]
+ gpio_defaults_block_31/gpio_defaults[11] gpio_defaults_block_31/gpio_defaults[12]
+ gpio_defaults_block_31/gpio_defaults[1] gpio_defaults_block_31/gpio_defaults[2]
+ gpio_defaults_block_31/gpio_defaults[3] gpio_defaults_block_31/gpio_defaults[4]
+ gpio_defaults_block_31/gpio_defaults[5] gpio_defaults_block_31/gpio_defaults[6]
+ gpio_defaults_block_31/gpio_defaults[7] gpio_defaults_block_31/gpio_defaults[8]
+ gpio_defaults_block_31/gpio_defaults[9] housekeeping/mgmt_gpio_in[31] gpio_control_in_2\[12\]/one
+ housekeeping/mgmt_gpio_in[31] gpio_control_in_2\[12\]/one padframe/mprj_io_analog_en[31]
+ padframe/mprj_io_analog_pol[31] padframe/mprj_io_analog_sel[31] padframe/mprj_io_dm[93]
+ padframe/mprj_io_dm[94] padframe/mprj_io_dm[95] padframe/mprj_io_holdover[31] padframe/mprj_io_ib_mode_sel[31]
+ padframe/mprj_io_in[31] padframe/mprj_io_inp_dis[31] padframe/mprj_io_out[31] padframe/mprj_io_oeb[31]
+ padframe/mprj_io_slow_sel[31] padframe/mprj_io_vtrip_sel[31] gpio_control_in_2\[12\]/resetn
+ gpio_control_in_2\[11\]/resetn gpio_control_in_2\[12\]/serial_clock gpio_control_in_2\[11\]/serial_clock
+ gpio_control_in_2\[12\]/serial_data_in gpio_control_in_2\[11\]/serial_data_in gpio_control_in_2\[12\]/serial_load
+ gpio_control_in_2\[11\]/serial_load mprj/io_in[31] mprj/io_oeb[31] mprj/io_out[31]
+ vccd1_core VSUBS gpio_control_in_2\[12\]/zero dw_8741_547738# vccd_core vssd1_core
+ gpio_control_block
Xgpio_control_in_1a\[1\] gpio_defaults_block_3/gpio_defaults[0] gpio_defaults_block_3/gpio_defaults[10]
+ gpio_defaults_block_3/gpio_defaults[11] gpio_defaults_block_3/gpio_defaults[12]
+ gpio_defaults_block_3/gpio_defaults[1] gpio_defaults_block_3/gpio_defaults[2] gpio_defaults_block_3/gpio_defaults[3]
+ gpio_defaults_block_3/gpio_defaults[4] gpio_defaults_block_3/gpio_defaults[5] gpio_defaults_block_3/gpio_defaults[6]
+ gpio_defaults_block_3/gpio_defaults[7] gpio_defaults_block_3/gpio_defaults[8] gpio_defaults_block_3/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[3] gpio_control_in_1a\[1\]/one housekeeping/mgmt_gpio_in[3]
+ gpio_control_in_1a\[1\]/one padframe/mprj_io_analog_en[3] padframe/mprj_io_analog_pol[3]
+ padframe/mprj_io_analog_sel[3] padframe/mprj_io_dm[9] padframe/mprj_io_dm[10] padframe/mprj_io_dm[11]
+ padframe/mprj_io_holdover[3] padframe/mprj_io_ib_mode_sel[3] padframe/mprj_io_in[3]
+ padframe/mprj_io_inp_dis[3] padframe/mprj_io_out[3] padframe/mprj_io_oeb[3] padframe/mprj_io_slow_sel[3]
+ padframe/mprj_io_vtrip_sel[3] gpio_control_in_1a\[1\]/resetn gpio_control_in_1a\[2\]/resetn
+ gpio_control_in_1a\[1\]/serial_clock gpio_control_in_1a\[2\]/serial_clock gpio_control_in_1a\[1\]/serial_data_in
+ gpio_control_in_1a\[2\]/serial_data_in gpio_control_in_1a\[1\]/serial_load gpio_control_in_1a\[2\]/serial_load
+ mprj/io_in[3] mprj/io_oeb[3] mprj/io_out[3] vccd1_core VSUBS gpio_control_in_1a\[1\]/zero
+ dw_707553_257938# vccd_core vssd1_core gpio_control_block
Xspare_logic_block_3 spare_logic_block_3/spare_xfq[0] spare_logic_block_3/spare_xfq[1]
+ spare_logic_block_3/spare_xfqn[0] spare_logic_block_3/spare_xfqn[1] spare_logic_block_3/spare_xi[0]
+ spare_logic_block_3/spare_xi[1] spare_logic_block_3/spare_xi[2] spare_logic_block_3/spare_xi[3]
+ spare_logic_block_3/spare_xib spare_logic_block_3/spare_xmx[0] spare_logic_block_3/spare_xmx[1]
+ spare_logic_block_3/spare_xna[0] spare_logic_block_3/spare_xna[1] spare_logic_block_3/spare_xno[0]
+ spare_logic_block_3/spare_xno[1] spare_logic_block_3/spare_xz[0] spare_logic_block_3/spare_xz[10]
+ spare_logic_block_3/spare_xz[11] spare_logic_block_3/spare_xz[12] spare_logic_block_3/spare_xz[13]
+ spare_logic_block_3/spare_xz[14] spare_logic_block_3/spare_xz[15] spare_logic_block_3/spare_xz[16]
+ spare_logic_block_3/spare_xz[17] spare_logic_block_3/spare_xz[18] spare_logic_block_3/spare_xz[19]
+ spare_logic_block_3/spare_xz[1] spare_logic_block_3/spare_xz[20] spare_logic_block_3/spare_xz[21]
+ spare_logic_block_3/spare_xz[22] spare_logic_block_3/spare_xz[23] spare_logic_block_3/spare_xz[24]
+ spare_logic_block_3/spare_xz[25] spare_logic_block_3/spare_xz[26] spare_logic_block_3/spare_xz[2]
+ spare_logic_block_3/spare_xz[3] spare_logic_block_3/spare_xz[4] spare_logic_block_3/spare_xz[5]
+ spare_logic_block_3/spare_xz[6] spare_logic_block_3/spare_xz[7] spare_logic_block_3/spare_xz[8]
+ spare_logic_block_3/spare_xz[9] VSUBS vccd_core spare_logic_block
Xgpio_defaults_block_17 VSUBS gpio_defaults_block_17/gpio_defaults[0] gpio_defaults_block_17/gpio_defaults[10]
+ gpio_defaults_block_17/gpio_defaults[11] gpio_defaults_block_17/gpio_defaults[12]
+ gpio_defaults_block_17/gpio_defaults[1] gpio_defaults_block_17/gpio_defaults[2]
+ gpio_defaults_block_17/gpio_defaults[3] gpio_defaults_block_17/gpio_defaults[4]
+ gpio_defaults_block_17/gpio_defaults[5] gpio_defaults_block_17/gpio_defaults[6]
+ gpio_defaults_block_17/gpio_defaults[7] gpio_defaults_block_17/gpio_defaults[8]
+ gpio_defaults_block_17/gpio_defaults[9] vccd_core gpio_defaults_block
Xgpio_control_in_2\[7\] gpio_defaults_block_26/gpio_defaults[0] gpio_defaults_block_26/gpio_defaults[10]
+ gpio_defaults_block_26/gpio_defaults[11] gpio_defaults_block_26/gpio_defaults[12]
+ gpio_defaults_block_26/gpio_defaults[1] gpio_defaults_block_26/gpio_defaults[2]
+ gpio_defaults_block_26/gpio_defaults[3] gpio_defaults_block_26/gpio_defaults[4]
+ gpio_defaults_block_26/gpio_defaults[5] gpio_defaults_block_26/gpio_defaults[6]
+ gpio_defaults_block_26/gpio_defaults[7] gpio_defaults_block_26/gpio_defaults[8]
+ gpio_defaults_block_26/gpio_defaults[9] housekeeping/mgmt_gpio_in[26] gpio_control_in_2\[7\]/one
+ housekeeping/mgmt_gpio_in[26] gpio_control_in_2\[7\]/one padframe/mprj_io_analog_en[26]
+ padframe/mprj_io_analog_pol[26] padframe/mprj_io_analog_sel[26] padframe/mprj_io_dm[78]
+ padframe/mprj_io_dm[79] padframe/mprj_io_dm[80] padframe/mprj_io_holdover[26] padframe/mprj_io_ib_mode_sel[26]
+ padframe/mprj_io_in[26] padframe/mprj_io_inp_dis[26] padframe/mprj_io_out[26] padframe/mprj_io_oeb[26]
+ padframe/mprj_io_slow_sel[26] padframe/mprj_io_vtrip_sel[26] gpio_control_in_2\[7\]/resetn
+ gpio_control_in_2\[6\]/resetn gpio_control_in_2\[7\]/serial_clock gpio_control_in_2\[6\]/serial_clock
+ gpio_control_in_2\[7\]/serial_data_in gpio_control_in_2\[6\]/serial_data_in gpio_control_in_2\[7\]/serial_load
+ gpio_control_in_2\[6\]/serial_load mprj/io_in[26] mprj/io_oeb[26] mprj/io_out[26]
+ vccd1_core VSUBS gpio_control_in_2\[7\]/zero dw_8741_763738# vccd_core vssd1_core
+ gpio_control_block
Xgpio_defaults_block_28 VSUBS gpio_defaults_block_28/gpio_defaults[0] gpio_defaults_block_28/gpio_defaults[10]
+ gpio_defaults_block_28/gpio_defaults[11] gpio_defaults_block_28/gpio_defaults[12]
+ gpio_defaults_block_28/gpio_defaults[1] gpio_defaults_block_28/gpio_defaults[2]
+ gpio_defaults_block_28/gpio_defaults[3] gpio_defaults_block_28/gpio_defaults[4]
+ gpio_defaults_block_28/gpio_defaults[5] gpio_defaults_block_28/gpio_defaults[6]
+ gpio_defaults_block_28/gpio_defaults[7] gpio_defaults_block_28/gpio_defaults[8]
+ gpio_defaults_block_28/gpio_defaults[9] vccd_core gpio_defaults_block
Xclocking soc/core_clk pll/osc clocking/ext_clk_sel housekeeping/reset pll/clockp[1]
+ pll/clockp[0] pll/resetb soc/core_rstn clocking/sel2[0] clocking/sel2[1] clocking/sel2[2]
+ clocking/sel[0] clocking/sel[1] clocking/sel[2] clocking/user_clk vccd_core VSUBS
+ caravel_clocking
Xgpio_defaults_block_18 VSUBS gpio_defaults_block_18/gpio_defaults[0] gpio_defaults_block_18/gpio_defaults[10]
+ gpio_defaults_block_18/gpio_defaults[11] gpio_defaults_block_18/gpio_defaults[12]
+ gpio_defaults_block_18/gpio_defaults[1] gpio_defaults_block_18/gpio_defaults[2]
+ gpio_defaults_block_18/gpio_defaults[3] gpio_defaults_block_18/gpio_defaults[4]
+ gpio_defaults_block_18/gpio_defaults[5] gpio_defaults_block_18/gpio_defaults[6]
+ gpio_defaults_block_18/gpio_defaults[7] gpio_defaults_block_18/gpio_defaults[8]
+ gpio_defaults_block_18/gpio_defaults[9] vccd_core gpio_defaults_block
Xgpio_defaults_block_19 VSUBS gpio_defaults_block_19/gpio_defaults[0] gpio_defaults_block_19/gpio_defaults[10]
+ gpio_defaults_block_19/gpio_defaults[11] gpio_defaults_block_19/gpio_defaults[12]
+ gpio_defaults_block_19/gpio_defaults[1] gpio_defaults_block_19/gpio_defaults[2]
+ gpio_defaults_block_19/gpio_defaults[3] gpio_defaults_block_19/gpio_defaults[4]
+ gpio_defaults_block_19/gpio_defaults[5] gpio_defaults_block_19/gpio_defaults[6]
+ gpio_defaults_block_19/gpio_defaults[7] gpio_defaults_block_19/gpio_defaults[8]
+ gpio_defaults_block_19/gpio_defaults[9] vccd_core gpio_defaults_block
Xgpio_control_in_1\[2\] gpio_defaults_block_10/gpio_defaults[0] gpio_defaults_block_10/gpio_defaults[10]
+ gpio_defaults_block_10/gpio_defaults[11] gpio_defaults_block_10/gpio_defaults[12]
+ gpio_defaults_block_10/gpio_defaults[1] gpio_defaults_block_10/gpio_defaults[2]
+ gpio_defaults_block_10/gpio_defaults[3] gpio_defaults_block_10/gpio_defaults[4]
+ gpio_defaults_block_10/gpio_defaults[5] gpio_defaults_block_10/gpio_defaults[6]
+ gpio_defaults_block_10/gpio_defaults[7] gpio_defaults_block_10/gpio_defaults[8]
+ gpio_defaults_block_10/gpio_defaults[9] housekeeping/mgmt_gpio_in[10] gpio_control_in_1\[2\]/one
+ housekeeping/mgmt_gpio_in[10] gpio_control_in_1\[2\]/one padframe/mprj_io_analog_en[10]
+ padframe/mprj_io_analog_pol[10] padframe/mprj_io_analog_sel[10] padframe/mprj_io_dm[30]
+ padframe/mprj_io_dm[31] padframe/mprj_io_dm[32] padframe/mprj_io_holdover[10] padframe/mprj_io_ib_mode_sel[10]
+ padframe/mprj_io_in[10] padframe/mprj_io_inp_dis[10] padframe/mprj_io_out[10] padframe/mprj_io_oeb[10]
+ padframe/mprj_io_slow_sel[10] padframe/mprj_io_vtrip_sel[10] gpio_control_in_1\[2\]/resetn
+ gpio_control_in_1\[3\]/resetn gpio_control_in_1\[2\]/serial_clock gpio_control_in_1\[3\]/serial_clock
+ gpio_control_in_1\[2\]/serial_data_in gpio_control_in_1\[3\]/serial_data_in gpio_control_in_1\[2\]/serial_load
+ gpio_control_in_1\[3\]/serial_load mprj/io_in[10] mprj/io_oeb[10] mprj/io_out[10]
+ vccd1_core VSUBS gpio_control_in_1\[2\]/zero dw_707553_615538# vccd_core vssd1_core
+ gpio_control_block
Xgpio_defaults_block_29 VSUBS gpio_defaults_block_29/gpio_defaults[0] gpio_defaults_block_29/gpio_defaults[10]
+ gpio_defaults_block_29/gpio_defaults[11] gpio_defaults_block_29/gpio_defaults[12]
+ gpio_defaults_block_29/gpio_defaults[1] gpio_defaults_block_29/gpio_defaults[2]
+ gpio_defaults_block_29/gpio_defaults[3] gpio_defaults_block_29/gpio_defaults[4]
+ gpio_defaults_block_29/gpio_defaults[5] gpio_defaults_block_29/gpio_defaults[6]
+ gpio_defaults_block_29/gpio_defaults[7] gpio_defaults_block_29/gpio_defaults[8]
+ gpio_defaults_block_29/gpio_defaults[9] vccd_core gpio_defaults_block
Xgpio_control_in_2\[10\] gpio_defaults_block_29/gpio_defaults[0] gpio_defaults_block_29/gpio_defaults[10]
+ gpio_defaults_block_29/gpio_defaults[11] gpio_defaults_block_29/gpio_defaults[12]
+ gpio_defaults_block_29/gpio_defaults[1] gpio_defaults_block_29/gpio_defaults[2]
+ gpio_defaults_block_29/gpio_defaults[3] gpio_defaults_block_29/gpio_defaults[4]
+ gpio_defaults_block_29/gpio_defaults[5] gpio_defaults_block_29/gpio_defaults[6]
+ gpio_defaults_block_29/gpio_defaults[7] gpio_defaults_block_29/gpio_defaults[8]
+ gpio_defaults_block_29/gpio_defaults[9] housekeeping/mgmt_gpio_in[29] gpio_control_in_2\[10\]/one
+ housekeeping/mgmt_gpio_in[29] gpio_control_in_2\[10\]/one padframe/mprj_io_analog_en[29]
+ padframe/mprj_io_analog_pol[29] padframe/mprj_io_analog_sel[29] padframe/mprj_io_dm[87]
+ padframe/mprj_io_dm[88] padframe/mprj_io_dm[89] padframe/mprj_io_holdover[29] padframe/mprj_io_ib_mode_sel[29]
+ padframe/mprj_io_in[29] padframe/mprj_io_inp_dis[29] padframe/mprj_io_out[29] padframe/mprj_io_oeb[29]
+ padframe/mprj_io_slow_sel[29] padframe/mprj_io_vtrip_sel[29] gpio_control_in_2\[10\]/resetn
+ gpio_control_in_2\[9\]/resetn gpio_control_in_2\[10\]/serial_clock gpio_control_in_2\[9\]/serial_clock
+ gpio_control_in_2\[10\]/serial_data_in gpio_control_in_2\[9\]/serial_data_in gpio_control_in_2\[10\]/serial_load
+ gpio_control_in_2\[9\]/serial_load mprj/io_in[29] mprj/io_oeb[29] mprj/io_out[29]
+ vccd1_core VSUBS gpio_control_in_2\[10\]/zero dw_8741_634138# vccd_core vssd1_core
+ gpio_control_block
Xgpio_control_in_1\[10\] gpio_defaults_block_18/gpio_defaults[0] gpio_defaults_block_18/gpio_defaults[10]
+ gpio_defaults_block_18/gpio_defaults[11] gpio_defaults_block_18/gpio_defaults[12]
+ gpio_defaults_block_18/gpio_defaults[1] gpio_defaults_block_18/gpio_defaults[2]
+ gpio_defaults_block_18/gpio_defaults[3] gpio_defaults_block_18/gpio_defaults[4]
+ gpio_defaults_block_18/gpio_defaults[5] gpio_defaults_block_18/gpio_defaults[6]
+ gpio_defaults_block_18/gpio_defaults[7] gpio_defaults_block_18/gpio_defaults[8]
+ gpio_defaults_block_18/gpio_defaults[9] housekeeping/mgmt_gpio_in[18] gpio_control_in_1\[10\]/one
+ housekeeping/mgmt_gpio_in[18] gpio_control_in_1\[10\]/one padframe/mprj_io_analog_en[18]
+ padframe/mprj_io_analog_pol[18] padframe/mprj_io_analog_sel[18] padframe/mprj_io_dm[54]
+ padframe/mprj_io_dm[55] padframe/mprj_io_dm[56] padframe/mprj_io_holdover[18] padframe/mprj_io_ib_mode_sel[18]
+ padframe/mprj_io_in[18] padframe/mprj_io_inp_dis[18] padframe/mprj_io_out[18] padframe/mprj_io_oeb[18]
+ padframe/mprj_io_slow_sel[18] padframe/mprj_io_vtrip_sel[18] gpio_control_in_1\[10\]/resetn
+ gpio_control_in_1\[10\]/resetn_out gpio_control_in_1\[10\]/serial_clock gpio_control_in_1\[10\]/serial_clock_out
+ gpio_control_in_1\[9\]/serial_data_out gpio_control_in_1\[10\]/serial_data_out gpio_control_in_1\[10\]/serial_load
+ gpio_control_in_1\[10\]/serial_load_out mprj/io_in[18] mprj/io_oeb[18] mprj/io_out[18]
+ vccd1_core VSUBS gpio_control_in_1\[10\]/zero dw_354938_1027427# vccd_core vssd1_core
+ gpio_control_block
Xgpio_control_in_2\[5\] gpio_defaults_block_24/gpio_defaults[0] gpio_defaults_block_24/gpio_defaults[10]
+ gpio_defaults_block_24/gpio_defaults[11] gpio_defaults_block_24/gpio_defaults[12]
+ gpio_defaults_block_24/gpio_defaults[1] gpio_defaults_block_24/gpio_defaults[2]
+ gpio_defaults_block_24/gpio_defaults[3] gpio_defaults_block_24/gpio_defaults[4]
+ gpio_defaults_block_24/gpio_defaults[5] gpio_defaults_block_24/gpio_defaults[6]
+ gpio_defaults_block_24/gpio_defaults[7] gpio_defaults_block_24/gpio_defaults[8]
+ gpio_defaults_block_24/gpio_defaults[9] housekeeping/mgmt_gpio_in[24] gpio_control_in_2\[5\]/one
+ housekeeping/mgmt_gpio_in[24] gpio_control_in_2\[5\]/one padframe/mprj_io_analog_en[24]
+ padframe/mprj_io_analog_pol[24] padframe/mprj_io_analog_sel[24] padframe/mprj_io_dm[72]
+ padframe/mprj_io_dm[73] padframe/mprj_io_dm[74] padframe/mprj_io_holdover[24] padframe/mprj_io_ib_mode_sel[24]
+ padframe/mprj_io_in[24] padframe/mprj_io_inp_dis[24] padframe/mprj_io_out[24] padframe/mprj_io_oeb[24]
+ padframe/mprj_io_slow_sel[24] padframe/mprj_io_vtrip_sel[24] gpio_control_in_2\[5\]/resetn
+ gpio_control_in_2\[4\]/resetn gpio_control_in_2\[5\]/serial_clock gpio_control_in_2\[4\]/serial_clock
+ gpio_control_in_2\[5\]/serial_data_in gpio_control_in_2\[4\]/serial_data_in gpio_control_in_2\[5\]/serial_load
+ gpio_control_in_2\[4\]/serial_load mprj/io_in[24] mprj/io_oeb[24] mprj/io_out[24]
+ vccd1_core VSUBS gpio_control_in_2\[5\]/zero dw_8741_932738# vccd_core vssd1_core
+ gpio_control_block
Xgpio_control_in_1\[0\] gpio_defaults_block_8/gpio_defaults[0] gpio_defaults_block_8/gpio_defaults[10]
+ gpio_defaults_block_8/gpio_defaults[11] gpio_defaults_block_8/gpio_defaults[12]
+ gpio_defaults_block_8/gpio_defaults[1] gpio_defaults_block_8/gpio_defaults[2] gpio_defaults_block_8/gpio_defaults[3]
+ gpio_defaults_block_8/gpio_defaults[4] gpio_defaults_block_8/gpio_defaults[5] gpio_defaults_block_8/gpio_defaults[6]
+ gpio_defaults_block_8/gpio_defaults[7] gpio_defaults_block_8/gpio_defaults[8] gpio_defaults_block_8/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[8] gpio_control_in_1\[0\]/one housekeeping/mgmt_gpio_in[8]
+ gpio_control_in_1\[0\]/one padframe/mprj_io_analog_en[8] padframe/mprj_io_analog_pol[8]
+ padframe/mprj_io_analog_sel[8] padframe/mprj_io_dm[24] padframe/mprj_io_dm[25] padframe/mprj_io_dm[26]
+ padframe/mprj_io_holdover[8] padframe/mprj_io_ib_mode_sel[8] padframe/mprj_io_in[8]
+ padframe/mprj_io_inp_dis[8] padframe/mprj_io_out[8] padframe/mprj_io_oeb[8] padframe/mprj_io_slow_sel[8]
+ padframe/mprj_io_vtrip_sel[8] gpio_control_in_1\[0\]/resetn gpio_control_in_1\[1\]/resetn
+ gpio_control_in_1\[0\]/serial_clock gpio_control_in_1\[1\]/serial_clock gpio_control_in_1\[0\]/serial_data_in
+ gpio_control_in_1\[1\]/serial_data_in gpio_control_in_1\[0\]/serial_load gpio_control_in_1\[1\]/serial_load
+ mprj/io_in[8] mprj/io_oeb[8] mprj/io_out[8] vccd1_core VSUBS gpio_control_in_1\[0\]/zero
+ dw_707553_525338# vccd_core vssd1_core gpio_control_block
Xgpio_defaults_block_0 VSUBS vccd_core gpio_defaults_block_0/gpio_defaults[0] gpio_defaults_block_0/gpio_defaults[10]
+ gpio_defaults_block_0/gpio_defaults[11] gpio_defaults_block_0/gpio_defaults[12]
+ gpio_defaults_block_0/gpio_defaults[1] gpio_defaults_block_0/gpio_defaults[2] gpio_defaults_block_0/gpio_defaults[3]
+ gpio_defaults_block_0/gpio_defaults[4] gpio_defaults_block_0/gpio_defaults[5] gpio_defaults_block_0/gpio_defaults[6]
+ gpio_defaults_block_0/gpio_defaults[7] gpio_defaults_block_0/gpio_defaults[8] gpio_defaults_block_0/gpio_defaults[9]
+ gpio_defaults_block_1803
Xgpio_defaults_block_1 VSUBS vccd_core gpio_defaults_block_1/gpio_defaults[0] gpio_defaults_block_1/gpio_defaults[10]
+ gpio_defaults_block_1/gpio_defaults[11] gpio_defaults_block_1/gpio_defaults[12]
+ gpio_defaults_block_1/gpio_defaults[1] gpio_defaults_block_1/gpio_defaults[2] gpio_defaults_block_1/gpio_defaults[3]
+ gpio_defaults_block_1/gpio_defaults[4] gpio_defaults_block_1/gpio_defaults[5] gpio_defaults_block_1/gpio_defaults[6]
+ gpio_defaults_block_1/gpio_defaults[7] gpio_defaults_block_1/gpio_defaults[8] gpio_defaults_block_1/gpio_defaults[9]
+ gpio_defaults_block_1803
Xuser_id_value user_id_value/mask_rev[0] user_id_value/mask_rev[10] user_id_value/mask_rev[11]
+ user_id_value/mask_rev[12] user_id_value/mask_rev[13] user_id_value/mask_rev[14]
+ user_id_value/mask_rev[15] user_id_value/mask_rev[16] user_id_value/mask_rev[17]
+ user_id_value/mask_rev[18] user_id_value/mask_rev[19] user_id_value/mask_rev[1]
+ user_id_value/mask_rev[20] user_id_value/mask_rev[21] user_id_value/mask_rev[22]
+ user_id_value/mask_rev[23] user_id_value/mask_rev[24] user_id_value/mask_rev[25]
+ user_id_value/mask_rev[26] user_id_value/mask_rev[27] user_id_value/mask_rev[28]
+ user_id_value/mask_rev[29] user_id_value/mask_rev[2] user_id_value/mask_rev[30]
+ user_id_value/mask_rev[31] user_id_value/mask_rev[3] user_id_value/mask_rev[4] user_id_value/mask_rev[5]
+ user_id_value/mask_rev[6] user_id_value/mask_rev[7] user_id_value/mask_rev[8] user_id_value/mask_rev[9]
+ VSUBS vccd_core user_id_programming
Xgpio_control_in_2\[3\] gpio_defaults_block_22/gpio_defaults[0] gpio_defaults_block_22/gpio_defaults[10]
+ gpio_defaults_block_22/gpio_defaults[11] gpio_defaults_block_22/gpio_defaults[12]
+ gpio_defaults_block_22/gpio_defaults[1] gpio_defaults_block_22/gpio_defaults[2]
+ gpio_defaults_block_22/gpio_defaults[3] gpio_defaults_block_22/gpio_defaults[4]
+ gpio_defaults_block_22/gpio_defaults[5] gpio_defaults_block_22/gpio_defaults[6]
+ gpio_defaults_block_22/gpio_defaults[7] gpio_defaults_block_22/gpio_defaults[8]
+ gpio_defaults_block_22/gpio_defaults[9] housekeeping/mgmt_gpio_in[22] gpio_control_in_2\[3\]/one
+ housekeeping/mgmt_gpio_in[22] gpio_control_in_2\[3\]/one padframe/mprj_io_analog_en[22]
+ padframe/mprj_io_analog_pol[22] padframe/mprj_io_analog_sel[22] padframe/mprj_io_dm[66]
+ padframe/mprj_io_dm[67] padframe/mprj_io_dm[68] padframe/mprj_io_holdover[22] padframe/mprj_io_ib_mode_sel[22]
+ padframe/mprj_io_in[22] padframe/mprj_io_inp_dis[22] padframe/mprj_io_out[22] padframe/mprj_io_oeb[22]
+ padframe/mprj_io_slow_sel[22] padframe/mprj_io_vtrip_sel[22] gpio_control_in_2\[3\]/resetn
+ gpio_control_in_2\[2\]/resetn gpio_control_in_2\[3\]/serial_clock gpio_control_in_2\[2\]/serial_clock
+ gpio_control_in_2\[3\]/serial_data_in gpio_control_in_2\[2\]/serial_data_in gpio_control_in_2\[3\]/serial_load
+ gpio_control_in_2\[2\]/serial_load mprj/io_in[22] mprj/io_oeb[22] mprj/io_out[22]
+ vccd1_core VSUBS gpio_control_in_2\[3\]/zero dw_150138_1027427# vccd_core vssd1_core
+ gpio_control_block
Xgpio_defaults_block_2 VSUBS vccd_core gpio_defaults_block_2/gpio_defaults[0] gpio_defaults_block_2/gpio_defaults[10]
+ gpio_defaults_block_2/gpio_defaults[11] gpio_defaults_block_2/gpio_defaults[12]
+ gpio_defaults_block_2/gpio_defaults[1] gpio_defaults_block_2/gpio_defaults[2] gpio_defaults_block_2/gpio_defaults[3]
+ gpio_defaults_block_2/gpio_defaults[4] gpio_defaults_block_2/gpio_defaults[5] gpio_defaults_block_2/gpio_defaults[6]
+ gpio_defaults_block_2/gpio_defaults[7] gpio_defaults_block_2/gpio_defaults[8] gpio_defaults_block_2/gpio_defaults[9]
+ gpio_defaults_block_0403
Xgpio_defaults_block_3 VSUBS vccd_core gpio_defaults_block_3/gpio_defaults[0] gpio_defaults_block_3/gpio_defaults[10]
+ gpio_defaults_block_3/gpio_defaults[11] gpio_defaults_block_3/gpio_defaults[12]
+ gpio_defaults_block_3/gpio_defaults[1] gpio_defaults_block_3/gpio_defaults[2] gpio_defaults_block_3/gpio_defaults[3]
+ gpio_defaults_block_3/gpio_defaults[4] gpio_defaults_block_3/gpio_defaults[5] gpio_defaults_block_3/gpio_defaults[6]
+ gpio_defaults_block_3/gpio_defaults[7] gpio_defaults_block_3/gpio_defaults[8] gpio_defaults_block_3/gpio_defaults[9]
+ gpio_defaults_block_0403
Xgpio_control_bidir_1\[0\] gpio_defaults_block_0/gpio_defaults[0] gpio_defaults_block_0/gpio_defaults[10]
+ gpio_defaults_block_0/gpio_defaults[11] gpio_defaults_block_0/gpio_defaults[12]
+ gpio_defaults_block_0/gpio_defaults[1] gpio_defaults_block_0/gpio_defaults[2] gpio_defaults_block_0/gpio_defaults[3]
+ gpio_defaults_block_0/gpio_defaults[4] gpio_defaults_block_0/gpio_defaults[5] gpio_defaults_block_0/gpio_defaults[6]
+ gpio_defaults_block_0/gpio_defaults[7] gpio_defaults_block_0/gpio_defaults[8] gpio_defaults_block_0/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[0] housekeeping/mgmt_gpio_oeb[0] housekeeping/mgmt_gpio_out[0]
+ gpio_control_bidir_1\[0\]/one padframe/mprj_io_analog_en[0] padframe/mprj_io_analog_pol[0]
+ padframe/mprj_io_analog_sel[0] padframe/mprj_io_dm[0] padframe/mprj_io_dm[1] padframe/mprj_io_dm[2]
+ padframe/mprj_io_holdover[0] padframe/mprj_io_ib_mode_sel[0] padframe/mprj_io_in[0]
+ padframe/mprj_io_inp_dis[0] padframe/mprj_io_out[0] padframe/mprj_io_oeb[0] padframe/mprj_io_slow_sel[0]
+ padframe/mprj_io_vtrip_sel[0] housekeeping/serial_resetn gpio_control_bidir_1\[1\]/resetn
+ housekeeping/serial_clock gpio_control_bidir_1\[1\]/serial_clock housekeeping/serial_data_1
+ gpio_control_bidir_1\[1\]/serial_data_in housekeeping/serial_load gpio_control_bidir_1\[1\]/serial_load
+ mprj/io_in[0] mprj/io_oeb[0] mprj/io_out[0] vccd1_core VSUBS gpio_control_bidir_1\[0\]/zero
+ dw_707553_122538# vccd_core vssd1_core gpio_control_block
Xgpio_control_in_1\[9\] gpio_defaults_block_17/gpio_defaults[0] gpio_defaults_block_17/gpio_defaults[10]
+ gpio_defaults_block_17/gpio_defaults[11] gpio_defaults_block_17/gpio_defaults[12]
+ gpio_defaults_block_17/gpio_defaults[1] gpio_defaults_block_17/gpio_defaults[2]
+ gpio_defaults_block_17/gpio_defaults[3] gpio_defaults_block_17/gpio_defaults[4]
+ gpio_defaults_block_17/gpio_defaults[5] gpio_defaults_block_17/gpio_defaults[6]
+ gpio_defaults_block_17/gpio_defaults[7] gpio_defaults_block_17/gpio_defaults[8]
+ gpio_defaults_block_17/gpio_defaults[9] housekeeping/mgmt_gpio_in[17] gpio_control_in_1\[9\]/one
+ housekeeping/mgmt_gpio_in[17] gpio_control_in_1\[9\]/one padframe/mprj_io_analog_en[17]
+ padframe/mprj_io_analog_pol[17] padframe/mprj_io_analog_sel[17] padframe/mprj_io_dm[51]
+ padframe/mprj_io_dm[52] padframe/mprj_io_dm[53] padframe/mprj_io_holdover[17] padframe/mprj_io_ib_mode_sel[17]
+ padframe/mprj_io_in[17] padframe/mprj_io_inp_dis[17] padframe/mprj_io_out[17] padframe/mprj_io_oeb[17]
+ padframe/mprj_io_slow_sel[17] padframe/mprj_io_vtrip_sel[17] gpio_control_in_1\[9\]/resetn
+ gpio_control_in_1\[10\]/resetn gpio_control_in_1\[9\]/serial_clock gpio_control_in_1\[10\]/serial_clock
+ gpio_control_in_1\[9\]/serial_data_in gpio_control_in_1\[9\]/serial_data_out gpio_control_in_1\[9\]/serial_load
+ gpio_control_in_1\[10\]/serial_load mprj/io_in[17] mprj/io_oeb[17] mprj/io_out[17]
+ vccd1_core VSUBS gpio_control_in_1\[9\]/zero dw_422338_1027427# vccd_core vssd1_core
+ gpio_control_block
Xgpio_defaults_block_5 VSUBS gpio_defaults_block_5/gpio_defaults[0] gpio_defaults_block_5/gpio_defaults[10]
+ gpio_defaults_block_5/gpio_defaults[11] gpio_defaults_block_5/gpio_defaults[12]
+ gpio_defaults_block_5/gpio_defaults[1] gpio_defaults_block_5/gpio_defaults[2] gpio_defaults_block_5/gpio_defaults[3]
+ gpio_defaults_block_5/gpio_defaults[4] gpio_defaults_block_5/gpio_defaults[5] gpio_defaults_block_5/gpio_defaults[6]
+ gpio_defaults_block_5/gpio_defaults[7] gpio_defaults_block_5/gpio_defaults[8] gpio_defaults_block_5/gpio_defaults[9]
+ vccd_core gpio_defaults_block
Xgpio_defaults_block_4 VSUBS vccd_core gpio_defaults_block_4/gpio_defaults[0] gpio_defaults_block_4/gpio_defaults[10]
+ gpio_defaults_block_4/gpio_defaults[11] gpio_defaults_block_4/gpio_defaults[12]
+ gpio_defaults_block_4/gpio_defaults[1] gpio_defaults_block_4/gpio_defaults[2] gpio_defaults_block_4/gpio_defaults[3]
+ gpio_defaults_block_4/gpio_defaults[4] gpio_defaults_block_4/gpio_defaults[5] gpio_defaults_block_4/gpio_defaults[6]
+ gpio_defaults_block_4/gpio_defaults[7] gpio_defaults_block_4/gpio_defaults[8] gpio_defaults_block_4/gpio_defaults[9]
+ gpio_defaults_block_0403
Xgpio_control_in_2\[1\] gpio_defaults_block_20/gpio_defaults[0] gpio_defaults_block_20/gpio_defaults[10]
+ gpio_defaults_block_20/gpio_defaults[11] gpio_defaults_block_20/gpio_defaults[12]
+ gpio_defaults_block_20/gpio_defaults[1] gpio_defaults_block_20/gpio_defaults[2]
+ gpio_defaults_block_20/gpio_defaults[3] gpio_defaults_block_20/gpio_defaults[4]
+ gpio_defaults_block_20/gpio_defaults[5] gpio_defaults_block_20/gpio_defaults[6]
+ gpio_defaults_block_20/gpio_defaults[7] gpio_defaults_block_20/gpio_defaults[8]
+ gpio_defaults_block_20/gpio_defaults[9] housekeeping/mgmt_gpio_in[20] gpio_control_in_2\[1\]/one
+ housekeeping/mgmt_gpio_in[20] gpio_control_in_2\[1\]/one padframe/mprj_io_analog_en[20]
+ padframe/mprj_io_analog_pol[20] padframe/mprj_io_analog_sel[20] padframe/mprj_io_dm[60]
+ padframe/mprj_io_dm[61] padframe/mprj_io_dm[62] padframe/mprj_io_holdover[20] padframe/mprj_io_ib_mode_sel[20]
+ padframe/mprj_io_in[20] padframe/mprj_io_inp_dis[20] padframe/mprj_io_out[20] padframe/mprj_io_oeb[20]
+ padframe/mprj_io_slow_sel[20] padframe/mprj_io_vtrip_sel[20] gpio_control_in_2\[1\]/resetn
+ gpio_control_in_2\[0\]/resetn gpio_control_in_2\[1\]/serial_clock gpio_control_in_2\[0\]/serial_clock
+ gpio_control_in_2\[1\]/serial_data_in gpio_control_in_2\[0\]/serial_data_in gpio_control_in_2\[1\]/serial_load
+ gpio_control_in_2\[0\]/serial_load mprj/io_in[20] mprj/io_oeb[20] mprj/io_out[20]
+ vccd1_core VSUBS gpio_control_in_2\[1\]/zero dw_252938_1027427# vccd_core vssd1_core
+ gpio_control_block
Xgpio_defaults_block_6 VSUBS gpio_defaults_block_6/gpio_defaults[0] gpio_defaults_block_6/gpio_defaults[10]
+ gpio_defaults_block_6/gpio_defaults[11] gpio_defaults_block_6/gpio_defaults[12]
+ gpio_defaults_block_6/gpio_defaults[1] gpio_defaults_block_6/gpio_defaults[2] gpio_defaults_block_6/gpio_defaults[3]
+ gpio_defaults_block_6/gpio_defaults[4] gpio_defaults_block_6/gpio_defaults[5] gpio_defaults_block_6/gpio_defaults[6]
+ gpio_defaults_block_6/gpio_defaults[7] gpio_defaults_block_6/gpio_defaults[8] gpio_defaults_block_6/gpio_defaults[9]
+ vccd_core gpio_defaults_block
Xgpio_defaults_block_7 VSUBS gpio_defaults_block_7/gpio_defaults[0] gpio_defaults_block_7/gpio_defaults[10]
+ gpio_defaults_block_7/gpio_defaults[11] gpio_defaults_block_7/gpio_defaults[12]
+ gpio_defaults_block_7/gpio_defaults[1] gpio_defaults_block_7/gpio_defaults[2] gpio_defaults_block_7/gpio_defaults[3]
+ gpio_defaults_block_7/gpio_defaults[4] gpio_defaults_block_7/gpio_defaults[5] gpio_defaults_block_7/gpio_defaults[6]
+ gpio_defaults_block_7/gpio_defaults[7] gpio_defaults_block_7/gpio_defaults[8] gpio_defaults_block_7/gpio_defaults[9]
+ vccd_core gpio_defaults_block
Xgpio_control_in_1\[7\] gpio_defaults_block_15/gpio_defaults[0] gpio_defaults_block_15/gpio_defaults[10]
+ gpio_defaults_block_15/gpio_defaults[11] gpio_defaults_block_15/gpio_defaults[12]
+ gpio_defaults_block_15/gpio_defaults[1] gpio_defaults_block_15/gpio_defaults[2]
+ gpio_defaults_block_15/gpio_defaults[3] gpio_defaults_block_15/gpio_defaults[4]
+ gpio_defaults_block_15/gpio_defaults[5] gpio_defaults_block_15/gpio_defaults[6]
+ gpio_defaults_block_15/gpio_defaults[7] gpio_defaults_block_15/gpio_defaults[8]
+ gpio_defaults_block_15/gpio_defaults[9] housekeeping/mgmt_gpio_in[15] gpio_control_in_1\[7\]/one
+ housekeeping/mgmt_gpio_in[15] gpio_control_in_1\[7\]/one padframe/mprj_io_analog_en[15]
+ padframe/mprj_io_analog_pol[15] padframe/mprj_io_analog_sel[15] padframe/mprj_io_dm[45]
+ padframe/mprj_io_dm[46] padframe/mprj_io_dm[47] padframe/mprj_io_holdover[15] padframe/mprj_io_ib_mode_sel[15]
+ padframe/mprj_io_in[15] padframe/mprj_io_inp_dis[15] padframe/mprj_io_out[15] padframe/mprj_io_oeb[15]
+ padframe/mprj_io_slow_sel[15] padframe/mprj_io_vtrip_sel[15] gpio_control_in_1\[7\]/resetn
+ gpio_control_in_1\[8\]/resetn gpio_control_in_1\[7\]/serial_clock gpio_control_in_1\[8\]/serial_clock
+ gpio_control_in_1\[7\]/serial_data_in gpio_control_in_1\[8\]/serial_data_in gpio_control_in_1\[7\]/serial_load
+ gpio_control_in_1\[8\]/serial_load mprj/io_in[15] mprj/io_oeb[15] mprj/io_out[15]
+ vccd1_core VSUBS gpio_control_in_1\[7\]/zero dw_550738_1027427# vccd_core vssd1_core
+ gpio_control_block
Xgpio_defaults_block_8 VSUBS gpio_defaults_block_8/gpio_defaults[0] gpio_defaults_block_8/gpio_defaults[10]
+ gpio_defaults_block_8/gpio_defaults[11] gpio_defaults_block_8/gpio_defaults[12]
+ gpio_defaults_block_8/gpio_defaults[1] gpio_defaults_block_8/gpio_defaults[2] gpio_defaults_block_8/gpio_defaults[3]
+ gpio_defaults_block_8/gpio_defaults[4] gpio_defaults_block_8/gpio_defaults[5] gpio_defaults_block_8/gpio_defaults[6]
+ gpio_defaults_block_8/gpio_defaults[7] gpio_defaults_block_8/gpio_defaults[8] gpio_defaults_block_8/gpio_defaults[9]
+ vccd_core gpio_defaults_block
Xgpio_control_in_1a\[4\] gpio_defaults_block_6/gpio_defaults[0] gpio_defaults_block_6/gpio_defaults[10]
+ gpio_defaults_block_6/gpio_defaults[11] gpio_defaults_block_6/gpio_defaults[12]
+ gpio_defaults_block_6/gpio_defaults[1] gpio_defaults_block_6/gpio_defaults[2] gpio_defaults_block_6/gpio_defaults[3]
+ gpio_defaults_block_6/gpio_defaults[4] gpio_defaults_block_6/gpio_defaults[5] gpio_defaults_block_6/gpio_defaults[6]
+ gpio_defaults_block_6/gpio_defaults[7] gpio_defaults_block_6/gpio_defaults[8] gpio_defaults_block_6/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[6] gpio_control_in_1a\[4\]/one housekeeping/mgmt_gpio_in[6]
+ gpio_control_in_1a\[4\]/one padframe/mprj_io_analog_en[6] padframe/mprj_io_analog_pol[6]
+ padframe/mprj_io_analog_sel[6] padframe/mprj_io_dm[18] padframe/mprj_io_dm[19] padframe/mprj_io_dm[20]
+ padframe/mprj_io_holdover[6] padframe/mprj_io_ib_mode_sel[6] padframe/mprj_io_in[6]
+ padframe/mprj_io_inp_dis[6] padframe/mprj_io_out[6] padframe/mprj_io_oeb[6] padframe/mprj_io_slow_sel[6]
+ padframe/mprj_io_vtrip_sel[6] gpio_control_in_1a\[4\]/resetn gpio_control_in_1a\[5\]/resetn
+ gpio_control_in_1a\[4\]/serial_clock gpio_control_in_1a\[5\]/serial_clock gpio_control_in_1a\[4\]/serial_data_in
+ gpio_control_in_1a\[5\]/serial_data_in gpio_control_in_1a\[4\]/serial_load gpio_control_in_1a\[5\]/serial_load
+ mprj/io_in[6] mprj/io_oeb[6] mprj/io_out[6] vccd1_core VSUBS gpio_control_in_1a\[4\]/zero
+ dw_707553_393138# vccd_core vssd1_core gpio_control_block
Xmgmt_buffers soc/core_clk clocking/user_clk soc/core_rstn mprj/la_data_in[0] mprj/la_data_in[100]
+ mprj/la_data_in[101] mprj/la_data_in[102] mprj/la_data_in[103] mprj/la_data_in[104]
+ mprj/la_data_in[105] mprj/la_data_in[106] mprj/la_data_in[107] mprj/la_data_in[108]
+ mprj/la_data_in[109] mprj/la_data_in[10] mprj/la_data_in[110] mprj/la_data_in[111]
+ mprj/la_data_in[112] mprj/la_data_in[113] mprj/la_data_in[114] mprj/la_data_in[115]
+ mprj/la_data_in[116] mprj/la_data_in[117] mprj/la_data_in[118] mprj/la_data_in[119]
+ mprj/la_data_in[11] mprj/la_data_in[120] mprj/la_data_in[121] mprj/la_data_in[122]
+ mprj/la_data_in[123] mprj/la_data_in[124] mprj/la_data_in[125] mprj/la_data_in[126]
+ mprj/la_data_in[127] mprj/la_data_in[12] mprj/la_data_in[13] mprj/la_data_in[14]
+ mprj/la_data_in[15] mprj/la_data_in[16] mprj/la_data_in[17] mprj/la_data_in[18]
+ mprj/la_data_in[19] mprj/la_data_in[1] mprj/la_data_in[20] mprj/la_data_in[21] mprj/la_data_in[22]
+ mprj/la_data_in[23] mprj/la_data_in[24] mprj/la_data_in[25] mprj/la_data_in[26]
+ mprj/la_data_in[27] mprj/la_data_in[28] mprj/la_data_in[29] mprj/la_data_in[2] mprj/la_data_in[30]
+ mprj/la_data_in[31] mprj/la_data_in[32] mprj/la_data_in[33] mprj/la_data_in[34]
+ mprj/la_data_in[35] mprj/la_data_in[36] mprj/la_data_in[37] mprj/la_data_in[38]
+ mprj/la_data_in[39] mprj/la_data_in[3] mprj/la_data_in[40] mprj/la_data_in[41] mprj/la_data_in[42]
+ mprj/la_data_in[43] mprj/la_data_in[44] mprj/la_data_in[45] mprj/la_data_in[46]
+ mprj/la_data_in[47] mprj/la_data_in[48] mprj/la_data_in[49] mprj/la_data_in[4] mprj/la_data_in[50]
+ mprj/la_data_in[51] mprj/la_data_in[52] mprj/la_data_in[53] mprj/la_data_in[54]
+ mprj/la_data_in[55] mprj/la_data_in[56] mprj/la_data_in[57] mprj/la_data_in[58]
+ mprj/la_data_in[59] mprj/la_data_in[5] mprj/la_data_in[60] mprj/la_data_in[61] mprj/la_data_in[62]
+ mprj/la_data_in[63] mprj/la_data_in[64] mprj/la_data_in[65] mprj/la_data_in[66]
+ mprj/la_data_in[67] mprj/la_data_in[68] mprj/la_data_in[69] mprj/la_data_in[6] mprj/la_data_in[70]
+ mprj/la_data_in[71] mprj/la_data_in[72] mprj/la_data_in[73] mprj/la_data_in[74]
+ mprj/la_data_in[75] mprj/la_data_in[76] mprj/la_data_in[77] mprj/la_data_in[78]
+ mprj/la_data_in[79] mprj/la_data_in[7] mprj/la_data_in[80] mprj/la_data_in[81] mprj/la_data_in[82]
+ mprj/la_data_in[83] mprj/la_data_in[84] mprj/la_data_in[85] mprj/la_data_in[86]
+ mprj/la_data_in[87] mprj/la_data_in[88] mprj/la_data_in[89] mprj/la_data_in[8] mprj/la_data_in[90]
+ mprj/la_data_in[91] mprj/la_data_in[92] mprj/la_data_in[93] mprj/la_data_in[94]
+ mprj/la_data_in[95] mprj/la_data_in[96] mprj/la_data_in[97] mprj/la_data_in[98]
+ mprj/la_data_in[99] mprj/la_data_in[9] soc/la_input[0] soc/la_input[100] soc/la_input[101]
+ soc/la_input[102] soc/la_input[103] soc/la_input[104] soc/la_input[105] soc/la_input[106]
+ soc/la_input[107] soc/la_input[108] soc/la_input[109] soc/la_input[10] soc/la_input[110]
+ soc/la_input[111] soc/la_input[112] soc/la_input[113] soc/la_input[114] soc/la_input[115]
+ soc/la_input[116] soc/la_input[117] soc/la_input[118] soc/la_input[119] soc/la_input[11]
+ soc/la_input[120] soc/la_input[121] soc/la_input[122] soc/la_input[123] soc/la_input[124]
+ soc/la_input[125] soc/la_input[126] soc/la_input[127] soc/la_input[12] soc/la_input[13]
+ soc/la_input[14] soc/la_input[15] soc/la_input[16] soc/la_input[17] soc/la_input[18]
+ soc/la_input[19] soc/la_input[1] soc/la_input[20] soc/la_input[21] soc/la_input[22]
+ soc/la_input[23] soc/la_input[24] soc/la_input[25] soc/la_input[26] soc/la_input[27]
+ soc/la_input[28] soc/la_input[29] soc/la_input[2] soc/la_input[30] soc/la_input[31]
+ soc/la_input[32] soc/la_input[33] soc/la_input[34] soc/la_input[35] soc/la_input[36]
+ soc/la_input[37] soc/la_input[38] soc/la_input[39] soc/la_input[3] soc/la_input[40]
+ soc/la_input[41] soc/la_input[42] soc/la_input[43] soc/la_input[44] soc/la_input[45]
+ soc/la_input[46] soc/la_input[47] soc/la_input[48] soc/la_input[49] soc/la_input[4]
+ soc/la_input[50] soc/la_input[51] soc/la_input[52] soc/la_input[53] soc/la_input[54]
+ soc/la_input[55] soc/la_input[56] soc/la_input[57] soc/la_input[58] soc/la_input[59]
+ soc/la_input[5] soc/la_input[60] soc/la_input[61] soc/la_input[62] soc/la_input[63]
+ soc/la_input[64] soc/la_input[65] soc/la_input[66] soc/la_input[67] soc/la_input[68]
+ soc/la_input[69] soc/la_input[6] soc/la_input[70] soc/la_input[71] soc/la_input[72]
+ soc/la_input[73] soc/la_input[74] soc/la_input[75] soc/la_input[76] soc/la_input[77]
+ soc/la_input[78] soc/la_input[79] soc/la_input[7] soc/la_input[80] soc/la_input[81]
+ soc/la_input[82] soc/la_input[83] soc/la_input[84] soc/la_input[85] soc/la_input[86]
+ soc/la_input[87] soc/la_input[88] soc/la_input[89] soc/la_input[8] soc/la_input[90]
+ soc/la_input[91] soc/la_input[92] soc/la_input[93] soc/la_input[94] soc/la_input[95]
+ soc/la_input[96] soc/la_input[97] soc/la_input[98] soc/la_input[99] soc/la_input[9]
+ mprj/la_data_out[0] mprj/la_data_out[100] mprj/la_data_out[101] mprj/la_data_out[102]
+ mprj/la_data_out[103] mprj/la_data_out[104] mprj/la_data_out[105] mprj/la_data_out[106]
+ mprj/la_data_out[107] mprj/la_data_out[108] mprj/la_data_out[109] mprj/la_data_out[10]
+ mprj/la_data_out[110] mprj/la_data_out[111] mprj/la_data_out[112] mprj/la_data_out[113]
+ mprj/la_data_out[114] mprj/la_data_out[115] mprj/la_data_out[116] mprj/la_data_out[117]
+ mprj/la_data_out[118] mprj/la_data_out[119] mprj/la_data_out[11] mprj/la_data_out[120]
+ mprj/la_data_out[121] mprj/la_data_out[122] mprj/la_data_out[123] mprj/la_data_out[124]
+ mprj/la_data_out[125] mprj/la_data_out[126] mprj/la_data_out[127] mprj/la_data_out[12]
+ mprj/la_data_out[13] mprj/la_data_out[14] mprj/la_data_out[15] mprj/la_data_out[16]
+ mprj/la_data_out[17] mprj/la_data_out[18] mprj/la_data_out[19] mprj/la_data_out[1]
+ mprj/la_data_out[20] mprj/la_data_out[21] mprj/la_data_out[22] mprj/la_data_out[23]
+ mprj/la_data_out[24] mprj/la_data_out[25] mprj/la_data_out[26] mprj/la_data_out[27]
+ mprj/la_data_out[28] mprj/la_data_out[29] mprj/la_data_out[2] mprj/la_data_out[30]
+ mprj/la_data_out[31] mprj/la_data_out[32] mprj/la_data_out[33] mprj/la_data_out[34]
+ mprj/la_data_out[35] mprj/la_data_out[36] mprj/la_data_out[37] mprj/la_data_out[38]
+ mprj/la_data_out[39] mprj/la_data_out[3] mprj/la_data_out[40] mprj/la_data_out[41]
+ mprj/la_data_out[42] mprj/la_data_out[43] mprj/la_data_out[44] mprj/la_data_out[45]
+ mprj/la_data_out[46] mprj/la_data_out[47] mprj/la_data_out[48] mprj/la_data_out[49]
+ mprj/la_data_out[4] mprj/la_data_out[50] mprj/la_data_out[51] mprj/la_data_out[52]
+ mprj/la_data_out[53] mprj/la_data_out[54] mprj/la_data_out[55] mprj/la_data_out[56]
+ mprj/la_data_out[57] mprj/la_data_out[58] mprj/la_data_out[59] mprj/la_data_out[5]
+ mprj/la_data_out[60] mprj/la_data_out[61] mprj/la_data_out[62] mprj/la_data_out[63]
+ mprj/la_data_out[64] mprj/la_data_out[65] mprj/la_data_out[66] mprj/la_data_out[67]
+ mprj/la_data_out[68] mprj/la_data_out[69] mprj/la_data_out[6] mprj/la_data_out[70]
+ mprj/la_data_out[71] mprj/la_data_out[72] mprj/la_data_out[73] mprj/la_data_out[74]
+ mprj/la_data_out[75] mprj/la_data_out[76] mprj/la_data_out[77] mprj/la_data_out[78]
+ mprj/la_data_out[79] mprj/la_data_out[7] mprj/la_data_out[80] mprj/la_data_out[81]
+ mprj/la_data_out[82] mprj/la_data_out[83] mprj/la_data_out[84] mprj/la_data_out[85]
+ mprj/la_data_out[86] mprj/la_data_out[87] mprj/la_data_out[88] mprj/la_data_out[89]
+ mprj/la_data_out[8] mprj/la_data_out[90] mprj/la_data_out[91] mprj/la_data_out[92]
+ mprj/la_data_out[93] mprj/la_data_out[94] mprj/la_data_out[95] mprj/la_data_out[96]
+ mprj/la_data_out[97] mprj/la_data_out[98] mprj/la_data_out[99] mprj/la_data_out[9]
+ soc/la_output[0] soc/la_output[100] soc/la_output[101] soc/la_output[102] soc/la_output[103]
+ soc/la_output[104] soc/la_output[105] soc/la_output[106] soc/la_output[107] soc/la_output[108]
+ soc/la_output[109] soc/la_output[10] soc/la_output[110] soc/la_output[111] soc/la_output[112]
+ soc/la_output[113] soc/la_output[114] soc/la_output[115] soc/la_output[116] soc/la_output[117]
+ soc/la_output[118] soc/la_output[119] soc/la_output[11] soc/la_output[120] soc/la_output[121]
+ soc/la_output[122] soc/la_output[123] soc/la_output[124] soc/la_output[125] soc/la_output[126]
+ soc/la_output[127] soc/la_output[12] soc/la_output[13] soc/la_output[14] soc/la_output[15]
+ soc/la_output[16] soc/la_output[17] soc/la_output[18] soc/la_output[19] soc/la_output[1]
+ soc/la_output[20] soc/la_output[21] soc/la_output[22] soc/la_output[23] soc/la_output[24]
+ soc/la_output[25] soc/la_output[26] soc/la_output[27] soc/la_output[28] soc/la_output[29]
+ soc/la_output[2] soc/la_output[30] soc/la_output[31] soc/la_output[32] soc/la_output[33]
+ soc/la_output[34] soc/la_output[35] soc/la_output[36] soc/la_output[37] soc/la_output[38]
+ soc/la_output[39] soc/la_output[3] soc/la_output[40] soc/la_output[41] soc/la_output[42]
+ soc/la_output[43] soc/la_output[44] soc/la_output[45] soc/la_output[46] soc/la_output[47]
+ soc/la_output[48] soc/la_output[49] soc/la_output[4] soc/la_output[50] soc/la_output[51]
+ soc/la_output[52] soc/la_output[53] soc/la_output[54] soc/la_output[55] soc/la_output[56]
+ soc/la_output[57] soc/la_output[58] soc/la_output[59] soc/la_output[5] soc/la_output[60]
+ soc/la_output[61] soc/la_output[62] soc/la_output[63] soc/la_output[64] soc/la_output[65]
+ soc/la_output[66] soc/la_output[67] soc/la_output[68] soc/la_output[69] soc/la_output[6]
+ soc/la_output[70] soc/la_output[71] soc/la_output[72] soc/la_output[73] soc/la_output[74]
+ soc/la_output[75] soc/la_output[76] soc/la_output[77] soc/la_output[78] soc/la_output[79]
+ soc/la_output[7] soc/la_output[80] soc/la_output[81] soc/la_output[82] soc/la_output[83]
+ soc/la_output[84] soc/la_output[85] soc/la_output[86] soc/la_output[87] soc/la_output[88]
+ soc/la_output[89] soc/la_output[8] soc/la_output[90] soc/la_output[91] soc/la_output[92]
+ soc/la_output[93] soc/la_output[94] soc/la_output[95] soc/la_output[96] soc/la_output[97]
+ soc/la_output[98] soc/la_output[99] soc/la_output[9] soc/la_iena[0] soc/la_iena[100]
+ soc/la_iena[101] soc/la_iena[102] soc/la_iena[103] soc/la_iena[104] soc/la_iena[105]
+ soc/la_iena[106] soc/la_iena[107] soc/la_iena[108] soc/la_iena[109] soc/la_iena[10]
+ soc/la_iena[110] soc/la_iena[111] soc/la_iena[112] soc/la_iena[113] soc/la_iena[114]
+ soc/la_iena[115] soc/la_iena[116] soc/la_iena[117] soc/la_iena[118] soc/la_iena[119]
+ soc/la_iena[11] soc/la_iena[120] soc/la_iena[121] soc/la_iena[122] soc/la_iena[123]
+ soc/la_iena[124] soc/la_iena[125] soc/la_iena[126] soc/la_iena[127] soc/la_iena[12]
+ soc/la_iena[13] soc/la_iena[14] soc/la_iena[15] soc/la_iena[16] soc/la_iena[17]
+ soc/la_iena[18] soc/la_iena[19] soc/la_iena[1] soc/la_iena[20] soc/la_iena[21] soc/la_iena[22]
+ soc/la_iena[23] soc/la_iena[24] soc/la_iena[25] soc/la_iena[26] soc/la_iena[27]
+ soc/la_iena[28] soc/la_iena[29] soc/la_iena[2] soc/la_iena[30] soc/la_iena[31] soc/la_iena[32]
+ soc/la_iena[33] soc/la_iena[34] soc/la_iena[35] soc/la_iena[36] soc/la_iena[37]
+ soc/la_iena[38] soc/la_iena[39] soc/la_iena[3] soc/la_iena[40] soc/la_iena[41] soc/la_iena[42]
+ soc/la_iena[43] soc/la_iena[44] soc/la_iena[45] soc/la_iena[46] soc/la_iena[47]
+ soc/la_iena[48] soc/la_iena[49] soc/la_iena[4] soc/la_iena[50] soc/la_iena[51] soc/la_iena[52]
+ soc/la_iena[53] soc/la_iena[54] soc/la_iena[55] soc/la_iena[56] soc/la_iena[57]
+ soc/la_iena[58] soc/la_iena[59] soc/la_iena[5] soc/la_iena[60] soc/la_iena[61] soc/la_iena[62]
+ soc/la_iena[63] soc/la_iena[64] soc/la_iena[65] soc/la_iena[66] soc/la_iena[67]
+ soc/la_iena[68] soc/la_iena[69] soc/la_iena[6] soc/la_iena[70] soc/la_iena[71] soc/la_iena[72]
+ soc/la_iena[73] soc/la_iena[74] soc/la_iena[75] soc/la_iena[76] soc/la_iena[77]
+ soc/la_iena[78] soc/la_iena[79] soc/la_iena[7] soc/la_iena[80] soc/la_iena[81] soc/la_iena[82]
+ soc/la_iena[83] soc/la_iena[84] soc/la_iena[85] soc/la_iena[86] soc/la_iena[87]
+ soc/la_iena[88] soc/la_iena[89] soc/la_iena[8] soc/la_iena[90] soc/la_iena[91] soc/la_iena[92]
+ soc/la_iena[93] soc/la_iena[94] soc/la_iena[95] soc/la_iena[96] soc/la_iena[97]
+ soc/la_iena[98] soc/la_iena[99] soc/la_iena[9] mprj/la_oenb[0] mprj/la_oenb[100]
+ mprj/la_oenb[101] mprj/la_oenb[102] mprj/la_oenb[103] mprj/la_oenb[104] mprj/la_oenb[105]
+ mprj/la_oenb[106] mprj/la_oenb[107] mprj/la_oenb[108] mprj/la_oenb[109] mprj/la_oenb[10]
+ mprj/la_oenb[110] mprj/la_oenb[111] mprj/la_oenb[112] mprj/la_oenb[113] mprj/la_oenb[114]
+ mprj/la_oenb[115] mprj/la_oenb[116] mprj/la_oenb[117] mprj/la_oenb[118] mprj/la_oenb[119]
+ mprj/la_oenb[11] mprj/la_oenb[120] mprj/la_oenb[121] mprj/la_oenb[122] mprj/la_oenb[123]
+ mprj/la_oenb[124] mprj/la_oenb[125] mprj/la_oenb[126] mprj/la_oenb[127] mprj/la_oenb[12]
+ mprj/la_oenb[13] mprj/la_oenb[14] mprj/la_oenb[15] mprj/la_oenb[16] mprj/la_oenb[17]
+ mprj/la_oenb[18] mprj/la_oenb[19] mprj/la_oenb[1] mprj/la_oenb[20] mprj/la_oenb[21]
+ mprj/la_oenb[22] mprj/la_oenb[23] mprj/la_oenb[24] mprj/la_oenb[25] mprj/la_oenb[26]
+ mprj/la_oenb[27] mprj/la_oenb[28] mprj/la_oenb[29] mprj/la_oenb[2] mprj/la_oenb[30]
+ mprj/la_oenb[31] mprj/la_oenb[32] mprj/la_oenb[33] mprj/la_oenb[34] mprj/la_oenb[35]
+ mprj/la_oenb[36] mprj/la_oenb[37] mprj/la_oenb[38] mprj/la_oenb[39] mprj/la_oenb[3]
+ mprj/la_oenb[40] mprj/la_oenb[41] mprj/la_oenb[42] mprj/la_oenb[43] mprj/la_oenb[44]
+ mprj/la_oenb[45] mprj/la_oenb[46] mprj/la_oenb[47] mprj/la_oenb[48] mprj/la_oenb[49]
+ mprj/la_oenb[4] mprj/la_oenb[50] mprj/la_oenb[51] mprj/la_oenb[52] mprj/la_oenb[53]
+ mprj/la_oenb[54] mprj/la_oenb[55] mprj/la_oenb[56] mprj/la_oenb[57] mprj/la_oenb[58]
+ mprj/la_oenb[59] mprj/la_oenb[5] mprj/la_oenb[60] mprj/la_oenb[61] mprj/la_oenb[62]
+ mprj/la_oenb[63] mprj/la_oenb[64] mprj/la_oenb[65] mprj/la_oenb[66] mprj/la_oenb[67]
+ mprj/la_oenb[68] mprj/la_oenb[69] mprj/la_oenb[6] mprj/la_oenb[70] mprj/la_oenb[71]
+ mprj/la_oenb[72] mprj/la_oenb[73] mprj/la_oenb[74] mprj/la_oenb[75] mprj/la_oenb[76]
+ mprj/la_oenb[77] mprj/la_oenb[78] mprj/la_oenb[79] mprj/la_oenb[7] mprj/la_oenb[80]
+ mprj/la_oenb[81] mprj/la_oenb[82] mprj/la_oenb[83] mprj/la_oenb[84] mprj/la_oenb[85]
+ mprj/la_oenb[86] mprj/la_oenb[87] mprj/la_oenb[88] mprj/la_oenb[89] mprj/la_oenb[8]
+ mprj/la_oenb[90] mprj/la_oenb[91] mprj/la_oenb[92] mprj/la_oenb[93] mprj/la_oenb[94]
+ mprj/la_oenb[95] mprj/la_oenb[96] mprj/la_oenb[97] mprj/la_oenb[98] mprj/la_oenb[99]
+ mprj/la_oenb[9] soc/la_oenb[0] soc/la_oenb[100] soc/la_oenb[101] soc/la_oenb[102]
+ soc/la_oenb[103] soc/la_oenb[104] soc/la_oenb[105] soc/la_oenb[106] soc/la_oenb[107]
+ soc/la_oenb[108] soc/la_oenb[109] soc/la_oenb[10] soc/la_oenb[110] soc/la_oenb[111]
+ soc/la_oenb[112] soc/la_oenb[113] soc/la_oenb[114] soc/la_oenb[115] soc/la_oenb[116]
+ soc/la_oenb[117] soc/la_oenb[118] soc/la_oenb[119] soc/la_oenb[11] soc/la_oenb[120]
+ soc/la_oenb[121] soc/la_oenb[122] soc/la_oenb[123] soc/la_oenb[124] soc/la_oenb[125]
+ soc/la_oenb[126] soc/la_oenb[127] soc/la_oenb[12] soc/la_oenb[13] soc/la_oenb[14]
+ soc/la_oenb[15] soc/la_oenb[16] soc/la_oenb[17] soc/la_oenb[18] soc/la_oenb[19]
+ soc/la_oenb[1] soc/la_oenb[20] soc/la_oenb[21] soc/la_oenb[22] soc/la_oenb[23] soc/la_oenb[24]
+ soc/la_oenb[25] soc/la_oenb[26] soc/la_oenb[27] soc/la_oenb[28] soc/la_oenb[29]
+ soc/la_oenb[2] soc/la_oenb[30] soc/la_oenb[31] soc/la_oenb[32] soc/la_oenb[33] soc/la_oenb[34]
+ soc/la_oenb[35] soc/la_oenb[36] soc/la_oenb[37] soc/la_oenb[38] soc/la_oenb[39]
+ soc/la_oenb[3] soc/la_oenb[40] soc/la_oenb[41] soc/la_oenb[42] soc/la_oenb[43] soc/la_oenb[44]
+ soc/la_oenb[45] soc/la_oenb[46] soc/la_oenb[47] soc/la_oenb[48] soc/la_oenb[49]
+ soc/la_oenb[4] soc/la_oenb[50] soc/la_oenb[51] soc/la_oenb[52] soc/la_oenb[53] soc/la_oenb[54]
+ soc/la_oenb[55] soc/la_oenb[56] soc/la_oenb[57] soc/la_oenb[58] soc/la_oenb[59]
+ soc/la_oenb[5] soc/la_oenb[60] soc/la_oenb[61] soc/la_oenb[62] soc/la_oenb[63] soc/la_oenb[64]
+ soc/la_oenb[65] soc/la_oenb[66] soc/la_oenb[67] soc/la_oenb[68] soc/la_oenb[69]
+ soc/la_oenb[6] soc/la_oenb[70] soc/la_oenb[71] soc/la_oenb[72] soc/la_oenb[73] soc/la_oenb[74]
+ soc/la_oenb[75] soc/la_oenb[76] soc/la_oenb[77] soc/la_oenb[78] soc/la_oenb[79]
+ soc/la_oenb[7] soc/la_oenb[80] soc/la_oenb[81] soc/la_oenb[82] soc/la_oenb[83] soc/la_oenb[84]
+ soc/la_oenb[85] soc/la_oenb[86] soc/la_oenb[87] soc/la_oenb[88] soc/la_oenb[89]
+ soc/la_oenb[8] soc/la_oenb[90] soc/la_oenb[91] soc/la_oenb[92] soc/la_oenb[93] soc/la_oenb[94]
+ soc/la_oenb[95] soc/la_oenb[96] soc/la_oenb[97] soc/la_oenb[98] soc/la_oenb[99]
+ soc/la_oenb[9] soc/mprj_ack_i mprj/wbs_ack_o soc/mprj_adr_o[0] soc/mprj_adr_o[10]
+ soc/mprj_adr_o[11] soc/mprj_adr_o[12] soc/mprj_adr_o[13] soc/mprj_adr_o[14] soc/mprj_adr_o[15]
+ soc/mprj_adr_o[16] soc/mprj_adr_o[17] soc/mprj_adr_o[18] soc/mprj_adr_o[19] soc/mprj_adr_o[1]
+ soc/mprj_adr_o[20] soc/mprj_adr_o[21] soc/mprj_adr_o[22] soc/mprj_adr_o[23] soc/mprj_adr_o[24]
+ soc/mprj_adr_o[25] soc/mprj_adr_o[26] soc/mprj_adr_o[27] soc/mprj_adr_o[28] soc/mprj_adr_o[29]
+ soc/mprj_adr_o[2] soc/mprj_adr_o[30] soc/mprj_adr_o[31] soc/mprj_adr_o[3] soc/mprj_adr_o[4]
+ soc/mprj_adr_o[5] soc/mprj_adr_o[6] soc/mprj_adr_o[7] soc/mprj_adr_o[8] soc/mprj_adr_o[9]
+ mprj/wbs_adr_i[0] mprj/wbs_adr_i[10] mprj/wbs_adr_i[11] mprj/wbs_adr_i[12] mprj/wbs_adr_i[13]
+ mprj/wbs_adr_i[14] mprj/wbs_adr_i[15] mprj/wbs_adr_i[16] mprj/wbs_adr_i[17] mprj/wbs_adr_i[18]
+ mprj/wbs_adr_i[19] mprj/wbs_adr_i[1] mprj/wbs_adr_i[20] mprj/wbs_adr_i[21] mprj/wbs_adr_i[22]
+ mprj/wbs_adr_i[23] mprj/wbs_adr_i[24] mprj/wbs_adr_i[25] mprj/wbs_adr_i[26] mprj/wbs_adr_i[27]
+ mprj/wbs_adr_i[28] mprj/wbs_adr_i[29] mprj/wbs_adr_i[2] mprj/wbs_adr_i[30] mprj/wbs_adr_i[31]
+ mprj/wbs_adr_i[3] mprj/wbs_adr_i[4] mprj/wbs_adr_i[5] mprj/wbs_adr_i[6] mprj/wbs_adr_i[7]
+ mprj/wbs_adr_i[8] mprj/wbs_adr_i[9] soc/mprj_cyc_o mprj/wbs_cyc_i soc/mprj_dat_i[0]
+ soc/mprj_dat_i[10] soc/mprj_dat_i[11] soc/mprj_dat_i[12] soc/mprj_dat_i[13] soc/mprj_dat_i[14]
+ soc/mprj_dat_i[15] soc/mprj_dat_i[16] soc/mprj_dat_i[17] soc/mprj_dat_i[18] soc/mprj_dat_i[19]
+ soc/mprj_dat_i[1] soc/mprj_dat_i[20] soc/mprj_dat_i[21] soc/mprj_dat_i[22] soc/mprj_dat_i[23]
+ soc/mprj_dat_i[24] soc/mprj_dat_i[25] soc/mprj_dat_i[26] soc/mprj_dat_i[27] soc/mprj_dat_i[28]
+ soc/mprj_dat_i[29] soc/mprj_dat_i[2] soc/mprj_dat_i[30] soc/mprj_dat_i[31] soc/mprj_dat_i[3]
+ soc/mprj_dat_i[4] soc/mprj_dat_i[5] soc/mprj_dat_i[6] soc/mprj_dat_i[7] soc/mprj_dat_i[8]
+ soc/mprj_dat_i[9] mprj/wbs_dat_o[0] mprj/wbs_dat_o[10] mprj/wbs_dat_o[11] mprj/wbs_dat_o[12]
+ mprj/wbs_dat_o[13] mprj/wbs_dat_o[14] mprj/wbs_dat_o[15] mprj/wbs_dat_o[16] mprj/wbs_dat_o[17]
+ mprj/wbs_dat_o[18] mprj/wbs_dat_o[19] mprj/wbs_dat_o[1] mprj/wbs_dat_o[20] mprj/wbs_dat_o[21]
+ mprj/wbs_dat_o[22] mprj/wbs_dat_o[23] mprj/wbs_dat_o[24] mprj/wbs_dat_o[25] mprj/wbs_dat_o[26]
+ mprj/wbs_dat_o[27] mprj/wbs_dat_o[28] mprj/wbs_dat_o[29] mprj/wbs_dat_o[2] mprj/wbs_dat_o[30]
+ mprj/wbs_dat_o[31] mprj/wbs_dat_o[3] mprj/wbs_dat_o[4] mprj/wbs_dat_o[5] mprj/wbs_dat_o[6]
+ mprj/wbs_dat_o[7] mprj/wbs_dat_o[8] mprj/wbs_dat_o[9] soc/mprj_dat_o[0] soc/mprj_dat_o[10]
+ soc/mprj_dat_o[11] soc/mprj_dat_o[12] soc/mprj_dat_o[13] soc/mprj_dat_o[14] soc/mprj_dat_o[15]
+ soc/mprj_dat_o[16] soc/mprj_dat_o[17] soc/mprj_dat_o[18] soc/mprj_dat_o[19] soc/mprj_dat_o[1]
+ soc/mprj_dat_o[20] soc/mprj_dat_o[21] soc/mprj_dat_o[22] soc/mprj_dat_o[23] soc/mprj_dat_o[24]
+ soc/mprj_dat_o[25] soc/mprj_dat_o[26] soc/mprj_dat_o[27] soc/mprj_dat_o[28] soc/mprj_dat_o[29]
+ soc/mprj_dat_o[2] soc/mprj_dat_o[30] soc/mprj_dat_o[31] soc/mprj_dat_o[3] soc/mprj_dat_o[4]
+ soc/mprj_dat_o[5] soc/mprj_dat_o[6] soc/mprj_dat_o[7] soc/mprj_dat_o[8] soc/mprj_dat_o[9]
+ mprj/wbs_dat_i[0] mprj/wbs_dat_i[10] mprj/wbs_dat_i[11] mprj/wbs_dat_i[12] mprj/wbs_dat_i[13]
+ mprj/wbs_dat_i[14] mprj/wbs_dat_i[15] mprj/wbs_dat_i[16] mprj/wbs_dat_i[17] mprj/wbs_dat_i[18]
+ mprj/wbs_dat_i[19] mprj/wbs_dat_i[1] mprj/wbs_dat_i[20] mprj/wbs_dat_i[21] mprj/wbs_dat_i[22]
+ mprj/wbs_dat_i[23] mprj/wbs_dat_i[24] mprj/wbs_dat_i[25] mprj/wbs_dat_i[26] mprj/wbs_dat_i[27]
+ mprj/wbs_dat_i[28] mprj/wbs_dat_i[29] mprj/wbs_dat_i[2] mprj/wbs_dat_i[30] mprj/wbs_dat_i[31]
+ mprj/wbs_dat_i[3] mprj/wbs_dat_i[4] mprj/wbs_dat_i[5] mprj/wbs_dat_i[6] mprj/wbs_dat_i[7]
+ mprj/wbs_dat_i[8] mprj/wbs_dat_i[9] soc/mprj_wb_iena soc/mprj_sel_o[0] soc/mprj_sel_o[1]
+ soc/mprj_sel_o[2] soc/mprj_sel_o[3] mprj/wbs_sel_i[0] mprj/wbs_sel_i[1] mprj/wbs_sel_i[2]
+ mprj/wbs_sel_i[3] soc/mprj_stb_o mprj/wbs_stb_i soc/mprj_we_o mprj/wbs_we_i housekeeping/usr1_vcc_pwrgood
+ housekeeping/usr1_vdd_pwrgood housekeeping/usr2_vcc_pwrgood housekeeping/usr2_vdd_pwrgood
+ mprj/wb_clk_i mprj/user_clock2 soc/irq[0] soc/irq[1] soc/irq[2] mprj/user_irq[0]
+ mprj/user_irq[1] mprj/user_irq[2] soc/user_irq_ena[0] soc/user_irq_ena[1] soc/user_irq_ena[2]
+ mprj/wb_rst_i vccd1_core vccd2_core vdda1_core vdda2_core VSUBS dw_394166_241200#
+ dw_386584_241220# vssa2_core vssd2_core vssa1_core dw_193956_239226# dw_263310_241106#
+ vccd_core vssd1_core mgmt_protect
Xrstb_level rstb_level/A pll/resetb por/vdd3v3 vccd_core VSUBS por/vss3v3 xres_buf
Xgpio_defaults_block_9 VSUBS gpio_defaults_block_9/gpio_defaults[0] gpio_defaults_block_9/gpio_defaults[10]
+ gpio_defaults_block_9/gpio_defaults[11] gpio_defaults_block_9/gpio_defaults[12]
+ gpio_defaults_block_9/gpio_defaults[1] gpio_defaults_block_9/gpio_defaults[2] gpio_defaults_block_9/gpio_defaults[3]
+ gpio_defaults_block_9/gpio_defaults[4] gpio_defaults_block_9/gpio_defaults[5] gpio_defaults_block_9/gpio_defaults[6]
+ gpio_defaults_block_9/gpio_defaults[7] gpio_defaults_block_9/gpio_defaults[8] gpio_defaults_block_9/gpio_defaults[9]
+ vccd_core gpio_defaults_block
Xgpio_control_in_2\[15\] gpio_control_in_2\[15\]/gpio_defaults[0] gpio_control_in_2\[15\]/gpio_defaults[10]
+ gpio_control_in_2\[15\]/gpio_defaults[11] gpio_control_in_2\[15\]/gpio_defaults[12]
+ gpio_control_in_2\[15\]/gpio_defaults[1] gpio_control_in_2\[15\]/gpio_defaults[2]
+ gpio_control_in_2\[15\]/gpio_defaults[3] gpio_control_in_2\[15\]/gpio_defaults[4]
+ gpio_control_in_2\[15\]/gpio_defaults[5] gpio_control_in_2\[15\]/gpio_defaults[6]
+ gpio_control_in_2\[15\]/gpio_defaults[7] gpio_control_in_2\[15\]/gpio_defaults[8]
+ gpio_control_in_2\[15\]/gpio_defaults[9] housekeeping/mgmt_gpio_in[34] gpio_control_in_2\[15\]/one
+ housekeeping/mgmt_gpio_in[34] gpio_control_in_2\[15\]/one padframe/mprj_io_analog_en[34]
+ padframe/mprj_io_analog_pol[34] padframe/mprj_io_analog_sel[34] padframe/mprj_io_dm[102]
+ padframe/mprj_io_dm[103] padframe/mprj_io_dm[104] padframe/mprj_io_holdover[34]
+ padframe/mprj_io_ib_mode_sel[34] padframe/mprj_io_in[34] padframe/mprj_io_inp_dis[34]
+ padframe/mprj_io_out[34] padframe/mprj_io_oeb[34] padframe/mprj_io_slow_sel[34]
+ padframe/mprj_io_vtrip_sel[34] gpio_control_in_2\[15\]/resetn gpio_control_in_2\[14\]/resetn
+ gpio_control_in_2\[15\]/serial_clock gpio_control_in_2\[14\]/serial_clock gpio_control_in_2\[15\]/serial_data_in
+ gpio_control_in_2\[14\]/serial_data_in gpio_control_in_2\[15\]/serial_load gpio_control_in_2\[14\]/serial_load
+ mprj/io_in[34] mprj/io_oeb[34] mprj/io_out[34] vccd1_core VSUBS gpio_control_in_2\[15\]/zero
+ dw_8741_333738# vccd_core vssd1_core gpio_control_block
Xgpio_control_bidir_2\[1\] gpio_defaults_block_36/gpio_defaults[0] gpio_defaults_block_36/gpio_defaults[10]
+ gpio_defaults_block_36/gpio_defaults[11] gpio_defaults_block_36/gpio_defaults[12]
+ gpio_defaults_block_36/gpio_defaults[1] gpio_defaults_block_36/gpio_defaults[2]
+ gpio_defaults_block_36/gpio_defaults[3] gpio_defaults_block_36/gpio_defaults[4]
+ gpio_defaults_block_36/gpio_defaults[5] gpio_defaults_block_36/gpio_defaults[6]
+ gpio_defaults_block_36/gpio_defaults[7] gpio_defaults_block_36/gpio_defaults[8]
+ gpio_defaults_block_36/gpio_defaults[9] housekeeping/mgmt_gpio_in[36] housekeeping/mgmt_gpio_oeb[36]
+ housekeeping/mgmt_gpio_out[36] gpio_control_bidir_2\[1\]/one padframe/mprj_io_analog_en[36]
+ padframe/mprj_io_analog_pol[36] padframe/mprj_io_analog_sel[36] padframe/mprj_io_dm[108]
+ padframe/mprj_io_dm[109] padframe/mprj_io_dm[110] padframe/mprj_io_holdover[36]
+ padframe/mprj_io_ib_mode_sel[36] padframe/mprj_io_in[36] padframe/mprj_io_inp_dis[36]
+ padframe/mprj_io_out[36] padframe/mprj_io_oeb[36] padframe/mprj_io_slow_sel[36]
+ padframe/mprj_io_vtrip_sel[36] gpio_control_bidir_2\[1\]/resetn gpio_control_bidir_2\[0\]/resetn
+ gpio_control_bidir_2\[1\]/serial_clock gpio_control_bidir_2\[0\]/serial_clock gpio_control_bidir_2\[1\]/serial_data_in
+ gpio_control_bidir_2\[0\]/serial_data_in gpio_control_bidir_2\[1\]/serial_load gpio_control_bidir_2\[0\]/serial_load
+ mprj/io_in[36] mprj/io_oeb[36] mprj/io_out[36] vccd1_core VSUBS gpio_control_bidir_2\[1\]/zero
+ dw_8741_247338# vccd_core vssd1_core gpio_control_block
Xgpio_control_in_1\[5\] gpio_defaults_block_13/gpio_defaults[0] gpio_defaults_block_13/gpio_defaults[10]
+ gpio_defaults_block_13/gpio_defaults[11] gpio_defaults_block_13/gpio_defaults[12]
+ gpio_defaults_block_13/gpio_defaults[1] gpio_defaults_block_13/gpio_defaults[2]
+ gpio_defaults_block_13/gpio_defaults[3] gpio_defaults_block_13/gpio_defaults[4]
+ gpio_defaults_block_13/gpio_defaults[5] gpio_defaults_block_13/gpio_defaults[6]
+ gpio_defaults_block_13/gpio_defaults[7] gpio_defaults_block_13/gpio_defaults[8]
+ gpio_defaults_block_13/gpio_defaults[9] housekeeping/mgmt_gpio_in[13] gpio_control_in_1\[5\]/one
+ housekeeping/mgmt_gpio_in[13] gpio_control_in_1\[5\]/one padframe/mprj_io_analog_en[13]
+ padframe/mprj_io_analog_pol[13] padframe/mprj_io_analog_sel[13] padframe/mprj_io_dm[39]
+ padframe/mprj_io_dm[40] padframe/mprj_io_dm[41] padframe/mprj_io_holdover[13] padframe/mprj_io_ib_mode_sel[13]
+ padframe/mprj_io_in[13] padframe/mprj_io_inp_dis[13] padframe/mprj_io_out[13] padframe/mprj_io_oeb[13]
+ padframe/mprj_io_slow_sel[13] padframe/mprj_io_vtrip_sel[13] gpio_control_in_1\[5\]/resetn
+ gpio_control_in_1\[6\]/resetn gpio_control_in_1\[5\]/serial_clock gpio_control_in_1\[6\]/serial_clock
+ gpio_control_in_1\[5\]/serial_data_in gpio_control_in_1\[6\]/serial_data_in gpio_control_in_1\[5\]/serial_load
+ gpio_control_in_1\[6\]/serial_load mprj/io_in[13] mprj/io_oeb[13] mprj/io_out[13]
+ vccd1_core VSUBS gpio_control_in_1\[5\]/zero dw_707553_750738# vccd_core vssd1_core
+ gpio_control_block
Xgpio_control_in_2\[13\] gpio_defaults_block_32/gpio_defaults[0] gpio_defaults_block_32/gpio_defaults[10]
+ gpio_defaults_block_32/gpio_defaults[11] gpio_defaults_block_32/gpio_defaults[12]
+ gpio_defaults_block_32/gpio_defaults[1] gpio_defaults_block_32/gpio_defaults[2]
+ gpio_defaults_block_32/gpio_defaults[3] gpio_defaults_block_32/gpio_defaults[4]
+ gpio_defaults_block_32/gpio_defaults[5] gpio_defaults_block_32/gpio_defaults[6]
+ gpio_defaults_block_32/gpio_defaults[7] gpio_defaults_block_32/gpio_defaults[8]
+ gpio_defaults_block_32/gpio_defaults[9] housekeeping/mgmt_gpio_in[32] gpio_control_in_2\[13\]/one
+ housekeeping/mgmt_gpio_in[32] gpio_control_in_2\[13\]/one padframe/mprj_io_analog_en[32]
+ padframe/mprj_io_analog_pol[32] padframe/mprj_io_analog_sel[32] padframe/mprj_io_dm[96]
+ padframe/mprj_io_dm[97] padframe/mprj_io_dm[98] padframe/mprj_io_holdover[32] padframe/mprj_io_ib_mode_sel[32]
+ padframe/mprj_io_in[32] padframe/mprj_io_inp_dis[32] padframe/mprj_io_out[32] padframe/mprj_io_oeb[32]
+ padframe/mprj_io_slow_sel[32] padframe/mprj_io_vtrip_sel[32] gpio_control_in_2\[13\]/resetn
+ gpio_control_in_2\[12\]/resetn gpio_control_in_2\[13\]/serial_clock gpio_control_in_2\[12\]/serial_clock
+ gpio_control_in_2\[13\]/serial_data_in gpio_control_in_2\[12\]/serial_data_in gpio_control_in_2\[13\]/serial_load
+ gpio_control_in_2\[12\]/serial_load mprj/io_in[32] mprj/io_oeb[32] mprj/io_out[32]
+ vccd1_core VSUBS gpio_control_in_2\[13\]/zero dw_8741_420138# vccd_core vssd1_core
+ gpio_control_block
Xgpio_control_in_1a\[2\] gpio_defaults_block_4/gpio_defaults[0] gpio_defaults_block_4/gpio_defaults[10]
+ gpio_defaults_block_4/gpio_defaults[11] gpio_defaults_block_4/gpio_defaults[12]
+ gpio_defaults_block_4/gpio_defaults[1] gpio_defaults_block_4/gpio_defaults[2] gpio_defaults_block_4/gpio_defaults[3]
+ gpio_defaults_block_4/gpio_defaults[4] gpio_defaults_block_4/gpio_defaults[5] gpio_defaults_block_4/gpio_defaults[6]
+ gpio_defaults_block_4/gpio_defaults[7] gpio_defaults_block_4/gpio_defaults[8] gpio_defaults_block_4/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[4] gpio_control_in_1a\[2\]/one housekeeping/mgmt_gpio_in[4]
+ gpio_control_in_1a\[2\]/one padframe/mprj_io_analog_en[4] padframe/mprj_io_analog_pol[4]
+ padframe/mprj_io_analog_sel[4] padframe/mprj_io_dm[12] padframe/mprj_io_dm[13] padframe/mprj_io_dm[14]
+ padframe/mprj_io_holdover[4] padframe/mprj_io_ib_mode_sel[4] padframe/mprj_io_in[4]
+ padframe/mprj_io_inp_dis[4] padframe/mprj_io_out[4] padframe/mprj_io_oeb[4] padframe/mprj_io_slow_sel[4]
+ padframe/mprj_io_vtrip_sel[4] gpio_control_in_1a\[2\]/resetn gpio_control_in_1a\[3\]/resetn
+ gpio_control_in_1a\[2\]/serial_clock gpio_control_in_1a\[3\]/serial_clock gpio_control_in_1a\[2\]/serial_data_in
+ gpio_control_in_1a\[3\]/serial_data_in gpio_control_in_1a\[2\]/serial_load gpio_control_in_1a\[3\]/serial_load
+ mprj/io_in[4] mprj/io_oeb[4] mprj/io_out[4] vccd1_core VSUBS gpio_control_in_1a\[2\]/zero
+ dw_707553_302938# vccd_core vssd1_core gpio_control_block
Xgpio_control_in_2\[8\] gpio_defaults_block_27/gpio_defaults[0] gpio_defaults_block_27/gpio_defaults[10]
+ gpio_defaults_block_27/gpio_defaults[11] gpio_defaults_block_27/gpio_defaults[12]
+ gpio_defaults_block_27/gpio_defaults[1] gpio_defaults_block_27/gpio_defaults[2]
+ gpio_defaults_block_27/gpio_defaults[3] gpio_defaults_block_27/gpio_defaults[4]
+ gpio_defaults_block_27/gpio_defaults[5] gpio_defaults_block_27/gpio_defaults[6]
+ gpio_defaults_block_27/gpio_defaults[7] gpio_defaults_block_27/gpio_defaults[8]
+ gpio_defaults_block_27/gpio_defaults[9] housekeeping/mgmt_gpio_in[27] gpio_control_in_2\[8\]/one
+ housekeeping/mgmt_gpio_in[27] gpio_control_in_2\[8\]/one padframe/mprj_io_analog_en[27]
+ padframe/mprj_io_analog_pol[27] padframe/mprj_io_analog_sel[27] padframe/mprj_io_dm[81]
+ padframe/mprj_io_dm[82] padframe/mprj_io_dm[83] padframe/mprj_io_holdover[27] padframe/mprj_io_ib_mode_sel[27]
+ padframe/mprj_io_in[27] padframe/mprj_io_inp_dis[27] padframe/mprj_io_out[27] padframe/mprj_io_oeb[27]
+ padframe/mprj_io_slow_sel[27] padframe/mprj_io_vtrip_sel[27] gpio_control_in_2\[8\]/resetn
+ gpio_control_in_2\[7\]/resetn gpio_control_in_2\[8\]/serial_clock gpio_control_in_2\[7\]/serial_clock
+ gpio_control_in_2\[8\]/serial_data_in gpio_control_in_2\[7\]/serial_data_in gpio_control_in_2\[8\]/serial_load
+ gpio_control_in_2\[7\]/serial_load mprj/io_in[27] mprj/io_oeb[27] mprj/io_out[27]
+ vccd1_core VSUBS gpio_control_in_2\[8\]/zero dw_8741_720538# vccd_core vssd1_core
+ gpio_control_block
Xgpio_control_in_1\[3\] gpio_defaults_block_11/gpio_defaults[0] gpio_defaults_block_11/gpio_defaults[10]
+ gpio_defaults_block_11/gpio_defaults[11] gpio_defaults_block_11/gpio_defaults[12]
+ gpio_defaults_block_11/gpio_defaults[1] gpio_defaults_block_11/gpio_defaults[2]
+ gpio_defaults_block_11/gpio_defaults[3] gpio_defaults_block_11/gpio_defaults[4]
+ gpio_defaults_block_11/gpio_defaults[5] gpio_defaults_block_11/gpio_defaults[6]
+ gpio_defaults_block_11/gpio_defaults[7] gpio_defaults_block_11/gpio_defaults[8]
+ gpio_defaults_block_11/gpio_defaults[9] housekeeping/mgmt_gpio_in[11] gpio_control_in_1\[3\]/one
+ housekeeping/mgmt_gpio_in[11] gpio_control_in_1\[3\]/one padframe/mprj_io_analog_en[11]
+ padframe/mprj_io_analog_pol[11] padframe/mprj_io_analog_sel[11] padframe/mprj_io_dm[33]
+ padframe/mprj_io_dm[34] padframe/mprj_io_dm[35] padframe/mprj_io_holdover[11] padframe/mprj_io_ib_mode_sel[11]
+ padframe/mprj_io_in[11] padframe/mprj_io_inp_dis[11] padframe/mprj_io_out[11] padframe/mprj_io_oeb[11]
+ padframe/mprj_io_slow_sel[11] padframe/mprj_io_vtrip_sel[11] gpio_control_in_1\[3\]/resetn
+ gpio_control_in_1\[4\]/resetn gpio_control_in_1\[3\]/serial_clock gpio_control_in_1\[4\]/serial_clock
+ gpio_control_in_1\[3\]/serial_data_in gpio_control_in_1\[4\]/serial_data_in gpio_control_in_1\[3\]/serial_load
+ gpio_control_in_1\[4\]/serial_load mprj/io_in[11] mprj/io_oeb[11] mprj/io_out[11]
+ vccd1_core VSUBS gpio_control_in_1\[3\]/zero dw_707553_660538# vccd_core vssd1_core
+ gpio_control_block
Xgpio_control_in_2\[11\] gpio_defaults_block_30/gpio_defaults[0] gpio_defaults_block_30/gpio_defaults[10]
+ gpio_defaults_block_30/gpio_defaults[11] gpio_defaults_block_30/gpio_defaults[12]
+ gpio_defaults_block_30/gpio_defaults[1] gpio_defaults_block_30/gpio_defaults[2]
+ gpio_defaults_block_30/gpio_defaults[3] gpio_defaults_block_30/gpio_defaults[4]
+ gpio_defaults_block_30/gpio_defaults[5] gpio_defaults_block_30/gpio_defaults[6]
+ gpio_defaults_block_30/gpio_defaults[7] gpio_defaults_block_30/gpio_defaults[8]
+ gpio_defaults_block_30/gpio_defaults[9] housekeeping/mgmt_gpio_in[30] gpio_control_in_2\[11\]/one
+ housekeeping/mgmt_gpio_in[30] gpio_control_in_2\[11\]/one padframe/mprj_io_analog_en[30]
+ padframe/mprj_io_analog_pol[30] padframe/mprj_io_analog_sel[30] padframe/mprj_io_dm[90]
+ padframe/mprj_io_dm[91] padframe/mprj_io_dm[92] padframe/mprj_io_holdover[30] padframe/mprj_io_ib_mode_sel[30]
+ padframe/mprj_io_in[30] padframe/mprj_io_inp_dis[30] padframe/mprj_io_out[30] padframe/mprj_io_oeb[30]
+ padframe/mprj_io_slow_sel[30] padframe/mprj_io_vtrip_sel[30] gpio_control_in_2\[11\]/resetn
+ gpio_control_in_2\[10\]/resetn gpio_control_in_2\[11\]/serial_clock gpio_control_in_2\[10\]/serial_clock
+ gpio_control_in_2\[11\]/serial_data_in gpio_control_in_2\[10\]/serial_data_in gpio_control_in_2\[11\]/serial_load
+ gpio_control_in_2\[10\]/serial_load mprj/io_in[30] mprj/io_oeb[30] mprj/io_out[30]
+ vccd1_core VSUBS gpio_control_in_2\[11\]/zero dw_8741_590938# vccd_core vssd1_core
+ gpio_control_block
Xgpio_control_in_1a\[0\] gpio_defaults_block_2/gpio_defaults[0] gpio_defaults_block_2/gpio_defaults[10]
+ gpio_defaults_block_2/gpio_defaults[11] gpio_defaults_block_2/gpio_defaults[12]
+ gpio_defaults_block_2/gpio_defaults[1] gpio_defaults_block_2/gpio_defaults[2] gpio_defaults_block_2/gpio_defaults[3]
+ gpio_defaults_block_2/gpio_defaults[4] gpio_defaults_block_2/gpio_defaults[5] gpio_defaults_block_2/gpio_defaults[6]
+ gpio_defaults_block_2/gpio_defaults[7] gpio_defaults_block_2/gpio_defaults[8] gpio_defaults_block_2/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[2] gpio_control_in_1a\[0\]/one housekeeping/mgmt_gpio_in[2]
+ gpio_control_in_1a\[0\]/one padframe/mprj_io_analog_en[2] padframe/mprj_io_analog_pol[2]
+ padframe/mprj_io_analog_sel[2] padframe/mprj_io_dm[6] padframe/mprj_io_dm[7] padframe/mprj_io_dm[8]
+ padframe/mprj_io_holdover[2] padframe/mprj_io_ib_mode_sel[2] padframe/mprj_io_in[2]
+ padframe/mprj_io_inp_dis[2] padframe/mprj_io_out[2] padframe/mprj_io_oeb[2] padframe/mprj_io_slow_sel[2]
+ padframe/mprj_io_vtrip_sel[2] gpio_control_in_1a\[0\]/resetn gpio_control_in_1a\[1\]/resetn
+ gpio_control_in_1a\[0\]/serial_clock gpio_control_in_1a\[1\]/serial_clock gpio_control_in_1a\[0\]/serial_data_in
+ gpio_control_in_1a\[1\]/serial_data_in gpio_control_in_1a\[0\]/serial_load gpio_control_in_1a\[1\]/serial_load
+ mprj/io_in[2] mprj/io_oeb[2] mprj/io_out[2] vccd1_core VSUBS gpio_control_in_1a\[0\]/zero
+ dw_707553_212738# vccd_core vssd1_core gpio_control_block
Xgpio_control_in_2\[6\] gpio_defaults_block_25/gpio_defaults[0] gpio_defaults_block_25/gpio_defaults[10]
+ gpio_defaults_block_25/gpio_defaults[11] gpio_defaults_block_25/gpio_defaults[12]
+ gpio_defaults_block_25/gpio_defaults[1] gpio_defaults_block_25/gpio_defaults[2]
+ gpio_defaults_block_25/gpio_defaults[3] gpio_defaults_block_25/gpio_defaults[4]
+ gpio_defaults_block_25/gpio_defaults[5] gpio_defaults_block_25/gpio_defaults[6]
+ gpio_defaults_block_25/gpio_defaults[7] gpio_defaults_block_25/gpio_defaults[8]
+ gpio_defaults_block_25/gpio_defaults[9] housekeeping/mgmt_gpio_in[25] gpio_control_in_2\[6\]/one
+ housekeeping/mgmt_gpio_in[25] gpio_control_in_2\[6\]/one padframe/mprj_io_analog_en[25]
+ padframe/mprj_io_analog_pol[25] padframe/mprj_io_analog_sel[25] padframe/mprj_io_dm[75]
+ padframe/mprj_io_dm[76] padframe/mprj_io_dm[77] padframe/mprj_io_holdover[25] padframe/mprj_io_ib_mode_sel[25]
+ padframe/mprj_io_in[25] padframe/mprj_io_inp_dis[25] padframe/mprj_io_out[25] padframe/mprj_io_oeb[25]
+ padframe/mprj_io_slow_sel[25] padframe/mprj_io_vtrip_sel[25] gpio_control_in_2\[6\]/resetn
+ gpio_control_in_2\[5\]/resetn gpio_control_in_2\[6\]/serial_clock gpio_control_in_2\[5\]/serial_clock
+ gpio_control_in_2\[6\]/serial_data_in gpio_control_in_2\[5\]/serial_data_in gpio_control_in_2\[6\]/serial_load
+ gpio_control_in_2\[5\]/serial_load mprj/io_in[25] mprj/io_oeb[25] mprj/io_out[25]
+ vccd1_core VSUBS gpio_control_in_2\[6\]/zero dw_8741_806938# vccd_core vssd1_core
+ gpio_control_block
Xgpio_control_in_1\[1\] gpio_defaults_block_9/gpio_defaults[0] gpio_defaults_block_9/gpio_defaults[10]
+ gpio_defaults_block_9/gpio_defaults[11] gpio_defaults_block_9/gpio_defaults[12]
+ gpio_defaults_block_9/gpio_defaults[1] gpio_defaults_block_9/gpio_defaults[2] gpio_defaults_block_9/gpio_defaults[3]
+ gpio_defaults_block_9/gpio_defaults[4] gpio_defaults_block_9/gpio_defaults[5] gpio_defaults_block_9/gpio_defaults[6]
+ gpio_defaults_block_9/gpio_defaults[7] gpio_defaults_block_9/gpio_defaults[8] gpio_defaults_block_9/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[9] gpio_control_in_1\[1\]/one housekeeping/mgmt_gpio_in[9]
+ gpio_control_in_1\[1\]/one padframe/mprj_io_analog_en[9] padframe/mprj_io_analog_pol[9]
+ padframe/mprj_io_analog_sel[9] padframe/mprj_io_dm[27] padframe/mprj_io_dm[28] padframe/mprj_io_dm[29]
+ padframe/mprj_io_holdover[9] padframe/mprj_io_ib_mode_sel[9] padframe/mprj_io_in[9]
+ padframe/mprj_io_inp_dis[9] padframe/mprj_io_out[9] padframe/mprj_io_oeb[9] padframe/mprj_io_slow_sel[9]
+ padframe/mprj_io_vtrip_sel[9] gpio_control_in_1\[1\]/resetn gpio_control_in_1\[2\]/resetn
+ gpio_control_in_1\[1\]/serial_clock gpio_control_in_1\[2\]/serial_clock gpio_control_in_1\[1\]/serial_data_in
+ gpio_control_in_1\[2\]/serial_data_in gpio_control_in_1\[1\]/serial_load gpio_control_in_1\[2\]/serial_load
+ mprj/io_in[9] mprj/io_oeb[9] mprj/io_out[9] vccd1_core VSUBS gpio_control_in_1\[1\]/zero
+ dw_707553_570338# vccd_core vssd1_core gpio_control_block
Xmprj mprj/analog_io[0] mprj/analog_io[10] mprj/analog_io[11] mprj/analog_io[12] mprj/analog_io[13]
+ mprj/analog_io[14] mprj/analog_io[15] mprj/analog_io[16] mprj/analog_io[17] mprj/analog_io[18]
+ mprj/analog_io[19] mprj/analog_io[1] mprj/analog_io[20] mprj/analog_io[21] mprj/analog_io[22]
+ mprj/analog_io[23] mprj/analog_io[24] mprj/analog_io[25] mprj/analog_io[26] mprj/analog_io[27]
+ mprj/analog_io[28] mprj/analog_io[2] mprj/analog_io[3] mprj/analog_io[4] mprj/analog_io[5]
+ mprj/analog_io[6] mprj/analog_io[7] mprj/analog_io[8] mprj/analog_io[9] mprj/io_in[0]
+ mprj/io_in[10] mprj/io_in[11] mprj/io_in[12] mprj/io_in[13] mprj/io_in[14] mprj/io_in[15]
+ mprj/io_in[16] mprj/io_in[17] mprj/io_in[18] mprj/io_in[19] mprj/io_in[1] mprj/io_in[20]
+ mprj/io_in[21] mprj/io_in[22] mprj/io_in[23] mprj/io_in[24] mprj/io_in[25] mprj/io_in[26]
+ mprj/io_in[27] mprj/io_in[28] mprj/io_in[29] mprj/io_in[2] mprj/io_in[30] mprj/io_in[31]
+ mprj/io_in[32] mprj/io_in[33] mprj/io_in[34] mprj/io_in[35] mprj/io_in[36] mprj/io_in[37]
+ mprj/io_in[3] mprj/io_in[4] mprj/io_in[5] mprj/io_in[6] mprj/io_in[7] mprj/io_in[8]
+ mprj/io_in[9] mprj/io_oeb[0] mprj/io_oeb[10] mprj/io_oeb[11] mprj/io_oeb[12] mprj/io_oeb[13]
+ mprj/io_oeb[14] mprj/io_oeb[15] mprj/io_oeb[16] mprj/io_oeb[17] mprj/io_oeb[18]
+ mprj/io_oeb[19] mprj/io_oeb[1] mprj/io_oeb[20] mprj/io_oeb[21] mprj/io_oeb[22] mprj/io_oeb[23]
+ mprj/io_oeb[24] mprj/io_oeb[25] mprj/io_oeb[26] mprj/io_oeb[27] mprj/io_oeb[28]
+ mprj/io_oeb[29] mprj/io_oeb[2] mprj/io_oeb[30] mprj/io_oeb[31] mprj/io_oeb[32] mprj/io_oeb[33]
+ mprj/io_oeb[34] mprj/io_oeb[35] mprj/io_oeb[36] mprj/io_oeb[37] mprj/io_oeb[3] mprj/io_oeb[4]
+ mprj/io_oeb[5] mprj/io_oeb[6] mprj/io_oeb[7] mprj/io_oeb[8] mprj/io_oeb[9] mprj/io_out[0]
+ mprj/io_out[10] mprj/io_out[11] mprj/io_out[12] mprj/io_out[13] mprj/io_out[14]
+ mprj/io_out[15] mprj/io_out[16] mprj/io_out[17] mprj/io_out[18] mprj/io_out[19]
+ mprj/io_out[1] mprj/io_out[20] mprj/io_out[21] mprj/io_out[22] mprj/io_out[23] mprj/io_out[24]
+ mprj/io_out[25] mprj/io_out[26] mprj/io_out[27] mprj/io_out[28] mprj/io_out[29]
+ mprj/io_out[2] mprj/io_out[30] mprj/io_out[31] mprj/io_out[32] mprj/io_out[33] mprj/io_out[34]
+ mprj/io_out[35] mprj/io_out[36] mprj/io_out[37] mprj/io_out[3] mprj/io_out[4] mprj/io_out[5]
+ mprj/io_out[6] mprj/io_out[7] mprj/io_out[8] mprj/io_out[9] mprj/la_data_in[0] mprj/la_data_in[100]
+ mprj/la_data_in[101] mprj/la_data_in[102] mprj/la_data_in[103] mprj/la_data_in[104]
+ mprj/la_data_in[105] mprj/la_data_in[106] mprj/la_data_in[107] mprj/la_data_in[108]
+ mprj/la_data_in[109] mprj/la_data_in[10] mprj/la_data_in[110] mprj/la_data_in[111]
+ mprj/la_data_in[112] mprj/la_data_in[113] mprj/la_data_in[114] mprj/la_data_in[115]
+ mprj/la_data_in[116] mprj/la_data_in[117] mprj/la_data_in[118] mprj/la_data_in[119]
+ mprj/la_data_in[11] mprj/la_data_in[120] mprj/la_data_in[121] mprj/la_data_in[122]
+ mprj/la_data_in[123] mprj/la_data_in[124] mprj/la_data_in[125] mprj/la_data_in[126]
+ mprj/la_data_in[127] mprj/la_data_in[12] mprj/la_data_in[13] mprj/la_data_in[14]
+ mprj/la_data_in[15] mprj/la_data_in[16] mprj/la_data_in[17] mprj/la_data_in[18]
+ mprj/la_data_in[19] mprj/la_data_in[1] mprj/la_data_in[20] mprj/la_data_in[21] mprj/la_data_in[22]
+ mprj/la_data_in[23] mprj/la_data_in[24] mprj/la_data_in[25] mprj/la_data_in[26]
+ mprj/la_data_in[27] mprj/la_data_in[28] mprj/la_data_in[29] mprj/la_data_in[2] mprj/la_data_in[30]
+ mprj/la_data_in[31] mprj/la_data_in[32] mprj/la_data_in[33] mprj/la_data_in[34]
+ mprj/la_data_in[35] mprj/la_data_in[36] mprj/la_data_in[37] mprj/la_data_in[38]
+ mprj/la_data_in[39] mprj/la_data_in[3] mprj/la_data_in[40] mprj/la_data_in[41] mprj/la_data_in[42]
+ mprj/la_data_in[43] mprj/la_data_in[44] mprj/la_data_in[45] mprj/la_data_in[46]
+ mprj/la_data_in[47] mprj/la_data_in[48] mprj/la_data_in[49] mprj/la_data_in[4] mprj/la_data_in[50]
+ mprj/la_data_in[51] mprj/la_data_in[52] mprj/la_data_in[53] mprj/la_data_in[54]
+ mprj/la_data_in[55] mprj/la_data_in[56] mprj/la_data_in[57] mprj/la_data_in[58]
+ mprj/la_data_in[59] mprj/la_data_in[5] mprj/la_data_in[60] mprj/la_data_in[61] mprj/la_data_in[62]
+ mprj/la_data_in[63] mprj/la_data_in[64] mprj/la_data_in[65] mprj/la_data_in[66]
+ mprj/la_data_in[67] mprj/la_data_in[68] mprj/la_data_in[69] mprj/la_data_in[6] mprj/la_data_in[70]
+ mprj/la_data_in[71] mprj/la_data_in[72] mprj/la_data_in[73] mprj/la_data_in[74]
+ mprj/la_data_in[75] mprj/la_data_in[76] mprj/la_data_in[77] mprj/la_data_in[78]
+ mprj/la_data_in[79] mprj/la_data_in[7] mprj/la_data_in[80] mprj/la_data_in[81] mprj/la_data_in[82]
+ mprj/la_data_in[83] mprj/la_data_in[84] mprj/la_data_in[85] mprj/la_data_in[86]
+ mprj/la_data_in[87] mprj/la_data_in[88] mprj/la_data_in[89] mprj/la_data_in[8] mprj/la_data_in[90]
+ mprj/la_data_in[91] mprj/la_data_in[92] mprj/la_data_in[93] mprj/la_data_in[94]
+ mprj/la_data_in[95] mprj/la_data_in[96] mprj/la_data_in[97] mprj/la_data_in[98]
+ mprj/la_data_in[99] mprj/la_data_in[9] mprj/la_data_out[0] mprj/la_data_out[100]
+ mprj/la_data_out[101] mprj/la_data_out[102] mprj/la_data_out[103] mprj/la_data_out[104]
+ mprj/la_data_out[105] mprj/la_data_out[106] mprj/la_data_out[107] mprj/la_data_out[108]
+ mprj/la_data_out[109] mprj/la_data_out[10] mprj/la_data_out[110] mprj/la_data_out[111]
+ mprj/la_data_out[112] mprj/la_data_out[113] mprj/la_data_out[114] mprj/la_data_out[115]
+ mprj/la_data_out[116] mprj/la_data_out[117] mprj/la_data_out[118] mprj/la_data_out[119]
+ mprj/la_data_out[11] mprj/la_data_out[120] mprj/la_data_out[121] mprj/la_data_out[122]
+ mprj/la_data_out[123] mprj/la_data_out[124] mprj/la_data_out[125] mprj/la_data_out[126]
+ mprj/la_data_out[127] mprj/la_data_out[12] mprj/la_data_out[13] mprj/la_data_out[14]
+ mprj/la_data_out[15] mprj/la_data_out[16] mprj/la_data_out[17] mprj/la_data_out[18]
+ mprj/la_data_out[19] mprj/la_data_out[1] mprj/la_data_out[20] mprj/la_data_out[21]
+ mprj/la_data_out[22] mprj/la_data_out[23] mprj/la_data_out[24] mprj/la_data_out[25]
+ mprj/la_data_out[26] mprj/la_data_out[27] mprj/la_data_out[28] mprj/la_data_out[29]
+ mprj/la_data_out[2] mprj/la_data_out[30] mprj/la_data_out[31] mprj/la_data_out[32]
+ mprj/la_data_out[33] mprj/la_data_out[34] mprj/la_data_out[35] mprj/la_data_out[36]
+ mprj/la_data_out[37] mprj/la_data_out[38] mprj/la_data_out[39] mprj/la_data_out[3]
+ mprj/la_data_out[40] mprj/la_data_out[41] mprj/la_data_out[42] mprj/la_data_out[43]
+ mprj/la_data_out[44] mprj/la_data_out[45] mprj/la_data_out[46] mprj/la_data_out[47]
+ mprj/la_data_out[48] mprj/la_data_out[49] mprj/la_data_out[4] mprj/la_data_out[50]
+ mprj/la_data_out[51] mprj/la_data_out[52] mprj/la_data_out[53] mprj/la_data_out[54]
+ mprj/la_data_out[55] mprj/la_data_out[56] mprj/la_data_out[57] mprj/la_data_out[58]
+ mprj/la_data_out[59] mprj/la_data_out[5] mprj/la_data_out[60] mprj/la_data_out[61]
+ mprj/la_data_out[62] mprj/la_data_out[63] mprj/la_data_out[64] mprj/la_data_out[65]
+ mprj/la_data_out[66] mprj/la_data_out[67] mprj/la_data_out[68] mprj/la_data_out[69]
+ mprj/la_data_out[6] mprj/la_data_out[70] mprj/la_data_out[71] mprj/la_data_out[72]
+ mprj/la_data_out[73] mprj/la_data_out[74] mprj/la_data_out[75] mprj/la_data_out[76]
+ mprj/la_data_out[77] mprj/la_data_out[78] mprj/la_data_out[79] mprj/la_data_out[7]
+ mprj/la_data_out[80] mprj/la_data_out[81] mprj/la_data_out[82] mprj/la_data_out[83]
+ mprj/la_data_out[84] mprj/la_data_out[85] mprj/la_data_out[86] mprj/la_data_out[87]
+ mprj/la_data_out[88] mprj/la_data_out[89] mprj/la_data_out[8] mprj/la_data_out[90]
+ mprj/la_data_out[91] mprj/la_data_out[92] mprj/la_data_out[93] mprj/la_data_out[94]
+ mprj/la_data_out[95] mprj/la_data_out[96] mprj/la_data_out[97] mprj/la_data_out[98]
+ mprj/la_data_out[99] mprj/la_data_out[9] mprj/la_oenb[0] mprj/la_oenb[100] mprj/la_oenb[101]
+ mprj/la_oenb[102] mprj/la_oenb[103] mprj/la_oenb[104] mprj/la_oenb[105] mprj/la_oenb[106]
+ mprj/la_oenb[107] mprj/la_oenb[108] mprj/la_oenb[109] mprj/la_oenb[10] mprj/la_oenb[110]
+ mprj/la_oenb[111] mprj/la_oenb[112] mprj/la_oenb[113] mprj/la_oenb[114] mprj/la_oenb[115]
+ mprj/la_oenb[116] mprj/la_oenb[117] mprj/la_oenb[118] mprj/la_oenb[119] mprj/la_oenb[11]
+ mprj/la_oenb[120] mprj/la_oenb[121] mprj/la_oenb[122] mprj/la_oenb[123] mprj/la_oenb[124]
+ mprj/la_oenb[125] mprj/la_oenb[126] mprj/la_oenb[127] mprj/la_oenb[12] mprj/la_oenb[13]
+ mprj/la_oenb[14] mprj/la_oenb[15] mprj/la_oenb[16] mprj/la_oenb[17] mprj/la_oenb[18]
+ mprj/la_oenb[19] mprj/la_oenb[1] mprj/la_oenb[20] mprj/la_oenb[21] mprj/la_oenb[22]
+ mprj/la_oenb[23] mprj/la_oenb[24] mprj/la_oenb[25] mprj/la_oenb[26] mprj/la_oenb[27]
+ mprj/la_oenb[28] mprj/la_oenb[29] mprj/la_oenb[2] mprj/la_oenb[30] mprj/la_oenb[31]
+ mprj/la_oenb[32] mprj/la_oenb[33] mprj/la_oenb[34] mprj/la_oenb[35] mprj/la_oenb[36]
+ mprj/la_oenb[37] mprj/la_oenb[38] mprj/la_oenb[39] mprj/la_oenb[3] mprj/la_oenb[40]
+ mprj/la_oenb[41] mprj/la_oenb[42] mprj/la_oenb[43] mprj/la_oenb[44] mprj/la_oenb[45]
+ mprj/la_oenb[46] mprj/la_oenb[47] mprj/la_oenb[48] mprj/la_oenb[49] mprj/la_oenb[4]
+ mprj/la_oenb[50] mprj/la_oenb[51] mprj/la_oenb[52] mprj/la_oenb[53] mprj/la_oenb[54]
+ mprj/la_oenb[55] mprj/la_oenb[56] mprj/la_oenb[57] mprj/la_oenb[58] mprj/la_oenb[59]
+ mprj/la_oenb[5] mprj/la_oenb[60] mprj/la_oenb[61] mprj/la_oenb[62] mprj/la_oenb[63]
+ mprj/la_oenb[64] mprj/la_oenb[65] mprj/la_oenb[66] mprj/la_oenb[67] mprj/la_oenb[68]
+ mprj/la_oenb[69] mprj/la_oenb[6] mprj/la_oenb[70] mprj/la_oenb[71] mprj/la_oenb[72]
+ mprj/la_oenb[73] mprj/la_oenb[74] mprj/la_oenb[75] mprj/la_oenb[76] mprj/la_oenb[77]
+ mprj/la_oenb[78] mprj/la_oenb[79] mprj/la_oenb[7] mprj/la_oenb[80] mprj/la_oenb[81]
+ mprj/la_oenb[82] mprj/la_oenb[83] mprj/la_oenb[84] mprj/la_oenb[85] mprj/la_oenb[86]
+ mprj/la_oenb[87] mprj/la_oenb[88] mprj/la_oenb[89] mprj/la_oenb[8] mprj/la_oenb[90]
+ mprj/la_oenb[91] mprj/la_oenb[92] mprj/la_oenb[93] mprj/la_oenb[94] mprj/la_oenb[95]
+ mprj/la_oenb[96] mprj/la_oenb[97] mprj/la_oenb[98] mprj/la_oenb[99] mprj/la_oenb[9]
+ mprj/user_clock2 mprj/user_irq[0] mprj/user_irq[1] mprj/user_irq[2] vccd1_core vccd2_core
+ vdda1_core vdda2_core vssa1_core vssa2_core vssd1_core vssd2_core mprj/wb_clk_i
+ mprj/wb_rst_i mprj/wbs_ack_o mprj/wbs_adr_i[0] mprj/wbs_adr_i[10] mprj/wbs_adr_i[11]
+ mprj/wbs_adr_i[12] mprj/wbs_adr_i[13] mprj/wbs_adr_i[14] mprj/wbs_adr_i[15] mprj/wbs_adr_i[16]
+ mprj/wbs_adr_i[17] mprj/wbs_adr_i[18] mprj/wbs_adr_i[19] mprj/wbs_adr_i[1] mprj/wbs_adr_i[20]
+ mprj/wbs_adr_i[21] mprj/wbs_adr_i[22] mprj/wbs_adr_i[23] mprj/wbs_adr_i[24] mprj/wbs_adr_i[25]
+ mprj/wbs_adr_i[26] mprj/wbs_adr_i[27] mprj/wbs_adr_i[28] mprj/wbs_adr_i[29] mprj/wbs_adr_i[2]
+ mprj/wbs_adr_i[30] mprj/wbs_adr_i[31] mprj/wbs_adr_i[3] mprj/wbs_adr_i[4] mprj/wbs_adr_i[5]
+ mprj/wbs_adr_i[6] mprj/wbs_adr_i[7] mprj/wbs_adr_i[8] mprj/wbs_adr_i[9] mprj/wbs_cyc_i
+ mprj/wbs_dat_i[0] mprj/wbs_dat_i[10] mprj/wbs_dat_i[11] mprj/wbs_dat_i[12] mprj/wbs_dat_i[13]
+ mprj/wbs_dat_i[14] mprj/wbs_dat_i[15] mprj/wbs_dat_i[16] mprj/wbs_dat_i[17] mprj/wbs_dat_i[18]
+ mprj/wbs_dat_i[19] mprj/wbs_dat_i[1] mprj/wbs_dat_i[20] mprj/wbs_dat_i[21] mprj/wbs_dat_i[22]
+ mprj/wbs_dat_i[23] mprj/wbs_dat_i[24] mprj/wbs_dat_i[25] mprj/wbs_dat_i[26] mprj/wbs_dat_i[27]
+ mprj/wbs_dat_i[28] mprj/wbs_dat_i[29] mprj/wbs_dat_i[2] mprj/wbs_dat_i[30] mprj/wbs_dat_i[31]
+ mprj/wbs_dat_i[3] mprj/wbs_dat_i[4] mprj/wbs_dat_i[5] mprj/wbs_dat_i[6] mprj/wbs_dat_i[7]
+ mprj/wbs_dat_i[8] mprj/wbs_dat_i[9] mprj/wbs_dat_o[0] mprj/wbs_dat_o[10] mprj/wbs_dat_o[11]
+ mprj/wbs_dat_o[12] mprj/wbs_dat_o[13] mprj/wbs_dat_o[14] mprj/wbs_dat_o[15] mprj/wbs_dat_o[16]
+ mprj/wbs_dat_o[17] mprj/wbs_dat_o[18] mprj/wbs_dat_o[19] mprj/wbs_dat_o[1] mprj/wbs_dat_o[20]
+ mprj/wbs_dat_o[21] mprj/wbs_dat_o[22] mprj/wbs_dat_o[23] mprj/wbs_dat_o[24] mprj/wbs_dat_o[25]
+ mprj/wbs_dat_o[26] mprj/wbs_dat_o[27] mprj/wbs_dat_o[28] mprj/wbs_dat_o[29] mprj/wbs_dat_o[2]
+ mprj/wbs_dat_o[30] mprj/wbs_dat_o[31] mprj/wbs_dat_o[3] mprj/wbs_dat_o[4] mprj/wbs_dat_o[5]
+ mprj/wbs_dat_o[6] mprj/wbs_dat_o[7] mprj/wbs_dat_o[8] mprj/wbs_dat_o[9] mprj/wbs_sel_i[0]
+ mprj/wbs_sel_i[1] mprj/wbs_sel_i[2] mprj/wbs_sel_i[3] mprj/wbs_stb_i mprj/wbs_we_i
+ user_project_wrapper
Xgpio_control_in_2\[4\] gpio_defaults_block_23/gpio_defaults[0] gpio_defaults_block_23/gpio_defaults[10]
+ gpio_defaults_block_23/gpio_defaults[11] gpio_defaults_block_23/gpio_defaults[12]
+ gpio_defaults_block_23/gpio_defaults[1] gpio_defaults_block_23/gpio_defaults[2]
+ gpio_defaults_block_23/gpio_defaults[3] gpio_defaults_block_23/gpio_defaults[4]
+ gpio_defaults_block_23/gpio_defaults[5] gpio_defaults_block_23/gpio_defaults[6]
+ gpio_defaults_block_23/gpio_defaults[7] gpio_defaults_block_23/gpio_defaults[8]
+ gpio_defaults_block_23/gpio_defaults[9] housekeeping/mgmt_gpio_in[23] gpio_control_in_2\[4\]/one
+ housekeeping/mgmt_gpio_in[23] gpio_control_in_2\[4\]/one padframe/mprj_io_analog_en[23]
+ padframe/mprj_io_analog_pol[23] padframe/mprj_io_analog_sel[23] padframe/mprj_io_dm[69]
+ padframe/mprj_io_dm[70] padframe/mprj_io_dm[71] padframe/mprj_io_holdover[23] padframe/mprj_io_ib_mode_sel[23]
+ padframe/mprj_io_in[23] padframe/mprj_io_inp_dis[23] padframe/mprj_io_out[23] padframe/mprj_io_oeb[23]
+ padframe/mprj_io_slow_sel[23] padframe/mprj_io_vtrip_sel[23] gpio_control_in_2\[4\]/resetn
+ gpio_control_in_2\[3\]/resetn gpio_control_in_2\[4\]/serial_clock gpio_control_in_2\[3\]/serial_clock
+ gpio_control_in_2\[4\]/serial_data_in gpio_control_in_2\[3\]/serial_data_in gpio_control_in_2\[4\]/serial_load
+ gpio_control_in_2\[3\]/serial_load mprj/io_in[23] mprj/io_oeb[23] mprj/io_out[23]
+ vccd1_core VSUBS gpio_control_in_2\[4\]/zero dw_98738_1027427# vccd_core vssd1_core
+ gpio_control_block
Xgpio_control_bidir_1\[1\] gpio_defaults_block_1/gpio_defaults[0] gpio_defaults_block_1/gpio_defaults[10]
+ gpio_defaults_block_1/gpio_defaults[11] gpio_defaults_block_1/gpio_defaults[12]
+ gpio_defaults_block_1/gpio_defaults[1] gpio_defaults_block_1/gpio_defaults[2] gpio_defaults_block_1/gpio_defaults[3]
+ gpio_defaults_block_1/gpio_defaults[4] gpio_defaults_block_1/gpio_defaults[5] gpio_defaults_block_1/gpio_defaults[6]
+ gpio_defaults_block_1/gpio_defaults[7] gpio_defaults_block_1/gpio_defaults[8] gpio_defaults_block_1/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[1] housekeeping/mgmt_gpio_oeb[1] housekeeping/mgmt_gpio_out[1]
+ gpio_control_bidir_1\[1\]/one padframe/mprj_io_analog_en[1] padframe/mprj_io_analog_pol[1]
+ padframe/mprj_io_analog_sel[1] padframe/mprj_io_dm[3] padframe/mprj_io_dm[4] padframe/mprj_io_dm[5]
+ padframe/mprj_io_holdover[1] padframe/mprj_io_ib_mode_sel[1] padframe/mprj_io_in[1]
+ padframe/mprj_io_inp_dis[1] padframe/mprj_io_out[1] padframe/mprj_io_oeb[1] padframe/mprj_io_slow_sel[1]
+ padframe/mprj_io_vtrip_sel[1] gpio_control_bidir_1\[1\]/resetn gpio_control_in_1a\[0\]/resetn
+ gpio_control_bidir_1\[1\]/serial_clock gpio_control_in_1a\[0\]/serial_clock gpio_control_bidir_1\[1\]/serial_data_in
+ gpio_control_in_1a\[0\]/serial_data_in gpio_control_bidir_1\[1\]/serial_load gpio_control_in_1a\[0\]/serial_load
+ mprj/io_in[1] mprj/io_oeb[1] mprj/io_out[1] vccd1_core VSUBS gpio_control_bidir_1\[1\]/zero
+ dw_707553_167738# vccd_core vssd1_core gpio_control_block
Xhousekeeping soc/debug_in soc/debug_mode soc/debug_oeb soc/debug_out soc/irq[3] soc/irq[4]
+ soc/irq[5] user_id_value/mask_rev[0] user_id_value/mask_rev[10] user_id_value/mask_rev[11]
+ user_id_value/mask_rev[12] user_id_value/mask_rev[13] user_id_value/mask_rev[14]
+ user_id_value/mask_rev[15] user_id_value/mask_rev[16] user_id_value/mask_rev[17]
+ user_id_value/mask_rev[18] user_id_value/mask_rev[19] user_id_value/mask_rev[1]
+ user_id_value/mask_rev[20] user_id_value/mask_rev[21] user_id_value/mask_rev[22]
+ user_id_value/mask_rev[23] user_id_value/mask_rev[24] user_id_value/mask_rev[25]
+ user_id_value/mask_rev[26] user_id_value/mask_rev[27] user_id_value/mask_rev[28]
+ user_id_value/mask_rev[29] user_id_value/mask_rev[2] user_id_value/mask_rev[30]
+ user_id_value/mask_rev[31] user_id_value/mask_rev[3] user_id_value/mask_rev[4] user_id_value/mask_rev[5]
+ user_id_value/mask_rev[6] user_id_value/mask_rev[7] user_id_value/mask_rev[8] user_id_value/mask_rev[9]
+ housekeeping/mgmt_gpio_in[0] housekeeping/mgmt_gpio_in[10] housekeeping/mgmt_gpio_in[11]
+ housekeeping/mgmt_gpio_in[12] housekeeping/mgmt_gpio_in[13] housekeeping/mgmt_gpio_in[14]
+ housekeeping/mgmt_gpio_in[15] housekeeping/mgmt_gpio_in[16] housekeeping/mgmt_gpio_in[17]
+ housekeeping/mgmt_gpio_in[18] housekeeping/mgmt_gpio_in[19] housekeeping/mgmt_gpio_in[1]
+ housekeeping/mgmt_gpio_in[20] housekeeping/mgmt_gpio_in[21] housekeeping/mgmt_gpio_in[22]
+ housekeeping/mgmt_gpio_in[23] housekeeping/mgmt_gpio_in[24] housekeeping/mgmt_gpio_in[25]
+ housekeeping/mgmt_gpio_in[26] housekeeping/mgmt_gpio_in[27] housekeeping/mgmt_gpio_in[28]
+ housekeeping/mgmt_gpio_in[29] housekeeping/mgmt_gpio_in[2] housekeeping/mgmt_gpio_in[30]
+ housekeeping/mgmt_gpio_in[31] housekeeping/mgmt_gpio_in[32] housekeeping/mgmt_gpio_in[33]
+ housekeeping/mgmt_gpio_in[34] housekeeping/mgmt_gpio_in[35] housekeeping/mgmt_gpio_in[36]
+ housekeeping/mgmt_gpio_in[37] housekeeping/mgmt_gpio_in[3] housekeeping/mgmt_gpio_in[4]
+ housekeeping/mgmt_gpio_in[5] housekeeping/mgmt_gpio_in[6] housekeeping/mgmt_gpio_in[7]
+ housekeeping/mgmt_gpio_in[8] housekeeping/mgmt_gpio_in[9] housekeeping/mgmt_gpio_oeb[0]
+ housekeeping/mgmt_gpio_oeb[10] housekeeping/mgmt_gpio_oeb[11] housekeeping/mgmt_gpio_oeb[12]
+ housekeeping/mgmt_gpio_oeb[13] housekeeping/mgmt_gpio_oeb[14] housekeeping/mgmt_gpio_oeb[15]
+ housekeeping/mgmt_gpio_oeb[16] housekeeping/mgmt_gpio_oeb[17] housekeeping/mgmt_gpio_oeb[18]
+ housekeeping/mgmt_gpio_oeb[19] housekeeping/mgmt_gpio_oeb[1] housekeeping/mgmt_gpio_oeb[20]
+ housekeeping/mgmt_gpio_oeb[21] housekeeping/mgmt_gpio_oeb[22] housekeeping/mgmt_gpio_oeb[23]
+ housekeeping/mgmt_gpio_oeb[24] housekeeping/mgmt_gpio_oeb[25] housekeeping/mgmt_gpio_oeb[26]
+ housekeeping/mgmt_gpio_oeb[27] housekeeping/mgmt_gpio_oeb[28] housekeeping/mgmt_gpio_oeb[29]
+ housekeeping/mgmt_gpio_oeb[2] housekeeping/mgmt_gpio_oeb[30] housekeeping/mgmt_gpio_oeb[31]
+ housekeeping/mgmt_gpio_oeb[32] housekeeping/mgmt_gpio_oeb[33] housekeeping/mgmt_gpio_oeb[34]
+ housekeeping/mgmt_gpio_oeb[35] housekeeping/mgmt_gpio_oeb[36] housekeeping/mgmt_gpio_oeb[37]
+ housekeeping/mgmt_gpio_oeb[3] housekeeping/mgmt_gpio_oeb[4] housekeeping/mgmt_gpio_oeb[5]
+ housekeeping/mgmt_gpio_oeb[6] housekeeping/mgmt_gpio_oeb[7] housekeeping/mgmt_gpio_oeb[8]
+ housekeeping/mgmt_gpio_oeb[9] housekeeping/mgmt_gpio_out[0] housekeeping/mgmt_gpio_in[10]
+ housekeeping/mgmt_gpio_in[11] housekeeping/mgmt_gpio_in[12] housekeeping/mgmt_gpio_in[13]
+ housekeeping/mgmt_gpio_in[14] housekeeping/mgmt_gpio_in[15] housekeeping/mgmt_gpio_in[16]
+ housekeeping/mgmt_gpio_in[17] housekeeping/mgmt_gpio_in[18] housekeeping/mgmt_gpio_in[19]
+ housekeeping/mgmt_gpio_out[1] housekeeping/mgmt_gpio_in[20] housekeeping/mgmt_gpio_in[21]
+ housekeeping/mgmt_gpio_in[22] housekeeping/mgmt_gpio_in[23] housekeeping/mgmt_gpio_in[24]
+ housekeeping/mgmt_gpio_in[25] housekeeping/mgmt_gpio_in[26] housekeeping/mgmt_gpio_in[27]
+ housekeeping/mgmt_gpio_in[28] housekeeping/mgmt_gpio_in[29] housekeeping/mgmt_gpio_in[2]
+ housekeeping/mgmt_gpio_in[30] housekeeping/mgmt_gpio_in[31] housekeeping/mgmt_gpio_in[32]
+ housekeeping/mgmt_gpio_in[33] housekeeping/mgmt_gpio_in[34] housekeeping/mgmt_gpio_out[35]
+ housekeeping/mgmt_gpio_out[36] housekeeping/mgmt_gpio_out[37] housekeeping/mgmt_gpio_in[3]
+ housekeeping/mgmt_gpio_in[4] housekeeping/mgmt_gpio_in[5] housekeeping/mgmt_gpio_in[6]
+ housekeeping/mgmt_gpio_in[7] housekeeping/mgmt_gpio_in[8] housekeeping/mgmt_gpio_in[9]
+ padframe/flash_clk_core padframe/flash_clk_oeb_core padframe/flash_csb_core padframe/flash_csb_oeb_core
+ padframe/flash_io0_di_core padframe/flash_io0_do_core padframe/flash_io0_ieb_core
+ padframe/flash_io0_oeb_core padframe/flash_io1_di_core padframe/flash_io1_do_core
+ padframe/flash_io1_ieb_core padframe/flash_io1_oeb_core clocking/sel2[0] clocking/sel2[1]
+ clocking/sel2[2] clocking/ext_clk_sel pll/dco pll/div[0] pll/div[1] pll/div[2] pll/div[3]
+ pll/div[4] pll/enable clocking/sel[0] clocking/sel[1] clocking/sel[2] pll/ext_trim[0]
+ pll/ext_trim[10] pll/ext_trim[11] pll/ext_trim[12] pll/ext_trim[13] pll/ext_trim[14]
+ pll/ext_trim[15] pll/ext_trim[16] pll/ext_trim[17] pll/ext_trim[18] pll/ext_trim[19]
+ pll/ext_trim[1] pll/ext_trim[20] pll/ext_trim[21] pll/ext_trim[22] pll/ext_trim[23]
+ pll/ext_trim[24] pll/ext_trim[25] pll/ext_trim[2] pll/ext_trim[3] pll/ext_trim[4]
+ pll/ext_trim[5] pll/ext_trim[6] pll/ext_trim[7] pll/ext_trim[8] pll/ext_trim[9]
+ por/porb_l housekeeping/pwr_ctrl_out[0] housekeeping/pwr_ctrl_out[1] housekeeping/pwr_ctrl_out[2]
+ housekeeping/pwr_ctrl_out[3] soc/qspi_enabled housekeeping/reset soc/ser_rx soc/ser_tx
+ housekeeping/serial_clock housekeeping/serial_data_1 housekeeping/serial_data_2
+ housekeeping/serial_load housekeeping/serial_resetn soc/spi_csb soc/spi_enabled
+ soc/spi_sck soc/spi_sdi soc/spi_sdo soc/spi_sdoenb soc/flash_clk soc/flash_csb soc/flash_io0_di
+ soc/flash_io0_do soc/flash_io0_oeb soc/flash_io1_di soc/flash_io1_do soc/flash_io1_oeb
+ soc/flash_io2_di soc/flash_io2_do soc/flash_io2_oeb soc/flash_io3_di soc/flash_io3_do
+ soc/flash_io3_oeb soc/sram_ro_addr[0] soc/sram_ro_addr[1] soc/sram_ro_addr[2] soc/sram_ro_addr[3]
+ soc/sram_ro_addr[4] soc/sram_ro_addr[5] soc/sram_ro_addr[6] soc/sram_ro_addr[7]
+ soc/sram_ro_clk soc/sram_ro_csb soc/sram_ro_data[0] soc/sram_ro_data[10] soc/sram_ro_data[11]
+ soc/sram_ro_data[12] soc/sram_ro_data[13] soc/sram_ro_data[14] soc/sram_ro_data[15]
+ soc/sram_ro_data[16] soc/sram_ro_data[17] soc/sram_ro_data[18] soc/sram_ro_data[19]
+ soc/sram_ro_data[1] soc/sram_ro_data[20] soc/sram_ro_data[21] soc/sram_ro_data[22]
+ soc/sram_ro_data[23] soc/sram_ro_data[24] soc/sram_ro_data[25] soc/sram_ro_data[26]
+ soc/sram_ro_data[27] soc/sram_ro_data[28] soc/sram_ro_data[29] soc/sram_ro_data[2]
+ soc/sram_ro_data[30] soc/sram_ro_data[31] soc/sram_ro_data[3] soc/sram_ro_data[4]
+ soc/sram_ro_data[5] soc/sram_ro_data[6] soc/sram_ro_data[7] soc/sram_ro_data[8]
+ soc/sram_ro_data[9] soc/trap soc/uart_enabled clocking/user_clk housekeeping/usr1_vcc_pwrgood
+ housekeeping/usr1_vdd_pwrgood housekeeping/usr2_vcc_pwrgood housekeeping/usr2_vdd_pwrgood
+ soc/hk_ack_i soc/mprj_adr_o[0] soc/mprj_adr_o[10] soc/mprj_adr_o[11] soc/mprj_adr_o[12]
+ soc/mprj_adr_o[13] soc/mprj_adr_o[14] soc/mprj_adr_o[15] soc/mprj_adr_o[16] soc/mprj_adr_o[17]
+ soc/mprj_adr_o[18] soc/mprj_adr_o[19] soc/mprj_adr_o[1] soc/mprj_adr_o[20] soc/mprj_adr_o[21]
+ soc/mprj_adr_o[22] soc/mprj_adr_o[23] soc/mprj_adr_o[24] soc/mprj_adr_o[25] soc/mprj_adr_o[26]
+ soc/mprj_adr_o[27] soc/mprj_adr_o[28] soc/mprj_adr_o[29] soc/mprj_adr_o[2] soc/mprj_adr_o[30]
+ soc/mprj_adr_o[31] soc/mprj_adr_o[3] soc/mprj_adr_o[4] soc/mprj_adr_o[5] soc/mprj_adr_o[6]
+ soc/mprj_adr_o[7] soc/mprj_adr_o[8] soc/mprj_adr_o[9] soc/core_clk soc/hk_cyc_o
+ soc/mprj_dat_o[0] soc/mprj_dat_o[10] soc/mprj_dat_o[11] soc/mprj_dat_o[12] soc/mprj_dat_o[13]
+ soc/mprj_dat_o[14] soc/mprj_dat_o[15] soc/mprj_dat_o[16] soc/mprj_dat_o[17] soc/mprj_dat_o[18]
+ soc/mprj_dat_o[19] soc/mprj_dat_o[1] soc/mprj_dat_o[20] soc/mprj_dat_o[21] soc/mprj_dat_o[22]
+ soc/mprj_dat_o[23] soc/mprj_dat_o[24] soc/mprj_dat_o[25] soc/mprj_dat_o[26] soc/mprj_dat_o[27]
+ soc/mprj_dat_o[28] soc/mprj_dat_o[29] soc/mprj_dat_o[2] soc/mprj_dat_o[30] soc/mprj_dat_o[31]
+ soc/mprj_dat_o[3] soc/mprj_dat_o[4] soc/mprj_dat_o[5] soc/mprj_dat_o[6] soc/mprj_dat_o[7]
+ soc/mprj_dat_o[8] soc/mprj_dat_o[9] soc/hk_dat_i[0] soc/hk_dat_i[10] soc/hk_dat_i[11]
+ soc/hk_dat_i[12] soc/hk_dat_i[13] soc/hk_dat_i[14] soc/hk_dat_i[15] soc/hk_dat_i[16]
+ soc/hk_dat_i[17] soc/hk_dat_i[18] soc/hk_dat_i[19] soc/hk_dat_i[1] soc/hk_dat_i[20]
+ soc/hk_dat_i[21] soc/hk_dat_i[22] soc/hk_dat_i[23] soc/hk_dat_i[24] soc/hk_dat_i[25]
+ soc/hk_dat_i[26] soc/hk_dat_i[27] soc/hk_dat_i[28] soc/hk_dat_i[29] soc/hk_dat_i[2]
+ soc/hk_dat_i[30] soc/hk_dat_i[31] soc/hk_dat_i[3] soc/hk_dat_i[4] soc/hk_dat_i[5]
+ soc/hk_dat_i[6] soc/hk_dat_i[7] soc/hk_dat_i[8] soc/hk_dat_i[9] soc/core_rstn soc/mprj_sel_o[0]
+ soc/mprj_sel_o[1] soc/mprj_sel_o[2] soc/mprj_sel_o[3] soc/hk_stb_o soc/mprj_we_o
+ VSUBS vccd_core housekeeping
Xgpio_control_in_2\[2\] gpio_defaults_block_21/gpio_defaults[0] gpio_defaults_block_21/gpio_defaults[10]
+ gpio_defaults_block_21/gpio_defaults[11] gpio_defaults_block_21/gpio_defaults[12]
+ gpio_defaults_block_21/gpio_defaults[1] gpio_defaults_block_21/gpio_defaults[2]
+ gpio_defaults_block_21/gpio_defaults[3] gpio_defaults_block_21/gpio_defaults[4]
+ gpio_defaults_block_21/gpio_defaults[5] gpio_defaults_block_21/gpio_defaults[6]
+ gpio_defaults_block_21/gpio_defaults[7] gpio_defaults_block_21/gpio_defaults[8]
+ gpio_defaults_block_21/gpio_defaults[9] housekeeping/mgmt_gpio_in[21] gpio_control_in_2\[2\]/one
+ housekeeping/mgmt_gpio_in[21] gpio_control_in_2\[2\]/one padframe/mprj_io_analog_en[21]
+ padframe/mprj_io_analog_pol[21] padframe/mprj_io_analog_sel[21] padframe/mprj_io_dm[63]
+ padframe/mprj_io_dm[64] padframe/mprj_io_dm[65] padframe/mprj_io_holdover[21] padframe/mprj_io_ib_mode_sel[21]
+ padframe/mprj_io_in[21] padframe/mprj_io_inp_dis[21] padframe/mprj_io_out[21] padframe/mprj_io_oeb[21]
+ padframe/mprj_io_slow_sel[21] padframe/mprj_io_vtrip_sel[21] gpio_control_in_2\[2\]/resetn
+ gpio_control_in_2\[1\]/resetn gpio_control_in_2\[2\]/serial_clock gpio_control_in_2\[1\]/serial_clock
+ gpio_control_in_2\[2\]/serial_data_in gpio_control_in_2\[1\]/serial_data_in gpio_control_in_2\[2\]/serial_load
+ gpio_control_in_2\[1\]/serial_load mprj/io_in[21] mprj/io_oeb[21] mprj/io_out[21]
+ vccd1_core VSUBS gpio_control_in_2\[2\]/zero dw_201538_1027427# vccd_core vssd1_core
+ gpio_control_block
Xgpio_control_in_1\[8\] gpio_defaults_block_16/gpio_defaults[0] gpio_defaults_block_16/gpio_defaults[10]
+ gpio_defaults_block_16/gpio_defaults[11] gpio_defaults_block_16/gpio_defaults[12]
+ gpio_defaults_block_16/gpio_defaults[1] gpio_defaults_block_16/gpio_defaults[2]
+ gpio_defaults_block_16/gpio_defaults[3] gpio_defaults_block_16/gpio_defaults[4]
+ gpio_defaults_block_16/gpio_defaults[5] gpio_defaults_block_16/gpio_defaults[6]
+ gpio_defaults_block_16/gpio_defaults[7] gpio_defaults_block_16/gpio_defaults[8]
+ gpio_defaults_block_16/gpio_defaults[9] housekeeping/mgmt_gpio_in[16] gpio_control_in_1\[8\]/one
+ housekeeping/mgmt_gpio_in[16] gpio_control_in_1\[8\]/one padframe/mprj_io_analog_en[16]
+ padframe/mprj_io_analog_pol[16] padframe/mprj_io_analog_sel[16] padframe/mprj_io_dm[48]
+ padframe/mprj_io_dm[49] padframe/mprj_io_dm[50] padframe/mprj_io_holdover[16] padframe/mprj_io_ib_mode_sel[16]
+ padframe/mprj_io_in[16] padframe/mprj_io_inp_dis[16] padframe/mprj_io_out[16] padframe/mprj_io_oeb[16]
+ padframe/mprj_io_slow_sel[16] padframe/mprj_io_vtrip_sel[16] gpio_control_in_1\[8\]/resetn
+ gpio_control_in_1\[9\]/resetn gpio_control_in_1\[8\]/serial_clock gpio_control_in_1\[9\]/serial_clock
+ gpio_control_in_1\[8\]/serial_data_in gpio_control_in_1\[9\]/serial_data_in gpio_control_in_1\[8\]/serial_load
+ gpio_control_in_1\[9\]/serial_load mprj/io_in[16] mprj/io_oeb[16] mprj/io_out[16]
+ vccd1_core VSUBS gpio_control_in_1\[8\]/zero dw_499338_1027427# vccd_core vssd1_core
+ gpio_control_block
Xgpio_defaults_block_30 VSUBS gpio_defaults_block_30/gpio_defaults[0] gpio_defaults_block_30/gpio_defaults[10]
+ gpio_defaults_block_30/gpio_defaults[11] gpio_defaults_block_30/gpio_defaults[12]
+ gpio_defaults_block_30/gpio_defaults[1] gpio_defaults_block_30/gpio_defaults[2]
+ gpio_defaults_block_30/gpio_defaults[3] gpio_defaults_block_30/gpio_defaults[4]
+ gpio_defaults_block_30/gpio_defaults[5] gpio_defaults_block_30/gpio_defaults[6]
+ gpio_defaults_block_30/gpio_defaults[7] gpio_defaults_block_30/gpio_defaults[8]
+ gpio_defaults_block_30/gpio_defaults[9] vccd_core gpio_defaults_block
Xgpio_defaults_block_20 VSUBS gpio_defaults_block_20/gpio_defaults[0] gpio_defaults_block_20/gpio_defaults[10]
+ gpio_defaults_block_20/gpio_defaults[11] gpio_defaults_block_20/gpio_defaults[12]
+ gpio_defaults_block_20/gpio_defaults[1] gpio_defaults_block_20/gpio_defaults[2]
+ gpio_defaults_block_20/gpio_defaults[3] gpio_defaults_block_20/gpio_defaults[4]
+ gpio_defaults_block_20/gpio_defaults[5] gpio_defaults_block_20/gpio_defaults[6]
+ gpio_defaults_block_20/gpio_defaults[7] gpio_defaults_block_20/gpio_defaults[8]
+ gpio_defaults_block_20/gpio_defaults[9] vccd_core gpio_defaults_block
Xgpio_defaults_block_21 VSUBS gpio_defaults_block_21/gpio_defaults[0] gpio_defaults_block_21/gpio_defaults[10]
+ gpio_defaults_block_21/gpio_defaults[11] gpio_defaults_block_21/gpio_defaults[12]
+ gpio_defaults_block_21/gpio_defaults[1] gpio_defaults_block_21/gpio_defaults[2]
+ gpio_defaults_block_21/gpio_defaults[3] gpio_defaults_block_21/gpio_defaults[4]
+ gpio_defaults_block_21/gpio_defaults[5] gpio_defaults_block_21/gpio_defaults[6]
+ gpio_defaults_block_21/gpio_defaults[7] gpio_defaults_block_21/gpio_defaults[8]
+ gpio_defaults_block_21/gpio_defaults[9] vccd_core gpio_defaults_block
Xgpio_defaults_block_10 VSUBS gpio_defaults_block_10/gpio_defaults[0] gpio_defaults_block_10/gpio_defaults[10]
+ gpio_defaults_block_10/gpio_defaults[11] gpio_defaults_block_10/gpio_defaults[12]
+ gpio_defaults_block_10/gpio_defaults[1] gpio_defaults_block_10/gpio_defaults[2]
+ gpio_defaults_block_10/gpio_defaults[3] gpio_defaults_block_10/gpio_defaults[4]
+ gpio_defaults_block_10/gpio_defaults[5] gpio_defaults_block_10/gpio_defaults[6]
+ gpio_defaults_block_10/gpio_defaults[7] gpio_defaults_block_10/gpio_defaults[8]
+ gpio_defaults_block_10/gpio_defaults[9] vccd_core gpio_defaults_block
Xgpio_defaults_block_31 VSUBS gpio_defaults_block_31/gpio_defaults[0] gpio_defaults_block_31/gpio_defaults[10]
+ gpio_defaults_block_31/gpio_defaults[11] gpio_defaults_block_31/gpio_defaults[12]
+ gpio_defaults_block_31/gpio_defaults[1] gpio_defaults_block_31/gpio_defaults[2]
+ gpio_defaults_block_31/gpio_defaults[3] gpio_defaults_block_31/gpio_defaults[4]
+ gpio_defaults_block_31/gpio_defaults[5] gpio_defaults_block_31/gpio_defaults[6]
+ gpio_defaults_block_31/gpio_defaults[7] gpio_defaults_block_31/gpio_defaults[8]
+ gpio_defaults_block_31/gpio_defaults[9] vccd_core gpio_defaults_block
Xgpio_control_in_1a\[5\] gpio_defaults_block_7/gpio_defaults[0] gpio_defaults_block_7/gpio_defaults[10]
+ gpio_defaults_block_7/gpio_defaults[11] gpio_defaults_block_7/gpio_defaults[12]
+ gpio_defaults_block_7/gpio_defaults[1] gpio_defaults_block_7/gpio_defaults[2] gpio_defaults_block_7/gpio_defaults[3]
+ gpio_defaults_block_7/gpio_defaults[4] gpio_defaults_block_7/gpio_defaults[5] gpio_defaults_block_7/gpio_defaults[6]
+ gpio_defaults_block_7/gpio_defaults[7] gpio_defaults_block_7/gpio_defaults[8] gpio_defaults_block_7/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[7] gpio_control_in_1a\[5\]/one housekeeping/mgmt_gpio_in[7]
+ gpio_control_in_1a\[5\]/one padframe/mprj_io_analog_en[7] padframe/mprj_io_analog_pol[7]
+ padframe/mprj_io_analog_sel[7] padframe/mprj_io_dm[21] padframe/mprj_io_dm[22] padframe/mprj_io_dm[23]
+ padframe/mprj_io_holdover[7] padframe/mprj_io_ib_mode_sel[7] padframe/mprj_io_in[7]
+ padframe/mprj_io_inp_dis[7] padframe/mprj_io_out[7] padframe/mprj_io_oeb[7] padframe/mprj_io_slow_sel[7]
+ padframe/mprj_io_vtrip_sel[7] gpio_control_in_1a\[5\]/resetn gpio_control_in_1\[0\]/resetn
+ gpio_control_in_1a\[5\]/serial_clock gpio_control_in_1\[0\]/serial_clock gpio_control_in_1a\[5\]/serial_data_in
+ gpio_control_in_1\[0\]/serial_data_in gpio_control_in_1a\[5\]/serial_load gpio_control_in_1\[0\]/serial_load
+ mprj/io_in[7] mprj/io_oeb[7] mprj/io_out[7] vccd1_core VSUBS gpio_control_in_1a\[5\]/zero
+ dw_707553_481338# vccd_core vssd1_core gpio_control_block
Xgpio_defaults_block_32 VSUBS gpio_defaults_block_32/gpio_defaults[0] gpio_defaults_block_32/gpio_defaults[10]
+ gpio_defaults_block_32/gpio_defaults[11] gpio_defaults_block_32/gpio_defaults[12]
+ gpio_defaults_block_32/gpio_defaults[1] gpio_defaults_block_32/gpio_defaults[2]
+ gpio_defaults_block_32/gpio_defaults[3] gpio_defaults_block_32/gpio_defaults[4]
+ gpio_defaults_block_32/gpio_defaults[5] gpio_defaults_block_32/gpio_defaults[6]
+ gpio_defaults_block_32/gpio_defaults[7] gpio_defaults_block_32/gpio_defaults[8]
+ gpio_defaults_block_32/gpio_defaults[9] vccd_core gpio_defaults_block
Xgpio_control_bidir_2\[2\] gpio_defaults_block_37/gpio_defaults[0] gpio_defaults_block_37/gpio_defaults[10]
+ gpio_defaults_block_37/gpio_defaults[11] gpio_defaults_block_37/gpio_defaults[12]
+ gpio_defaults_block_37/gpio_defaults[1] gpio_defaults_block_37/gpio_defaults[2]
+ gpio_defaults_block_37/gpio_defaults[3] gpio_defaults_block_37/gpio_defaults[4]
+ gpio_defaults_block_37/gpio_defaults[5] gpio_defaults_block_37/gpio_defaults[6]
+ gpio_defaults_block_37/gpio_defaults[7] gpio_defaults_block_37/gpio_defaults[8]
+ gpio_defaults_block_37/gpio_defaults[9] housekeeping/mgmt_gpio_in[37] housekeeping/mgmt_gpio_oeb[37]
+ housekeeping/mgmt_gpio_out[37] gpio_control_bidir_2\[2\]/one padframe/mprj_io_analog_en[37]
+ padframe/mprj_io_analog_pol[37] padframe/mprj_io_analog_sel[37] padframe/mprj_io_dm[111]
+ padframe/mprj_io_dm[112] padframe/mprj_io_dm[113] padframe/mprj_io_holdover[37]
+ padframe/mprj_io_ib_mode_sel[37] padframe/mprj_io_in[37] padframe/mprj_io_inp_dis[37]
+ padframe/mprj_io_out[37] padframe/mprj_io_oeb[37] padframe/mprj_io_slow_sel[37]
+ padframe/mprj_io_vtrip_sel[37] housekeeping/serial_resetn gpio_control_bidir_2\[1\]/resetn
+ housekeeping/serial_clock gpio_control_bidir_2\[1\]/serial_clock housekeeping/serial_data_2
+ gpio_control_bidir_2\[1\]/serial_data_in housekeeping/serial_load gpio_control_bidir_2\[1\]/serial_load
+ mprj/io_in[37] mprj/io_oeb[37] mprj/io_out[37] vccd1_core VSUBS gpio_control_bidir_2\[2\]/zero
+ dw_8741_204138# vccd_core vssd1_core gpio_control_block
.ends

