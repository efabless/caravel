* NGSPICE file created from caravan.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__dfbbn_1 abstract view
.subckt sky130_fd_sc_hd__dfbbn_1 CLK_N D RESET_B SET_B VGND VNB VPB VPWR Q Q_N
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1#0 abstract view
.subckt sky130_fd_sc_hd__fill_1#0 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2#0 abstract view
.subckt sky130_fd_sc_hd__fill_2#0 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12#0 abstract view
.subckt sky130_fd_sc_hd__decap_12#0 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3#0 abstract view
.subckt sky130_fd_sc_hd__decap_3#0 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1#0 abstract view
.subckt sky130_fd_sc_hd__conb_1#0 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__einvp_2 abstract view
.subckt sky130_fd_sc_hd__einvp_2 A TE VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6#0 abstract view
.subckt sky130_fd_sc_hd__decap_6#0 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1#0 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1#0 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_1 abstract view
.subckt sky130_fd_sc_hd__ebufn_1 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

.subckt sky130_fd_sc_hd__decap_6 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
.ends

.subckt sky130_fd_sc_hd__decap_8 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
.ends

.subckt sky130_fd_sc_hd__decap_3 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
.ends

.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
R0 HI VPWR sky130_fd_pr__res_generic_po w=480000u l=45000u
R1 VGND LO sky130_fd_pr__res_generic_po w=480000u l=45000u
.ends

.subckt gpio_logic_high gpio_logic1 vccd1 vssd1
XFILLER_3_3 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_3 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_0 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_5 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_6 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_7 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_8 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_9 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_3 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_3 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_4
Xgpio_logic_high vssd1 vssd1 vccd1 vccd1 gpio_logic1 gpio_logic_high/LO sky130_fd_sc_hd__conb_1
XFILLER_4_9 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_9 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8#0 abstract view
.subckt sky130_fd_sc_hd__decap_8#0 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for gpio_control_block abstract view
.subckt gpio_control_block gpio_defaults[0] gpio_defaults[10] gpio_defaults[11] gpio_defaults[12]
+ gpio_defaults[1] gpio_defaults[2] gpio_defaults[3] gpio_defaults[4] gpio_defaults[5]
+ gpio_defaults[6] gpio_defaults[7] gpio_defaults[8] gpio_defaults[9] mgmt_gpio_in
+ mgmt_gpio_oeb mgmt_gpio_out one pad_gpio_ana_en pad_gpio_ana_pol pad_gpio_ana_sel
+ pad_gpio_dm[0] pad_gpio_dm[1] pad_gpio_dm[2] pad_gpio_holdover pad_gpio_ib_mode_sel
+ pad_gpio_in pad_gpio_inenb pad_gpio_out pad_gpio_outenb pad_gpio_slow_sel pad_gpio_vtrip_sel
+ resetn resetn_out serial_clock serial_clock_out serial_data_in serial_data_out serial_load
+ serial_load_out user_gpio_in user_gpio_oeb user_gpio_out vccd vccd1 vssd vssd1 zero
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4#0 abstract view
.subckt sky130_fd_sc_hd__decap_4#0 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for gpio_defaults_block abstract view
.subckt gpio_defaults_block VGND VPWR gpio_defaults[0] gpio_defaults[10] gpio_defaults[11]
+ gpio_defaults[12] gpio_defaults[1] gpio_defaults[2] gpio_defaults[3] gpio_defaults[4]
+ gpio_defaults[5] gpio_defaults[6] gpio_defaults[7] gpio_defaults[8] gpio_defaults[9]
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_1 abstract view
.subckt sky130_fd_sc_hd__clkinv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__einvn_8 abstract view
.subckt sky130_fd_sc_hd__einvn_8 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__einvn_4 abstract view
.subckt sky130_fd_sc_hd__einvn_4 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__einvp_1 abstract view
.subckt sky130_fd_sc_hd__einvp_1 A TE VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for digital_pll abstract view
.subckt digital_pll VGND VPWR clockp[0] clockp[1] dco div[0] div[1] div[2] div[3]
+ div[4] enable ext_trim[0] ext_trim[10] ext_trim[11] ext_trim[12] ext_trim[13] ext_trim[14]
+ ext_trim[15] ext_trim[16] ext_trim[17] ext_trim[18] ext_trim[19] ext_trim[1] ext_trim[20]
+ ext_trim[21] ext_trim[22] ext_trim[23] ext_trim[24] ext_trim[25] ext_trim[2] ext_trim[3]
+ ext_trim[4] ext_trim[5] ext_trim[6] ext_trim[7] ext_trim[8] ext_trim[9] osc resetb
.ends

* Black-box entry subcircuit for sky130_ef_io__com_bus_slice_20um abstract view
.subckt sky130_ef_io__com_bus_slice_20um AMUXBUS_A AMUXBUS_B VSSA VDDA VSWITCH VDDIO_Q
+ VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
.ends

* Black-box entry subcircuit for sky130_ef_io__gpiov2_pad_wrapped abstract view
.subckt sky130_ef_io__gpiov2_pad_wrapped IN_H PAD_A_NOESD_H PAD_A_ESD_0_H PAD_A_ESD_1_H
+ PAD DM[2] DM[1] DM[0] HLD_H_N IN INP_DIS IB_MODE_SEL ENABLE_H ENABLE_VDDA_H ENABLE_INP_H
+ OE_N TIE_HI_ESD TIE_LO_ESD SLOW VTRIP_SEL HLD_OVR ANALOG_EN ANALOG_SEL ENABLE_VDDIO
+ ENABLE_VSWITCH_H ANALOG_POL OUT AMUXBUS_A AMUXBUS_B VSSA VDDA VSWITCH VDDIO_Q VCCHIB
+ VDDIO VCCD VSSIO VSSD VSSIO_Q
.ends

* Black-box entry subcircuit for sky130_ef_io__com_bus_slice_1um abstract view
.subckt sky130_ef_io__com_bus_slice_1um AMUXBUS_A AMUXBUS_B VSSA VDDA VSWITCH VDDIO_Q
+ VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
.ends

* Black-box entry subcircuit for sky130_ef_io__com_bus_slice_10um abstract view
.subckt sky130_ef_io__com_bus_slice_10um AMUXBUS_A AMUXBUS_B VSSA VDDA VSWITCH VDDIO_Q
+ VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
.ends

* Black-box entry subcircuit for sky130_ef_io__vccd_lvc_clamped_pad abstract view
.subckt sky130_ef_io__vccd_lvc_clamped_pad AMUXBUS_A AMUXBUS_B VCCD_PAD VSSA VDDA
+ VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
.ends

* Black-box entry subcircuit for sky130_ef_io__com_bus_slice_5um abstract view
.subckt sky130_ef_io__com_bus_slice_5um AMUXBUS_A AMUXBUS_B VSSA VDDA VSWITCH VDDIO_Q
+ VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
.ends

* Black-box entry subcircuit for sky130_ef_io__analog_pad abstract view
.subckt sky130_ef_io__analog_pad P_CORE VSSA VSSD AMUXBUS_B AMUXBUS_A VDDIO_Q VDDIO
+ VSWITCH VSSIO VDDA VCCD VCCHIB VSSIO_Q P_PAD
.ends

* Black-box entry subcircuit for sky130_ef_io__disconnect_vdda_slice_5um abstract view
.subckt sky130_ef_io__disconnect_vdda_slice_5um AMUXBUS_A AMUXBUS_B VSWITCH VDDIO_Q
+ VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
.ends

* Black-box entry subcircuit for sky130_ef_io__corner_pad abstract view
.subckt sky130_ef_io__corner_pad AMUXBUS_A AMUXBUS_B VSSA VDDA VSWITCH VDDIO_Q VCCHIB
+ VDDIO VCCD VSSIO VSSD VSSIO_Q
.ends

* Black-box entry subcircuit for sky130_ef_io__vddio_hvc_clamped_pad abstract view
.subckt sky130_ef_io__vddio_hvc_clamped_pad AMUXBUS_A AMUXBUS_B VDDIO_PAD VSSA VDDA
+ VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
.ends

* Black-box entry subcircuit for sky130_ef_io__vssio_hvc_clamped_pad abstract view
.subckt sky130_ef_io__vssio_hvc_clamped_pad AMUXBUS_A AMUXBUS_B VSSIO_PAD VSSA VDDA
+ VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
.ends

* Black-box entry subcircuit for sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um abstract view
.subckt sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um AMUXBUS_A AMUXBUS_B
+ VSSA VDDA VDDIO_Q VDDIO VCCD VSSIO VSSD VSSIO_Q VSWITCH VCCHIB
.ends

* Black-box entry subcircuit for sky130_ef_io__vdda_hvc_clamped_pad abstract view
.subckt sky130_ef_io__vdda_hvc_clamped_pad AMUXBUS_A AMUXBUS_B VDDA_PAD VSSA VDDA
+ VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
.ends

* Black-box entry subcircuit for sky130_ef_io__top_power_hvc abstract view
.subckt sky130_ef_io__top_power_hvc AMUXBUS_A AMUXBUS_B DRN_HVC P_CORE P_PAD SRC_BDY_HVC
+ VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
.ends

* Black-box entry subcircuit for sky130_ef_io__vssd_lvc_clamped3_pad abstract view
.subckt sky130_ef_io__vssd_lvc_clamped3_pad AMUXBUS_A AMUXBUS_B VSSD_PAD VSSA VDDA
+ VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q VCCD1 VSSD1
.ends

* Black-box entry subcircuit for sky130_ef_io__vssd_lvc_clamped_pad abstract view
.subckt sky130_ef_io__vssd_lvc_clamped_pad AMUXBUS_A AMUXBUS_B VSSD_PAD VSSA VDDA
+ VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
.ends

* Black-box entry subcircuit for sky130_ef_io__vccd_lvc_clamped3_pad abstract view
.subckt sky130_ef_io__vccd_lvc_clamped3_pad AMUXBUS_A AMUXBUS_B VCCD_PAD VSSA VDDA
+ VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q VCCD1 VSSD1
.ends

* Black-box entry subcircuit for sky130_ef_io__vssa_hvc_clamped_pad abstract view
.subckt sky130_ef_io__vssa_hvc_clamped_pad AMUXBUS_A AMUXBUS_B VSSA_PAD VSSA VDDA
+ VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
.ends

* Black-box entry subcircuit for sky130_fd_io__top_xres4v2 abstract view
.subckt sky130_fd_io__top_xres4v2 PAD_A_ESD_H XRES_H_N FILT_IN_H ENABLE_VDDIO TIE_WEAK_HI_H
+ ENABLE_H PULLUP_H EN_VDDIO_SIG_H TIE_LO_ESD TIE_HI_ESD DISABLE_PULLUP_H INP_SEL_H
+ VSSIO VSSA VSSD AMUXBUS_B AMUXBUS_A VDDIO_Q VDDIO VSWITCH VDDA VCCD VCCHIB VSSIO_Q
+ PAD
.ends

* Black-box entry subcircuit for chip_io_alt abstract view
.subckt chip_io_alt clock clock_core por flash_clk flash_csb flash_io0 flash_io0_di_core
+ flash_io0_do_core flash_io0_ieb_core flash_io0_oeb_core flash_io1 flash_io1_di_core
+ flash_io1_do_core flash_io1_ieb_core flash_io1_oeb_core gpio gpio_in_core gpio_inenb_core
+ gpio_mode0_core gpio_mode1_core gpio_out_core gpio_outenb_core vccd_pad vdda_pad
+ vddio_pad vddio_pad2 vssa_pad vssd_pad vssio_pad vssio_pad2 mprj_io[0] mprj_io_analog_en[0]
+ mprj_io_analog_pol[0] mprj_io_analog_sel[0] mprj_io_dm[0] mprj_io_dm[1] mprj_io_dm[2]
+ mprj_io_holdover[0] mprj_io_ib_mode_sel[0] mprj_io_inp_dis[0] mprj_io_oeb[0] mprj_io_out[0]
+ mprj_io_slow_sel[0] mprj_io_vtrip_sel[0] mprj_io_in[0] mprj_io_in_3v3[0] mprj_gpio_analog[3]
+ mprj_gpio_noesd[3] mprj_io[10] mprj_io_analog_en[10] mprj_io_analog_pol[10] mprj_io_analog_sel[10]
+ mprj_io_dm[30] mprj_io_dm[31] mprj_io_dm[32] mprj_io_holdover[10] mprj_io_ib_mode_sel[10]
+ mprj_io_inp_dis[10] mprj_io_oeb[10] mprj_io_out[10] mprj_io_slow_sel[10] mprj_io_vtrip_sel[10]
+ mprj_io_in[10] mprj_io_in_3v3[10] mprj_gpio_analog[4] mprj_gpio_noesd[4] mprj_io[11]
+ mprj_io_analog_en[11] mprj_io_analog_pol[11] mprj_io_analog_sel[11] mprj_io_dm[33]
+ mprj_io_dm[34] mprj_io_dm[35] mprj_io_holdover[11] mprj_io_ib_mode_sel[11] mprj_io_inp_dis[11]
+ mprj_io_oeb[11] mprj_io_out[11] mprj_io_slow_sel[11] mprj_io_vtrip_sel[11] mprj_io_in[11]
+ mprj_io_in_3v3[11] mprj_gpio_analog[5] mprj_gpio_noesd[5] mprj_io[12] mprj_io_analog_en[12]
+ mprj_io_analog_pol[12] mprj_io_analog_sel[12] mprj_io_dm[36] mprj_io_dm[37] mprj_io_dm[38]
+ mprj_io_holdover[12] mprj_io_ib_mode_sel[12] mprj_io_inp_dis[12] mprj_io_oeb[12]
+ mprj_io_out[12] mprj_io_slow_sel[12] mprj_io_vtrip_sel[12] mprj_io_in[12] mprj_io_in_3v3[12]
+ mprj_gpio_analog[6] mprj_gpio_noesd[6] mprj_io[13] mprj_io_analog_en[13] mprj_io_analog_pol[13]
+ mprj_io_analog_sel[13] mprj_io_dm[39] mprj_io_dm[40] mprj_io_dm[41] mprj_io_holdover[13]
+ mprj_io_ib_mode_sel[13] mprj_io_inp_dis[13] mprj_io_oeb[13] mprj_io_out[13] mprj_io_slow_sel[13]
+ mprj_io_vtrip_sel[13] mprj_io_in[13] mprj_io_in_3v3[13] mprj_io[1] mprj_io_analog_en[1]
+ mprj_io_analog_pol[1] mprj_io_analog_sel[1] mprj_io_dm[3] mprj_io_dm[4] mprj_io_dm[5]
+ mprj_io_holdover[1] mprj_io_ib_mode_sel[1] mprj_io_inp_dis[1] mprj_io_oeb[1] mprj_io_out[1]
+ mprj_io_slow_sel[1] mprj_io_vtrip_sel[1] mprj_io_in[1] mprj_io_in_3v3[1] mprj_io[2]
+ mprj_io_analog_en[2] mprj_io_analog_pol[2] mprj_io_analog_sel[2] mprj_io_dm[6] mprj_io_dm[7]
+ mprj_io_dm[8] mprj_io_holdover[2] mprj_io_ib_mode_sel[2] mprj_io_inp_dis[2] mprj_io_oeb[2]
+ mprj_io_out[2] mprj_io_slow_sel[2] mprj_io_vtrip_sel[2] mprj_io_in[2] mprj_io_in_3v3[2]
+ mprj_io[3] mprj_io_analog_en[3] mprj_io_analog_pol[3] mprj_io_analog_sel[3] mprj_io_dm[10]
+ mprj_io_dm[11] mprj_io_dm[9] mprj_io_holdover[3] mprj_io_ib_mode_sel[3] mprj_io_inp_dis[3]
+ mprj_io_oeb[3] mprj_io_out[3] mprj_io_slow_sel[3] mprj_io_vtrip_sel[3] mprj_io_in[3]
+ mprj_io_in_3v3[3] mprj_io[4] mprj_io_analog_en[4] mprj_io_analog_pol[4] mprj_io_analog_sel[4]
+ mprj_io_dm[12] mprj_io_dm[13] mprj_io_dm[14] mprj_io_holdover[4] mprj_io_ib_mode_sel[4]
+ mprj_io_inp_dis[4] mprj_io_oeb[4] mprj_io_out[4] mprj_io_slow_sel[4] mprj_io_vtrip_sel[4]
+ mprj_io_in[4] mprj_io_in_3v3[4] mprj_io[5] mprj_io_analog_en[5] mprj_io_analog_pol[5]
+ mprj_io_analog_sel[5] mprj_io_dm[15] mprj_io_dm[16] mprj_io_dm[17] mprj_io_holdover[5]
+ mprj_io_ib_mode_sel[5] mprj_io_inp_dis[5] mprj_io_oeb[5] mprj_io_out[5] mprj_io_slow_sel[5]
+ mprj_io_vtrip_sel[5] mprj_io_in[5] mprj_io_in_3v3[5] mprj_io[6] mprj_io_analog_en[6]
+ mprj_io_analog_pol[6] mprj_io_analog_sel[6] mprj_io_dm[18] mprj_io_dm[19] mprj_io_dm[20]
+ mprj_io_holdover[6] mprj_io_ib_mode_sel[6] mprj_io_inp_dis[6] mprj_io_oeb[6] mprj_io_out[6]
+ mprj_io_slow_sel[6] mprj_io_vtrip_sel[6] mprj_io_in[6] mprj_io_in_3v3[6] mprj_gpio_analog[0]
+ mprj_gpio_noesd[0] mprj_io[7] mprj_io_analog_en[7] mprj_io_analog_pol[7] mprj_io_analog_sel[7]
+ mprj_io_dm[21] mprj_io_dm[22] mprj_io_dm[23] mprj_io_holdover[7] mprj_io_ib_mode_sel[7]
+ mprj_io_inp_dis[7] mprj_io_oeb[7] mprj_io_out[7] mprj_io_slow_sel[7] mprj_io_vtrip_sel[7]
+ mprj_io_in[7] mprj_io_in_3v3[7] mprj_gpio_analog[1] mprj_gpio_noesd[1] mprj_io[8]
+ mprj_io_analog_en[8] mprj_io_analog_pol[8] mprj_io_analog_sel[8] mprj_io_dm[24]
+ mprj_io_dm[25] mprj_io_dm[26] mprj_io_holdover[8] mprj_io_ib_mode_sel[8] mprj_io_inp_dis[8]
+ mprj_io_oeb[8] mprj_io_out[8] mprj_io_slow_sel[8] mprj_io_vtrip_sel[8] mprj_io_in[8]
+ mprj_io_in_3v3[8] mprj_gpio_analog[2] mprj_gpio_noesd[2] mprj_io[9] mprj_io_analog_en[9]
+ mprj_io_analog_pol[9] mprj_io_analog_sel[9] mprj_io_dm[27] mprj_io_dm[28] mprj_io_dm[29]
+ mprj_io_holdover[9] mprj_io_ib_mode_sel[9] mprj_io_inp_dis[9] mprj_io_oeb[9] mprj_io_out[9]
+ mprj_io_slow_sel[9] mprj_io_vtrip_sel[9] mprj_io_in[9] mprj_io_in_3v3[9] mprj_gpio_analog[7]
+ mprj_gpio_noesd[7] mprj_io[25] mprj_io_analog_en[14] mprj_io_analog_pol[14] mprj_io_analog_sel[14]
+ mprj_io_dm[42] mprj_io_dm[43] mprj_io_dm[44] mprj_io_holdover[14] mprj_io_ib_mode_sel[14]
+ mprj_io_inp_dis[14] mprj_io_oeb[14] mprj_io_out[14] mprj_io_slow_sel[14] mprj_io_vtrip_sel[14]
+ mprj_io_in[14] mprj_io_in_3v3[14] mprj_gpio_analog[17] mprj_gpio_noesd[17] mprj_io[35]
+ mprj_io_analog_en[24] mprj_io_analog_pol[24] mprj_io_analog_sel[24] mprj_io_dm[72]
+ mprj_io_dm[73] mprj_io_dm[74] mprj_io_holdover[24] mprj_io_ib_mode_sel[24] mprj_io_inp_dis[24]
+ mprj_io_oeb[24] mprj_io_out[24] mprj_io_slow_sel[24] mprj_io_vtrip_sel[24] mprj_io_in[24]
+ mprj_io_in_3v3[24] mprj_io[36] mprj_io_analog_en[25] mprj_io_analog_pol[25] mprj_io_analog_sel[25]
+ mprj_io_dm[75] mprj_io_dm[76] mprj_io_dm[77] mprj_io_holdover[25] mprj_io_ib_mode_sel[25]
+ mprj_io_inp_dis[25] mprj_io_oeb[25] mprj_io_out[25] mprj_io_slow_sel[25] mprj_io_vtrip_sel[25]
+ mprj_io_in[25] mprj_io_in_3v3[25] mprj_io[37] mprj_io_analog_en[26] mprj_io_analog_pol[26]
+ mprj_io_analog_sel[26] mprj_io_dm[78] mprj_io_dm[79] mprj_io_dm[80] mprj_io_holdover[26]
+ mprj_io_ib_mode_sel[26] mprj_io_inp_dis[26] mprj_io_oeb[26] mprj_io_out[26] mprj_io_slow_sel[26]
+ mprj_io_vtrip_sel[26] mprj_io_in[26] mprj_io_in_3v3[26] mprj_gpio_analog[8] mprj_gpio_noesd[8]
+ mprj_io[26] mprj_io_analog_en[15] mprj_io_analog_pol[15] mprj_io_analog_sel[15]
+ mprj_io_dm[45] mprj_io_dm[46] mprj_io_dm[47] mprj_io_holdover[15] mprj_io_ib_mode_sel[15]
+ mprj_io_inp_dis[15] mprj_io_oeb[15] mprj_io_out[15] mprj_io_slow_sel[15] mprj_io_vtrip_sel[15]
+ mprj_io_in[15] mprj_io_in_3v3[15] mprj_gpio_analog[9] mprj_gpio_noesd[9] mprj_io[27]
+ mprj_io_analog_en[16] mprj_io_analog_pol[16] mprj_io_analog_sel[16] mprj_io_dm[48]
+ mprj_io_dm[49] mprj_io_dm[50] mprj_io_holdover[16] mprj_io_ib_mode_sel[16] mprj_io_inp_dis[16]
+ mprj_io_oeb[16] mprj_io_out[16] mprj_io_slow_sel[16] mprj_io_vtrip_sel[16] mprj_io_in[16]
+ mprj_io_in_3v3[16] mprj_gpio_analog[10] mprj_gpio_noesd[10] mprj_io[28] mprj_io_analog_en[17]
+ mprj_io_analog_pol[17] mprj_io_analog_sel[17] mprj_io_dm[51] mprj_io_dm[52] mprj_io_dm[53]
+ mprj_io_holdover[17] mprj_io_ib_mode_sel[17] mprj_io_inp_dis[17] mprj_io_oeb[17]
+ mprj_io_out[17] mprj_io_slow_sel[17] mprj_io_vtrip_sel[17] mprj_io_in[17] mprj_io_in_3v3[17]
+ mprj_gpio_analog[11] mprj_gpio_noesd[11] mprj_io[29] mprj_io_analog_en[18] mprj_io_analog_pol[18]
+ mprj_io_analog_sel[18] mprj_io_dm[54] mprj_io_dm[55] mprj_io_dm[56] mprj_io_holdover[18]
+ mprj_io_ib_mode_sel[18] mprj_io_inp_dis[18] mprj_io_oeb[18] mprj_io_out[18] mprj_io_slow_sel[18]
+ mprj_io_vtrip_sel[18] mprj_io_in[18] mprj_io_in_3v3[18] mprj_gpio_analog[12] mprj_gpio_noesd[12]
+ mprj_io[30] mprj_io_analog_en[19] mprj_io_analog_pol[19] mprj_io_analog_sel[19]
+ mprj_io_dm[57] mprj_io_dm[58] mprj_io_dm[59] mprj_io_holdover[19] mprj_io_ib_mode_sel[19]
+ mprj_io_inp_dis[19] mprj_io_oeb[19] mprj_io_out[19] mprj_io_slow_sel[19] mprj_io_vtrip_sel[19]
+ mprj_io_in[19] mprj_io_in_3v3[19] mprj_gpio_analog[13] mprj_gpio_noesd[13] mprj_io[31]
+ mprj_io_analog_en[20] mprj_io_analog_pol[20] mprj_io_analog_sel[20] mprj_io_dm[60]
+ mprj_io_dm[61] mprj_io_dm[62] mprj_io_holdover[20] mprj_io_ib_mode_sel[20] mprj_io_inp_dis[20]
+ mprj_io_oeb[20] mprj_io_out[20] mprj_io_slow_sel[20] mprj_io_vtrip_sel[20] mprj_io_in[20]
+ mprj_io_in_3v3[20] mprj_gpio_analog[14] mprj_gpio_noesd[14] mprj_io[32] mprj_io_analog_en[21]
+ mprj_io_analog_pol[21] mprj_io_analog_sel[21] mprj_io_dm[63] mprj_io_dm[64] mprj_io_dm[65]
+ mprj_io_holdover[21] mprj_io_ib_mode_sel[21] mprj_io_inp_dis[21] mprj_io_oeb[21]
+ mprj_io_out[21] mprj_io_slow_sel[21] mprj_io_vtrip_sel[21] mprj_io_in[21] mprj_io_in_3v3[21]
+ mprj_gpio_analog[15] mprj_gpio_noesd[15] mprj_io[33] mprj_io_analog_en[22] mprj_io_analog_pol[22]
+ mprj_io_analog_sel[22] mprj_io_dm[66] mprj_io_dm[67] mprj_io_dm[68] mprj_io_holdover[22]
+ mprj_io_ib_mode_sel[22] mprj_io_inp_dis[22] mprj_io_oeb[22] mprj_io_out[22] mprj_io_slow_sel[22]
+ mprj_io_vtrip_sel[22] mprj_io_in[22] mprj_io_in_3v3[22] mprj_gpio_analog[16] mprj_gpio_noesd[16]
+ mprj_io[34] mprj_io_analog_en[23] mprj_io_analog_pol[23] mprj_io_analog_sel[23]
+ mprj_io_dm[69] mprj_io_dm[70] mprj_io_dm[71] mprj_io_holdover[23] mprj_io_ib_mode_sel[23]
+ mprj_io_inp_dis[23] mprj_io_oeb[23] mprj_io_out[23] mprj_io_slow_sel[23] mprj_io_vtrip_sel[23]
+ mprj_io_in[23] mprj_io_in_3v3[23] porb_h resetb resetb_core_h vdda vssa vssd mprj_analog[1]
+ mprj_io[15] mprj_analog[2] mprj_io[16] mprj_analog[3] mprj_io[17] mprj_analog[0]
+ mprj_io[14] mprj_analog[4] mprj_clamp_high[0] mprj_clamp_low[0] mprj_io[18] vccd1_pad
+ vdda1_pad vdda1_pad2 vssa1_pad vssa1_pad2 vccd1 vdda1 vssa1 vssd1 vssd1_pad mprj_analog[7]
+ mprj_io[21] mprj_analog[8] mprj_io[22] mprj_analog[9] mprj_io[23] mprj_analog[10]
+ mprj_io[24] mprj_analog[5] mprj_clamp_high[1] mprj_clamp_low[1] mprj_io[19] mprj_analog[6]
+ mprj_clamp_high[2] mprj_clamp_low[2] mprj_io[20] vccd2_pad vdda2_pad vssa2_pad vccd
+ vccd2 vdda2 vddio vssa2 vssd2 vssd2_pad vssio flash_csb_core flash_clk_ieb_core
+ flash_clk_oeb_core flash_clk_core flash_csb_oeb_core flash_csb_ieb_core
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfbbp_1 abstract view
.subckt sky130_fd_sc_hd__dfbbp_1 CLK D RESET_B SET_B VGND VNB VPB VPWR Q Q_N
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for spare_logic_block abstract view
.subckt spare_logic_block spare_xfq[0] spare_xfq[1] spare_xfqn[0] spare_xfqn[1] spare_xi[0]
+ spare_xi[1] spare_xi[2] spare_xi[3] spare_xib spare_xmx[0] spare_xmx[1] spare_xna[0]
+ spare_xna[1] spare_xno[0] spare_xno[1] spare_xz[0] spare_xz[10] spare_xz[11] spare_xz[12]
+ spare_xz[13] spare_xz[14] spare_xz[15] spare_xz[16] spare_xz[17] spare_xz[18] spare_xz[19]
+ spare_xz[1] spare_xz[20] spare_xz[21] spare_xz[22] spare_xz[23] spare_xz[24] spare_xz[25]
+ spare_xz[26] spare_xz[2] spare_xz[3] spare_xz[4] spare_xz[5] spare_xz[6] spare_xz[7]
+ spare_xz[8] spare_xz[9] vccd vssd
.ends

* Black-box entry subcircuit for mgmt_core_wrapper abstract view
.subckt mgmt_core_wrapper VGND VPWR core_clk core_rstn debug_in debug_mode debug_oeb
+ debug_out flash_clk flash_csb flash_io0_di flash_io0_do flash_io0_oeb flash_io1_di
+ flash_io1_do flash_io1_oeb flash_io2_di flash_io2_do flash_io2_oeb flash_io3_di
+ flash_io3_do flash_io3_oeb gpio_in_pad gpio_inenb_pad gpio_mode0_pad gpio_mode1_pad
+ gpio_out_pad gpio_outenb_pad hk_ack_i hk_cyc_o hk_dat_i[0] hk_dat_i[10] hk_dat_i[11]
+ hk_dat_i[12] hk_dat_i[13] hk_dat_i[14] hk_dat_i[15] hk_dat_i[16] hk_dat_i[17] hk_dat_i[18]
+ hk_dat_i[19] hk_dat_i[1] hk_dat_i[20] hk_dat_i[21] hk_dat_i[22] hk_dat_i[23] hk_dat_i[24]
+ hk_dat_i[25] hk_dat_i[26] hk_dat_i[27] hk_dat_i[28] hk_dat_i[29] hk_dat_i[2] hk_dat_i[30]
+ hk_dat_i[31] hk_dat_i[3] hk_dat_i[4] hk_dat_i[5] hk_dat_i[6] hk_dat_i[7] hk_dat_i[8]
+ hk_dat_i[9] hk_stb_o irq[0] irq[1] irq[2] irq[3] irq[4] irq[5] la_iena[0] la_iena[100]
+ la_iena[101] la_iena[102] la_iena[103] la_iena[104] la_iena[105] la_iena[106] la_iena[107]
+ la_iena[108] la_iena[109] la_iena[10] la_iena[110] la_iena[111] la_iena[112] la_iena[113]
+ la_iena[114] la_iena[115] la_iena[116] la_iena[117] la_iena[118] la_iena[119] la_iena[11]
+ la_iena[120] la_iena[121] la_iena[122] la_iena[123] la_iena[124] la_iena[125] la_iena[126]
+ la_iena[127] la_iena[12] la_iena[13] la_iena[14] la_iena[15] la_iena[16] la_iena[17]
+ la_iena[18] la_iena[19] la_iena[1] la_iena[20] la_iena[21] la_iena[22] la_iena[23]
+ la_iena[24] la_iena[25] la_iena[26] la_iena[27] la_iena[28] la_iena[29] la_iena[2]
+ la_iena[30] la_iena[31] la_iena[32] la_iena[33] la_iena[34] la_iena[35] la_iena[36]
+ la_iena[37] la_iena[38] la_iena[39] la_iena[3] la_iena[40] la_iena[41] la_iena[42]
+ la_iena[43] la_iena[44] la_iena[45] la_iena[46] la_iena[47] la_iena[48] la_iena[49]
+ la_iena[4] la_iena[50] la_iena[51] la_iena[52] la_iena[53] la_iena[54] la_iena[55]
+ la_iena[56] la_iena[57] la_iena[58] la_iena[59] la_iena[5] la_iena[60] la_iena[61]
+ la_iena[62] la_iena[63] la_iena[64] la_iena[65] la_iena[66] la_iena[67] la_iena[68]
+ la_iena[69] la_iena[6] la_iena[70] la_iena[71] la_iena[72] la_iena[73] la_iena[74]
+ la_iena[75] la_iena[76] la_iena[77] la_iena[78] la_iena[79] la_iena[7] la_iena[80]
+ la_iena[81] la_iena[82] la_iena[83] la_iena[84] la_iena[85] la_iena[86] la_iena[87]
+ la_iena[88] la_iena[89] la_iena[8] la_iena[90] la_iena[91] la_iena[92] la_iena[93]
+ la_iena[94] la_iena[95] la_iena[96] la_iena[97] la_iena[98] la_iena[99] la_iena[9]
+ la_input[0] la_input[100] la_input[101] la_input[102] la_input[103] la_input[104]
+ la_input[105] la_input[106] la_input[107] la_input[108] la_input[109] la_input[10]
+ la_input[110] la_input[111] la_input[112] la_input[113] la_input[114] la_input[115]
+ la_input[116] la_input[117] la_input[118] la_input[119] la_input[11] la_input[120]
+ la_input[121] la_input[122] la_input[123] la_input[124] la_input[125] la_input[126]
+ la_input[127] la_input[12] la_input[13] la_input[14] la_input[15] la_input[16] la_input[17]
+ la_input[18] la_input[19] la_input[1] la_input[20] la_input[21] la_input[22] la_input[23]
+ la_input[24] la_input[25] la_input[26] la_input[27] la_input[28] la_input[29] la_input[2]
+ la_input[30] la_input[31] la_input[32] la_input[33] la_input[34] la_input[35] la_input[36]
+ la_input[37] la_input[38] la_input[39] la_input[3] la_input[40] la_input[41] la_input[42]
+ la_input[43] la_input[44] la_input[45] la_input[46] la_input[47] la_input[48] la_input[49]
+ la_input[4] la_input[50] la_input[51] la_input[52] la_input[53] la_input[54] la_input[55]
+ la_input[56] la_input[57] la_input[58] la_input[59] la_input[5] la_input[60] la_input[61]
+ la_input[62] la_input[63] la_input[64] la_input[65] la_input[66] la_input[67] la_input[68]
+ la_input[69] la_input[6] la_input[70] la_input[71] la_input[72] la_input[73] la_input[74]
+ la_input[75] la_input[76] la_input[77] la_input[78] la_input[79] la_input[7] la_input[80]
+ la_input[81] la_input[82] la_input[83] la_input[84] la_input[85] la_input[86] la_input[87]
+ la_input[88] la_input[89] la_input[8] la_input[90] la_input[91] la_input[92] la_input[93]
+ la_input[94] la_input[95] la_input[96] la_input[97] la_input[98] la_input[99] la_input[9]
+ la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104] la_oenb[105]
+ la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109] la_oenb[10] la_oenb[110] la_oenb[111]
+ la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117] la_oenb[118]
+ la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121] la_oenb[122] la_oenb[123] la_oenb[124]
+ la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12] la_oenb[13] la_oenb[14] la_oenb[15]
+ la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20] la_oenb[21]
+ la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27] la_oenb[28]
+ la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33] la_oenb[34]
+ la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3] la_oenb[40]
+ la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46] la_oenb[47]
+ la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52] la_oenb[53]
+ la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59] la_oenb[5]
+ la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65] la_oenb[66]
+ la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6] la_oenb[70] la_oenb[71] la_oenb[72]
+ la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76] la_oenb[77] la_oenb[78] la_oenb[79]
+ la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84] la_oenb[85]
+ la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89] la_oenb[8] la_oenb[90] la_oenb[91]
+ la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97] la_oenb[98]
+ la_oenb[99] la_oenb[9] la_output[0] la_output[100] la_output[101] la_output[102]
+ la_output[103] la_output[104] la_output[105] la_output[106] la_output[107] la_output[108]
+ la_output[109] la_output[10] la_output[110] la_output[111] la_output[112] la_output[113]
+ la_output[114] la_output[115] la_output[116] la_output[117] la_output[118] la_output[119]
+ la_output[11] la_output[120] la_output[121] la_output[122] la_output[123] la_output[124]
+ la_output[125] la_output[126] la_output[127] la_output[12] la_output[13] la_output[14]
+ la_output[15] la_output[16] la_output[17] la_output[18] la_output[19] la_output[1]
+ la_output[20] la_output[21] la_output[22] la_output[23] la_output[24] la_output[25]
+ la_output[26] la_output[27] la_output[28] la_output[29] la_output[2] la_output[30]
+ la_output[31] la_output[32] la_output[33] la_output[34] la_output[35] la_output[36]
+ la_output[37] la_output[38] la_output[39] la_output[3] la_output[40] la_output[41]
+ la_output[42] la_output[43] la_output[44] la_output[45] la_output[46] la_output[47]
+ la_output[48] la_output[49] la_output[4] la_output[50] la_output[51] la_output[52]
+ la_output[53] la_output[54] la_output[55] la_output[56] la_output[57] la_output[58]
+ la_output[59] la_output[5] la_output[60] la_output[61] la_output[62] la_output[63]
+ la_output[64] la_output[65] la_output[66] la_output[67] la_output[68] la_output[69]
+ la_output[6] la_output[70] la_output[71] la_output[72] la_output[73] la_output[74]
+ la_output[75] la_output[76] la_output[77] la_output[78] la_output[79] la_output[7]
+ la_output[80] la_output[81] la_output[82] la_output[83] la_output[84] la_output[85]
+ la_output[86] la_output[87] la_output[88] la_output[89] la_output[8] la_output[90]
+ la_output[91] la_output[92] la_output[93] la_output[94] la_output[95] la_output[96]
+ la_output[97] la_output[98] la_output[99] la_output[9] mprj_ack_i mprj_adr_o[0]
+ mprj_adr_o[10] mprj_adr_o[11] mprj_adr_o[12] mprj_adr_o[13] mprj_adr_o[14] mprj_adr_o[15]
+ mprj_adr_o[16] mprj_adr_o[17] mprj_adr_o[18] mprj_adr_o[19] mprj_adr_o[1] mprj_adr_o[20]
+ mprj_adr_o[21] mprj_adr_o[22] mprj_adr_o[23] mprj_adr_o[24] mprj_adr_o[25] mprj_adr_o[26]
+ mprj_adr_o[27] mprj_adr_o[28] mprj_adr_o[29] mprj_adr_o[2] mprj_adr_o[30] mprj_adr_o[31]
+ mprj_adr_o[3] mprj_adr_o[4] mprj_adr_o[5] mprj_adr_o[6] mprj_adr_o[7] mprj_adr_o[8]
+ mprj_adr_o[9] mprj_cyc_o mprj_dat_i[0] mprj_dat_i[10] mprj_dat_i[11] mprj_dat_i[12]
+ mprj_dat_i[13] mprj_dat_i[14] mprj_dat_i[15] mprj_dat_i[16] mprj_dat_i[17] mprj_dat_i[18]
+ mprj_dat_i[19] mprj_dat_i[1] mprj_dat_i[20] mprj_dat_i[21] mprj_dat_i[22] mprj_dat_i[23]
+ mprj_dat_i[24] mprj_dat_i[25] mprj_dat_i[26] mprj_dat_i[27] mprj_dat_i[28] mprj_dat_i[29]
+ mprj_dat_i[2] mprj_dat_i[30] mprj_dat_i[31] mprj_dat_i[3] mprj_dat_i[4] mprj_dat_i[5]
+ mprj_dat_i[6] mprj_dat_i[7] mprj_dat_i[8] mprj_dat_i[9] mprj_dat_o[0] mprj_dat_o[10]
+ mprj_dat_o[11] mprj_dat_o[12] mprj_dat_o[13] mprj_dat_o[14] mprj_dat_o[15] mprj_dat_o[16]
+ mprj_dat_o[17] mprj_dat_o[18] mprj_dat_o[19] mprj_dat_o[1] mprj_dat_o[20] mprj_dat_o[21]
+ mprj_dat_o[22] mprj_dat_o[23] mprj_dat_o[24] mprj_dat_o[25] mprj_dat_o[26] mprj_dat_o[27]
+ mprj_dat_o[28] mprj_dat_o[29] mprj_dat_o[2] mprj_dat_o[30] mprj_dat_o[31] mprj_dat_o[3]
+ mprj_dat_o[4] mprj_dat_o[5] mprj_dat_o[6] mprj_dat_o[7] mprj_dat_o[8] mprj_dat_o[9]
+ mprj_sel_o[0] mprj_sel_o[1] mprj_sel_o[2] mprj_sel_o[3] mprj_stb_o mprj_wb_iena
+ mprj_we_o qspi_enabled ser_rx ser_tx spi_csb spi_enabled spi_sck spi_sdi spi_sdo
+ spi_sdoenb sram_ro_addr[0] sram_ro_addr[1] sram_ro_addr[2] sram_ro_addr[3] sram_ro_addr[4]
+ sram_ro_addr[5] sram_ro_addr[6] sram_ro_addr[7] sram_ro_clk sram_ro_csb sram_ro_data[0]
+ sram_ro_data[10] sram_ro_data[11] sram_ro_data[12] sram_ro_data[13] sram_ro_data[14]
+ sram_ro_data[15] sram_ro_data[16] sram_ro_data[17] sram_ro_data[18] sram_ro_data[19]
+ sram_ro_data[1] sram_ro_data[20] sram_ro_data[21] sram_ro_data[22] sram_ro_data[23]
+ sram_ro_data[24] sram_ro_data[25] sram_ro_data[26] sram_ro_data[27] sram_ro_data[28]
+ sram_ro_data[29] sram_ro_data[2] sram_ro_data[30] sram_ro_data[31] sram_ro_data[3]
+ sram_ro_data[4] sram_ro_data[5] sram_ro_data[6] sram_ro_data[7] sram_ro_data[8]
+ sram_ro_data[9] trap uart_enabled user_irq_ena[0] user_irq_ena[1] user_irq_ena[2]
.ends

* Black-box entry subcircuit for user_id_textblock abstract view
.subckt user_id_textblock
.ends

.subckt sky130_fd_pr__cap_mim_m3_2_W5U4AW c2_n3079_n3000# m4_n3179_n3100#
X0 c2_n3079_n3000# m4_n3179_n3100# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
.ends

* Black-box entry subcircuit for sky130_fd_sc_hvl__buf_8 abstract view
.subckt sky130_fd_sc_hvl__buf_8 A VGND VNB VPB VPWR X
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_ZEUEFZ a_n683_n200# a_n189_n297# a_29_n297# a_189_n200#
+ a_n901_n200# a_247_n297# a_n407_n297# a_465_n297# a_407_n200# a_n625_n297# a_683_n297#
+ a_625_n200# a_n843_n297# w_n1101_n497# a_843_n200# a_n29_n200# a_n247_n200# a_n465_n200#
X0 a_n247_n200# a_n407_n297# a_n465_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X1 a_843_n200# a_683_n297# a_625_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X2 a_407_n200# a_247_n297# a_189_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X3 a_189_n200# a_29_n297# a_n29_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X4 a_n465_n200# a_n625_n297# a_n683_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X5 a_625_n200# a_465_n297# a_407_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X6 a_n29_n200# a_n189_n297# a_n247_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X7 a_n683_n200# a_n843_n297# a_n901_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_TGFUGS a_n792_n200# a_298_n200# a_516_n200# a_734_n200#
+ w_n962_n458# a_138_n288# a_n298_n288# a_80_n200# a_356_n288# a_n516_n288# a_574_n288#
+ a_n734_n288# a_n138_n200# a_n356_n200# a_n574_n200# a_n80_n288#
X0 a_80_n200# a_n80_n288# a_n138_n200# w_n962_n458# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X1 a_n574_n200# a_n734_n288# a_n792_n200# w_n962_n458# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X2 a_734_n200# a_574_n288# a_516_n200# w_n962_n458# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X3 a_298_n200# a_138_n288# a_80_n200# w_n962_n458# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X4 a_n138_n200# a_n298_n288# a_n356_n200# w_n962_n458# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X5 a_n356_n200# a_n516_n288# a_n574_n200# w_n962_n458# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X6 a_516_n200# a_356_n288# a_298_n200# w_n962_n458# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p69_S5N9F3 a_n1806_2500# a_n4122_n2932# a_n5280_2500#
+ a_2054_n2932# a_896_n2932# a_4756_2500# a_3598_n2932# a_3212_2500# a_n3736_n2932#
+ a_1668_n2932# a_n1806_n2932# a_5142_n2932# a_896_2500# a_510_n2932# a_n3350_2500#
+ a_n4508_2500# a_3212_n2932# a_n4894_2500# a_1282_2500# w_n5446_n3098# a_4756_n2932#
+ a_2826_2500# a_2826_n2932# a_n2192_n2932# a_n1034_2500# a_n2578_2500# a_n1420_2500#
+ a_n2964_2500# a_n648_n2932# a_n648_2500# a_n5280_n2932# a_n3350_n2932# a_4370_2500#
+ a_1282_n2932# a_124_n2932# a_n1420_n2932# a_n4894_n2932# a_124_2500# a_n2964_n2932#
+ a_n4122_2500# a_2054_2500# a_510_2500# a_n4508_n2932# a_4370_n2932# a_3598_2500#
+ a_3984_2500# a_2440_n2932# a_2440_2500# a_3984_n2932# a_n2192_2500# a_n3736_2500#
+ a_1668_2500# a_n262_n2932# a_n262_2500# a_n1034_n2932# a_5142_2500# a_n2578_n2932#
X0 a_n2578_n2932# a_n2578_2500# w_n5446_n3098# sky130_fd_pr__res_xhigh_po_0p69 l=2.5e+07u
X1 a_n1420_n2932# a_n1420_2500# w_n5446_n3098# sky130_fd_pr__res_xhigh_po_0p69 l=2.5e+07u
X2 a_n1806_n2932# a_n1806_2500# w_n5446_n3098# sky130_fd_pr__res_xhigh_po_0p69 l=2.5e+07u
X3 a_3212_n2932# a_3212_2500# w_n5446_n3098# sky130_fd_pr__res_xhigh_po_0p69 l=2.5e+07u
X4 a_3598_n2932# a_3598_2500# w_n5446_n3098# sky130_fd_pr__res_xhigh_po_0p69 l=2.5e+07u
X5 a_n2964_n2932# a_n2964_2500# w_n5446_n3098# sky130_fd_pr__res_xhigh_po_0p69 l=2.5e+07u
X6 a_2826_n2932# a_2826_2500# w_n5446_n3098# sky130_fd_pr__res_xhigh_po_0p69 l=2.5e+07u
X7 a_4370_n2932# a_4370_2500# w_n5446_n3098# sky130_fd_pr__res_xhigh_po_0p69 l=2.5e+07u
X8 a_3984_n2932# a_3984_2500# w_n5446_n3098# sky130_fd_pr__res_xhigh_po_0p69 l=2.5e+07u
X9 a_n262_n2932# a_n262_2500# w_n5446_n3098# sky130_fd_pr__res_xhigh_po_0p69 l=2.5e+07u
X10 a_n3350_n2932# a_n3350_2500# w_n5446_n3098# sky130_fd_pr__res_xhigh_po_0p69 l=2.5e+07u
X11 a_n4122_n2932# a_n4122_2500# w_n5446_n3098# sky130_fd_pr__res_xhigh_po_0p69 l=2.5e+07u
X12 a_n3736_n2932# a_n3736_2500# w_n5446_n3098# sky130_fd_pr__res_xhigh_po_0p69 l=2.5e+07u
X13 a_5142_n2932# a_5142_2500# w_n5446_n3098# sky130_fd_pr__res_xhigh_po_0p69 l=2.5e+07u
X14 a_n4894_n2932# a_n4894_2500# w_n5446_n3098# sky130_fd_pr__res_xhigh_po_0p69 l=2.5e+07u
X15 a_1282_n2932# a_1282_2500# w_n5446_n3098# sky130_fd_pr__res_xhigh_po_0p69 l=2.5e+07u
X16 a_4756_n2932# a_4756_2500# w_n5446_n3098# sky130_fd_pr__res_xhigh_po_0p69 l=2.5e+07u
X17 a_124_n2932# a_124_2500# w_n5446_n3098# sky130_fd_pr__res_xhigh_po_0p69 l=2.5e+07u
X18 a_510_n2932# a_510_2500# w_n5446_n3098# sky130_fd_pr__res_xhigh_po_0p69 l=2.5e+07u
X19 a_896_n2932# a_896_2500# w_n5446_n3098# sky130_fd_pr__res_xhigh_po_0p69 l=2.5e+07u
X20 a_n648_n2932# a_n648_2500# w_n5446_n3098# sky130_fd_pr__res_xhigh_po_0p69 l=2.5e+07u
X21 a_n5280_n2932# a_n5280_2500# w_n5446_n3098# sky130_fd_pr__res_xhigh_po_0p69 l=2.5e+07u
X22 a_n4508_n2932# a_n4508_2500# w_n5446_n3098# sky130_fd_pr__res_xhigh_po_0p69 l=2.5e+07u
X23 a_n1034_n2932# a_n1034_2500# w_n5446_n3098# sky130_fd_pr__res_xhigh_po_0p69 l=2.5e+07u
X24 a_n2192_n2932# a_n2192_2500# w_n5446_n3098# sky130_fd_pr__res_xhigh_po_0p69 l=2.5e+07u
X25 a_2054_n2932# a_2054_2500# w_n5446_n3098# sky130_fd_pr__res_xhigh_po_0p69 l=2.5e+07u
X26 a_1668_n2932# a_1668_2500# w_n5446_n3098# sky130_fd_pr__res_xhigh_po_0p69 l=2.5e+07u
X27 a_2440_n2932# a_2440_2500# w_n5446_n3098# sky130_fd_pr__res_xhigh_po_0p69 l=2.5e+07u
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_3YBPVB a_n80_n297# a_80_n200# w_n338_n497# a_n138_n200#
X0 a_80_n200# a_n80_n297# a_n138_n200# w_n338_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
.ends

* Black-box entry subcircuit for sky130_fd_sc_hvl__schmittbuf_1 abstract view
.subckt sky130_fd_sc_hvl__schmittbuf_1 A VGND VNB VPB VPWR X
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_PKVMTM w_n308_n458# a_80_n200# a_n138_n200# a_n80_n288#
X0 a_80_n200# a_n80_n288# a_n138_n200# w_n308_n458# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_YUHPXE a_n80_n297# a_80_n200# w_n338_n497# a_n138_n200#
X0 a_80_n200# a_n80_n297# a_n138_n200# w_n338_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_ZK8HQC w_n308_n458# a_80_n200# a_n138_n200# a_n80_n288#
X0 a_80_n200# a_n80_n288# a_n138_n200# w_n308_n458# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_WRT4AW c1_n3036_n3000# m3_n3136_n3100#
X0 c1_n3036_n3000# m3_n3136_n3100# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_YEUEBV a_n792_n200# a_138_n297# a_n298_n297#
+ a_298_n200# a_356_n297# a_n516_n297# a_574_n297# a_516_n200# a_n734_n297# a_734_n200#
+ a_n80_n297# a_80_n200# a_n138_n200# a_n356_n200# a_n574_n200# w_n992_n497#
X0 a_80_n200# a_n80_n297# a_n138_n200# w_n992_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X1 a_n574_n200# a_n734_n297# a_n792_n200# w_n992_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X2 a_734_n200# a_574_n297# a_516_n200# w_n992_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X3 a_298_n200# a_138_n297# a_80_n200# w_n992_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X4 a_n138_n200# a_n298_n297# a_n356_n200# w_n992_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X5 a_n356_n200# a_n516_n297# a_n574_n200# w_n992_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X6 a_516_n200# a_356_n297# a_298_n200# w_n992_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_YUHPBG a_n80_n297# a_80_n200# w_n338_n497# a_n138_n200#
X0 a_80_n200# a_n80_n297# a_n138_n200# w_n338_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
.ends

* Black-box entry subcircuit for sky130_fd_sc_hvl__fill_4 abstract view
.subckt sky130_fd_sc_hvl__fill_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hvl__inv_8 abstract view
.subckt sky130_fd_sc_hvl__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for simple_por abstract view
.subckt simple_por vdd3v3 vdd1v8 vss3v3 porb_h por_l porb_l vss1v8
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtn_1 abstract view
.subckt sky130_fd_sc_hd__dfrtn_1 CLK_N D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_4 abstract view
.subckt sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd1_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd1_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for caravel_clocking abstract view
.subckt caravel_clocking VGND VPWR core_clk ext_clk ext_clk_sel ext_reset pll_clk
+ pll_clk90 resetb resetb_sync sel2[0] sel2[1] sel2[2] sel[0] sel[1] sel[2] user_clk
.ends

* Black-box entry subcircuit for gpio_defaults_block_1803 abstract view
.subckt gpio_defaults_block_1803 VGND VPWR gpio_defaults[0] gpio_defaults[10] gpio_defaults[11]
+ gpio_defaults[12] gpio_defaults[1] gpio_defaults[2] gpio_defaults[3] gpio_defaults[4]
+ gpio_defaults[5] gpio_defaults[6] gpio_defaults[7] gpio_defaults[8] gpio_defaults[9]
.ends

* Black-box entry subcircuit for user_id_programming abstract view
.subckt user_id_programming mask_rev[0] mask_rev[10] mask_rev[11] mask_rev[12] mask_rev[13]
+ mask_rev[14] mask_rev[15] mask_rev[16] mask_rev[17] mask_rev[18] mask_rev[19] mask_rev[1]
+ mask_rev[20] mask_rev[21] mask_rev[22] mask_rev[23] mask_rev[24] mask_rev[25] mask_rev[26]
+ mask_rev[27] mask_rev[28] mask_rev[29] mask_rev[2] mask_rev[30] mask_rev[31] mask_rev[3]
+ mask_rev[4] mask_rev[5] mask_rev[6] mask_rev[7] mask_rev[8] mask_rev[9] VPWR VGND
.ends

* Black-box entry subcircuit for gpio_defaults_block_0403 abstract view
.subckt gpio_defaults_block_0403 VGND VPWR gpio_defaults[0] gpio_defaults[10] gpio_defaults[11]
+ gpio_defaults[12] gpio_defaults[1] gpio_defaults[2] gpio_defaults[3] gpio_defaults[4]
+ gpio_defaults[5] gpio_defaults[6] gpio_defaults[7] gpio_defaults[8] gpio_defaults[9]
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__einvp_8 abstract view
.subckt sky130_fd_sc_hd__einvp_8 A TE VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_12 abstract view
.subckt sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__einvp_4 abstract view
.subckt sky130_fd_sc_hd__einvp_4 A TE VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

.subckt sky130_fd_sc_hd__decap_12 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
.ends

.subckt mprj2_logic_high HI vccd2 vssd2
XFILLER_0_57 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_209 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_69 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_15 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_81 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_1_181 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_29 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_3 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_193 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_1_95 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XPHY_0 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_1 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_1_85 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_1_41 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_53 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_2 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_3 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_1_141 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_197 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_153 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_165 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_209 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_1_57 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_113 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_69 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_169 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_125 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_15 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_181 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_137 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_193 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_1_29 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_107 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_141 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_197 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_153 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_165 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_113 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_3 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_169 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_125 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_137 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_81 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_3
Xinst vssd2 vssd2 vccd2 vccd2 HI inst/LO sky130_fd_sc_hd__conb_1
XFILLER_0_85 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_41 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_109 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_97 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_53 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_3
.ends

.subckt mprj_logic_high HI[0] HI[100] HI[101] HI[102] HI[103] HI[104] HI[105] HI[106]
+ HI[107] HI[108] HI[109] HI[10] HI[110] HI[111] HI[112] HI[113] HI[114] HI[115] HI[116]
+ HI[117] HI[118] HI[119] HI[11] HI[120] HI[121] HI[122] HI[123] HI[124] HI[125] HI[126]
+ HI[127] HI[128] HI[129] HI[12] HI[130] HI[131] HI[132] HI[133] HI[134] HI[135] HI[136]
+ HI[137] HI[138] HI[139] HI[13] HI[140] HI[141] HI[142] HI[143] HI[144] HI[145] HI[146]
+ HI[147] HI[148] HI[149] HI[14] HI[150] HI[151] HI[152] HI[153] HI[154] HI[155] HI[156]
+ HI[157] HI[158] HI[159] HI[15] HI[160] HI[161] HI[162] HI[163] HI[164] HI[165] HI[166]
+ HI[167] HI[168] HI[169] HI[16] HI[170] HI[171] HI[172] HI[173] HI[174] HI[175] HI[176]
+ HI[177] HI[178] HI[179] HI[17] HI[180] HI[181] HI[182] HI[183] HI[184] HI[185] HI[186]
+ HI[187] HI[188] HI[189] HI[18] HI[190] HI[191] HI[192] HI[193] HI[194] HI[195] HI[196]
+ HI[197] HI[198] HI[199] HI[19] HI[1] HI[200] HI[201] HI[202] HI[203] HI[204] HI[205]
+ HI[206] HI[207] HI[208] HI[209] HI[20] HI[210] HI[211] HI[212] HI[213] HI[214] HI[215]
+ HI[216] HI[217] HI[218] HI[219] HI[21] HI[220] HI[221] HI[222] HI[223] HI[224] HI[225]
+ HI[226] HI[227] HI[228] HI[229] HI[22] HI[230] HI[231] HI[232] HI[233] HI[234] HI[235]
+ HI[236] HI[237] HI[238] HI[239] HI[23] HI[240] HI[241] HI[242] HI[243] HI[244] HI[245]
+ HI[246] HI[247] HI[248] HI[249] HI[24] HI[250] HI[251] HI[252] HI[253] HI[254] HI[255]
+ HI[256] HI[257] HI[258] HI[259] HI[25] HI[260] HI[261] HI[262] HI[263] HI[264] HI[265]
+ HI[266] HI[267] HI[268] HI[269] HI[26] HI[270] HI[271] HI[272] HI[273] HI[274] HI[275]
+ HI[276] HI[277] HI[278] HI[279] HI[27] HI[280] HI[281] HI[282] HI[283] HI[284] HI[285]
+ HI[286] HI[287] HI[288] HI[289] HI[28] HI[290] HI[291] HI[292] HI[293] HI[294] HI[295]
+ HI[296] HI[297] HI[298] HI[299] HI[29] HI[2] HI[300] HI[301] HI[302] HI[303] HI[304]
+ HI[305] HI[306] HI[307] HI[308] HI[309] HI[30] HI[310] HI[311] HI[312] HI[313] HI[314]
+ HI[315] HI[316] HI[317] HI[318] HI[319] HI[31] HI[320] HI[321] HI[322] HI[323] HI[324]
+ HI[325] HI[326] HI[327] HI[328] HI[329] HI[32] HI[330] HI[331] HI[332] HI[333] HI[334]
+ HI[335] HI[336] HI[337] HI[338] HI[339] HI[33] HI[340] HI[341] HI[342] HI[343] HI[344]
+ HI[345] HI[346] HI[347] HI[348] HI[349] HI[34] HI[350] HI[351] HI[352] HI[353] HI[354]
+ HI[355] HI[356] HI[357] HI[358] HI[359] HI[35] HI[360] HI[361] HI[362] HI[363] HI[364]
+ HI[365] HI[366] HI[367] HI[368] HI[369] HI[36] HI[370] HI[371] HI[372] HI[373] HI[374]
+ HI[375] HI[376] HI[377] HI[378] HI[379] HI[37] HI[380] HI[381] HI[382] HI[383] HI[384]
+ HI[385] HI[386] HI[387] HI[388] HI[389] HI[38] HI[390] HI[391] HI[392] HI[393] HI[394]
+ HI[395] HI[396] HI[397] HI[398] HI[399] HI[39] HI[3] HI[400] HI[401] HI[402] HI[403]
+ HI[404] HI[405] HI[406] HI[407] HI[408] HI[409] HI[40] HI[410] HI[411] HI[412] HI[413]
+ HI[414] HI[415] HI[416] HI[417] HI[418] HI[419] HI[41] HI[420] HI[421] HI[422] HI[423]
+ HI[424] HI[425] HI[426] HI[427] HI[428] HI[429] HI[42] HI[430] HI[431] HI[432] HI[433]
+ HI[434] HI[435] HI[436] HI[437] HI[438] HI[439] HI[43] HI[440] HI[441] HI[442] HI[443]
+ HI[444] HI[445] HI[446] HI[447] HI[448] HI[449] HI[44] HI[450] HI[451] HI[452] HI[453]
+ HI[454] HI[455] HI[456] HI[457] HI[458] HI[459] HI[45] HI[460] HI[461] HI[462] HI[46]
+ HI[47] HI[48] HI[49] HI[4] HI[50] HI[51] HI[52] HI[53] HI[54] HI[55] HI[56] HI[57]
+ HI[58] HI[59] HI[5] HI[60] HI[61] HI[62] HI[63] HI[64] HI[65] HI[66] HI[67] HI[68]
+ HI[69] HI[6] HI[70] HI[71] HI[72] HI[73] HI[74] HI[75] HI[76] HI[77] HI[78] HI[79]
+ HI[7] HI[80] HI[81] HI[82] HI[83] HI[84] HI[85] HI[86] HI[87] HI[88] HI[89] HI[8]
+ HI[90] HI[91] HI[92] HI[93] HI[94] HI[95] HI[96] HI[97] HI[98] HI[99] HI[9] vccd1
+ vssd1
Xinsts\[210\] vssd1 vssd1 vccd1 vccd1 HI[210] insts\[210\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[308\] vssd1 vssd1 vccd1 vccd1 HI[308] insts\[308\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[425\] vssd1 vssd1 vccd1 vccd1 HI[425] insts\[425\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[160\] vssd1 vssd1 vccd1 vccd1 HI[160] insts\[160\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_357 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_302 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[258\] vssd1 vssd1 vccd1 vccd1 HI[258] insts\[258\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[40\] vssd1 vssd1 vccd1 vccd1 HI[40] insts\[40\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[375\] vssd1 vssd1 vccd1 vccd1 HI[375] insts\[375\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[88\] vssd1 vssd1 vccd1 vccd1 HI[88] insts\[88\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_165 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[123\] vssd1 vssd1 vccd1 vccd1 HI[123] insts\[123\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_669 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[338\] vssd1 vssd1 vccd1 vccd1 HI[338] insts\[338\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[240\] vssd1 vssd1 vccd1 vccd1 HI[240] insts\[240\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[9\] vssd1 vssd1 vccd1 vccd1 HI[9] insts\[9\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[455\] vssd1 vssd1 vccd1 vccd1 HI[455] insts\[455\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[288\] vssd1 vssd1 vccd1 vccd1 HI[288] insts\[288\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[190\] vssd1 vssd1 vccd1 vccd1 HI[190] insts\[190\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[70\] vssd1 vssd1 vccd1 vccd1 HI[70] insts\[70\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[203\] vssd1 vssd1 vccd1 vccd1 HI[203] insts\[203\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_561 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[418\] vssd1 vssd1 vccd1 vccd1 HI[418] insts\[418\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[153\] vssd1 vssd1 vccd1 vccd1 HI[153] insts\[153\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[320\] vssd1 vssd1 vccd1 vccd1 HI[320] insts\[320\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[33\] vssd1 vssd1 vccd1 vccd1 HI[33] insts\[33\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[368\] vssd1 vssd1 vccd1 vccd1 HI[368] insts\[368\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[270\] vssd1 vssd1 vccd1 vccd1 HI[270] insts\[270\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_177 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_486 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[116\] vssd1 vssd1 vccd1 vccd1 HI[116] insts\[116\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[400\] vssd1 vssd1 vccd1 vccd1 HI[400] insts\[400\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[233\] vssd1 vssd1 vccd1 vccd1 HI[233] insts\[233\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_209 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[183\] vssd1 vssd1 vccd1 vccd1 HI[183] insts\[183\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[350\] vssd1 vssd1 vccd1 vccd1 HI[350] insts\[350\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[448\] vssd1 vssd1 vccd1 vccd1 HI[448] insts\[448\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_721 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[63\] vssd1 vssd1 vccd1 vccd1 HI[63] insts\[63\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[398\] vssd1 vssd1 vccd1 vccd1 HI[398] insts\[398\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_573 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[146\] vssd1 vssd1 vccd1 vccd1 HI[146] insts\[146\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[313\] vssd1 vssd1 vccd1 vccd1 HI[313] insts\[313\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[26\] vssd1 vssd1 vccd1 vccd1 HI[26] insts\[26\]/LO sky130_fd_sc_hd__conb_1
XFILLER_3_3 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[430\] vssd1 vssd1 vccd1 vccd1 HI[430] insts\[430\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_189 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[263\] vssd1 vssd1 vccd1 vccd1 HI[263] insts\[263\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[380\] vssd1 vssd1 vccd1 vccd1 HI[380] insts\[380\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[109\] vssd1 vssd1 vccd1 vccd1 HI[109] insts\[109\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[93\] vssd1 vssd1 vccd1 vccd1 HI[93] insts\[93\]/LO sky130_fd_sc_hd__conb_1
XFILLER_3_498 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_80 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[226\] vssd1 vssd1 vccd1 vccd1 HI[226] insts\[226\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[343\] vssd1 vssd1 vccd1 vccd1 HI[343] insts\[343\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[176\] vssd1 vssd1 vccd1 vccd1 HI[176] insts\[176\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[56\] vssd1 vssd1 vccd1 vccd1 HI[56] insts\[56\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[460\] vssd1 vssd1 vccd1 vccd1 HI[460] insts\[460\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[293\] vssd1 vssd1 vccd1 vccd1 HI[293] insts\[293\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_541 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_585 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[139\] vssd1 vssd1 vccd1 vccd1 HI[139] insts\[139\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[306\] vssd1 vssd1 vccd1 vccd1 HI[306] insts\[306\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[19\] vssd1 vssd1 vccd1 vccd1 HI[19] insts\[19\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_393 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[423\] vssd1 vssd1 vccd1 vccd1 HI[423] insts\[423\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[256\] vssd1 vssd1 vccd1 vccd1 HI[256] insts\[256\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[373\] vssd1 vssd1 vccd1 vccd1 HI[373] insts\[373\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_617 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[86\] vssd1 vssd1 vccd1 vccd1 HI[86] insts\[86\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[121\] vssd1 vssd1 vccd1 vccd1 HI[121] insts\[121\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[219\] vssd1 vssd1 vccd1 vccd1 HI[219] insts\[219\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[336\] vssd1 vssd1 vccd1 vccd1 HI[336] insts\[336\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[169\] vssd1 vssd1 vccd1 vccd1 HI[169] insts\[169\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[49\] vssd1 vssd1 vccd1 vccd1 HI[49] insts\[49\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[286\] vssd1 vssd1 vccd1 vccd1 HI[286] insts\[286\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[7\] vssd1 vssd1 vccd1 vccd1 HI[7] insts\[7\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[453\] vssd1 vssd1 vccd1 vccd1 HI[453] insts\[453\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_597 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[201\] vssd1 vssd1 vccd1 vccd1 HI[201] insts\[201\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[416\] vssd1 vssd1 vccd1 vccd1 HI[416] insts\[416\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[151\] vssd1 vssd1 vccd1 vccd1 HI[151] insts\[151\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[249\] vssd1 vssd1 vccd1 vccd1 HI[249] insts\[249\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_681 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_8
Xinsts\[31\] vssd1 vssd1 vccd1 vccd1 HI[31] insts\[31\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_629 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[366\] vssd1 vssd1 vccd1 vccd1 HI[366] insts\[366\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[199\] vssd1 vssd1 vccd1 vccd1 HI[199] insts\[199\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[79\] vssd1 vssd1 vccd1 vccd1 HI[79] insts\[79\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[114\] vssd1 vssd1 vccd1 vccd1 HI[114] insts\[114\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[329\] vssd1 vssd1 vccd1 vccd1 HI[329] insts\[329\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[231\] vssd1 vssd1 vccd1 vccd1 HI[231] insts\[231\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[446\] vssd1 vssd1 vccd1 vccd1 HI[446] insts\[446\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[181\] vssd1 vssd1 vccd1 vccd1 HI[181] insts\[181\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[279\] vssd1 vssd1 vccd1 vccd1 HI[279] insts\[279\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[61\] vssd1 vssd1 vccd1 vccd1 HI[61] insts\[61\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[396\] vssd1 vssd1 vccd1 vccd1 HI[396] insts\[396\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[144\] vssd1 vssd1 vccd1 vccd1 HI[144] insts\[144\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[409\] vssd1 vssd1 vccd1 vccd1 HI[409] insts\[409\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[311\] vssd1 vssd1 vccd1 vccd1 HI[311] insts\[311\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[24\] vssd1 vssd1 vccd1 vccd1 HI[24] insts\[24\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[359\] vssd1 vssd1 vccd1 vccd1 HI[359] insts\[359\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_3 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[261\] vssd1 vssd1 vccd1 vccd1 HI[261] insts\[261\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[107\] vssd1 vssd1 vccd1 vccd1 HI[107] insts\[107\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[91\] vssd1 vssd1 vccd1 vccd1 HI[91] insts\[91\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[224\] vssd1 vssd1 vccd1 vccd1 HI[224] insts\[224\]/LO sky130_fd_sc_hd__conb_1
XPHY_0 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[439\] vssd1 vssd1 vccd1 vccd1 HI[439] insts\[439\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[174\] vssd1 vssd1 vccd1 vccd1 HI[174] insts\[174\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[341\] vssd1 vssd1 vccd1 vccd1 HI[341] insts\[341\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[54\] vssd1 vssd1 vccd1 vccd1 HI[54] insts\[54\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[389\] vssd1 vssd1 vccd1 vccd1 HI[389] insts\[389\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[291\] vssd1 vssd1 vccd1 vccd1 HI[291] insts\[291\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[137\] vssd1 vssd1 vccd1 vccd1 HI[137] insts\[137\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[304\] vssd1 vssd1 vccd1 vccd1 HI[304] insts\[304\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[17\] vssd1 vssd1 vccd1 vccd1 HI[17] insts\[17\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[421\] vssd1 vssd1 vccd1 vccd1 HI[421] insts\[421\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[254\] vssd1 vssd1 vccd1 vccd1 HI[254] insts\[254\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[371\] vssd1 vssd1 vccd1 vccd1 HI[371] insts\[371\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[84\] vssd1 vssd1 vccd1 vccd1 HI[84] insts\[84\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[217\] vssd1 vssd1 vccd1 vccd1 HI[217] insts\[217\]/LO sky130_fd_sc_hd__conb_1
XPHY_1 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[334\] vssd1 vssd1 vccd1 vccd1 HI[334] insts\[334\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[167\] vssd1 vssd1 vccd1 vccd1 HI[167] insts\[167\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[47\] vssd1 vssd1 vccd1 vccd1 HI[47] insts\[47\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_309 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[5\] vssd1 vssd1 vccd1 vccd1 HI[5] insts\[5\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[451\] vssd1 vssd1 vccd1 vccd1 HI[451] insts\[451\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[284\] vssd1 vssd1 vccd1 vccd1 HI[284] insts\[284\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_331 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_172 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[247\] vssd1 vssd1 vccd1 vccd1 HI[247] insts\[247\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[414\] vssd1 vssd1 vccd1 vccd1 HI[414] insts\[414\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_470 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_96 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[364\] vssd1 vssd1 vccd1 vccd1 HI[364] insts\[364\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[197\] vssd1 vssd1 vccd1 vccd1 HI[197] insts\[197\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[77\] vssd1 vssd1 vccd1 vccd1 HI[77] insts\[77\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[112\] vssd1 vssd1 vccd1 vccd1 HI[112] insts\[112\]/LO sky130_fd_sc_hd__conb_1
XPHY_2 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[327\] vssd1 vssd1 vccd1 vccd1 HI[327] insts\[327\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_557 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[444\] vssd1 vssd1 vccd1 vccd1 HI[444] insts\[444\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[277\] vssd1 vssd1 vccd1 vccd1 HI[277] insts\[277\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_343 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[394\] vssd1 vssd1 vccd1 vccd1 HI[394] insts\[394\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_118 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_184 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[407\] vssd1 vssd1 vccd1 vccd1 HI[407] insts\[407\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[142\] vssd1 vssd1 vccd1 vccd1 HI[142] insts\[142\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[22\] vssd1 vssd1 vccd1 vccd1 HI[22] insts\[22\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[357\] vssd1 vssd1 vccd1 vccd1 HI[357] insts\[357\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[105\] vssd1 vssd1 vccd1 vccd1 HI[105] insts\[105\]/LO sky130_fd_sc_hd__conb_1
XPHY_3 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[222\] vssd1 vssd1 vccd1 vccd1 HI[222] insts\[222\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[437\] vssd1 vssd1 vccd1 vccd1 HI[437] insts\[437\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[172\] vssd1 vssd1 vccd1 vccd1 HI[172] insts\[172\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_355 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[52\] vssd1 vssd1 vccd1 vccd1 HI[52] insts\[52\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[387\] vssd1 vssd1 vccd1 vccd1 HI[387] insts\[387\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_196 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_8
Xinsts\[135\] vssd1 vssd1 vccd1 vccd1 HI[135] insts\[135\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[302\] vssd1 vssd1 vccd1 vccd1 HI[302] insts\[302\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[15\] vssd1 vssd1 vccd1 vccd1 HI[15] insts\[15\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[252\] vssd1 vssd1 vccd1 vccd1 HI[252] insts\[252\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[82\] vssd1 vssd1 vccd1 vccd1 HI[82] insts\[82\]/LO sky130_fd_sc_hd__conb_1
XPHY_4 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[215\] vssd1 vssd1 vccd1 vccd1 HI[215] insts\[215\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[165\] vssd1 vssd1 vccd1 vccd1 HI[165] insts\[165\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[332\] vssd1 vssd1 vccd1 vccd1 HI[332] insts\[332\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_301 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_367 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[45\] vssd1 vssd1 vccd1 vccd1 HI[45] insts\[45\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_109 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[3\] vssd1 vssd1 vccd1 vccd1 HI[3] insts\[3\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_142 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[282\] vssd1 vssd1 vccd1 vccd1 HI[282] insts\[282\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[128\] vssd1 vssd1 vccd1 vccd1 HI[128] insts\[128\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[412\] vssd1 vssd1 vccd1 vccd1 HI[412] insts\[412\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[245\] vssd1 vssd1 vccd1 vccd1 HI[245] insts\[245\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[362\] vssd1 vssd1 vccd1 vccd1 HI[362] insts\[362\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[195\] vssd1 vssd1 vccd1 vccd1 HI[195] insts\[195\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[75\] vssd1 vssd1 vccd1 vccd1 HI[75] insts\[75\]/LO sky130_fd_sc_hd__conb_1
XPHY_5 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[110\] vssd1 vssd1 vccd1 vccd1 HI[110] insts\[110\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[208\] vssd1 vssd1 vccd1 vccd1 HI[208] insts\[208\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_505 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[158\] vssd1 vssd1 vccd1 vccd1 HI[158] insts\[158\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[325\] vssd1 vssd1 vccd1 vccd1 HI[325] insts\[325\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_379 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[38\] vssd1 vssd1 vccd1 vccd1 HI[38] insts\[38\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[442\] vssd1 vssd1 vccd1 vccd1 HI[442] insts\[442\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[275\] vssd1 vssd1 vccd1 vccd1 HI[275] insts\[275\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_154 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_121 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[392\] vssd1 vssd1 vccd1 vccd1 HI[392] insts\[392\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[405\] vssd1 vssd1 vccd1 vccd1 HI[405] insts\[405\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[140\] vssd1 vssd1 vccd1 vccd1 HI[140] insts\[140\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[238\] vssd1 vssd1 vccd1 vccd1 HI[238] insts\[238\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[20\] vssd1 vssd1 vccd1 vccd1 HI[20] insts\[20\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[355\] vssd1 vssd1 vccd1 vccd1 HI[355] insts\[355\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[188\] vssd1 vssd1 vccd1 vccd1 HI[188] insts\[188\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_709 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[68\] vssd1 vssd1 vccd1 vccd1 HI[68] insts\[68\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_517 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[103\] vssd1 vssd1 vccd1 vccd1 HI[103] insts\[103\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[318\] vssd1 vssd1 vccd1 vccd1 HI[318] insts\[318\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[220\] vssd1 vssd1 vccd1 vccd1 HI[220] insts\[220\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[170\] vssd1 vssd1 vccd1 vccd1 HI[170] insts\[170\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[435\] vssd1 vssd1 vccd1 vccd1 HI[435] insts\[435\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_689 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_645 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_601 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_133 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[268\] vssd1 vssd1 vccd1 vccd1 HI[268] insts\[268\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[50\] vssd1 vssd1 vccd1 vccd1 HI[50] insts\[50\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[385\] vssd1 vssd1 vccd1 vccd1 HI[385] insts\[385\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[98\] vssd1 vssd1 vccd1 vccd1 HI[98] insts\[98\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_442 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_68 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[133\] vssd1 vssd1 vccd1 vccd1 HI[133] insts\[133\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[300\] vssd1 vssd1 vccd1 vccd1 HI[300] insts\[300\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[13\] vssd1 vssd1 vccd1 vccd1 HI[13] insts\[13\]/LO sky130_fd_sc_hd__conb_1
XPHY_7 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[348\] vssd1 vssd1 vccd1 vccd1 HI[348] insts\[348\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[250\] vssd1 vssd1 vccd1 vccd1 HI[250] insts\[250\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[298\] vssd1 vssd1 vccd1 vccd1 HI[298] insts\[298\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_529 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[80\] vssd1 vssd1 vccd1 vccd1 HI[80] insts\[80\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[213\] vssd1 vssd1 vccd1 vccd1 HI[213] insts\[213\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_337 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[428\] vssd1 vssd1 vccd1 vccd1 HI[428] insts\[428\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_657 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_613 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[330\] vssd1 vssd1 vccd1 vccd1 HI[330] insts\[330\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[163\] vssd1 vssd1 vccd1 vccd1 HI[163] insts\[163\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[43\] vssd1 vssd1 vccd1 vccd1 HI[43] insts\[43\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[378\] vssd1 vssd1 vccd1 vccd1 HI[378] insts\[378\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[280\] vssd1 vssd1 vccd1 vccd1 HI[280] insts\[280\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[1\] vssd1 vssd1 vccd1 vccd1 HI[1] insts\[1\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_454 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_421 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_410 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_8
Xinsts\[126\] vssd1 vssd1 vccd1 vccd1 HI[126] insts\[126\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[410\] vssd1 vssd1 vccd1 vccd1 HI[410] insts\[410\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[243\] vssd1 vssd1 vccd1 vccd1 HI[243] insts\[243\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[458\] vssd1 vssd1 vccd1 vccd1 HI[458] insts\[458\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[360\] vssd1 vssd1 vccd1 vccd1 HI[360] insts\[360\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[193\] vssd1 vssd1 vccd1 vccd1 HI[193] insts\[193\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[73\] vssd1 vssd1 vccd1 vccd1 HI[73] insts\[73\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[206\] vssd1 vssd1 vccd1 vccd1 HI[206] insts\[206\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_669 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_625 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_113 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[156\] vssd1 vssd1 vccd1 vccd1 HI[156] insts\[156\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[323\] vssd1 vssd1 vccd1 vccd1 HI[323] insts\[323\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[36\] vssd1 vssd1 vccd1 vccd1 HI[36] insts\[36\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[273\] vssd1 vssd1 vccd1 vccd1 HI[273] insts\[273\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[440\] vssd1 vssd1 vccd1 vccd1 HI[440] insts\[440\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_433 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[390\] vssd1 vssd1 vccd1 vccd1 HI[390] insts\[390\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[119\] vssd1 vssd1 vccd1 vccd1 HI[119] insts\[119\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[403\] vssd1 vssd1 vccd1 vccd1 HI[403] insts\[403\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[236\] vssd1 vssd1 vccd1 vccd1 HI[236] insts\[236\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_701 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[353\] vssd1 vssd1 vccd1 vccd1 HI[353] insts\[353\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[186\] vssd1 vssd1 vccd1 vccd1 HI[186] insts\[186\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[66\] vssd1 vssd1 vccd1 vccd1 HI[66] insts\[66\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[101\] vssd1 vssd1 vccd1 vccd1 HI[101] insts\[101\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[149\] vssd1 vssd1 vccd1 vccd1 HI[149] insts\[149\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_637 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[316\] vssd1 vssd1 vccd1 vccd1 HI[316] insts\[316\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[29\] vssd1 vssd1 vccd1 vccd1 HI[29] insts\[29\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[433\] vssd1 vssd1 vccd1 vccd1 HI[433] insts\[433\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[266\] vssd1 vssd1 vccd1 vccd1 HI[266] insts\[266\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[383\] vssd1 vssd1 vccd1 vccd1 HI[383] insts\[383\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[96\] vssd1 vssd1 vccd1 vccd1 HI[96] insts\[96\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_253 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[131\] vssd1 vssd1 vccd1 vccd1 HI[131] insts\[131\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[229\] vssd1 vssd1 vccd1 vccd1 HI[229] insts\[229\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_713 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[11\] vssd1 vssd1 vccd1 vccd1 HI[11] insts\[11\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[346\] vssd1 vssd1 vccd1 vccd1 HI[346] insts\[346\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[179\] vssd1 vssd1 vccd1 vccd1 HI[179] insts\[179\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[59\] vssd1 vssd1 vccd1 vccd1 HI[59] insts\[59\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_307 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[296\] vssd1 vssd1 vccd1 vccd1 HI[296] insts\[296\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[309\] vssd1 vssd1 vccd1 vccd1 HI[309] insts\[309\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[211\] vssd1 vssd1 vccd1 vccd1 HI[211] insts\[211\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[426\] vssd1 vssd1 vccd1 vccd1 HI[426] insts\[426\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[161\] vssd1 vssd1 vccd1 vccd1 HI[161] insts\[161\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[259\] vssd1 vssd1 vccd1 vccd1 HI[259] insts\[259\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[41\] vssd1 vssd1 vccd1 vccd1 HI[41] insts\[41\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_490 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_722 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[376\] vssd1 vssd1 vccd1 vccd1 HI[376] insts\[376\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_265 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_221 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[89\] vssd1 vssd1 vccd1 vccd1 HI[89] insts\[89\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_60 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[124\] vssd1 vssd1 vccd1 vccd1 HI[124] insts\[124\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_725 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[241\] vssd1 vssd1 vccd1 vccd1 HI[241] insts\[241\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[339\] vssd1 vssd1 vccd1 vccd1 HI[339] insts\[339\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_319 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_8
Xinsts\[456\] vssd1 vssd1 vccd1 vccd1 HI[456] insts\[456\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[289\] vssd1 vssd1 vccd1 vccd1 HI[289] insts\[289\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[191\] vssd1 vssd1 vccd1 vccd1 HI[191] insts\[191\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[71\] vssd1 vssd1 vccd1 vccd1 HI[71] insts\[71\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[204\] vssd1 vssd1 vccd1 vccd1 HI[204] insts\[204\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[419\] vssd1 vssd1 vccd1 vccd1 HI[419] insts\[419\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[154\] vssd1 vssd1 vccd1 vccd1 HI[154] insts\[154\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[321\] vssd1 vssd1 vccd1 vccd1 HI[321] insts\[321\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[34\] vssd1 vssd1 vccd1 vccd1 HI[34] insts\[34\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[369\] vssd1 vssd1 vccd1 vccd1 HI[369] insts\[369\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_277 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_233 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[271\] vssd1 vssd1 vccd1 vccd1 HI[271] insts\[271\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_72 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[117\] vssd1 vssd1 vccd1 vccd1 HI[117] insts\[117\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[234\] vssd1 vssd1 vccd1 vccd1 HI[234] insts\[234\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[401\] vssd1 vssd1 vccd1 vccd1 HI[401] insts\[401\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[351\] vssd1 vssd1 vccd1 vccd1 HI[351] insts\[351\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[449\] vssd1 vssd1 vccd1 vccd1 HI[449] insts\[449\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[184\] vssd1 vssd1 vccd1 vccd1 HI[184] insts\[184\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[64\] vssd1 vssd1 vccd1 vccd1 HI[64] insts\[64\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[399\] vssd1 vssd1 vccd1 vccd1 HI[399] insts\[399\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_673 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[147\] vssd1 vssd1 vccd1 vccd1 HI[147] insts\[147\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[314\] vssd1 vssd1 vccd1 vccd1 HI[314] insts\[314\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[27\] vssd1 vssd1 vccd1 vccd1 HI[27] insts\[27\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[431\] vssd1 vssd1 vccd1 vccd1 HI[431] insts\[431\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_289 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_245 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[264\] vssd1 vssd1 vccd1 vccd1 HI[264] insts\[264\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[381\] vssd1 vssd1 vccd1 vccd1 HI[381] insts\[381\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[94\] vssd1 vssd1 vccd1 vccd1 HI[94] insts\[94\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[227\] vssd1 vssd1 vccd1 vccd1 HI[227] insts\[227\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[344\] vssd1 vssd1 vccd1 vccd1 HI[344] insts\[344\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[177\] vssd1 vssd1 vccd1 vccd1 HI[177] insts\[177\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[57\] vssd1 vssd1 vccd1 vccd1 HI[57] insts\[57\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[461\] vssd1 vssd1 vccd1 vccd1 HI[461] insts\[461\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[294\] vssd1 vssd1 vccd1 vccd1 HI[294] insts\[294\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_641 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_685 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[307\] vssd1 vssd1 vccd1 vccd1 HI[307] insts\[307\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_471 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_8
Xinsts\[424\] vssd1 vssd1 vccd1 vccd1 HI[424] insts\[424\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[257\] vssd1 vssd1 vccd1 vccd1 HI[257] insts\[257\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_85 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_511 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[374\] vssd1 vssd1 vccd1 vccd1 HI[374] insts\[374\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[87\] vssd1 vssd1 vccd1 vccd1 HI[87] insts\[87\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[122\] vssd1 vssd1 vccd1 vccd1 HI[122] insts\[122\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[337\] vssd1 vssd1 vccd1 vccd1 HI[337] insts\[337\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_108 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[8\] vssd1 vssd1 vccd1 vccd1 HI[8] insts\[8\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[454\] vssd1 vssd1 vccd1 vccd1 HI[454] insts\[454\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[287\] vssd1 vssd1 vccd1 vccd1 HI[287] insts\[287\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_653 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_697 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[202\] vssd1 vssd1 vccd1 vccd1 HI[202] insts\[202\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_461 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[417\] vssd1 vssd1 vccd1 vccd1 HI[417] insts\[417\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[152\] vssd1 vssd1 vccd1 vccd1 HI[152] insts\[152\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_97 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[32\] vssd1 vssd1 vccd1 vccd1 HI[32] insts\[32\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[367\] vssd1 vssd1 vccd1 vccd1 HI[367] insts\[367\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[115\] vssd1 vssd1 vccd1 vccd1 HI[115] insts\[115\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[232\] vssd1 vssd1 vccd1 vccd1 HI[232] insts\[232\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[447\] vssd1 vssd1 vccd1 vccd1 HI[447] insts\[447\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[182\] vssd1 vssd1 vccd1 vccd1 HI[182] insts\[182\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[62\] vssd1 vssd1 vccd1 vccd1 HI[62] insts\[62\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_665 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[397\] vssd1 vssd1 vccd1 vccd1 HI[397] insts\[397\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_484 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[145\] vssd1 vssd1 vccd1 vccd1 HI[145] insts\[145\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[312\] vssd1 vssd1 vccd1 vccd1 HI[312] insts\[312\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[25\] vssd1 vssd1 vccd1 vccd1 HI[25] insts\[25\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_281 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[262\] vssd1 vssd1 vccd1 vccd1 HI[262] insts\[262\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_3 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_8
Xinsts\[108\] vssd1 vssd1 vccd1 vccd1 HI[108] insts\[108\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[92\] vssd1 vssd1 vccd1 vccd1 HI[92] insts\[92\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[225\] vssd1 vssd1 vccd1 vccd1 HI[225] insts\[225\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[342\] vssd1 vssd1 vccd1 vccd1 HI[342] insts\[342\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[175\] vssd1 vssd1 vccd1 vccd1 HI[175] insts\[175\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[55\] vssd1 vssd1 vccd1 vccd1 HI[55] insts\[55\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[292\] vssd1 vssd1 vccd1 vccd1 HI[292] insts\[292\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_441 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[138\] vssd1 vssd1 vccd1 vccd1 HI[138] insts\[138\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[305\] vssd1 vssd1 vccd1 vccd1 HI[305] insts\[305\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[18\] vssd1 vssd1 vccd1 vccd1 HI[18] insts\[18\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_293 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_8
Xinsts\[422\] vssd1 vssd1 vccd1 vccd1 HI[422] insts\[422\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[255\] vssd1 vssd1 vccd1 vccd1 HI[255] insts\[255\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[372\] vssd1 vssd1 vccd1 vccd1 HI[372] insts\[372\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[85\] vssd1 vssd1 vccd1 vccd1 HI[85] insts\[85\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[120\] vssd1 vssd1 vccd1 vccd1 HI[120] insts\[120\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[218\] vssd1 vssd1 vccd1 vccd1 HI[218] insts\[218\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[335\] vssd1 vssd1 vccd1 vccd1 HI[335] insts\[335\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[168\] vssd1 vssd1 vccd1 vccd1 HI[168] insts\[168\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[48\] vssd1 vssd1 vccd1 vccd1 HI[48] insts\[48\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[6\] vssd1 vssd1 vccd1 vccd1 HI[6] insts\[6\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[452\] vssd1 vssd1 vccd1 vccd1 HI[452] insts\[452\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[285\] vssd1 vssd1 vccd1 vccd1 HI[285] insts\[285\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[200\] vssd1 vssd1 vccd1 vccd1 HI[200] insts\[200\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_261 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[415\] vssd1 vssd1 vccd1 vccd1 HI[415] insts\[415\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[150\] vssd1 vssd1 vccd1 vccd1 HI[150] insts\[150\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[248\] vssd1 vssd1 vccd1 vccd1 HI[248] insts\[248\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_581 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[30\] vssd1 vssd1 vccd1 vccd1 HI[30] insts\[30\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[365\] vssd1 vssd1 vccd1 vccd1 HI[365] insts\[365\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[198\] vssd1 vssd1 vccd1 vccd1 HI[198] insts\[198\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[78\] vssd1 vssd1 vccd1 vccd1 HI[78] insts\[78\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[113\] vssd1 vssd1 vccd1 vccd1 HI[113] insts\[113\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[230\] vssd1 vssd1 vccd1 vccd1 HI[230] insts\[230\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[328\] vssd1 vssd1 vccd1 vccd1 HI[328] insts\[328\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[445\] vssd1 vssd1 vccd1 vccd1 HI[445] insts\[445\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[278\] vssd1 vssd1 vccd1 vccd1 HI[278] insts\[278\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[180\] vssd1 vssd1 vccd1 vccd1 HI[180] insts\[180\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[60\] vssd1 vssd1 vccd1 vccd1 HI[60] insts\[60\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[395\] vssd1 vssd1 vccd1 vccd1 HI[395] insts\[395\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_273 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[408\] vssd1 vssd1 vccd1 vccd1 HI[408] insts\[408\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[143\] vssd1 vssd1 vccd1 vccd1 HI[143] insts\[143\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[310\] vssd1 vssd1 vccd1 vccd1 HI[310] insts\[310\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[23\] vssd1 vssd1 vccd1 vccd1 HI[23] insts\[23\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[358\] vssd1 vssd1 vccd1 vccd1 HI[358] insts\[358\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[260\] vssd1 vssd1 vccd1 vccd1 HI[260] insts\[260\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[106\] vssd1 vssd1 vccd1 vccd1 HI[106] insts\[106\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[90\] vssd1 vssd1 vccd1 vccd1 HI[90] insts\[90\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[223\] vssd1 vssd1 vccd1 vccd1 HI[223] insts\[223\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[438\] vssd1 vssd1 vccd1 vccd1 HI[438] insts\[438\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[340\] vssd1 vssd1 vccd1 vccd1 HI[340] insts\[340\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[173\] vssd1 vssd1 vccd1 vccd1 HI[173] insts\[173\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[53\] vssd1 vssd1 vccd1 vccd1 HI[53] insts\[53\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[388\] vssd1 vssd1 vccd1 vccd1 HI[388] insts\[388\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[290\] vssd1 vssd1 vccd1 vccd1 HI[290] insts\[290\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_230 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[136\] vssd1 vssd1 vccd1 vccd1 HI[136] insts\[136\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[303\] vssd1 vssd1 vccd1 vccd1 HI[303] insts\[303\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[16\] vssd1 vssd1 vccd1 vccd1 HI[16] insts\[16\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[420\] vssd1 vssd1 vccd1 vccd1 HI[420] insts\[420\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[253\] vssd1 vssd1 vccd1 vccd1 HI[253] insts\[253\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[370\] vssd1 vssd1 vccd1 vccd1 HI[370] insts\[370\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[83\] vssd1 vssd1 vccd1 vccd1 HI[83] insts\[83\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[216\] vssd1 vssd1 vccd1 vccd1 HI[216] insts\[216\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[166\] vssd1 vssd1 vccd1 vccd1 HI[166] insts\[166\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[333\] vssd1 vssd1 vccd1 vccd1 HI[333] insts\[333\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[46\] vssd1 vssd1 vccd1 vccd1 HI[46] insts\[46\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[450\] vssd1 vssd1 vccd1 vccd1 HI[450] insts\[450\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_209 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[283\] vssd1 vssd1 vccd1 vccd1 HI[283] insts\[283\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[4\] vssd1 vssd1 vccd1 vccd1 HI[4] insts\[4\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_710 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_242 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[129\] vssd1 vssd1 vccd1 vccd1 HI[129] insts\[129\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[413\] vssd1 vssd1 vccd1 vccd1 HI[413] insts\[413\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[246\] vssd1 vssd1 vccd1 vccd1 HI[246] insts\[246\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[196\] vssd1 vssd1 vccd1 vccd1 HI[196] insts\[196\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[363\] vssd1 vssd1 vccd1 vccd1 HI[363] insts\[363\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[76\] vssd1 vssd1 vccd1 vccd1 HI[76] insts\[76\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[209\] vssd1 vssd1 vccd1 vccd1 HI[209] insts\[209\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[111\] vssd1 vssd1 vccd1 vccd1 HI[111] insts\[111\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[326\] vssd1 vssd1 vccd1 vccd1 HI[326] insts\[326\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[159\] vssd1 vssd1 vccd1 vccd1 HI[159] insts\[159\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[39\] vssd1 vssd1 vccd1 vccd1 HI[39] insts\[39\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_722 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_8
Xinsts\[443\] vssd1 vssd1 vccd1 vccd1 HI[443] insts\[443\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_221 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_254 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[276\] vssd1 vssd1 vccd1 vccd1 HI[276] insts\[276\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[393\] vssd1 vssd1 vccd1 vccd1 HI[393] insts\[393\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[406\] vssd1 vssd1 vccd1 vccd1 HI[406] insts\[406\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[141\] vssd1 vssd1 vccd1 vccd1 HI[141] insts\[141\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[239\] vssd1 vssd1 vccd1 vccd1 HI[239] insts\[239\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[21\] vssd1 vssd1 vccd1 vccd1 HI[21] insts\[21\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[356\] vssd1 vssd1 vccd1 vccd1 HI[356] insts\[356\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[189\] vssd1 vssd1 vccd1 vccd1 HI[189] insts\[189\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[69\] vssd1 vssd1 vccd1 vccd1 HI[69] insts\[69\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[104\] vssd1 vssd1 vccd1 vccd1 HI[104] insts\[104\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_617 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[221\] vssd1 vssd1 vccd1 vccd1 HI[221] insts\[221\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[319\] vssd1 vssd1 vccd1 vccd1 HI[319] insts\[319\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[436\] vssd1 vssd1 vccd1 vccd1 HI[436] insts\[436\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[171\] vssd1 vssd1 vccd1 vccd1 HI[171] insts\[171\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[269\] vssd1 vssd1 vccd1 vccd1 HI[269] insts\[269\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[51\] vssd1 vssd1 vccd1 vccd1 HI[51] insts\[51\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[386\] vssd1 vssd1 vccd1 vccd1 HI[386] insts\[386\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[99\] vssd1 vssd1 vccd1 vccd1 HI[99] insts\[99\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[134\] vssd1 vssd1 vccd1 vccd1 HI[134] insts\[134\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[301\] vssd1 vssd1 vccd1 vccd1 HI[301] insts\[301\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[14\] vssd1 vssd1 vccd1 vccd1 HI[14] insts\[14\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[349\] vssd1 vssd1 vccd1 vccd1 HI[349] insts\[349\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[251\] vssd1 vssd1 vccd1 vccd1 HI[251] insts\[251\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[299\] vssd1 vssd1 vccd1 vccd1 HI[299] insts\[299\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_629 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_673 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[81\] vssd1 vssd1 vccd1 vccd1 HI[81] insts\[81\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[214\] vssd1 vssd1 vccd1 vccd1 HI[214] insts\[214\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[429\] vssd1 vssd1 vccd1 vccd1 HI[429] insts\[429\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[164\] vssd1 vssd1 vccd1 vccd1 HI[164] insts\[164\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[331\] vssd1 vssd1 vccd1 vccd1 HI[331] insts\[331\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[44\] vssd1 vssd1 vccd1 vccd1 HI[44] insts\[44\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[379\] vssd1 vssd1 vccd1 vccd1 HI[379] insts\[379\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[2\] vssd1 vssd1 vccd1 vccd1 HI[2] insts\[2\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[281\] vssd1 vssd1 vccd1 vccd1 HI[281] insts\[281\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[127\] vssd1 vssd1 vccd1 vccd1 HI[127] insts\[127\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[411\] vssd1 vssd1 vccd1 vccd1 HI[411] insts\[411\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[244\] vssd1 vssd1 vccd1 vccd1 HI[244] insts\[244\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[459\] vssd1 vssd1 vccd1 vccd1 HI[459] insts\[459\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[361\] vssd1 vssd1 vccd1 vccd1 HI[361] insts\[361\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[194\] vssd1 vssd1 vccd1 vccd1 HI[194] insts\[194\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_641 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_685 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[74\] vssd1 vssd1 vccd1 vccd1 HI[74] insts\[74\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_405 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_449 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[207\] vssd1 vssd1 vccd1 vccd1 HI[207] insts\[207\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[157\] vssd1 vssd1 vccd1 vccd1 HI[157] insts\[157\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[324\] vssd1 vssd1 vccd1 vccd1 HI[324] insts\[324\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[37\] vssd1 vssd1 vccd1 vccd1 HI[37] insts\[37\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[441\] vssd1 vssd1 vccd1 vccd1 HI[441] insts\[441\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_533 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[274\] vssd1 vssd1 vccd1 vccd1 HI[274] insts\[274\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[391\] vssd1 vssd1 vccd1 vccd1 HI[391] insts\[391\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[404\] vssd1 vssd1 vccd1 vccd1 HI[404] insts\[404\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[237\] vssd1 vssd1 vccd1 vccd1 HI[237] insts\[237\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_609 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[354\] vssd1 vssd1 vccd1 vccd1 HI[354] insts\[354\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[187\] vssd1 vssd1 vccd1 vccd1 HI[187] insts\[187\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[67\] vssd1 vssd1 vccd1 vccd1 HI[67] insts\[67\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_697 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[102\] vssd1 vssd1 vccd1 vccd1 HI[102] insts\[102\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_417 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[317\] vssd1 vssd1 vccd1 vccd1 HI[317] insts\[317\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[434\] vssd1 vssd1 vccd1 vccd1 HI[434] insts\[434\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_545 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[267\] vssd1 vssd1 vccd1 vccd1 HI[267] insts\[267\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_589 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[384\] vssd1 vssd1 vccd1 vccd1 HI[384] insts\[384\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_386 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[97\] vssd1 vssd1 vccd1 vccd1 HI[97] insts\[97\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[132\] vssd1 vssd1 vccd1 vccd1 HI[132] insts\[132\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[12\] vssd1 vssd1 vccd1 vccd1 HI[12] insts\[12\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[347\] vssd1 vssd1 vccd1 vccd1 HI[347] insts\[347\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_429 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[297\] vssd1 vssd1 vccd1 vccd1 HI[297] insts\[297\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[212\] vssd1 vssd1 vccd1 vccd1 HI[212] insts\[212\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[162\] vssd1 vssd1 vccd1 vccd1 HI[162] insts\[162\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[427\] vssd1 vssd1 vccd1 vccd1 HI[427] insts\[427\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_557 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_502 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[42\] vssd1 vssd1 vccd1 vccd1 HI[42] insts\[42\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[377\] vssd1 vssd1 vccd1 vccd1 HI[377] insts\[377\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_398 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_365 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_321 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[0\] vssd1 vssd1 vccd1 vccd1 HI[0] insts\[0\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[125\] vssd1 vssd1 vccd1 vccd1 HI[125] insts\[125\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[242\] vssd1 vssd1 vccd1 vccd1 HI[242] insts\[242\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[457\] vssd1 vssd1 vccd1 vccd1 HI[457] insts\[457\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[192\] vssd1 vssd1 vccd1 vccd1 HI[192] insts\[192\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[72\] vssd1 vssd1 vccd1 vccd1 HI[72] insts\[72\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[205\] vssd1 vssd1 vccd1 vccd1 HI[205] insts\[205\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_569 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_514 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[155\] vssd1 vssd1 vccd1 vccd1 HI[155] insts\[155\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[322\] vssd1 vssd1 vccd1 vccd1 HI[322] insts\[322\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[35\] vssd1 vssd1 vccd1 vccd1 HI[35] insts\[35\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[272\] vssd1 vssd1 vccd1 vccd1 HI[272] insts\[272\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_377 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_333 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[118\] vssd1 vssd1 vccd1 vccd1 HI[118] insts\[118\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_130 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_141 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[402\] vssd1 vssd1 vccd1 vccd1 HI[402] insts\[402\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[235\] vssd1 vssd1 vccd1 vccd1 HI[235] insts\[235\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_601 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_645 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[352\] vssd1 vssd1 vccd1 vccd1 HI[352] insts\[352\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[185\] vssd1 vssd1 vccd1 vccd1 HI[185] insts\[185\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[65\] vssd1 vssd1 vccd1 vccd1 HI[65] insts\[65\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[100\] vssd1 vssd1 vccd1 vccd1 HI[100] insts\[100\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[148\] vssd1 vssd1 vccd1 vccd1 HI[148] insts\[148\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_526 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[315\] vssd1 vssd1 vccd1 vccd1 HI[315] insts\[315\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[28\] vssd1 vssd1 vccd1 vccd1 HI[28] insts\[28\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[265\] vssd1 vssd1 vccd1 vccd1 HI[265] insts\[265\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[432\] vssd1 vssd1 vccd1 vccd1 HI[432] insts\[432\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_345 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[382\] vssd1 vssd1 vccd1 vccd1 HI[382] insts\[382\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_197 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_153 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[95\] vssd1 vssd1 vccd1 vccd1 HI[95] insts\[95\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[130\] vssd1 vssd1 vccd1 vccd1 HI[130] insts\[130\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[228\] vssd1 vssd1 vccd1 vccd1 HI[228] insts\[228\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_613 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_657 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[10\] vssd1 vssd1 vccd1 vccd1 HI[10] insts\[10\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[178\] vssd1 vssd1 vccd1 vccd1 HI[178] insts\[178\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[345\] vssd1 vssd1 vccd1 vccd1 HI[345] insts\[345\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[58\] vssd1 vssd1 vccd1 vccd1 HI[58] insts\[58\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[462\] vssd1 vssd1 vccd1 vccd1 HI[462] insts\[462\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[295\] vssd1 vssd1 vccd1 vccd1 HI[295] insts\[295\]/LO sky130_fd_sc_hd__conb_1
.ends

.subckt sky130_fd_sc_hvl__conb_1 VGND VNB VPB VPWR HI LO
R0 VGND LO sky130_fd_pr__res_generic_po w=510000u l=45000u
R1 HI VPWR sky130_fd_pr__res_generic_po w=510000u l=45000u
.ends

.subckt sky130_fd_sc_hvl__lsbufhv2lv_1 A VGND VPWR X VPWR_uq0 VGND_uq0 VNB VPB LVPWR
X0 a_30_1337# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X1 VGND_uq0 a_30_1337# a_30_207# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X2 VGND_uq0 a_30_207# a_389_141# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X3 VGND_uq0 a_30_207# a_389_141# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X4 a_389_1337# a_30_1337# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X5 VGND_uq0 a_30_207# a_389_141# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X6 VGND A a_30_1337# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X7 VGND a_30_1337# a_389_1337# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X8 a_389_141# a_30_207# VGND_uq0 VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X9 VGND a_30_1337# a_389_1337# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X10 LVPWR a_389_141# X LVPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X11 VGND_uq0 a_389_141# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X12 a_389_1337# a_30_1337# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X13 LVPWR a_389_1337# a_389_141# LVPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X14 a_30_207# a_30_1337# VPWR_uq0 VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X15 a_389_1337# a_389_141# LVPWR LVPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
.ends

.subckt mgmt_protect_hv vccd vssd vdda1 vdda2 mprj2_vdd_logic1 mprj_vdd_logic1 dw_6116_1496#
+ vssa1 dw_13698_1476# vssa2
Xmprj2_logic_high_hvl vssa2 vssa2 vdda2 vdda2 mprj2_logic_high_lv/A mprj2_logic_high_hvl/LO
+ sky130_fd_sc_hvl__conb_1
Xmprj_logic_high_hvl vssa1 vssa1 vdda1 vdda1 mprj_logic_high_lv/A mprj_logic_high_hvl/LO
+ sky130_fd_sc_hvl__conb_1
Xmprj_logic_high_lv mprj_logic_high_lv/A vssd vdda1 mprj_vdd_logic1 vdda1 vssd vssd
+ vdda1 vccd sky130_fd_sc_hvl__lsbufhv2lv_1
Xmprj2_logic_high_lv mprj2_logic_high_lv/A vssd vdda2 mprj2_vdd_logic1 vdda2 vssd
+ vssd vdda2 vccd sky130_fd_sc_hvl__lsbufhv2lv_1
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for mgmt_protect abstract view
.subckt mgmt_protect caravel_clk caravel_clk2 caravel_rstn la_data_in_core[0] la_data_in_core[100]
+ la_data_in_core[101] la_data_in_core[102] la_data_in_core[103] la_data_in_core[104]
+ la_data_in_core[105] la_data_in_core[106] la_data_in_core[107] la_data_in_core[108]
+ la_data_in_core[109] la_data_in_core[10] la_data_in_core[110] la_data_in_core[111]
+ la_data_in_core[112] la_data_in_core[113] la_data_in_core[114] la_data_in_core[115]
+ la_data_in_core[116] la_data_in_core[117] la_data_in_core[118] la_data_in_core[119]
+ la_data_in_core[11] la_data_in_core[120] la_data_in_core[121] la_data_in_core[122]
+ la_data_in_core[123] la_data_in_core[124] la_data_in_core[125] la_data_in_core[126]
+ la_data_in_core[127] la_data_in_core[12] la_data_in_core[13] la_data_in_core[14]
+ la_data_in_core[15] la_data_in_core[16] la_data_in_core[17] la_data_in_core[18]
+ la_data_in_core[19] la_data_in_core[1] la_data_in_core[20] la_data_in_core[21] la_data_in_core[22]
+ la_data_in_core[23] la_data_in_core[24] la_data_in_core[25] la_data_in_core[26]
+ la_data_in_core[27] la_data_in_core[28] la_data_in_core[29] la_data_in_core[2] la_data_in_core[30]
+ la_data_in_core[31] la_data_in_core[32] la_data_in_core[33] la_data_in_core[34]
+ la_data_in_core[35] la_data_in_core[36] la_data_in_core[37] la_data_in_core[38]
+ la_data_in_core[39] la_data_in_core[3] la_data_in_core[40] la_data_in_core[41] la_data_in_core[42]
+ la_data_in_core[43] la_data_in_core[44] la_data_in_core[45] la_data_in_core[46]
+ la_data_in_core[47] la_data_in_core[48] la_data_in_core[49] la_data_in_core[4] la_data_in_core[50]
+ la_data_in_core[51] la_data_in_core[52] la_data_in_core[53] la_data_in_core[54]
+ la_data_in_core[55] la_data_in_core[56] la_data_in_core[57] la_data_in_core[58]
+ la_data_in_core[59] la_data_in_core[5] la_data_in_core[60] la_data_in_core[61] la_data_in_core[62]
+ la_data_in_core[63] la_data_in_core[64] la_data_in_core[65] la_data_in_core[66]
+ la_data_in_core[67] la_data_in_core[68] la_data_in_core[69] la_data_in_core[6] la_data_in_core[70]
+ la_data_in_core[71] la_data_in_core[72] la_data_in_core[73] la_data_in_core[74]
+ la_data_in_core[75] la_data_in_core[76] la_data_in_core[77] la_data_in_core[78]
+ la_data_in_core[79] la_data_in_core[7] la_data_in_core[80] la_data_in_core[81] la_data_in_core[82]
+ la_data_in_core[83] la_data_in_core[84] la_data_in_core[85] la_data_in_core[86]
+ la_data_in_core[87] la_data_in_core[88] la_data_in_core[89] la_data_in_core[8] la_data_in_core[90]
+ la_data_in_core[91] la_data_in_core[92] la_data_in_core[93] la_data_in_core[94]
+ la_data_in_core[95] la_data_in_core[96] la_data_in_core[97] la_data_in_core[98]
+ la_data_in_core[99] la_data_in_core[9] la_data_in_mprj[0] la_data_in_mprj[100] la_data_in_mprj[101]
+ la_data_in_mprj[102] la_data_in_mprj[103] la_data_in_mprj[104] la_data_in_mprj[105]
+ la_data_in_mprj[106] la_data_in_mprj[107] la_data_in_mprj[108] la_data_in_mprj[109]
+ la_data_in_mprj[10] la_data_in_mprj[110] la_data_in_mprj[111] la_data_in_mprj[112]
+ la_data_in_mprj[113] la_data_in_mprj[114] la_data_in_mprj[115] la_data_in_mprj[116]
+ la_data_in_mprj[117] la_data_in_mprj[118] la_data_in_mprj[119] la_data_in_mprj[11]
+ la_data_in_mprj[120] la_data_in_mprj[121] la_data_in_mprj[122] la_data_in_mprj[123]
+ la_data_in_mprj[124] la_data_in_mprj[125] la_data_in_mprj[126] la_data_in_mprj[127]
+ la_data_in_mprj[12] la_data_in_mprj[13] la_data_in_mprj[14] la_data_in_mprj[15]
+ la_data_in_mprj[16] la_data_in_mprj[17] la_data_in_mprj[18] la_data_in_mprj[19]
+ la_data_in_mprj[1] la_data_in_mprj[20] la_data_in_mprj[21] la_data_in_mprj[22] la_data_in_mprj[23]
+ la_data_in_mprj[24] la_data_in_mprj[25] la_data_in_mprj[26] la_data_in_mprj[27]
+ la_data_in_mprj[28] la_data_in_mprj[29] la_data_in_mprj[2] la_data_in_mprj[30] la_data_in_mprj[31]
+ la_data_in_mprj[32] la_data_in_mprj[33] la_data_in_mprj[34] la_data_in_mprj[35]
+ la_data_in_mprj[36] la_data_in_mprj[37] la_data_in_mprj[38] la_data_in_mprj[39]
+ la_data_in_mprj[3] la_data_in_mprj[40] la_data_in_mprj[41] la_data_in_mprj[42] la_data_in_mprj[43]
+ la_data_in_mprj[44] la_data_in_mprj[45] la_data_in_mprj[46] la_data_in_mprj[47]
+ la_data_in_mprj[48] la_data_in_mprj[49] la_data_in_mprj[4] la_data_in_mprj[50] la_data_in_mprj[51]
+ la_data_in_mprj[52] la_data_in_mprj[53] la_data_in_mprj[54] la_data_in_mprj[55]
+ la_data_in_mprj[56] la_data_in_mprj[57] la_data_in_mprj[58] la_data_in_mprj[59]
+ la_data_in_mprj[5] la_data_in_mprj[60] la_data_in_mprj[61] la_data_in_mprj[62] la_data_in_mprj[63]
+ la_data_in_mprj[64] la_data_in_mprj[65] la_data_in_mprj[66] la_data_in_mprj[67]
+ la_data_in_mprj[68] la_data_in_mprj[69] la_data_in_mprj[6] la_data_in_mprj[70] la_data_in_mprj[71]
+ la_data_in_mprj[72] la_data_in_mprj[73] la_data_in_mprj[74] la_data_in_mprj[75]
+ la_data_in_mprj[76] la_data_in_mprj[77] la_data_in_mprj[78] la_data_in_mprj[79]
+ la_data_in_mprj[7] la_data_in_mprj[80] la_data_in_mprj[81] la_data_in_mprj[82] la_data_in_mprj[83]
+ la_data_in_mprj[84] la_data_in_mprj[85] la_data_in_mprj[86] la_data_in_mprj[87]
+ la_data_in_mprj[88] la_data_in_mprj[89] la_data_in_mprj[8] la_data_in_mprj[90] la_data_in_mprj[91]
+ la_data_in_mprj[92] la_data_in_mprj[93] la_data_in_mprj[94] la_data_in_mprj[95]
+ la_data_in_mprj[96] la_data_in_mprj[97] la_data_in_mprj[98] la_data_in_mprj[99]
+ la_data_in_mprj[9] la_data_out_core[0] la_data_out_core[100] la_data_out_core[101]
+ la_data_out_core[102] la_data_out_core[103] la_data_out_core[104] la_data_out_core[105]
+ la_data_out_core[106] la_data_out_core[107] la_data_out_core[108] la_data_out_core[109]
+ la_data_out_core[10] la_data_out_core[110] la_data_out_core[111] la_data_out_core[112]
+ la_data_out_core[113] la_data_out_core[114] la_data_out_core[115] la_data_out_core[116]
+ la_data_out_core[117] la_data_out_core[118] la_data_out_core[119] la_data_out_core[11]
+ la_data_out_core[120] la_data_out_core[121] la_data_out_core[122] la_data_out_core[123]
+ la_data_out_core[124] la_data_out_core[125] la_data_out_core[126] la_data_out_core[127]
+ la_data_out_core[12] la_data_out_core[13] la_data_out_core[14] la_data_out_core[15]
+ la_data_out_core[16] la_data_out_core[17] la_data_out_core[18] la_data_out_core[19]
+ la_data_out_core[1] la_data_out_core[20] la_data_out_core[21] la_data_out_core[22]
+ la_data_out_core[23] la_data_out_core[24] la_data_out_core[25] la_data_out_core[26]
+ la_data_out_core[27] la_data_out_core[28] la_data_out_core[29] la_data_out_core[2]
+ la_data_out_core[30] la_data_out_core[31] la_data_out_core[32] la_data_out_core[33]
+ la_data_out_core[34] la_data_out_core[35] la_data_out_core[36] la_data_out_core[37]
+ la_data_out_core[38] la_data_out_core[39] la_data_out_core[3] la_data_out_core[40]
+ la_data_out_core[41] la_data_out_core[42] la_data_out_core[43] la_data_out_core[44]
+ la_data_out_core[45] la_data_out_core[46] la_data_out_core[47] la_data_out_core[48]
+ la_data_out_core[49] la_data_out_core[4] la_data_out_core[50] la_data_out_core[51]
+ la_data_out_core[52] la_data_out_core[53] la_data_out_core[54] la_data_out_core[55]
+ la_data_out_core[56] la_data_out_core[57] la_data_out_core[58] la_data_out_core[59]
+ la_data_out_core[5] la_data_out_core[60] la_data_out_core[61] la_data_out_core[62]
+ la_data_out_core[63] la_data_out_core[64] la_data_out_core[65] la_data_out_core[66]
+ la_data_out_core[67] la_data_out_core[68] la_data_out_core[69] la_data_out_core[6]
+ la_data_out_core[70] la_data_out_core[71] la_data_out_core[72] la_data_out_core[73]
+ la_data_out_core[74] la_data_out_core[75] la_data_out_core[76] la_data_out_core[77]
+ la_data_out_core[78] la_data_out_core[79] la_data_out_core[7] la_data_out_core[80]
+ la_data_out_core[81] la_data_out_core[82] la_data_out_core[83] la_data_out_core[84]
+ la_data_out_core[85] la_data_out_core[86] la_data_out_core[87] la_data_out_core[88]
+ la_data_out_core[89] la_data_out_core[8] la_data_out_core[90] la_data_out_core[91]
+ la_data_out_core[92] la_data_out_core[93] la_data_out_core[94] la_data_out_core[95]
+ la_data_out_core[96] la_data_out_core[97] la_data_out_core[98] la_data_out_core[99]
+ la_data_out_core[9] la_data_out_mprj[0] la_data_out_mprj[100] la_data_out_mprj[101]
+ la_data_out_mprj[102] la_data_out_mprj[103] la_data_out_mprj[104] la_data_out_mprj[105]
+ la_data_out_mprj[106] la_data_out_mprj[107] la_data_out_mprj[108] la_data_out_mprj[109]
+ la_data_out_mprj[10] la_data_out_mprj[110] la_data_out_mprj[111] la_data_out_mprj[112]
+ la_data_out_mprj[113] la_data_out_mprj[114] la_data_out_mprj[115] la_data_out_mprj[116]
+ la_data_out_mprj[117] la_data_out_mprj[118] la_data_out_mprj[119] la_data_out_mprj[11]
+ la_data_out_mprj[120] la_data_out_mprj[121] la_data_out_mprj[122] la_data_out_mprj[123]
+ la_data_out_mprj[124] la_data_out_mprj[125] la_data_out_mprj[126] la_data_out_mprj[127]
+ la_data_out_mprj[12] la_data_out_mprj[13] la_data_out_mprj[14] la_data_out_mprj[15]
+ la_data_out_mprj[16] la_data_out_mprj[17] la_data_out_mprj[18] la_data_out_mprj[19]
+ la_data_out_mprj[1] la_data_out_mprj[20] la_data_out_mprj[21] la_data_out_mprj[22]
+ la_data_out_mprj[23] la_data_out_mprj[24] la_data_out_mprj[25] la_data_out_mprj[26]
+ la_data_out_mprj[27] la_data_out_mprj[28] la_data_out_mprj[29] la_data_out_mprj[2]
+ la_data_out_mprj[30] la_data_out_mprj[31] la_data_out_mprj[32] la_data_out_mprj[33]
+ la_data_out_mprj[34] la_data_out_mprj[35] la_data_out_mprj[36] la_data_out_mprj[37]
+ la_data_out_mprj[38] la_data_out_mprj[39] la_data_out_mprj[3] la_data_out_mprj[40]
+ la_data_out_mprj[41] la_data_out_mprj[42] la_data_out_mprj[43] la_data_out_mprj[44]
+ la_data_out_mprj[45] la_data_out_mprj[46] la_data_out_mprj[47] la_data_out_mprj[48]
+ la_data_out_mprj[49] la_data_out_mprj[4] la_data_out_mprj[50] la_data_out_mprj[51]
+ la_data_out_mprj[52] la_data_out_mprj[53] la_data_out_mprj[54] la_data_out_mprj[55]
+ la_data_out_mprj[56] la_data_out_mprj[57] la_data_out_mprj[58] la_data_out_mprj[59]
+ la_data_out_mprj[5] la_data_out_mprj[60] la_data_out_mprj[61] la_data_out_mprj[62]
+ la_data_out_mprj[63] la_data_out_mprj[64] la_data_out_mprj[65] la_data_out_mprj[66]
+ la_data_out_mprj[67] la_data_out_mprj[68] la_data_out_mprj[69] la_data_out_mprj[6]
+ la_data_out_mprj[70] la_data_out_mprj[71] la_data_out_mprj[72] la_data_out_mprj[73]
+ la_data_out_mprj[74] la_data_out_mprj[75] la_data_out_mprj[76] la_data_out_mprj[77]
+ la_data_out_mprj[78] la_data_out_mprj[79] la_data_out_mprj[7] la_data_out_mprj[80]
+ la_data_out_mprj[81] la_data_out_mprj[82] la_data_out_mprj[83] la_data_out_mprj[84]
+ la_data_out_mprj[85] la_data_out_mprj[86] la_data_out_mprj[87] la_data_out_mprj[88]
+ la_data_out_mprj[89] la_data_out_mprj[8] la_data_out_mprj[90] la_data_out_mprj[91]
+ la_data_out_mprj[92] la_data_out_mprj[93] la_data_out_mprj[94] la_data_out_mprj[95]
+ la_data_out_mprj[96] la_data_out_mprj[97] la_data_out_mprj[98] la_data_out_mprj[99]
+ la_data_out_mprj[9] la_iena_mprj[0] la_iena_mprj[100] la_iena_mprj[101] la_iena_mprj[102]
+ la_iena_mprj[103] la_iena_mprj[104] la_iena_mprj[105] la_iena_mprj[106] la_iena_mprj[107]
+ la_iena_mprj[108] la_iena_mprj[109] la_iena_mprj[10] la_iena_mprj[110] la_iena_mprj[111]
+ la_iena_mprj[112] la_iena_mprj[113] la_iena_mprj[114] la_iena_mprj[115] la_iena_mprj[116]
+ la_iena_mprj[117] la_iena_mprj[118] la_iena_mprj[119] la_iena_mprj[11] la_iena_mprj[120]
+ la_iena_mprj[121] la_iena_mprj[122] la_iena_mprj[123] la_iena_mprj[124] la_iena_mprj[125]
+ la_iena_mprj[126] la_iena_mprj[127] la_iena_mprj[12] la_iena_mprj[13] la_iena_mprj[14]
+ la_iena_mprj[15] la_iena_mprj[16] la_iena_mprj[17] la_iena_mprj[18] la_iena_mprj[19]
+ la_iena_mprj[1] la_iena_mprj[20] la_iena_mprj[21] la_iena_mprj[22] la_iena_mprj[23]
+ la_iena_mprj[24] la_iena_mprj[25] la_iena_mprj[26] la_iena_mprj[27] la_iena_mprj[28]
+ la_iena_mprj[29] la_iena_mprj[2] la_iena_mprj[30] la_iena_mprj[31] la_iena_mprj[32]
+ la_iena_mprj[33] la_iena_mprj[34] la_iena_mprj[35] la_iena_mprj[36] la_iena_mprj[37]
+ la_iena_mprj[38] la_iena_mprj[39] la_iena_mprj[3] la_iena_mprj[40] la_iena_mprj[41]
+ la_iena_mprj[42] la_iena_mprj[43] la_iena_mprj[44] la_iena_mprj[45] la_iena_mprj[46]
+ la_iena_mprj[47] la_iena_mprj[48] la_iena_mprj[49] la_iena_mprj[4] la_iena_mprj[50]
+ la_iena_mprj[51] la_iena_mprj[52] la_iena_mprj[53] la_iena_mprj[54] la_iena_mprj[55]
+ la_iena_mprj[56] la_iena_mprj[57] la_iena_mprj[58] la_iena_mprj[59] la_iena_mprj[5]
+ la_iena_mprj[60] la_iena_mprj[61] la_iena_mprj[62] la_iena_mprj[63] la_iena_mprj[64]
+ la_iena_mprj[65] la_iena_mprj[66] la_iena_mprj[67] la_iena_mprj[68] la_iena_mprj[69]
+ la_iena_mprj[6] la_iena_mprj[70] la_iena_mprj[71] la_iena_mprj[72] la_iena_mprj[73]
+ la_iena_mprj[74] la_iena_mprj[75] la_iena_mprj[76] la_iena_mprj[77] la_iena_mprj[78]
+ la_iena_mprj[79] la_iena_mprj[7] la_iena_mprj[80] la_iena_mprj[81] la_iena_mprj[82]
+ la_iena_mprj[83] la_iena_mprj[84] la_iena_mprj[85] la_iena_mprj[86] la_iena_mprj[87]
+ la_iena_mprj[88] la_iena_mprj[89] la_iena_mprj[8] la_iena_mprj[90] la_iena_mprj[91]
+ la_iena_mprj[92] la_iena_mprj[93] la_iena_mprj[94] la_iena_mprj[95] la_iena_mprj[96]
+ la_iena_mprj[97] la_iena_mprj[98] la_iena_mprj[99] la_iena_mprj[9] la_oenb_core[0]
+ la_oenb_core[100] la_oenb_core[101] la_oenb_core[102] la_oenb_core[103] la_oenb_core[104]
+ la_oenb_core[105] la_oenb_core[106] la_oenb_core[107] la_oenb_core[108] la_oenb_core[109]
+ la_oenb_core[10] la_oenb_core[110] la_oenb_core[111] la_oenb_core[112] la_oenb_core[113]
+ la_oenb_core[114] la_oenb_core[115] la_oenb_core[116] la_oenb_core[117] la_oenb_core[118]
+ la_oenb_core[119] la_oenb_core[11] la_oenb_core[120] la_oenb_core[121] la_oenb_core[122]
+ la_oenb_core[123] la_oenb_core[124] la_oenb_core[125] la_oenb_core[126] la_oenb_core[127]
+ la_oenb_core[12] la_oenb_core[13] la_oenb_core[14] la_oenb_core[15] la_oenb_core[16]
+ la_oenb_core[17] la_oenb_core[18] la_oenb_core[19] la_oenb_core[1] la_oenb_core[20]
+ la_oenb_core[21] la_oenb_core[22] la_oenb_core[23] la_oenb_core[24] la_oenb_core[25]
+ la_oenb_core[26] la_oenb_core[27] la_oenb_core[28] la_oenb_core[29] la_oenb_core[2]
+ la_oenb_core[30] la_oenb_core[31] la_oenb_core[32] la_oenb_core[33] la_oenb_core[34]
+ la_oenb_core[35] la_oenb_core[36] la_oenb_core[37] la_oenb_core[38] la_oenb_core[39]
+ la_oenb_core[3] la_oenb_core[40] la_oenb_core[41] la_oenb_core[42] la_oenb_core[43]
+ la_oenb_core[44] la_oenb_core[45] la_oenb_core[46] la_oenb_core[47] la_oenb_core[48]
+ la_oenb_core[49] la_oenb_core[4] la_oenb_core[50] la_oenb_core[51] la_oenb_core[52]
+ la_oenb_core[53] la_oenb_core[54] la_oenb_core[55] la_oenb_core[56] la_oenb_core[57]
+ la_oenb_core[58] la_oenb_core[59] la_oenb_core[5] la_oenb_core[60] la_oenb_core[61]
+ la_oenb_core[62] la_oenb_core[63] la_oenb_core[64] la_oenb_core[65] la_oenb_core[66]
+ la_oenb_core[67] la_oenb_core[68] la_oenb_core[69] la_oenb_core[6] la_oenb_core[70]
+ la_oenb_core[71] la_oenb_core[72] la_oenb_core[73] la_oenb_core[74] la_oenb_core[75]
+ la_oenb_core[76] la_oenb_core[77] la_oenb_core[78] la_oenb_core[79] la_oenb_core[7]
+ la_oenb_core[80] la_oenb_core[81] la_oenb_core[82] la_oenb_core[83] la_oenb_core[84]
+ la_oenb_core[85] la_oenb_core[86] la_oenb_core[87] la_oenb_core[88] la_oenb_core[89]
+ la_oenb_core[8] la_oenb_core[90] la_oenb_core[91] la_oenb_core[92] la_oenb_core[93]
+ la_oenb_core[94] la_oenb_core[95] la_oenb_core[96] la_oenb_core[97] la_oenb_core[98]
+ la_oenb_core[99] la_oenb_core[9] la_oenb_mprj[0] la_oenb_mprj[100] la_oenb_mprj[101]
+ la_oenb_mprj[102] la_oenb_mprj[103] la_oenb_mprj[104] la_oenb_mprj[105] la_oenb_mprj[106]
+ la_oenb_mprj[107] la_oenb_mprj[108] la_oenb_mprj[109] la_oenb_mprj[10] la_oenb_mprj[110]
+ la_oenb_mprj[111] la_oenb_mprj[112] la_oenb_mprj[113] la_oenb_mprj[114] la_oenb_mprj[115]
+ la_oenb_mprj[116] la_oenb_mprj[117] la_oenb_mprj[118] la_oenb_mprj[119] la_oenb_mprj[11]
+ la_oenb_mprj[120] la_oenb_mprj[121] la_oenb_mprj[122] la_oenb_mprj[123] la_oenb_mprj[124]
+ la_oenb_mprj[125] la_oenb_mprj[126] la_oenb_mprj[127] la_oenb_mprj[12] la_oenb_mprj[13]
+ la_oenb_mprj[14] la_oenb_mprj[15] la_oenb_mprj[16] la_oenb_mprj[17] la_oenb_mprj[18]
+ la_oenb_mprj[19] la_oenb_mprj[1] la_oenb_mprj[20] la_oenb_mprj[21] la_oenb_mprj[22]
+ la_oenb_mprj[23] la_oenb_mprj[24] la_oenb_mprj[25] la_oenb_mprj[26] la_oenb_mprj[27]
+ la_oenb_mprj[28] la_oenb_mprj[29] la_oenb_mprj[2] la_oenb_mprj[30] la_oenb_mprj[31]
+ la_oenb_mprj[32] la_oenb_mprj[33] la_oenb_mprj[34] la_oenb_mprj[35] la_oenb_mprj[36]
+ la_oenb_mprj[37] la_oenb_mprj[38] la_oenb_mprj[39] la_oenb_mprj[3] la_oenb_mprj[40]
+ la_oenb_mprj[41] la_oenb_mprj[42] la_oenb_mprj[43] la_oenb_mprj[44] la_oenb_mprj[45]
+ la_oenb_mprj[46] la_oenb_mprj[47] la_oenb_mprj[48] la_oenb_mprj[49] la_oenb_mprj[4]
+ la_oenb_mprj[50] la_oenb_mprj[51] la_oenb_mprj[52] la_oenb_mprj[53] la_oenb_mprj[54]
+ la_oenb_mprj[55] la_oenb_mprj[56] la_oenb_mprj[57] la_oenb_mprj[58] la_oenb_mprj[59]
+ la_oenb_mprj[5] la_oenb_mprj[60] la_oenb_mprj[61] la_oenb_mprj[62] la_oenb_mprj[63]
+ la_oenb_mprj[64] la_oenb_mprj[65] la_oenb_mprj[66] la_oenb_mprj[67] la_oenb_mprj[68]
+ la_oenb_mprj[69] la_oenb_mprj[6] la_oenb_mprj[70] la_oenb_mprj[71] la_oenb_mprj[72]
+ la_oenb_mprj[73] la_oenb_mprj[74] la_oenb_mprj[75] la_oenb_mprj[76] la_oenb_mprj[77]
+ la_oenb_mprj[78] la_oenb_mprj[79] la_oenb_mprj[7] la_oenb_mprj[80] la_oenb_mprj[81]
+ la_oenb_mprj[82] la_oenb_mprj[83] la_oenb_mprj[84] la_oenb_mprj[85] la_oenb_mprj[86]
+ la_oenb_mprj[87] la_oenb_mprj[88] la_oenb_mprj[89] la_oenb_mprj[8] la_oenb_mprj[90]
+ la_oenb_mprj[91] la_oenb_mprj[92] la_oenb_mprj[93] la_oenb_mprj[94] la_oenb_mprj[95]
+ la_oenb_mprj[96] la_oenb_mprj[97] la_oenb_mprj[98] la_oenb_mprj[99] la_oenb_mprj[9]
+ mprj_ack_i_core mprj_ack_i_user mprj_adr_o_core[0] mprj_adr_o_core[10] mprj_adr_o_core[11]
+ mprj_adr_o_core[12] mprj_adr_o_core[13] mprj_adr_o_core[14] mprj_adr_o_core[15]
+ mprj_adr_o_core[16] mprj_adr_o_core[17] mprj_adr_o_core[18] mprj_adr_o_core[19]
+ mprj_adr_o_core[1] mprj_adr_o_core[20] mprj_adr_o_core[21] mprj_adr_o_core[22] mprj_adr_o_core[23]
+ mprj_adr_o_core[24] mprj_adr_o_core[25] mprj_adr_o_core[26] mprj_adr_o_core[27]
+ mprj_adr_o_core[28] mprj_adr_o_core[29] mprj_adr_o_core[2] mprj_adr_o_core[30] mprj_adr_o_core[31]
+ mprj_adr_o_core[3] mprj_adr_o_core[4] mprj_adr_o_core[5] mprj_adr_o_core[6] mprj_adr_o_core[7]
+ mprj_adr_o_core[8] mprj_adr_o_core[9] mprj_adr_o_user[0] mprj_adr_o_user[10] mprj_adr_o_user[11]
+ mprj_adr_o_user[12] mprj_adr_o_user[13] mprj_adr_o_user[14] mprj_adr_o_user[15]
+ mprj_adr_o_user[16] mprj_adr_o_user[17] mprj_adr_o_user[18] mprj_adr_o_user[19]
+ mprj_adr_o_user[1] mprj_adr_o_user[20] mprj_adr_o_user[21] mprj_adr_o_user[22] mprj_adr_o_user[23]
+ mprj_adr_o_user[24] mprj_adr_o_user[25] mprj_adr_o_user[26] mprj_adr_o_user[27]
+ mprj_adr_o_user[28] mprj_adr_o_user[29] mprj_adr_o_user[2] mprj_adr_o_user[30] mprj_adr_o_user[31]
+ mprj_adr_o_user[3] mprj_adr_o_user[4] mprj_adr_o_user[5] mprj_adr_o_user[6] mprj_adr_o_user[7]
+ mprj_adr_o_user[8] mprj_adr_o_user[9] mprj_cyc_o_core mprj_cyc_o_user mprj_dat_i_core[0]
+ mprj_dat_i_core[10] mprj_dat_i_core[11] mprj_dat_i_core[12] mprj_dat_i_core[13]
+ mprj_dat_i_core[14] mprj_dat_i_core[15] mprj_dat_i_core[16] mprj_dat_i_core[17]
+ mprj_dat_i_core[18] mprj_dat_i_core[19] mprj_dat_i_core[1] mprj_dat_i_core[20] mprj_dat_i_core[21]
+ mprj_dat_i_core[22] mprj_dat_i_core[23] mprj_dat_i_core[24] mprj_dat_i_core[25]
+ mprj_dat_i_core[26] mprj_dat_i_core[27] mprj_dat_i_core[28] mprj_dat_i_core[29]
+ mprj_dat_i_core[2] mprj_dat_i_core[30] mprj_dat_i_core[31] mprj_dat_i_core[3] mprj_dat_i_core[4]
+ mprj_dat_i_core[5] mprj_dat_i_core[6] mprj_dat_i_core[7] mprj_dat_i_core[8] mprj_dat_i_core[9]
+ mprj_dat_i_user[0] mprj_dat_i_user[10] mprj_dat_i_user[11] mprj_dat_i_user[12] mprj_dat_i_user[13]
+ mprj_dat_i_user[14] mprj_dat_i_user[15] mprj_dat_i_user[16] mprj_dat_i_user[17]
+ mprj_dat_i_user[18] mprj_dat_i_user[19] mprj_dat_i_user[1] mprj_dat_i_user[20] mprj_dat_i_user[21]
+ mprj_dat_i_user[22] mprj_dat_i_user[23] mprj_dat_i_user[24] mprj_dat_i_user[25]
+ mprj_dat_i_user[26] mprj_dat_i_user[27] mprj_dat_i_user[28] mprj_dat_i_user[29]
+ mprj_dat_i_user[2] mprj_dat_i_user[30] mprj_dat_i_user[31] mprj_dat_i_user[3] mprj_dat_i_user[4]
+ mprj_dat_i_user[5] mprj_dat_i_user[6] mprj_dat_i_user[7] mprj_dat_i_user[8] mprj_dat_i_user[9]
+ mprj_dat_o_core[0] mprj_dat_o_core[10] mprj_dat_o_core[11] mprj_dat_o_core[12] mprj_dat_o_core[13]
+ mprj_dat_o_core[14] mprj_dat_o_core[15] mprj_dat_o_core[16] mprj_dat_o_core[17]
+ mprj_dat_o_core[18] mprj_dat_o_core[19] mprj_dat_o_core[1] mprj_dat_o_core[20] mprj_dat_o_core[21]
+ mprj_dat_o_core[22] mprj_dat_o_core[23] mprj_dat_o_core[24] mprj_dat_o_core[25]
+ mprj_dat_o_core[26] mprj_dat_o_core[27] mprj_dat_o_core[28] mprj_dat_o_core[29]
+ mprj_dat_o_core[2] mprj_dat_o_core[30] mprj_dat_o_core[31] mprj_dat_o_core[3] mprj_dat_o_core[4]
+ mprj_dat_o_core[5] mprj_dat_o_core[6] mprj_dat_o_core[7] mprj_dat_o_core[8] mprj_dat_o_core[9]
+ mprj_dat_o_user[0] mprj_dat_o_user[10] mprj_dat_o_user[11] mprj_dat_o_user[12] mprj_dat_o_user[13]
+ mprj_dat_o_user[14] mprj_dat_o_user[15] mprj_dat_o_user[16] mprj_dat_o_user[17]
+ mprj_dat_o_user[18] mprj_dat_o_user[19] mprj_dat_o_user[1] mprj_dat_o_user[20] mprj_dat_o_user[21]
+ mprj_dat_o_user[22] mprj_dat_o_user[23] mprj_dat_o_user[24] mprj_dat_o_user[25]
+ mprj_dat_o_user[26] mprj_dat_o_user[27] mprj_dat_o_user[28] mprj_dat_o_user[29]
+ mprj_dat_o_user[2] mprj_dat_o_user[30] mprj_dat_o_user[31] mprj_dat_o_user[3] mprj_dat_o_user[4]
+ mprj_dat_o_user[5] mprj_dat_o_user[6] mprj_dat_o_user[7] mprj_dat_o_user[8] mprj_dat_o_user[9]
+ mprj_iena_wb mprj_sel_o_core[0] mprj_sel_o_core[1] mprj_sel_o_core[2] mprj_sel_o_core[3]
+ mprj_sel_o_user[0] mprj_sel_o_user[1] mprj_sel_o_user[2] mprj_sel_o_user[3] mprj_stb_o_core
+ mprj_stb_o_user mprj_we_o_core mprj_we_o_user user1_vcc_powergood user1_vdd_powergood
+ user2_vcc_powergood user2_vdd_powergood user_clock user_clock2 user_irq[0] user_irq[1]
+ user_irq[2] user_irq_core[0] user_irq_core[1] user_irq_core[2] user_irq_ena[0] user_irq_ena[1]
+ user_irq_ena[2] user_reset vccd vccd1 vccd2 vdda1 vdda2 vssa1 vssa2 vssd vssd1 vssd2
.ends

* Black-box entry subcircuit for sky130_fd_sc_hvl__decap_4 abstract view
.subckt sky130_fd_sc_hvl__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hvl__decap_8 abstract view
.subckt sky130_fd_sc_hvl__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hvl__fill_2#0 abstract view
.subckt sky130_fd_sc_hvl__fill_2#0 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hvl__fill_1#0 abstract view
.subckt sky130_fd_sc_hvl__fill_1#0 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hvl__diode_2 abstract view
.subckt sky130_fd_sc_hvl__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hvl__lsbufhv2lv_1#0 abstract view
.subckt sky130_fd_sc_hvl__lsbufhv2lv_1#0 A LVPWR VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for xres_buf abstract view
.subckt xres_buf A X VPWR VGND LVPWR LVGND
.ends

* Black-box entry subcircuit for copyright_block_a abstract view
.subckt copyright_block_a
.ends

* Black-box entry subcircuit for caravan_power_routing abstract view
.subckt caravan_power_routing
.ends

* Black-box entry subcircuit for user_analog_project_wrapper abstract view
.subckt user_analog_project_wrapper gpio_analog[0] gpio_analog[10] gpio_analog[11]
+ gpio_analog[12] gpio_analog[13] gpio_analog[14] gpio_analog[15] gpio_analog[16]
+ gpio_analog[17] gpio_analog[1] gpio_analog[2] gpio_analog[3] gpio_analog[4] gpio_analog[5]
+ gpio_analog[6] gpio_analog[7] gpio_analog[8] gpio_analog[9] gpio_noesd[0] gpio_noesd[10]
+ gpio_noesd[11] gpio_noesd[12] gpio_noesd[13] gpio_noesd[14] gpio_noesd[15] gpio_noesd[16]
+ gpio_noesd[17] gpio_noesd[1] gpio_noesd[2] gpio_noesd[3] gpio_noesd[4] gpio_noesd[5]
+ gpio_noesd[6] gpio_noesd[7] gpio_noesd[8] gpio_noesd[9] io_analog[0] io_analog[10]
+ io_analog[1] io_analog[2] io_analog[3] io_analog[7] io_analog[8] io_analog[9] io_analog[4]
+ io_analog[5] io_analog[6] io_clamp_high[0] io_clamp_high[1] io_clamp_high[2] io_clamp_low[0]
+ io_clamp_low[1] io_clamp_low[2] io_in[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21]
+ io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_in[8] io_in[9] io_in_3v3[0] io_in_3v3[10] io_in_3v3[11] io_in_3v3[12]
+ io_in_3v3[13] io_in_3v3[14] io_in_3v3[15] io_in_3v3[16] io_in_3v3[17] io_in_3v3[18]
+ io_in_3v3[19] io_in_3v3[1] io_in_3v3[20] io_in_3v3[21] io_in_3v3[22] io_in_3v3[23]
+ io_in_3v3[24] io_in_3v3[25] io_in_3v3[26] io_in_3v3[2] io_in_3v3[3] io_in_3v3[4]
+ io_in_3v3[5] io_in_3v3[6] io_in_3v3[7] io_in_3v3[8] io_in_3v3[9] io_oeb[0] io_oeb[10]
+ io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18]
+ io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25]
+ io_oeb[26] io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8]
+ io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15]
+ io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22]
+ io_out[23] io_out[24] io_out[25] io_out[26] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100] la_data_in[101]
+ la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105] la_data_in[106]
+ la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110] la_data_in[111]
+ la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115] la_data_in[116]
+ la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120] la_data_in[121]
+ la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125] la_data_in[126]
+ la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15] la_data_in[16]
+ la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20] la_data_in[21]
+ la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26] la_data_in[27]
+ la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31] la_data_in[32]
+ la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37] la_data_in[38]
+ la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42] la_data_in[43]
+ la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48] la_data_in[49]
+ la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53] la_data_in[54]
+ la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59] la_data_in[5]
+ la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64] la_data_in[65]
+ la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6] la_data_in[70]
+ la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75] la_data_in[76]
+ la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80] la_data_in[81]
+ la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86] la_data_in[87]
+ la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91] la_data_in[92]
+ la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97] la_data_in[98]
+ la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101] la_data_out[102]
+ la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106] la_data_out[107]
+ la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110] la_data_out[111]
+ la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115] la_data_out[116]
+ la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11] la_data_out[120]
+ la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124] la_data_out[125]
+ la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24]
+ la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29]
+ la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34]
+ la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39]
+ la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44]
+ la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49]
+ la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54]
+ la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59]
+ la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[64]
+ la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68] la_data_out[69]
+ la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73] la_data_out[74]
+ la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78] la_data_out[79]
+ la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83] la_data_out[84]
+ la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88] la_data_out[89]
+ la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93] la_data_out[94]
+ la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98] la_data_out[99]
+ la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104]
+ la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109] la_oenb[10] la_oenb[110]
+ la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117]
+ la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121] la_oenb[122] la_oenb[123]
+ la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65]
+ la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6] la_oenb[70] la_oenb[71]
+ la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76] la_oenb[77] la_oenb[78]
+ la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84]
+ la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89] la_oenb[8] la_oenb[90]
+ la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97]
+ la_oenb[98] la_oenb[99] la_oenb[9] user_clock2 user_irq[0] user_irq[1] user_irq[2]
+ vccd1 vccd2 vdda1 vdda2 vssa1 vssa2 vssd1 vssd2 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0]
+ wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15]
+ wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20]
+ wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26]
+ wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31]
+ wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9]
+ wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13]
+ wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19]
+ wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24]
+ wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2]
+ wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6]
+ wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3]
+ wbs_stb_i wbs_we_i
.ends

* Black-box entry subcircuit for caravan_motto abstract view
.subckt caravan_motto
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_8 abstract view
.subckt sky130_fd_sc_hd__ebufn_8 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_2 abstract view
.subckt sky130_fd_sc_hd__ebufn_2 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_2 abstract view
.subckt sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_2 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_4 abstract view
.subckt sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4bb_1 abstract view
.subckt sky130_fd_sc_hd__nand4bb_1 A_N B_N C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for housekeeping abstract view
.subckt housekeeping VGND VPWR debug_in debug_mode debug_oeb debug_out irq[0] irq[1]
+ irq[2] mask_rev_in[0] mask_rev_in[10] mask_rev_in[11] mask_rev_in[12] mask_rev_in[13]
+ mask_rev_in[14] mask_rev_in[15] mask_rev_in[16] mask_rev_in[17] mask_rev_in[18]
+ mask_rev_in[19] mask_rev_in[1] mask_rev_in[20] mask_rev_in[21] mask_rev_in[22] mask_rev_in[23]
+ mask_rev_in[24] mask_rev_in[25] mask_rev_in[26] mask_rev_in[27] mask_rev_in[28]
+ mask_rev_in[29] mask_rev_in[2] mask_rev_in[30] mask_rev_in[31] mask_rev_in[3] mask_rev_in[4]
+ mask_rev_in[5] mask_rev_in[6] mask_rev_in[7] mask_rev_in[8] mask_rev_in[9] mgmt_gpio_in[0]
+ mgmt_gpio_in[10] mgmt_gpio_in[11] mgmt_gpio_in[12] mgmt_gpio_in[13] mgmt_gpio_in[14]
+ mgmt_gpio_in[15] mgmt_gpio_in[16] mgmt_gpio_in[17] mgmt_gpio_in[18] mgmt_gpio_in[19]
+ mgmt_gpio_in[1] mgmt_gpio_in[20] mgmt_gpio_in[21] mgmt_gpio_in[22] mgmt_gpio_in[23]
+ mgmt_gpio_in[24] mgmt_gpio_in[25] mgmt_gpio_in[26] mgmt_gpio_in[27] mgmt_gpio_in[28]
+ mgmt_gpio_in[29] mgmt_gpio_in[2] mgmt_gpio_in[30] mgmt_gpio_in[31] mgmt_gpio_in[32]
+ mgmt_gpio_in[33] mgmt_gpio_in[34] mgmt_gpio_in[35] mgmt_gpio_in[36] mgmt_gpio_in[37]
+ mgmt_gpio_in[3] mgmt_gpio_in[4] mgmt_gpio_in[5] mgmt_gpio_in[6] mgmt_gpio_in[7]
+ mgmt_gpio_in[8] mgmt_gpio_in[9] mgmt_gpio_oeb[0] mgmt_gpio_oeb[10] mgmt_gpio_oeb[11]
+ mgmt_gpio_oeb[12] mgmt_gpio_oeb[13] mgmt_gpio_oeb[14] mgmt_gpio_oeb[15] mgmt_gpio_oeb[16]
+ mgmt_gpio_oeb[17] mgmt_gpio_oeb[18] mgmt_gpio_oeb[19] mgmt_gpio_oeb[1] mgmt_gpio_oeb[20]
+ mgmt_gpio_oeb[21] mgmt_gpio_oeb[22] mgmt_gpio_oeb[23] mgmt_gpio_oeb[24] mgmt_gpio_oeb[25]
+ mgmt_gpio_oeb[26] mgmt_gpio_oeb[27] mgmt_gpio_oeb[28] mgmt_gpio_oeb[29] mgmt_gpio_oeb[2]
+ mgmt_gpio_oeb[30] mgmt_gpio_oeb[31] mgmt_gpio_oeb[32] mgmt_gpio_oeb[33] mgmt_gpio_oeb[34]
+ mgmt_gpio_oeb[35] mgmt_gpio_oeb[36] mgmt_gpio_oeb[37] mgmt_gpio_oeb[3] mgmt_gpio_oeb[4]
+ mgmt_gpio_oeb[5] mgmt_gpio_oeb[6] mgmt_gpio_oeb[7] mgmt_gpio_oeb[8] mgmt_gpio_oeb[9]
+ mgmt_gpio_out[0] mgmt_gpio_out[10] mgmt_gpio_out[11] mgmt_gpio_out[12] mgmt_gpio_out[13]
+ mgmt_gpio_out[14] mgmt_gpio_out[15] mgmt_gpio_out[16] mgmt_gpio_out[17] mgmt_gpio_out[18]
+ mgmt_gpio_out[19] mgmt_gpio_out[1] mgmt_gpio_out[20] mgmt_gpio_out[21] mgmt_gpio_out[22]
+ mgmt_gpio_out[23] mgmt_gpio_out[24] mgmt_gpio_out[25] mgmt_gpio_out[26] mgmt_gpio_out[27]
+ mgmt_gpio_out[28] mgmt_gpio_out[29] mgmt_gpio_out[2] mgmt_gpio_out[30] mgmt_gpio_out[31]
+ mgmt_gpio_out[32] mgmt_gpio_out[33] mgmt_gpio_out[34] mgmt_gpio_out[35] mgmt_gpio_out[36]
+ mgmt_gpio_out[37] mgmt_gpio_out[3] mgmt_gpio_out[4] mgmt_gpio_out[5] mgmt_gpio_out[6]
+ mgmt_gpio_out[7] mgmt_gpio_out[8] mgmt_gpio_out[9] pad_flash_clk pad_flash_clk_oeb
+ pad_flash_csb pad_flash_csb_oeb pad_flash_io0_di pad_flash_io0_do pad_flash_io0_ieb
+ pad_flash_io0_oeb pad_flash_io1_di pad_flash_io1_do pad_flash_io1_ieb pad_flash_io1_oeb
+ pll90_sel[0] pll90_sel[1] pll90_sel[2] pll_bypass pll_dco_ena pll_div[0] pll_div[1]
+ pll_div[2] pll_div[3] pll_div[4] pll_ena pll_sel[0] pll_sel[1] pll_sel[2] pll_trim[0]
+ pll_trim[10] pll_trim[11] pll_trim[12] pll_trim[13] pll_trim[14] pll_trim[15] pll_trim[16]
+ pll_trim[17] pll_trim[18] pll_trim[19] pll_trim[1] pll_trim[20] pll_trim[21] pll_trim[22]
+ pll_trim[23] pll_trim[24] pll_trim[25] pll_trim[2] pll_trim[3] pll_trim[4] pll_trim[5]
+ pll_trim[6] pll_trim[7] pll_trim[8] pll_trim[9] porb pwr_ctrl_out[0] pwr_ctrl_out[1]
+ pwr_ctrl_out[2] pwr_ctrl_out[3] qspi_enabled reset ser_rx ser_tx serial_clock serial_data_1
+ serial_data_2 serial_load serial_resetn spi_csb spi_enabled spi_sck spi_sdi spi_sdo
+ spi_sdoenb spimemio_flash_clk spimemio_flash_csb spimemio_flash_io0_di spimemio_flash_io0_do
+ spimemio_flash_io0_oeb spimemio_flash_io1_di spimemio_flash_io1_do spimemio_flash_io1_oeb
+ spimemio_flash_io2_di spimemio_flash_io2_do spimemio_flash_io2_oeb spimemio_flash_io3_di
+ spimemio_flash_io3_do spimemio_flash_io3_oeb sram_ro_addr[0] sram_ro_addr[1] sram_ro_addr[2]
+ sram_ro_addr[3] sram_ro_addr[4] sram_ro_addr[5] sram_ro_addr[6] sram_ro_addr[7]
+ sram_ro_clk sram_ro_csb sram_ro_data[0] sram_ro_data[10] sram_ro_data[11] sram_ro_data[12]
+ sram_ro_data[13] sram_ro_data[14] sram_ro_data[15] sram_ro_data[16] sram_ro_data[17]
+ sram_ro_data[18] sram_ro_data[19] sram_ro_data[1] sram_ro_data[20] sram_ro_data[21]
+ sram_ro_data[22] sram_ro_data[23] sram_ro_data[24] sram_ro_data[25] sram_ro_data[26]
+ sram_ro_data[27] sram_ro_data[28] sram_ro_data[29] sram_ro_data[2] sram_ro_data[30]
+ sram_ro_data[31] sram_ro_data[3] sram_ro_data[4] sram_ro_data[5] sram_ro_data[6]
+ sram_ro_data[7] sram_ro_data[8] sram_ro_data[9] trap uart_enabled user_clock usr1_vcc_pwrgood
+ usr1_vdd_pwrgood usr2_vcc_pwrgood usr2_vdd_pwrgood wb_ack_o wb_adr_i[0] wb_adr_i[10]
+ wb_adr_i[11] wb_adr_i[12] wb_adr_i[13] wb_adr_i[14] wb_adr_i[15] wb_adr_i[16] wb_adr_i[17]
+ wb_adr_i[18] wb_adr_i[19] wb_adr_i[1] wb_adr_i[20] wb_adr_i[21] wb_adr_i[22] wb_adr_i[23]
+ wb_adr_i[24] wb_adr_i[25] wb_adr_i[26] wb_adr_i[27] wb_adr_i[28] wb_adr_i[29] wb_adr_i[2]
+ wb_adr_i[30] wb_adr_i[31] wb_adr_i[3] wb_adr_i[4] wb_adr_i[5] wb_adr_i[6] wb_adr_i[7]
+ wb_adr_i[8] wb_adr_i[9] wb_clk_i wb_cyc_i wb_dat_i[0] wb_dat_i[10] wb_dat_i[11]
+ wb_dat_i[12] wb_dat_i[13] wb_dat_i[14] wb_dat_i[15] wb_dat_i[16] wb_dat_i[17] wb_dat_i[18]
+ wb_dat_i[19] wb_dat_i[1] wb_dat_i[20] wb_dat_i[21] wb_dat_i[22] wb_dat_i[23] wb_dat_i[24]
+ wb_dat_i[25] wb_dat_i[26] wb_dat_i[27] wb_dat_i[28] wb_dat_i[29] wb_dat_i[2] wb_dat_i[30]
+ wb_dat_i[31] wb_dat_i[3] wb_dat_i[4] wb_dat_i[5] wb_dat_i[6] wb_dat_i[7] wb_dat_i[8]
+ wb_dat_i[9] wb_dat_o[0] wb_dat_o[10] wb_dat_o[11] wb_dat_o[12] wb_dat_o[13] wb_dat_o[14]
+ wb_dat_o[15] wb_dat_o[16] wb_dat_o[17] wb_dat_o[18] wb_dat_o[19] wb_dat_o[1] wb_dat_o[20]
+ wb_dat_o[21] wb_dat_o[22] wb_dat_o[23] wb_dat_o[24] wb_dat_o[25] wb_dat_o[26] wb_dat_o[27]
+ wb_dat_o[28] wb_dat_o[29] wb_dat_o[2] wb_dat_o[30] wb_dat_o[31] wb_dat_o[3] wb_dat_o[4]
+ wb_dat_o[5] wb_dat_o[6] wb_dat_o[7] wb_dat_o[8] wb_dat_o[9] wb_rstn_i wb_sel_i[0]
+ wb_sel_i[1] wb_sel_i[2] wb_sel_i[3] wb_stb_i wb_we_i
.ends

.subckt caravan clock flash_clk flash_csb flash_io0 flash_io1 gpio mprj_io[0] mprj_io[10]
+ mprj_io[11] mprj_io[12] mprj_io[13] mprj_io[14] mprj_io[15] mprj_io[16] mprj_io[17]
+ mprj_io[18] mprj_io[19] mprj_io[1] mprj_io[20] mprj_io[21] mprj_io[22] mprj_io[23]
+ mprj_io[24] mprj_io[25] mprj_io[26] mprj_io[27] mprj_io[28] mprj_io[29] mprj_io[2]
+ mprj_io[30] mprj_io[31] mprj_io[32] mprj_io[33] mprj_io[34] mprj_io[35] mprj_io[36]
+ mprj_io[37] mprj_io[3] mprj_io[4] mprj_io[5] mprj_io[6] mprj_io[7] mprj_io[8] mprj_io[9]
+ resetb vccd vccd1 vccd2 vdda vdda1 vdda1_2 vdda2 vddio vddio_2 vssa vssa1 vssa1_2
+ vssa2 vssd vssd1 vssd2 vssio vssio_2
Xgpio_control_in_2\[0\] gpio_defaults_block_14/gpio_defaults[0] gpio_defaults_block_14/gpio_defaults[10]
+ gpio_defaults_block_14/gpio_defaults[11] gpio_defaults_block_14/gpio_defaults[12]
+ gpio_defaults_block_14/gpio_defaults[1] gpio_defaults_block_14/gpio_defaults[2]
+ gpio_defaults_block_14/gpio_defaults[3] gpio_defaults_block_14/gpio_defaults[4]
+ gpio_defaults_block_14/gpio_defaults[5] gpio_defaults_block_14/gpio_defaults[6]
+ gpio_defaults_block_14/gpio_defaults[7] gpio_defaults_block_14/gpio_defaults[8]
+ gpio_defaults_block_14/gpio_defaults[9] housekeeping/mgmt_gpio_in[25] gpio_control_in_2\[0\]/one
+ housekeeping/mgmt_gpio_in[25] gpio_control_in_2\[0\]/one padframe/mprj_io_analog_en[14]
+ padframe/mprj_io_analog_pol[14] padframe/mprj_io_analog_sel[14] padframe/mprj_io_dm[42]
+ padframe/mprj_io_dm[43] padframe/mprj_io_dm[44] padframe/mprj_io_holdover[14] padframe/mprj_io_ib_mode_sel[14]
+ padframe/mprj_io_in[14] padframe/mprj_io_inp_dis[14] padframe/mprj_io_out[14] padframe/mprj_io_oeb[14]
+ padframe/mprj_io_slow_sel[14] padframe/mprj_io_vtrip_sel[14] gpio_control_in_2\[0\]/resetn
+ gpio_control_in_2\[0\]/resetn_out gpio_control_in_2\[0\]/serial_clock gpio_control_in_2\[0\]/serial_clock_out
+ gpio_control_in_2\[0\]/serial_data_in gpio_control_in_2\[0\]/serial_data_out gpio_control_in_2\[0\]/serial_load
+ gpio_control_in_2\[0\]/serial_load_out mprj/io_in[14] mprj/io_oeb[14] mprj/io_out[14]
+ vccd_core vccd1_core VSUBS vssd1_core gpio_control_in_2\[0\]/zero gpio_control_block
Xgpio_defaults_block_11 VSUBS vccd_core gpio_defaults_block_11/gpio_defaults[0] gpio_defaults_block_11/gpio_defaults[10]
+ gpio_defaults_block_11/gpio_defaults[11] gpio_defaults_block_11/gpio_defaults[12]
+ gpio_defaults_block_11/gpio_defaults[1] gpio_defaults_block_11/gpio_defaults[2]
+ gpio_defaults_block_11/gpio_defaults[3] gpio_defaults_block_11/gpio_defaults[4]
+ gpio_defaults_block_11/gpio_defaults[5] gpio_defaults_block_11/gpio_defaults[6]
+ gpio_defaults_block_11/gpio_defaults[7] gpio_defaults_block_11/gpio_defaults[8]
+ gpio_defaults_block_11/gpio_defaults[9] gpio_defaults_block
Xgpio_defaults_block_33 VSUBS vccd_core gpio_defaults_block_33/gpio_defaults[0] gpio_defaults_block_33/gpio_defaults[10]
+ gpio_defaults_block_33/gpio_defaults[11] gpio_defaults_block_33/gpio_defaults[12]
+ gpio_defaults_block_33/gpio_defaults[1] gpio_defaults_block_33/gpio_defaults[2]
+ gpio_defaults_block_33/gpio_defaults[3] gpio_defaults_block_33/gpio_defaults[4]
+ gpio_defaults_block_33/gpio_defaults[5] gpio_defaults_block_33/gpio_defaults[6]
+ gpio_defaults_block_33/gpio_defaults[7] gpio_defaults_block_33/gpio_defaults[8]
+ gpio_defaults_block_33/gpio_defaults[9] gpio_defaults_block
Xgpio_defaults_block_12 VSUBS vccd_core gpio_defaults_block_12/gpio_defaults[0] gpio_defaults_block_12/gpio_defaults[10]
+ gpio_defaults_block_12/gpio_defaults[11] gpio_defaults_block_12/gpio_defaults[12]
+ gpio_defaults_block_12/gpio_defaults[1] gpio_defaults_block_12/gpio_defaults[2]
+ gpio_defaults_block_12/gpio_defaults[3] gpio_defaults_block_12/gpio_defaults[4]
+ gpio_defaults_block_12/gpio_defaults[5] gpio_defaults_block_12/gpio_defaults[6]
+ gpio_defaults_block_12/gpio_defaults[7] gpio_defaults_block_12/gpio_defaults[8]
+ gpio_defaults_block_12/gpio_defaults[9] gpio_defaults_block
Xgpio_defaults_block_34 VSUBS vccd_core gpio_defaults_block_34/gpio_defaults[0] gpio_defaults_block_34/gpio_defaults[10]
+ gpio_defaults_block_34/gpio_defaults[11] gpio_defaults_block_34/gpio_defaults[12]
+ gpio_defaults_block_34/gpio_defaults[1] gpio_defaults_block_34/gpio_defaults[2]
+ gpio_defaults_block_34/gpio_defaults[3] gpio_defaults_block_34/gpio_defaults[4]
+ gpio_defaults_block_34/gpio_defaults[5] gpio_defaults_block_34/gpio_defaults[6]
+ gpio_defaults_block_34/gpio_defaults[7] gpio_defaults_block_34/gpio_defaults[8]
+ gpio_defaults_block_34/gpio_defaults[9] gpio_defaults_block
Xpll VSUBS vccd_core pll/clockp[0] pll/clockp[1] pll/dco pll/div[0] pll/div[1] pll/div[2]
+ pll/div[3] pll/div[4] pll/enable pll/ext_trim[0] pll/ext_trim[10] pll/ext_trim[11]
+ pll/ext_trim[12] pll/ext_trim[13] pll/ext_trim[14] pll/ext_trim[15] pll/ext_trim[16]
+ pll/ext_trim[17] pll/ext_trim[18] pll/ext_trim[19] pll/ext_trim[1] pll/ext_trim[20]
+ pll/ext_trim[21] pll/ext_trim[22] pll/ext_trim[23] pll/ext_trim[24] pll/ext_trim[25]
+ pll/ext_trim[2] pll/ext_trim[3] pll/ext_trim[4] pll/ext_trim[5] pll/ext_trim[6]
+ pll/ext_trim[7] pll/ext_trim[8] pll/ext_trim[9] pll/osc pll/resetb digital_pll
Xpadframe clock pll/osc por/por_l flash_clk flash_csb flash_io0 padframe/flash_io0_di_core
+ padframe/flash_io0_do_core padframe/flash_io0_ieb_core padframe/flash_io0_oeb_core
+ flash_io1 padframe/flash_io1_di_core padframe/flash_io1_do_core padframe/flash_io1_ieb_core
+ padframe/flash_io1_oeb_core gpio soc/gpio_in_pad soc/gpio_inenb_pad soc/gpio_mode0_pad
+ soc/gpio_mode1_pad soc/gpio_out_pad soc/gpio_outenb_pad vccd vdda vddio vddio_2
+ vssa vssd vssio vssio_2 mprj_io[0] padframe/mprj_io_analog_en[0] padframe/mprj_io_analog_pol[0]
+ padframe/mprj_io_analog_sel[0] padframe/mprj_io_dm[0] padframe/mprj_io_dm[1] padframe/mprj_io_dm[2]
+ padframe/mprj_io_holdover[0] padframe/mprj_io_ib_mode_sel[0] padframe/mprj_io_inp_dis[0]
+ padframe/mprj_io_oeb[0] padframe/mprj_io_out[0] padframe/mprj_io_slow_sel[0] padframe/mprj_io_vtrip_sel[0]
+ padframe/mprj_io_in[0] mprj/io_in_3v3[0] mprj/gpio_analog[3] mprj/gpio_noesd[3]
+ mprj_io[10] padframe/mprj_io_analog_en[10] padframe/mprj_io_analog_pol[10] padframe/mprj_io_analog_sel[10]
+ padframe/mprj_io_dm[30] padframe/mprj_io_dm[31] padframe/mprj_io_dm[32] padframe/mprj_io_holdover[10]
+ padframe/mprj_io_ib_mode_sel[10] padframe/mprj_io_inp_dis[10] padframe/mprj_io_oeb[10]
+ padframe/mprj_io_out[10] padframe/mprj_io_slow_sel[10] padframe/mprj_io_vtrip_sel[10]
+ padframe/mprj_io_in[10] mprj/io_in_3v3[10] mprj/gpio_analog[4] mprj/gpio_noesd[4]
+ mprj_io[11] padframe/mprj_io_analog_en[11] padframe/mprj_io_analog_pol[11] padframe/mprj_io_analog_sel[11]
+ padframe/mprj_io_dm[33] padframe/mprj_io_dm[34] padframe/mprj_io_dm[35] padframe/mprj_io_holdover[11]
+ padframe/mprj_io_ib_mode_sel[11] padframe/mprj_io_inp_dis[11] padframe/mprj_io_oeb[11]
+ padframe/mprj_io_out[11] padframe/mprj_io_slow_sel[11] padframe/mprj_io_vtrip_sel[11]
+ padframe/mprj_io_in[11] mprj/io_in_3v3[11] mprj/gpio_analog[5] mprj/gpio_noesd[5]
+ mprj_io[12] padframe/mprj_io_analog_en[12] padframe/mprj_io_analog_pol[12] padframe/mprj_io_analog_sel[12]
+ padframe/mprj_io_dm[36] padframe/mprj_io_dm[37] padframe/mprj_io_dm[38] padframe/mprj_io_holdover[12]
+ padframe/mprj_io_ib_mode_sel[12] padframe/mprj_io_inp_dis[12] padframe/mprj_io_oeb[12]
+ padframe/mprj_io_out[12] padframe/mprj_io_slow_sel[12] padframe/mprj_io_vtrip_sel[12]
+ padframe/mprj_io_in[12] mprj/io_in_3v3[12] mprj/gpio_analog[6] mprj/gpio_noesd[6]
+ mprj_io[13] padframe/mprj_io_analog_en[13] padframe/mprj_io_analog_pol[13] padframe/mprj_io_analog_sel[13]
+ padframe/mprj_io_dm[39] padframe/mprj_io_dm[40] padframe/mprj_io_dm[41] padframe/mprj_io_holdover[13]
+ padframe/mprj_io_ib_mode_sel[13] padframe/mprj_io_inp_dis[13] padframe/mprj_io_oeb[13]
+ padframe/mprj_io_out[13] padframe/mprj_io_slow_sel[13] padframe/mprj_io_vtrip_sel[13]
+ padframe/mprj_io_in[13] mprj/io_in_3v3[13] mprj_io[1] padframe/mprj_io_analog_en[1]
+ padframe/mprj_io_analog_pol[1] padframe/mprj_io_analog_sel[1] padframe/mprj_io_dm[3]
+ padframe/mprj_io_dm[4] padframe/mprj_io_dm[5] padframe/mprj_io_holdover[1] padframe/mprj_io_ib_mode_sel[1]
+ padframe/mprj_io_inp_dis[1] padframe/mprj_io_oeb[1] padframe/mprj_io_out[1] padframe/mprj_io_slow_sel[1]
+ padframe/mprj_io_vtrip_sel[1] padframe/mprj_io_in[1] mprj/io_in_3v3[1] mprj_io[2]
+ padframe/mprj_io_analog_en[2] padframe/mprj_io_analog_pol[2] padframe/mprj_io_analog_sel[2]
+ padframe/mprj_io_dm[6] padframe/mprj_io_dm[7] padframe/mprj_io_dm[8] padframe/mprj_io_holdover[2]
+ padframe/mprj_io_ib_mode_sel[2] padframe/mprj_io_inp_dis[2] padframe/mprj_io_oeb[2]
+ padframe/mprj_io_out[2] padframe/mprj_io_slow_sel[2] padframe/mprj_io_vtrip_sel[2]
+ padframe/mprj_io_in[2] mprj/io_in_3v3[2] mprj_io[3] padframe/mprj_io_analog_en[3]
+ padframe/mprj_io_analog_pol[3] padframe/mprj_io_analog_sel[3] padframe/mprj_io_dm[10]
+ padframe/mprj_io_dm[11] padframe/mprj_io_dm[9] padframe/mprj_io_holdover[3] padframe/mprj_io_ib_mode_sel[3]
+ padframe/mprj_io_inp_dis[3] padframe/mprj_io_oeb[3] padframe/mprj_io_out[3] padframe/mprj_io_slow_sel[3]
+ padframe/mprj_io_vtrip_sel[3] padframe/mprj_io_in[3] mprj/io_in_3v3[3] mprj_io[4]
+ padframe/mprj_io_analog_en[4] padframe/mprj_io_analog_pol[4] padframe/mprj_io_analog_sel[4]
+ padframe/mprj_io_dm[12] padframe/mprj_io_dm[13] padframe/mprj_io_dm[14] padframe/mprj_io_holdover[4]
+ padframe/mprj_io_ib_mode_sel[4] padframe/mprj_io_inp_dis[4] padframe/mprj_io_oeb[4]
+ padframe/mprj_io_out[4] padframe/mprj_io_slow_sel[4] padframe/mprj_io_vtrip_sel[4]
+ padframe/mprj_io_in[4] mprj/io_in_3v3[4] mprj_io[5] padframe/mprj_io_analog_en[5]
+ padframe/mprj_io_analog_pol[5] padframe/mprj_io_analog_sel[5] padframe/mprj_io_dm[15]
+ padframe/mprj_io_dm[16] padframe/mprj_io_dm[17] padframe/mprj_io_holdover[5] padframe/mprj_io_ib_mode_sel[5]
+ padframe/mprj_io_inp_dis[5] padframe/mprj_io_oeb[5] padframe/mprj_io_out[5] padframe/mprj_io_slow_sel[5]
+ padframe/mprj_io_vtrip_sel[5] padframe/mprj_io_in[5] mprj/io_in_3v3[5] mprj_io[6]
+ padframe/mprj_io_analog_en[6] padframe/mprj_io_analog_pol[6] padframe/mprj_io_analog_sel[6]
+ padframe/mprj_io_dm[18] padframe/mprj_io_dm[19] padframe/mprj_io_dm[20] padframe/mprj_io_holdover[6]
+ padframe/mprj_io_ib_mode_sel[6] padframe/mprj_io_inp_dis[6] padframe/mprj_io_oeb[6]
+ padframe/mprj_io_out[6] padframe/mprj_io_slow_sel[6] padframe/mprj_io_vtrip_sel[6]
+ padframe/mprj_io_in[6] mprj/io_in_3v3[6] mprj/gpio_analog[0] mprj/gpio_noesd[0]
+ mprj_io[7] padframe/mprj_io_analog_en[7] padframe/mprj_io_analog_pol[7] padframe/mprj_io_analog_sel[7]
+ padframe/mprj_io_dm[21] padframe/mprj_io_dm[22] padframe/mprj_io_dm[23] padframe/mprj_io_holdover[7]
+ padframe/mprj_io_ib_mode_sel[7] padframe/mprj_io_inp_dis[7] padframe/mprj_io_oeb[7]
+ padframe/mprj_io_out[7] padframe/mprj_io_slow_sel[7] padframe/mprj_io_vtrip_sel[7]
+ padframe/mprj_io_in[7] mprj/io_in_3v3[7] mprj/gpio_analog[1] mprj/gpio_noesd[1]
+ mprj_io[8] padframe/mprj_io_analog_en[8] padframe/mprj_io_analog_pol[8] padframe/mprj_io_analog_sel[8]
+ padframe/mprj_io_dm[24] padframe/mprj_io_dm[25] padframe/mprj_io_dm[26] padframe/mprj_io_holdover[8]
+ padframe/mprj_io_ib_mode_sel[8] padframe/mprj_io_inp_dis[8] padframe/mprj_io_oeb[8]
+ padframe/mprj_io_out[8] padframe/mprj_io_slow_sel[8] padframe/mprj_io_vtrip_sel[8]
+ padframe/mprj_io_in[8] mprj/io_in_3v3[8] mprj/gpio_analog[2] mprj/gpio_noesd[2]
+ mprj_io[9] padframe/mprj_io_analog_en[9] padframe/mprj_io_analog_pol[9] padframe/mprj_io_analog_sel[9]
+ padframe/mprj_io_dm[27] padframe/mprj_io_dm[28] padframe/mprj_io_dm[29] padframe/mprj_io_holdover[9]
+ padframe/mprj_io_ib_mode_sel[9] padframe/mprj_io_inp_dis[9] padframe/mprj_io_oeb[9]
+ padframe/mprj_io_out[9] padframe/mprj_io_slow_sel[9] padframe/mprj_io_vtrip_sel[9]
+ padframe/mprj_io_in[9] mprj/io_in_3v3[9] mprj/gpio_analog[7] mprj/gpio_noesd[7]
+ mprj_io[25] padframe/mprj_io_analog_en[14] padframe/mprj_io_analog_pol[14] padframe/mprj_io_analog_sel[14]
+ padframe/mprj_io_dm[42] padframe/mprj_io_dm[43] padframe/mprj_io_dm[44] padframe/mprj_io_holdover[14]
+ padframe/mprj_io_ib_mode_sel[14] padframe/mprj_io_inp_dis[14] padframe/mprj_io_oeb[14]
+ padframe/mprj_io_out[14] padframe/mprj_io_slow_sel[14] padframe/mprj_io_vtrip_sel[14]
+ padframe/mprj_io_in[14] mprj/io_in_3v3[14] mprj/gpio_analog[17] mprj/gpio_noesd[17]
+ mprj_io[35] padframe/mprj_io_analog_en[24] padframe/mprj_io_analog_pol[24] padframe/mprj_io_analog_sel[24]
+ padframe/mprj_io_dm[72] padframe/mprj_io_dm[73] padframe/mprj_io_dm[74] padframe/mprj_io_holdover[24]
+ padframe/mprj_io_ib_mode_sel[24] padframe/mprj_io_inp_dis[24] padframe/mprj_io_oeb[24]
+ padframe/mprj_io_out[24] padframe/mprj_io_slow_sel[24] padframe/mprj_io_vtrip_sel[24]
+ padframe/mprj_io_in[24] mprj/io_in_3v3[24] mprj_io[36] padframe/mprj_io_analog_en[25]
+ padframe/mprj_io_analog_pol[25] padframe/mprj_io_analog_sel[25] padframe/mprj_io_dm[75]
+ padframe/mprj_io_dm[76] padframe/mprj_io_dm[77] padframe/mprj_io_holdover[25] padframe/mprj_io_ib_mode_sel[25]
+ padframe/mprj_io_inp_dis[25] padframe/mprj_io_oeb[25] padframe/mprj_io_out[25] padframe/mprj_io_slow_sel[25]
+ padframe/mprj_io_vtrip_sel[25] padframe/mprj_io_in[25] mprj/io_in_3v3[25] mprj_io[37]
+ padframe/mprj_io_analog_en[26] padframe/mprj_io_analog_pol[26] padframe/mprj_io_analog_sel[26]
+ padframe/mprj_io_dm[78] padframe/mprj_io_dm[79] padframe/mprj_io_dm[80] padframe/mprj_io_holdover[26]
+ padframe/mprj_io_ib_mode_sel[26] padframe/mprj_io_inp_dis[26] padframe/mprj_io_oeb[26]
+ padframe/mprj_io_out[26] padframe/mprj_io_slow_sel[26] padframe/mprj_io_vtrip_sel[26]
+ padframe/mprj_io_in[26] mprj/io_in_3v3[26] mprj/gpio_analog[8] mprj/gpio_noesd[8]
+ mprj_io[26] padframe/mprj_io_analog_en[15] padframe/mprj_io_analog_pol[15] padframe/mprj_io_analog_sel[15]
+ padframe/mprj_io_dm[45] padframe/mprj_io_dm[46] padframe/mprj_io_dm[47] padframe/mprj_io_holdover[15]
+ padframe/mprj_io_ib_mode_sel[15] padframe/mprj_io_inp_dis[15] padframe/mprj_io_oeb[15]
+ padframe/mprj_io_out[15] padframe/mprj_io_slow_sel[15] padframe/mprj_io_vtrip_sel[15]
+ padframe/mprj_io_in[15] mprj/io_in_3v3[15] mprj/gpio_analog[9] mprj/gpio_noesd[9]
+ mprj_io[27] padframe/mprj_io_analog_en[16] padframe/mprj_io_analog_pol[16] padframe/mprj_io_analog_sel[16]
+ padframe/mprj_io_dm[48] padframe/mprj_io_dm[49] padframe/mprj_io_dm[50] padframe/mprj_io_holdover[16]
+ padframe/mprj_io_ib_mode_sel[16] padframe/mprj_io_inp_dis[16] padframe/mprj_io_oeb[16]
+ padframe/mprj_io_out[16] padframe/mprj_io_slow_sel[16] padframe/mprj_io_vtrip_sel[16]
+ padframe/mprj_io_in[16] mprj/io_in_3v3[16] mprj/gpio_analog[10] mprj/gpio_noesd[10]
+ mprj_io[28] padframe/mprj_io_analog_en[17] padframe/mprj_io_analog_pol[17] padframe/mprj_io_analog_sel[17]
+ padframe/mprj_io_dm[51] padframe/mprj_io_dm[52] padframe/mprj_io_dm[53] padframe/mprj_io_holdover[17]
+ padframe/mprj_io_ib_mode_sel[17] padframe/mprj_io_inp_dis[17] padframe/mprj_io_oeb[17]
+ padframe/mprj_io_out[17] padframe/mprj_io_slow_sel[17] padframe/mprj_io_vtrip_sel[17]
+ padframe/mprj_io_in[17] mprj/io_in_3v3[17] mprj/gpio_analog[11] mprj/gpio_noesd[11]
+ mprj_io[29] padframe/mprj_io_analog_en[18] padframe/mprj_io_analog_pol[18] padframe/mprj_io_analog_sel[18]
+ padframe/mprj_io_dm[54] padframe/mprj_io_dm[55] padframe/mprj_io_dm[56] padframe/mprj_io_holdover[18]
+ padframe/mprj_io_ib_mode_sel[18] padframe/mprj_io_inp_dis[18] padframe/mprj_io_oeb[18]
+ padframe/mprj_io_out[18] padframe/mprj_io_slow_sel[18] padframe/mprj_io_vtrip_sel[18]
+ padframe/mprj_io_in[18] mprj/io_in_3v3[18] mprj/gpio_analog[12] mprj/gpio_noesd[12]
+ mprj_io[30] padframe/mprj_io_analog_en[19] padframe/mprj_io_analog_pol[19] padframe/mprj_io_analog_sel[19]
+ padframe/mprj_io_dm[57] padframe/mprj_io_dm[58] padframe/mprj_io_dm[59] padframe/mprj_io_holdover[19]
+ padframe/mprj_io_ib_mode_sel[19] padframe/mprj_io_inp_dis[19] padframe/mprj_io_oeb[19]
+ padframe/mprj_io_out[19] padframe/mprj_io_slow_sel[19] padframe/mprj_io_vtrip_sel[19]
+ padframe/mprj_io_in[19] mprj/io_in_3v3[19] mprj/gpio_analog[13] mprj/gpio_noesd[13]
+ mprj_io[31] padframe/mprj_io_analog_en[20] padframe/mprj_io_analog_pol[20] padframe/mprj_io_analog_sel[20]
+ padframe/mprj_io_dm[60] padframe/mprj_io_dm[61] padframe/mprj_io_dm[62] padframe/mprj_io_holdover[20]
+ padframe/mprj_io_ib_mode_sel[20] padframe/mprj_io_inp_dis[20] padframe/mprj_io_oeb[20]
+ padframe/mprj_io_out[20] padframe/mprj_io_slow_sel[20] padframe/mprj_io_vtrip_sel[20]
+ padframe/mprj_io_in[20] mprj/io_in_3v3[20] mprj/gpio_analog[14] mprj/gpio_noesd[14]
+ mprj_io[32] padframe/mprj_io_analog_en[21] padframe/mprj_io_analog_pol[21] padframe/mprj_io_analog_sel[21]
+ padframe/mprj_io_dm[63] padframe/mprj_io_dm[64] padframe/mprj_io_dm[65] padframe/mprj_io_holdover[21]
+ padframe/mprj_io_ib_mode_sel[21] padframe/mprj_io_inp_dis[21] padframe/mprj_io_oeb[21]
+ padframe/mprj_io_out[21] padframe/mprj_io_slow_sel[21] padframe/mprj_io_vtrip_sel[21]
+ padframe/mprj_io_in[21] mprj/io_in_3v3[21] mprj/gpio_analog[15] mprj/gpio_noesd[15]
+ mprj_io[33] padframe/mprj_io_analog_en[22] padframe/mprj_io_analog_pol[22] padframe/mprj_io_analog_sel[22]
+ padframe/mprj_io_dm[66] padframe/mprj_io_dm[67] padframe/mprj_io_dm[68] padframe/mprj_io_holdover[22]
+ padframe/mprj_io_ib_mode_sel[22] padframe/mprj_io_inp_dis[22] padframe/mprj_io_oeb[22]
+ padframe/mprj_io_out[22] padframe/mprj_io_slow_sel[22] padframe/mprj_io_vtrip_sel[22]
+ padframe/mprj_io_in[22] mprj/io_in_3v3[22] mprj/gpio_analog[16] mprj/gpio_noesd[16]
+ mprj_io[34] padframe/mprj_io_analog_en[23] padframe/mprj_io_analog_pol[23] padframe/mprj_io_analog_sel[23]
+ padframe/mprj_io_dm[69] padframe/mprj_io_dm[70] padframe/mprj_io_dm[71] padframe/mprj_io_holdover[23]
+ padframe/mprj_io_ib_mode_sel[23] padframe/mprj_io_inp_dis[23] padframe/mprj_io_oeb[23]
+ padframe/mprj_io_out[23] padframe/mprj_io_slow_sel[23] padframe/mprj_io_vtrip_sel[23]
+ padframe/mprj_io_in[23] mprj/io_in_3v3[23] por/porb_h resetb rstb_level/A padframe/vdda
+ padframe/vssa VSUBS mprj/io_analog[1] mprj_io[15] mprj/io_analog[2] mprj_io[16]
+ mprj/io_analog[3] mprj_io[17] mprj/io_analog[0] mprj_io[14] mprj/io_analog[4] mprj/io_clamp_high[0]
+ mprj/io_clamp_low[0] mprj_io[18] vccd1 vdda1 vdda1_2 vssa1 vssa1_2 vccd1_core vdda1_core
+ vssa1_core vssd1_core vssd1 mprj/io_analog[7] mprj_io[21] mprj/io_analog[8] mprj_io[22]
+ mprj/io_analog[9] mprj_io[23] mprj/io_analog[10] mprj_io[24] mprj/io_analog[5] mprj/io_clamp_high[1]
+ mprj/io_clamp_low[1] mprj_io[19] mprj/io_analog[6] mprj/io_clamp_high[2] mprj/io_clamp_low[2]
+ mprj_io[20] vccd2 vdda2 vssa2 vccd_core vccd2_core vdda2_core por/vdd3v3 vssa2_core
+ vssd2_core vssd2 por/vss3v3 padframe/flash_csb_core padframe/flash_clk_ieb_core
+ padframe/flash_clk_oeb_core padframe/flash_clk_core padframe/flash_csb_oeb_core
+ padframe/flash_csb_ieb_core chip_io_alt
Xgpio_defaults_block_13 VSUBS vccd_core gpio_defaults_block_13/gpio_defaults[0] gpio_defaults_block_13/gpio_defaults[10]
+ gpio_defaults_block_13/gpio_defaults[11] gpio_defaults_block_13/gpio_defaults[12]
+ gpio_defaults_block_13/gpio_defaults[1] gpio_defaults_block_13/gpio_defaults[2]
+ gpio_defaults_block_13/gpio_defaults[3] gpio_defaults_block_13/gpio_defaults[4]
+ gpio_defaults_block_13/gpio_defaults[5] gpio_defaults_block_13/gpio_defaults[6]
+ gpio_defaults_block_13/gpio_defaults[7] gpio_defaults_block_13/gpio_defaults[8]
+ gpio_defaults_block_13/gpio_defaults[9] gpio_defaults_block
Xgpio_control_in_1a\[3\] gpio_defaults_block_5/gpio_defaults[0] gpio_defaults_block_5/gpio_defaults[10]
+ gpio_defaults_block_5/gpio_defaults[11] gpio_defaults_block_5/gpio_defaults[12]
+ gpio_defaults_block_5/gpio_defaults[1] gpio_defaults_block_5/gpio_defaults[2] gpio_defaults_block_5/gpio_defaults[3]
+ gpio_defaults_block_5/gpio_defaults[4] gpio_defaults_block_5/gpio_defaults[5] gpio_defaults_block_5/gpio_defaults[6]
+ gpio_defaults_block_5/gpio_defaults[7] gpio_defaults_block_5/gpio_defaults[8] gpio_defaults_block_5/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[5] gpio_control_in_1a\[3\]/one housekeeping/mgmt_gpio_in[5]
+ gpio_control_in_1a\[3\]/one padframe/mprj_io_analog_en[5] padframe/mprj_io_analog_pol[5]
+ padframe/mprj_io_analog_sel[5] padframe/mprj_io_dm[15] padframe/mprj_io_dm[16] padframe/mprj_io_dm[17]
+ padframe/mprj_io_holdover[5] padframe/mprj_io_ib_mode_sel[5] padframe/mprj_io_in[5]
+ padframe/mprj_io_inp_dis[5] padframe/mprj_io_out[5] padframe/mprj_io_oeb[5] padframe/mprj_io_slow_sel[5]
+ padframe/mprj_io_vtrip_sel[5] gpio_control_in_1a\[3\]/resetn gpio_control_in_1a\[4\]/resetn
+ gpio_control_in_1a\[3\]/serial_clock gpio_control_in_1a\[4\]/serial_clock gpio_control_in_1a\[3\]/serial_data_in
+ gpio_control_in_1a\[4\]/serial_data_in gpio_control_in_1a\[3\]/serial_load gpio_control_in_1a\[4\]/serial_load
+ mprj/io_in[5] mprj/io_oeb[5] mprj/io_out[5] vccd_core vccd1_core VSUBS vssd1_core
+ gpio_control_in_1a\[3\]/zero gpio_control_block
Xgpio_defaults_block_35 VSUBS vccd_core gpio_defaults_block_35/gpio_defaults[0] gpio_defaults_block_35/gpio_defaults[10]
+ gpio_defaults_block_35/gpio_defaults[11] gpio_defaults_block_35/gpio_defaults[12]
+ gpio_defaults_block_35/gpio_defaults[1] gpio_defaults_block_35/gpio_defaults[2]
+ gpio_defaults_block_35/gpio_defaults[3] gpio_defaults_block_35/gpio_defaults[4]
+ gpio_defaults_block_35/gpio_defaults[5] gpio_defaults_block_35/gpio_defaults[6]
+ gpio_defaults_block_35/gpio_defaults[7] gpio_defaults_block_35/gpio_defaults[8]
+ gpio_defaults_block_35/gpio_defaults[9] gpio_defaults_block
Xgpio_control_bidir_2\[0\] gpio_defaults_block_35/gpio_defaults[0] gpio_defaults_block_35/gpio_defaults[10]
+ gpio_defaults_block_35/gpio_defaults[11] gpio_defaults_block_35/gpio_defaults[12]
+ gpio_defaults_block_35/gpio_defaults[1] gpio_defaults_block_35/gpio_defaults[2]
+ gpio_defaults_block_35/gpio_defaults[3] gpio_defaults_block_35/gpio_defaults[4]
+ gpio_defaults_block_35/gpio_defaults[5] gpio_defaults_block_35/gpio_defaults[6]
+ gpio_defaults_block_35/gpio_defaults[7] gpio_defaults_block_35/gpio_defaults[8]
+ gpio_defaults_block_35/gpio_defaults[9] housekeeping/mgmt_gpio_in[35] housekeeping/mgmt_gpio_oeb[35]
+ housekeeping/mgmt_gpio_out[35] gpio_control_bidir_2\[0\]/one padframe/mprj_io_analog_en[24]
+ padframe/mprj_io_analog_pol[24] padframe/mprj_io_analog_sel[24] padframe/mprj_io_dm[72]
+ padframe/mprj_io_dm[73] padframe/mprj_io_dm[74] padframe/mprj_io_holdover[24] padframe/mprj_io_ib_mode_sel[24]
+ padframe/mprj_io_in[24] padframe/mprj_io_inp_dis[24] padframe/mprj_io_out[24] padframe/mprj_io_oeb[24]
+ padframe/mprj_io_slow_sel[24] padframe/mprj_io_vtrip_sel[24] gpio_control_bidir_2\[0\]/resetn
+ gpio_control_in_2\[9\]/resetn gpio_control_bidir_2\[0\]/serial_clock gpio_control_in_2\[9\]/serial_clock
+ gpio_control_bidir_2\[0\]/serial_data_in gpio_control_in_2\[9\]/serial_data_in gpio_control_bidir_2\[0\]/serial_load
+ gpio_control_in_2\[9\]/serial_load mprj/io_in[24] mprj/io_oeb[24] mprj/io_out[24]
+ vccd_core vccd1_core VSUBS vssd1_core gpio_control_bidir_2\[0\]/zero gpio_control_block
Xspare_logic_block_0 spare_logic_block_0/spare_xfq[0] spare_logic_block_0/spare_xfq[1]
+ spare_logic_block_0/spare_xfqn[0] spare_logic_block_0/spare_xfqn[1] spare_logic_block_0/spare_xi[0]
+ spare_logic_block_0/spare_xi[1] spare_logic_block_0/spare_xi[2] spare_logic_block_0/spare_xi[3]
+ spare_logic_block_0/spare_xib spare_logic_block_0/spare_xmx[0] spare_logic_block_0/spare_xmx[1]
+ spare_logic_block_0/spare_xna[0] spare_logic_block_0/spare_xna[1] spare_logic_block_0/spare_xno[0]
+ spare_logic_block_0/spare_xno[1] spare_logic_block_0/spare_xz[0] spare_logic_block_0/spare_xz[10]
+ spare_logic_block_0/spare_xz[11] spare_logic_block_0/spare_xz[12] spare_logic_block_0/spare_xz[13]
+ spare_logic_block_0/spare_xz[14] spare_logic_block_0/spare_xz[15] spare_logic_block_0/spare_xz[16]
+ spare_logic_block_0/spare_xz[17] spare_logic_block_0/spare_xz[18] spare_logic_block_0/spare_xz[19]
+ spare_logic_block_0/spare_xz[1] spare_logic_block_0/spare_xz[20] spare_logic_block_0/spare_xz[21]
+ spare_logic_block_0/spare_xz[22] spare_logic_block_0/spare_xz[23] spare_logic_block_0/spare_xz[24]
+ spare_logic_block_0/spare_xz[25] spare_logic_block_0/spare_xz[26] spare_logic_block_0/spare_xz[2]
+ spare_logic_block_0/spare_xz[3] spare_logic_block_0/spare_xz[4] spare_logic_block_0/spare_xz[5]
+ spare_logic_block_0/spare_xz[6] spare_logic_block_0/spare_xz[7] spare_logic_block_0/spare_xz[8]
+ spare_logic_block_0/spare_xz[9] vccd_core VSUBS spare_logic_block
Xsoc VSUBS vccd_core soc/core_clk soc/core_rstn soc/debug_in soc/debug_mode soc/debug_oeb
+ soc/debug_out soc/flash_clk soc/flash_csb soc/flash_io0_di soc/flash_io0_do soc/flash_io0_oeb
+ soc/flash_io1_di soc/flash_io1_do soc/flash_io1_oeb soc/flash_io2_di soc/flash_io2_do
+ soc/flash_io2_oeb soc/flash_io3_di soc/flash_io3_do soc/flash_io3_oeb soc/gpio_in_pad
+ soc/gpio_inenb_pad soc/gpio_mode0_pad soc/gpio_mode1_pad soc/gpio_out_pad soc/gpio_outenb_pad
+ soc/hk_ack_i soc/hk_cyc_o soc/hk_dat_i[0] soc/hk_dat_i[10] soc/hk_dat_i[11] soc/hk_dat_i[12]
+ soc/hk_dat_i[13] soc/hk_dat_i[14] soc/hk_dat_i[15] soc/hk_dat_i[16] soc/hk_dat_i[17]
+ soc/hk_dat_i[18] soc/hk_dat_i[19] soc/hk_dat_i[1] soc/hk_dat_i[20] soc/hk_dat_i[21]
+ soc/hk_dat_i[22] soc/hk_dat_i[23] soc/hk_dat_i[24] soc/hk_dat_i[25] soc/hk_dat_i[26]
+ soc/hk_dat_i[27] soc/hk_dat_i[28] soc/hk_dat_i[29] soc/hk_dat_i[2] soc/hk_dat_i[30]
+ soc/hk_dat_i[31] soc/hk_dat_i[3] soc/hk_dat_i[4] soc/hk_dat_i[5] soc/hk_dat_i[6]
+ soc/hk_dat_i[7] soc/hk_dat_i[8] soc/hk_dat_i[9] soc/hk_stb_o soc/irq[0] soc/irq[1]
+ soc/irq[2] soc/irq[3] soc/irq[4] soc/irq[5] soc/la_iena[0] soc/la_iena[100] soc/la_iena[101]
+ soc/la_iena[102] soc/la_iena[103] soc/la_iena[104] soc/la_iena[105] soc/la_iena[106]
+ soc/la_iena[107] soc/la_iena[108] soc/la_iena[109] soc/la_iena[10] soc/la_iena[110]
+ soc/la_iena[111] soc/la_iena[112] soc/la_iena[113] soc/la_iena[114] soc/la_iena[115]
+ soc/la_iena[116] soc/la_iena[117] soc/la_iena[118] soc/la_iena[119] soc/la_iena[11]
+ soc/la_iena[120] soc/la_iena[121] soc/la_iena[122] soc/la_iena[123] soc/la_iena[124]
+ soc/la_iena[125] soc/la_iena[126] soc/la_iena[127] soc/la_iena[12] soc/la_iena[13]
+ soc/la_iena[14] soc/la_iena[15] soc/la_iena[16] soc/la_iena[17] soc/la_iena[18]
+ soc/la_iena[19] soc/la_iena[1] soc/la_iena[20] soc/la_iena[21] soc/la_iena[22] soc/la_iena[23]
+ soc/la_iena[24] soc/la_iena[25] soc/la_iena[26] soc/la_iena[27] soc/la_iena[28]
+ soc/la_iena[29] soc/la_iena[2] soc/la_iena[30] soc/la_iena[31] soc/la_iena[32] soc/la_iena[33]
+ soc/la_iena[34] soc/la_iena[35] soc/la_iena[36] soc/la_iena[37] soc/la_iena[38]
+ soc/la_iena[39] soc/la_iena[3] soc/la_iena[40] soc/la_iena[41] soc/la_iena[42] soc/la_iena[43]
+ soc/la_iena[44] soc/la_iena[45] soc/la_iena[46] soc/la_iena[47] soc/la_iena[48]
+ soc/la_iena[49] soc/la_iena[4] soc/la_iena[50] soc/la_iena[51] soc/la_iena[52] soc/la_iena[53]
+ soc/la_iena[54] soc/la_iena[55] soc/la_iena[56] soc/la_iena[57] soc/la_iena[58]
+ soc/la_iena[59] soc/la_iena[5] soc/la_iena[60] soc/la_iena[61] soc/la_iena[62] soc/la_iena[63]
+ soc/la_iena[64] soc/la_iena[65] soc/la_iena[66] soc/la_iena[67] soc/la_iena[68]
+ soc/la_iena[69] soc/la_iena[6] soc/la_iena[70] soc/la_iena[71] soc/la_iena[72] soc/la_iena[73]
+ soc/la_iena[74] soc/la_iena[75] soc/la_iena[76] soc/la_iena[77] soc/la_iena[78]
+ soc/la_iena[79] soc/la_iena[7] soc/la_iena[80] soc/la_iena[81] soc/la_iena[82] soc/la_iena[83]
+ soc/la_iena[84] soc/la_iena[85] soc/la_iena[86] soc/la_iena[87] soc/la_iena[88]
+ soc/la_iena[89] soc/la_iena[8] soc/la_iena[90] soc/la_iena[91] soc/la_iena[92] soc/la_iena[93]
+ soc/la_iena[94] soc/la_iena[95] soc/la_iena[96] soc/la_iena[97] soc/la_iena[98]
+ soc/la_iena[99] soc/la_iena[9] soc/la_input[0] soc/la_input[100] soc/la_input[101]
+ soc/la_input[102] soc/la_input[103] soc/la_input[104] soc/la_input[105] soc/la_input[106]
+ soc/la_input[107] soc/la_input[108] soc/la_input[109] soc/la_input[10] soc/la_input[110]
+ soc/la_input[111] soc/la_input[112] soc/la_input[113] soc/la_input[114] soc/la_input[115]
+ soc/la_input[116] soc/la_input[117] soc/la_input[118] soc/la_input[119] soc/la_input[11]
+ soc/la_input[120] soc/la_input[121] soc/la_input[122] soc/la_input[123] soc/la_input[124]
+ soc/la_input[125] soc/la_input[126] soc/la_input[127] soc/la_input[12] soc/la_input[13]
+ soc/la_input[14] soc/la_input[15] soc/la_input[16] soc/la_input[17] soc/la_input[18]
+ soc/la_input[19] soc/la_input[1] soc/la_input[20] soc/la_input[21] soc/la_input[22]
+ soc/la_input[23] soc/la_input[24] soc/la_input[25] soc/la_input[26] soc/la_input[27]
+ soc/la_input[28] soc/la_input[29] soc/la_input[2] soc/la_input[30] soc/la_input[31]
+ soc/la_input[32] soc/la_input[33] soc/la_input[34] soc/la_input[35] soc/la_input[36]
+ soc/la_input[37] soc/la_input[38] soc/la_input[39] soc/la_input[3] soc/la_input[40]
+ soc/la_input[41] soc/la_input[42] soc/la_input[43] soc/la_input[44] soc/la_input[45]
+ soc/la_input[46] soc/la_input[47] soc/la_input[48] soc/la_input[49] soc/la_input[4]
+ soc/la_input[50] soc/la_input[51] soc/la_input[52] soc/la_input[53] soc/la_input[54]
+ soc/la_input[55] soc/la_input[56] soc/la_input[57] soc/la_input[58] soc/la_input[59]
+ soc/la_input[5] soc/la_input[60] soc/la_input[61] soc/la_input[62] soc/la_input[63]
+ soc/la_input[64] soc/la_input[65] soc/la_input[66] soc/la_input[67] soc/la_input[68]
+ soc/la_input[69] soc/la_input[6] soc/la_input[70] soc/la_input[71] soc/la_input[72]
+ soc/la_input[73] soc/la_input[74] soc/la_input[75] soc/la_input[76] soc/la_input[77]
+ soc/la_input[78] soc/la_input[79] soc/la_input[7] soc/la_input[80] soc/la_input[81]
+ soc/la_input[82] soc/la_input[83] soc/la_input[84] soc/la_input[85] soc/la_input[86]
+ soc/la_input[87] soc/la_input[88] soc/la_input[89] soc/la_input[8] soc/la_input[90]
+ soc/la_input[91] soc/la_input[92] soc/la_input[93] soc/la_input[94] soc/la_input[95]
+ soc/la_input[96] soc/la_input[97] soc/la_input[98] soc/la_input[99] soc/la_input[9]
+ soc/la_oenb[0] soc/la_oenb[100] soc/la_oenb[101] soc/la_oenb[102] soc/la_oenb[103]
+ soc/la_oenb[104] soc/la_oenb[105] soc/la_oenb[106] soc/la_oenb[107] soc/la_oenb[108]
+ soc/la_oenb[109] soc/la_oenb[10] soc/la_oenb[110] soc/la_oenb[111] soc/la_oenb[112]
+ soc/la_oenb[113] soc/la_oenb[114] soc/la_oenb[115] soc/la_oenb[116] soc/la_oenb[117]
+ soc/la_oenb[118] soc/la_oenb[119] soc/la_oenb[11] soc/la_oenb[120] soc/la_oenb[121]
+ soc/la_oenb[122] soc/la_oenb[123] soc/la_oenb[124] soc/la_oenb[125] soc/la_oenb[126]
+ soc/la_oenb[127] soc/la_oenb[12] soc/la_oenb[13] soc/la_oenb[14] soc/la_oenb[15]
+ soc/la_oenb[16] soc/la_oenb[17] soc/la_oenb[18] soc/la_oenb[19] soc/la_oenb[1] soc/la_oenb[20]
+ soc/la_oenb[21] soc/la_oenb[22] soc/la_oenb[23] soc/la_oenb[24] soc/la_oenb[25]
+ soc/la_oenb[26] soc/la_oenb[27] soc/la_oenb[28] soc/la_oenb[29] soc/la_oenb[2] soc/la_oenb[30]
+ soc/la_oenb[31] soc/la_oenb[32] soc/la_oenb[33] soc/la_oenb[34] soc/la_oenb[35]
+ soc/la_oenb[36] soc/la_oenb[37] soc/la_oenb[38] soc/la_oenb[39] soc/la_oenb[3] soc/la_oenb[40]
+ soc/la_oenb[41] soc/la_oenb[42] soc/la_oenb[43] soc/la_oenb[44] soc/la_oenb[45]
+ soc/la_oenb[46] soc/la_oenb[47] soc/la_oenb[48] soc/la_oenb[49] soc/la_oenb[4] soc/la_oenb[50]
+ soc/la_oenb[51] soc/la_oenb[52] soc/la_oenb[53] soc/la_oenb[54] soc/la_oenb[55]
+ soc/la_oenb[56] soc/la_oenb[57] soc/la_oenb[58] soc/la_oenb[59] soc/la_oenb[5] soc/la_oenb[60]
+ soc/la_oenb[61] soc/la_oenb[62] soc/la_oenb[63] soc/la_oenb[64] soc/la_oenb[65]
+ soc/la_oenb[66] soc/la_oenb[67] soc/la_oenb[68] soc/la_oenb[69] soc/la_oenb[6] soc/la_oenb[70]
+ soc/la_oenb[71] soc/la_oenb[72] soc/la_oenb[73] soc/la_oenb[74] soc/la_oenb[75]
+ soc/la_oenb[76] soc/la_oenb[77] soc/la_oenb[78] soc/la_oenb[79] soc/la_oenb[7] soc/la_oenb[80]
+ soc/la_oenb[81] soc/la_oenb[82] soc/la_oenb[83] soc/la_oenb[84] soc/la_oenb[85]
+ soc/la_oenb[86] soc/la_oenb[87] soc/la_oenb[88] soc/la_oenb[89] soc/la_oenb[8] soc/la_oenb[90]
+ soc/la_oenb[91] soc/la_oenb[92] soc/la_oenb[93] soc/la_oenb[94] soc/la_oenb[95]
+ soc/la_oenb[96] soc/la_oenb[97] soc/la_oenb[98] soc/la_oenb[99] soc/la_oenb[9] soc/la_output[0]
+ soc/la_output[100] soc/la_output[101] soc/la_output[102] soc/la_output[103] soc/la_output[104]
+ soc/la_output[105] soc/la_output[106] soc/la_output[107] soc/la_output[108] soc/la_output[109]
+ soc/la_output[10] soc/la_output[110] soc/la_output[111] soc/la_output[112] soc/la_output[113]
+ soc/la_output[114] soc/la_output[115] soc/la_output[116] soc/la_output[117] soc/la_output[118]
+ soc/la_output[119] soc/la_output[11] soc/la_output[120] soc/la_output[121] soc/la_output[122]
+ soc/la_output[123] soc/la_output[124] soc/la_output[125] soc/la_output[126] soc/la_output[127]
+ soc/la_output[12] soc/la_output[13] soc/la_output[14] soc/la_output[15] soc/la_output[16]
+ soc/la_output[17] soc/la_output[18] soc/la_output[19] soc/la_output[1] soc/la_output[20]
+ soc/la_output[21] soc/la_output[22] soc/la_output[23] soc/la_output[24] soc/la_output[25]
+ soc/la_output[26] soc/la_output[27] soc/la_output[28] soc/la_output[29] soc/la_output[2]
+ soc/la_output[30] soc/la_output[31] soc/la_output[32] soc/la_output[33] soc/la_output[34]
+ soc/la_output[35] soc/la_output[36] soc/la_output[37] soc/la_output[38] soc/la_output[39]
+ soc/la_output[3] soc/la_output[40] soc/la_output[41] soc/la_output[42] soc/la_output[43]
+ soc/la_output[44] soc/la_output[45] soc/la_output[46] soc/la_output[47] soc/la_output[48]
+ soc/la_output[49] soc/la_output[4] soc/la_output[50] soc/la_output[51] soc/la_output[52]
+ soc/la_output[53] soc/la_output[54] soc/la_output[55] soc/la_output[56] soc/la_output[57]
+ soc/la_output[58] soc/la_output[59] soc/la_output[5] soc/la_output[60] soc/la_output[61]
+ soc/la_output[62] soc/la_output[63] soc/la_output[64] soc/la_output[65] soc/la_output[66]
+ soc/la_output[67] soc/la_output[68] soc/la_output[69] soc/la_output[6] soc/la_output[70]
+ soc/la_output[71] soc/la_output[72] soc/la_output[73] soc/la_output[74] soc/la_output[75]
+ soc/la_output[76] soc/la_output[77] soc/la_output[78] soc/la_output[79] soc/la_output[7]
+ soc/la_output[80] soc/la_output[81] soc/la_output[82] soc/la_output[83] soc/la_output[84]
+ soc/la_output[85] soc/la_output[86] soc/la_output[87] soc/la_output[88] soc/la_output[89]
+ soc/la_output[8] soc/la_output[90] soc/la_output[91] soc/la_output[92] soc/la_output[93]
+ soc/la_output[94] soc/la_output[95] soc/la_output[96] soc/la_output[97] soc/la_output[98]
+ soc/la_output[99] soc/la_output[9] soc/mprj_ack_i soc/mprj_adr_o[0] soc/mprj_adr_o[10]
+ soc/mprj_adr_o[11] soc/mprj_adr_o[12] soc/mprj_adr_o[13] soc/mprj_adr_o[14] soc/mprj_adr_o[15]
+ soc/mprj_adr_o[16] soc/mprj_adr_o[17] soc/mprj_adr_o[18] soc/mprj_adr_o[19] soc/mprj_adr_o[1]
+ soc/mprj_adr_o[20] soc/mprj_adr_o[21] soc/mprj_adr_o[22] soc/mprj_adr_o[23] soc/mprj_adr_o[24]
+ soc/mprj_adr_o[25] soc/mprj_adr_o[26] soc/mprj_adr_o[27] soc/mprj_adr_o[28] soc/mprj_adr_o[29]
+ soc/mprj_adr_o[2] soc/mprj_adr_o[30] soc/mprj_adr_o[31] soc/mprj_adr_o[3] soc/mprj_adr_o[4]
+ soc/mprj_adr_o[5] soc/mprj_adr_o[6] soc/mprj_adr_o[7] soc/mprj_adr_o[8] soc/mprj_adr_o[9]
+ soc/mprj_cyc_o soc/mprj_dat_i[0] soc/mprj_dat_i[10] soc/mprj_dat_i[11] soc/mprj_dat_i[12]
+ soc/mprj_dat_i[13] soc/mprj_dat_i[14] soc/mprj_dat_i[15] soc/mprj_dat_i[16] soc/mprj_dat_i[17]
+ soc/mprj_dat_i[18] soc/mprj_dat_i[19] soc/mprj_dat_i[1] soc/mprj_dat_i[20] soc/mprj_dat_i[21]
+ soc/mprj_dat_i[22] soc/mprj_dat_i[23] soc/mprj_dat_i[24] soc/mprj_dat_i[25] soc/mprj_dat_i[26]
+ soc/mprj_dat_i[27] soc/mprj_dat_i[28] soc/mprj_dat_i[29] soc/mprj_dat_i[2] soc/mprj_dat_i[30]
+ soc/mprj_dat_i[31] soc/mprj_dat_i[3] soc/mprj_dat_i[4] soc/mprj_dat_i[5] soc/mprj_dat_i[6]
+ soc/mprj_dat_i[7] soc/mprj_dat_i[8] soc/mprj_dat_i[9] soc/mprj_dat_o[0] soc/mprj_dat_o[10]
+ soc/mprj_dat_o[11] soc/mprj_dat_o[12] soc/mprj_dat_o[13] soc/mprj_dat_o[14] soc/mprj_dat_o[15]
+ soc/mprj_dat_o[16] soc/mprj_dat_o[17] soc/mprj_dat_o[18] soc/mprj_dat_o[19] soc/mprj_dat_o[1]
+ soc/mprj_dat_o[20] soc/mprj_dat_o[21] soc/mprj_dat_o[22] soc/mprj_dat_o[23] soc/mprj_dat_o[24]
+ soc/mprj_dat_o[25] soc/mprj_dat_o[26] soc/mprj_dat_o[27] soc/mprj_dat_o[28] soc/mprj_dat_o[29]
+ soc/mprj_dat_o[2] soc/mprj_dat_o[30] soc/mprj_dat_o[31] soc/mprj_dat_o[3] soc/mprj_dat_o[4]
+ soc/mprj_dat_o[5] soc/mprj_dat_o[6] soc/mprj_dat_o[7] soc/mprj_dat_o[8] soc/mprj_dat_o[9]
+ soc/mprj_sel_o[0] soc/mprj_sel_o[1] soc/mprj_sel_o[2] soc/mprj_sel_o[3] soc/mprj_stb_o
+ soc/mprj_wb_iena soc/mprj_we_o soc/qspi_enabled soc/ser_rx soc/ser_tx soc/spi_csb
+ soc/spi_enabled soc/spi_sck soc/spi_sdi soc/spi_sdo soc/spi_sdoenb soc/sram_ro_addr[0]
+ soc/sram_ro_addr[1] soc/sram_ro_addr[2] soc/sram_ro_addr[3] soc/sram_ro_addr[4]
+ soc/sram_ro_addr[5] soc/sram_ro_addr[6] soc/sram_ro_addr[7] soc/sram_ro_clk soc/sram_ro_csb
+ soc/sram_ro_data[0] soc/sram_ro_data[10] soc/sram_ro_data[11] soc/sram_ro_data[12]
+ soc/sram_ro_data[13] soc/sram_ro_data[14] soc/sram_ro_data[15] soc/sram_ro_data[16]
+ soc/sram_ro_data[17] soc/sram_ro_data[18] soc/sram_ro_data[19] soc/sram_ro_data[1]
+ soc/sram_ro_data[20] soc/sram_ro_data[21] soc/sram_ro_data[22] soc/sram_ro_data[23]
+ soc/sram_ro_data[24] soc/sram_ro_data[25] soc/sram_ro_data[26] soc/sram_ro_data[27]
+ soc/sram_ro_data[28] soc/sram_ro_data[29] soc/sram_ro_data[2] soc/sram_ro_data[30]
+ soc/sram_ro_data[31] soc/sram_ro_data[3] soc/sram_ro_data[4] soc/sram_ro_data[5]
+ soc/sram_ro_data[6] soc/sram_ro_data[7] soc/sram_ro_data[8] soc/sram_ro_data[9]
+ soc/trap soc/uart_enabled soc/user_irq_ena[0] soc/user_irq_ena[1] soc/user_irq_ena[2]
+ mgmt_core_wrapper
Xgpio_defaults_block_14 VSUBS vccd_core gpio_defaults_block_14/gpio_defaults[0] gpio_defaults_block_14/gpio_defaults[10]
+ gpio_defaults_block_14/gpio_defaults[11] gpio_defaults_block_14/gpio_defaults[12]
+ gpio_defaults_block_14/gpio_defaults[1] gpio_defaults_block_14/gpio_defaults[2]
+ gpio_defaults_block_14/gpio_defaults[3] gpio_defaults_block_14/gpio_defaults[4]
+ gpio_defaults_block_14/gpio_defaults[5] gpio_defaults_block_14/gpio_defaults[6]
+ gpio_defaults_block_14/gpio_defaults[7] gpio_defaults_block_14/gpio_defaults[8]
+ gpio_defaults_block_14/gpio_defaults[9] gpio_defaults_block
Xgpio_control_in_2\[9\] gpio_defaults_block_34/gpio_defaults[0] gpio_defaults_block_34/gpio_defaults[10]
+ gpio_defaults_block_34/gpio_defaults[11] gpio_defaults_block_34/gpio_defaults[12]
+ gpio_defaults_block_34/gpio_defaults[1] gpio_defaults_block_34/gpio_defaults[2]
+ gpio_defaults_block_34/gpio_defaults[3] gpio_defaults_block_34/gpio_defaults[4]
+ gpio_defaults_block_34/gpio_defaults[5] gpio_defaults_block_34/gpio_defaults[6]
+ gpio_defaults_block_34/gpio_defaults[7] gpio_defaults_block_34/gpio_defaults[8]
+ gpio_defaults_block_34/gpio_defaults[9] housekeeping/mgmt_gpio_in[34] gpio_control_in_2\[9\]/one
+ housekeeping/mgmt_gpio_in[34] gpio_control_in_2\[9\]/one padframe/mprj_io_analog_en[23]
+ padframe/mprj_io_analog_pol[23] padframe/mprj_io_analog_sel[23] padframe/mprj_io_dm[69]
+ padframe/mprj_io_dm[70] padframe/mprj_io_dm[71] padframe/mprj_io_holdover[23] padframe/mprj_io_ib_mode_sel[23]
+ padframe/mprj_io_in[23] padframe/mprj_io_inp_dis[23] padframe/mprj_io_out[23] padframe/mprj_io_oeb[23]
+ padframe/mprj_io_slow_sel[23] padframe/mprj_io_vtrip_sel[23] gpio_control_in_2\[9\]/resetn
+ gpio_control_in_2\[8\]/resetn gpio_control_in_2\[9\]/serial_clock gpio_control_in_2\[8\]/serial_clock
+ gpio_control_in_2\[9\]/serial_data_in gpio_control_in_2\[8\]/serial_data_in gpio_control_in_2\[9\]/serial_load
+ gpio_control_in_2\[8\]/serial_load mprj/io_in[23] mprj/io_oeb[23] mprj/io_out[23]
+ vccd_core vccd1_core VSUBS vssd1_core gpio_control_in_2\[9\]/zero gpio_control_block
Xgpio_defaults_block_36 VSUBS vccd_core gpio_defaults_block_36/gpio_defaults[0] gpio_defaults_block_36/gpio_defaults[10]
+ gpio_defaults_block_36/gpio_defaults[11] gpio_defaults_block_36/gpio_defaults[12]
+ gpio_defaults_block_36/gpio_defaults[1] gpio_defaults_block_36/gpio_defaults[2]
+ gpio_defaults_block_36/gpio_defaults[3] gpio_defaults_block_36/gpio_defaults[4]
+ gpio_defaults_block_36/gpio_defaults[5] gpio_defaults_block_36/gpio_defaults[6]
+ gpio_defaults_block_36/gpio_defaults[7] gpio_defaults_block_36/gpio_defaults[8]
+ gpio_defaults_block_36/gpio_defaults[9] gpio_defaults_block
Xspare_logic_block_1 spare_logic_block_1/spare_xfq[0] spare_logic_block_1/spare_xfq[1]
+ spare_logic_block_1/spare_xfqn[0] spare_logic_block_1/spare_xfqn[1] spare_logic_block_1/spare_xi[0]
+ spare_logic_block_1/spare_xi[1] spare_logic_block_1/spare_xi[2] spare_logic_block_1/spare_xi[3]
+ spare_logic_block_1/spare_xib spare_logic_block_1/spare_xmx[0] spare_logic_block_1/spare_xmx[1]
+ spare_logic_block_1/spare_xna[0] spare_logic_block_1/spare_xna[1] spare_logic_block_1/spare_xno[0]
+ spare_logic_block_1/spare_xno[1] spare_logic_block_1/spare_xz[0] spare_logic_block_1/spare_xz[10]
+ spare_logic_block_1/spare_xz[11] spare_logic_block_1/spare_xz[12] spare_logic_block_1/spare_xz[13]
+ spare_logic_block_1/spare_xz[14] spare_logic_block_1/spare_xz[15] spare_logic_block_1/spare_xz[16]
+ spare_logic_block_1/spare_xz[17] spare_logic_block_1/spare_xz[18] spare_logic_block_1/spare_xz[19]
+ spare_logic_block_1/spare_xz[1] spare_logic_block_1/spare_xz[20] spare_logic_block_1/spare_xz[21]
+ spare_logic_block_1/spare_xz[22] spare_logic_block_1/spare_xz[23] spare_logic_block_1/spare_xz[24]
+ spare_logic_block_1/spare_xz[25] spare_logic_block_1/spare_xz[26] spare_logic_block_1/spare_xz[2]
+ spare_logic_block_1/spare_xz[3] spare_logic_block_1/spare_xz[4] spare_logic_block_1/spare_xz[5]
+ spare_logic_block_1/spare_xz[6] spare_logic_block_1/spare_xz[7] spare_logic_block_1/spare_xz[8]
+ spare_logic_block_1/spare_xz[9] vccd_core VSUBS spare_logic_block
Xgpio_defaults_block_26 VSUBS vccd_core gpio_defaults_block_26/gpio_defaults[0] gpio_defaults_block_26/gpio_defaults[10]
+ gpio_defaults_block_26/gpio_defaults[11] gpio_defaults_block_26/gpio_defaults[12]
+ gpio_defaults_block_26/gpio_defaults[1] gpio_defaults_block_26/gpio_defaults[2]
+ gpio_defaults_block_26/gpio_defaults[3] gpio_defaults_block_26/gpio_defaults[4]
+ gpio_defaults_block_26/gpio_defaults[5] gpio_defaults_block_26/gpio_defaults[6]
+ gpio_defaults_block_26/gpio_defaults[7] gpio_defaults_block_26/gpio_defaults[8]
+ gpio_defaults_block_26/gpio_defaults[9] gpio_defaults_block
Xgpio_control_in_1\[4\] gpio_defaults_block_12/gpio_defaults[0] gpio_defaults_block_12/gpio_defaults[10]
+ gpio_defaults_block_12/gpio_defaults[11] gpio_defaults_block_12/gpio_defaults[12]
+ gpio_defaults_block_12/gpio_defaults[1] gpio_defaults_block_12/gpio_defaults[2]
+ gpio_defaults_block_12/gpio_defaults[3] gpio_defaults_block_12/gpio_defaults[4]
+ gpio_defaults_block_12/gpio_defaults[5] gpio_defaults_block_12/gpio_defaults[6]
+ gpio_defaults_block_12/gpio_defaults[7] gpio_defaults_block_12/gpio_defaults[8]
+ gpio_defaults_block_12/gpio_defaults[9] housekeeping/mgmt_gpio_in[12] gpio_control_in_1\[4\]/one
+ housekeeping/mgmt_gpio_in[12] gpio_control_in_1\[4\]/one padframe/mprj_io_analog_en[12]
+ padframe/mprj_io_analog_pol[12] padframe/mprj_io_analog_sel[12] padframe/mprj_io_dm[36]
+ padframe/mprj_io_dm[37] padframe/mprj_io_dm[38] padframe/mprj_io_holdover[12] padframe/mprj_io_ib_mode_sel[12]
+ padframe/mprj_io_in[12] padframe/mprj_io_inp_dis[12] padframe/mprj_io_out[12] padframe/mprj_io_oeb[12]
+ padframe/mprj_io_slow_sel[12] padframe/mprj_io_vtrip_sel[12] gpio_control_in_1\[4\]/resetn
+ gpio_control_in_1\[5\]/resetn gpio_control_in_1\[4\]/serial_clock gpio_control_in_1\[5\]/serial_clock
+ gpio_control_in_1\[4\]/serial_data_in gpio_control_in_1\[5\]/serial_data_in gpio_control_in_1\[4\]/serial_load
+ gpio_control_in_1\[5\]/serial_load mprj/io_in[12] mprj/io_oeb[12] mprj/io_out[12]
+ vccd_core vccd1_core VSUBS vssd1_core gpio_control_in_1\[4\]/zero gpio_control_block
Xspare_logic_block_2 spare_logic_block_2/spare_xfq[0] spare_logic_block_2/spare_xfq[1]
+ spare_logic_block_2/spare_xfqn[0] spare_logic_block_2/spare_xfqn[1] spare_logic_block_2/spare_xi[0]
+ spare_logic_block_2/spare_xi[1] spare_logic_block_2/spare_xi[2] spare_logic_block_2/spare_xi[3]
+ spare_logic_block_2/spare_xib spare_logic_block_2/spare_xmx[0] spare_logic_block_2/spare_xmx[1]
+ spare_logic_block_2/spare_xna[0] spare_logic_block_2/spare_xna[1] spare_logic_block_2/spare_xno[0]
+ spare_logic_block_2/spare_xno[1] spare_logic_block_2/spare_xz[0] spare_logic_block_2/spare_xz[10]
+ spare_logic_block_2/spare_xz[11] spare_logic_block_2/spare_xz[12] spare_logic_block_2/spare_xz[13]
+ spare_logic_block_2/spare_xz[14] spare_logic_block_2/spare_xz[15] spare_logic_block_2/spare_xz[16]
+ spare_logic_block_2/spare_xz[17] spare_logic_block_2/spare_xz[18] spare_logic_block_2/spare_xz[19]
+ spare_logic_block_2/spare_xz[1] spare_logic_block_2/spare_xz[20] spare_logic_block_2/spare_xz[21]
+ spare_logic_block_2/spare_xz[22] spare_logic_block_2/spare_xz[23] spare_logic_block_2/spare_xz[24]
+ spare_logic_block_2/spare_xz[25] spare_logic_block_2/spare_xz[26] spare_logic_block_2/spare_xz[2]
+ spare_logic_block_2/spare_xz[3] spare_logic_block_2/spare_xz[4] spare_logic_block_2/spare_xz[5]
+ spare_logic_block_2/spare_xz[6] spare_logic_block_2/spare_xz[7] spare_logic_block_2/spare_xz[8]
+ spare_logic_block_2/spare_xz[9] vccd_core VSUBS spare_logic_block
Xgpio_defaults_block_37 VSUBS vccd_core gpio_defaults_block_37/gpio_defaults[0] gpio_defaults_block_37/gpio_defaults[10]
+ gpio_defaults_block_37/gpio_defaults[11] gpio_defaults_block_37/gpio_defaults[12]
+ gpio_defaults_block_37/gpio_defaults[1] gpio_defaults_block_37/gpio_defaults[2]
+ gpio_defaults_block_37/gpio_defaults[3] gpio_defaults_block_37/gpio_defaults[4]
+ gpio_defaults_block_37/gpio_defaults[5] gpio_defaults_block_37/gpio_defaults[6]
+ gpio_defaults_block_37/gpio_defaults[7] gpio_defaults_block_37/gpio_defaults[8]
+ gpio_defaults_block_37/gpio_defaults[9] gpio_defaults_block
Xpor por/vdd3v3 vccd_core por/vss3v3 por/porb_h por/por_l por/porb_l VSUBS simple_por
Xgpio_defaults_block_27 VSUBS vccd_core gpio_defaults_block_27/gpio_defaults[0] gpio_defaults_block_27/gpio_defaults[10]
+ gpio_defaults_block_27/gpio_defaults[11] gpio_defaults_block_27/gpio_defaults[12]
+ gpio_defaults_block_27/gpio_defaults[1] gpio_defaults_block_27/gpio_defaults[2]
+ gpio_defaults_block_27/gpio_defaults[3] gpio_defaults_block_27/gpio_defaults[4]
+ gpio_defaults_block_27/gpio_defaults[5] gpio_defaults_block_27/gpio_defaults[6]
+ gpio_defaults_block_27/gpio_defaults[7] gpio_defaults_block_27/gpio_defaults[8]
+ gpio_defaults_block_27/gpio_defaults[9] gpio_defaults_block
Xgpio_control_in_1a\[1\] gpio_defaults_block_3/gpio_defaults[0] gpio_defaults_block_3/gpio_defaults[10]
+ gpio_defaults_block_3/gpio_defaults[11] gpio_defaults_block_3/gpio_defaults[12]
+ gpio_defaults_block_3/gpio_defaults[1] gpio_defaults_block_3/gpio_defaults[2] gpio_defaults_block_3/gpio_defaults[3]
+ gpio_defaults_block_3/gpio_defaults[4] gpio_defaults_block_3/gpio_defaults[5] gpio_defaults_block_3/gpio_defaults[6]
+ gpio_defaults_block_3/gpio_defaults[7] gpio_defaults_block_3/gpio_defaults[8] gpio_defaults_block_3/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[3] gpio_control_in_1a\[1\]/one housekeeping/mgmt_gpio_in[3]
+ gpio_control_in_1a\[1\]/one padframe/mprj_io_analog_en[3] padframe/mprj_io_analog_pol[3]
+ padframe/mprj_io_analog_sel[3] padframe/mprj_io_dm[9] padframe/mprj_io_dm[10] padframe/mprj_io_dm[11]
+ padframe/mprj_io_holdover[3] padframe/mprj_io_ib_mode_sel[3] padframe/mprj_io_in[3]
+ padframe/mprj_io_inp_dis[3] padframe/mprj_io_out[3] padframe/mprj_io_oeb[3] padframe/mprj_io_slow_sel[3]
+ padframe/mprj_io_vtrip_sel[3] gpio_control_in_1a\[1\]/resetn gpio_control_in_1a\[2\]/resetn
+ gpio_control_in_1a\[1\]/serial_clock gpio_control_in_1a\[2\]/serial_clock gpio_control_in_1a\[1\]/serial_data_in
+ gpio_control_in_1a\[2\]/serial_data_in gpio_control_in_1a\[1\]/serial_load gpio_control_in_1a\[2\]/serial_load
+ mprj/io_in[3] mprj/io_oeb[3] mprj/io_out[3] vccd_core vccd1_core VSUBS vssd1_core
+ gpio_control_in_1a\[1\]/zero gpio_control_block
Xspare_logic_block_3 spare_logic_block_3/spare_xfq[0] spare_logic_block_3/spare_xfq[1]
+ spare_logic_block_3/spare_xfqn[0] spare_logic_block_3/spare_xfqn[1] spare_logic_block_3/spare_xi[0]
+ spare_logic_block_3/spare_xi[1] spare_logic_block_3/spare_xi[2] spare_logic_block_3/spare_xi[3]
+ spare_logic_block_3/spare_xib spare_logic_block_3/spare_xmx[0] spare_logic_block_3/spare_xmx[1]
+ spare_logic_block_3/spare_xna[0] spare_logic_block_3/spare_xna[1] spare_logic_block_3/spare_xno[0]
+ spare_logic_block_3/spare_xno[1] spare_logic_block_3/spare_xz[0] spare_logic_block_3/spare_xz[10]
+ spare_logic_block_3/spare_xz[11] spare_logic_block_3/spare_xz[12] spare_logic_block_3/spare_xz[13]
+ spare_logic_block_3/spare_xz[14] spare_logic_block_3/spare_xz[15] spare_logic_block_3/spare_xz[16]
+ spare_logic_block_3/spare_xz[17] spare_logic_block_3/spare_xz[18] spare_logic_block_3/spare_xz[19]
+ spare_logic_block_3/spare_xz[1] spare_logic_block_3/spare_xz[20] spare_logic_block_3/spare_xz[21]
+ spare_logic_block_3/spare_xz[22] spare_logic_block_3/spare_xz[23] spare_logic_block_3/spare_xz[24]
+ spare_logic_block_3/spare_xz[25] spare_logic_block_3/spare_xz[26] spare_logic_block_3/spare_xz[2]
+ spare_logic_block_3/spare_xz[3] spare_logic_block_3/spare_xz[4] spare_logic_block_3/spare_xz[5]
+ spare_logic_block_3/spare_xz[6] spare_logic_block_3/spare_xz[7] spare_logic_block_3/spare_xz[8]
+ spare_logic_block_3/spare_xz[9] vccd_core VSUBS spare_logic_block
Xgpio_defaults_block_28 VSUBS vccd_core gpio_defaults_block_28/gpio_defaults[0] gpio_defaults_block_28/gpio_defaults[10]
+ gpio_defaults_block_28/gpio_defaults[11] gpio_defaults_block_28/gpio_defaults[12]
+ gpio_defaults_block_28/gpio_defaults[1] gpio_defaults_block_28/gpio_defaults[2]
+ gpio_defaults_block_28/gpio_defaults[3] gpio_defaults_block_28/gpio_defaults[4]
+ gpio_defaults_block_28/gpio_defaults[5] gpio_defaults_block_28/gpio_defaults[6]
+ gpio_defaults_block_28/gpio_defaults[7] gpio_defaults_block_28/gpio_defaults[8]
+ gpio_defaults_block_28/gpio_defaults[9] gpio_defaults_block
Xgpio_control_in_2\[7\] gpio_defaults_block_32/gpio_defaults[0] gpio_defaults_block_32/gpio_defaults[10]
+ gpio_defaults_block_32/gpio_defaults[11] gpio_defaults_block_32/gpio_defaults[12]
+ gpio_defaults_block_32/gpio_defaults[1] gpio_defaults_block_32/gpio_defaults[2]
+ gpio_defaults_block_32/gpio_defaults[3] gpio_defaults_block_32/gpio_defaults[4]
+ gpio_defaults_block_32/gpio_defaults[5] gpio_defaults_block_32/gpio_defaults[6]
+ gpio_defaults_block_32/gpio_defaults[7] gpio_defaults_block_32/gpio_defaults[8]
+ gpio_defaults_block_32/gpio_defaults[9] housekeeping/mgmt_gpio_in[32] gpio_control_in_2\[7\]/one
+ housekeeping/mgmt_gpio_in[32] gpio_control_in_2\[7\]/one padframe/mprj_io_analog_en[21]
+ padframe/mprj_io_analog_pol[21] padframe/mprj_io_analog_sel[21] padframe/mprj_io_dm[63]
+ padframe/mprj_io_dm[64] padframe/mprj_io_dm[65] padframe/mprj_io_holdover[21] padframe/mprj_io_ib_mode_sel[21]
+ padframe/mprj_io_in[21] padframe/mprj_io_inp_dis[21] padframe/mprj_io_out[21] padframe/mprj_io_oeb[21]
+ padframe/mprj_io_slow_sel[21] padframe/mprj_io_vtrip_sel[21] gpio_control_in_2\[7\]/resetn
+ gpio_control_in_2\[6\]/resetn gpio_control_in_2\[7\]/serial_clock gpio_control_in_2\[6\]/serial_clock
+ gpio_control_in_2\[7\]/serial_data_in gpio_control_in_2\[6\]/serial_data_in gpio_control_in_2\[7\]/serial_load
+ gpio_control_in_2\[6\]/serial_load mprj/io_in[21] mprj/io_oeb[21] mprj/io_out[21]
+ vccd_core vccd1_core VSUBS vssd1_core gpio_control_in_2\[7\]/zero gpio_control_block
Xclocking VSUBS vccd_core soc/core_clk pll/osc clocking/ext_clk_sel housekeeping/reset
+ pll/clockp[1] pll/clockp[0] pll/resetb soc/core_rstn clocking/sel2[0] clocking/sel2[1]
+ clocking/sel2[2] clocking/sel[0] clocking/sel[1] clocking/sel[2] clocking/user_clk
+ caravel_clocking
Xgpio_defaults_block_29 VSUBS vccd_core gpio_defaults_block_29/gpio_defaults[0] gpio_defaults_block_29/gpio_defaults[10]
+ gpio_defaults_block_29/gpio_defaults[11] gpio_defaults_block_29/gpio_defaults[12]
+ gpio_defaults_block_29/gpio_defaults[1] gpio_defaults_block_29/gpio_defaults[2]
+ gpio_defaults_block_29/gpio_defaults[3] gpio_defaults_block_29/gpio_defaults[4]
+ gpio_defaults_block_29/gpio_defaults[5] gpio_defaults_block_29/gpio_defaults[6]
+ gpio_defaults_block_29/gpio_defaults[7] gpio_defaults_block_29/gpio_defaults[8]
+ gpio_defaults_block_29/gpio_defaults[9] gpio_defaults_block
Xgpio_control_in_1\[2\] gpio_defaults_block_10/gpio_defaults[0] gpio_defaults_block_10/gpio_defaults[10]
+ gpio_defaults_block_10/gpio_defaults[11] gpio_defaults_block_10/gpio_defaults[12]
+ gpio_defaults_block_10/gpio_defaults[1] gpio_defaults_block_10/gpio_defaults[2]
+ gpio_defaults_block_10/gpio_defaults[3] gpio_defaults_block_10/gpio_defaults[4]
+ gpio_defaults_block_10/gpio_defaults[5] gpio_defaults_block_10/gpio_defaults[6]
+ gpio_defaults_block_10/gpio_defaults[7] gpio_defaults_block_10/gpio_defaults[8]
+ gpio_defaults_block_10/gpio_defaults[9] housekeeping/mgmt_gpio_in[10] gpio_control_in_1\[2\]/one
+ housekeeping/mgmt_gpio_in[10] gpio_control_in_1\[2\]/one padframe/mprj_io_analog_en[10]
+ padframe/mprj_io_analog_pol[10] padframe/mprj_io_analog_sel[10] padframe/mprj_io_dm[30]
+ padframe/mprj_io_dm[31] padframe/mprj_io_dm[32] padframe/mprj_io_holdover[10] padframe/mprj_io_ib_mode_sel[10]
+ padframe/mprj_io_in[10] padframe/mprj_io_inp_dis[10] padframe/mprj_io_out[10] padframe/mprj_io_oeb[10]
+ padframe/mprj_io_slow_sel[10] padframe/mprj_io_vtrip_sel[10] gpio_control_in_1\[2\]/resetn
+ gpio_control_in_1\[3\]/resetn gpio_control_in_1\[2\]/serial_clock gpio_control_in_1\[3\]/serial_clock
+ gpio_control_in_1\[2\]/serial_data_in gpio_control_in_1\[3\]/serial_data_in gpio_control_in_1\[2\]/serial_load
+ gpio_control_in_1\[3\]/serial_load mprj/io_in[10] mprj/io_oeb[10] mprj/io_out[10]
+ vccd_core vccd1_core VSUBS vssd1_core gpio_control_in_1\[2\]/zero gpio_control_block
Xgpio_control_in_1\[0\] gpio_defaults_block_8/gpio_defaults[0] gpio_defaults_block_8/gpio_defaults[10]
+ gpio_defaults_block_8/gpio_defaults[11] gpio_defaults_block_8/gpio_defaults[12]
+ gpio_defaults_block_8/gpio_defaults[1] gpio_defaults_block_8/gpio_defaults[2] gpio_defaults_block_8/gpio_defaults[3]
+ gpio_defaults_block_8/gpio_defaults[4] gpio_defaults_block_8/gpio_defaults[5] gpio_defaults_block_8/gpio_defaults[6]
+ gpio_defaults_block_8/gpio_defaults[7] gpio_defaults_block_8/gpio_defaults[8] gpio_defaults_block_8/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[8] gpio_control_in_1\[0\]/one housekeeping/mgmt_gpio_in[8]
+ gpio_control_in_1\[0\]/one padframe/mprj_io_analog_en[8] padframe/mprj_io_analog_pol[8]
+ padframe/mprj_io_analog_sel[8] padframe/mprj_io_dm[24] padframe/mprj_io_dm[25] padframe/mprj_io_dm[26]
+ padframe/mprj_io_holdover[8] padframe/mprj_io_ib_mode_sel[8] padframe/mprj_io_in[8]
+ padframe/mprj_io_inp_dis[8] padframe/mprj_io_out[8] padframe/mprj_io_oeb[8] padframe/mprj_io_slow_sel[8]
+ padframe/mprj_io_vtrip_sel[8] gpio_control_in_1\[0\]/resetn gpio_control_in_1\[1\]/resetn
+ gpio_control_in_1\[0\]/serial_clock gpio_control_in_1\[1\]/serial_clock gpio_control_in_1\[0\]/serial_data_in
+ gpio_control_in_1\[1\]/serial_data_in gpio_control_in_1\[0\]/serial_load gpio_control_in_1\[1\]/serial_load
+ mprj/io_in[8] mprj/io_oeb[8] mprj/io_out[8] vccd_core vccd1_core VSUBS vssd1_core
+ gpio_control_in_1\[0\]/zero gpio_control_block
Xgpio_control_in_2\[5\] gpio_defaults_block_30/gpio_defaults[0] gpio_defaults_block_30/gpio_defaults[10]
+ gpio_defaults_block_30/gpio_defaults[11] gpio_defaults_block_30/gpio_defaults[12]
+ gpio_defaults_block_30/gpio_defaults[1] gpio_defaults_block_30/gpio_defaults[2]
+ gpio_defaults_block_30/gpio_defaults[3] gpio_defaults_block_30/gpio_defaults[4]
+ gpio_defaults_block_30/gpio_defaults[5] gpio_defaults_block_30/gpio_defaults[6]
+ gpio_defaults_block_30/gpio_defaults[7] gpio_defaults_block_30/gpio_defaults[8]
+ gpio_defaults_block_30/gpio_defaults[9] housekeeping/mgmt_gpio_in[30] gpio_control_in_2\[5\]/one
+ housekeeping/mgmt_gpio_in[30] gpio_control_in_2\[5\]/one padframe/mprj_io_analog_en[19]
+ padframe/mprj_io_analog_pol[19] padframe/mprj_io_analog_sel[19] padframe/mprj_io_dm[57]
+ padframe/mprj_io_dm[58] padframe/mprj_io_dm[59] padframe/mprj_io_holdover[19] padframe/mprj_io_ib_mode_sel[19]
+ padframe/mprj_io_in[19] padframe/mprj_io_inp_dis[19] padframe/mprj_io_out[19] padframe/mprj_io_oeb[19]
+ padframe/mprj_io_slow_sel[19] padframe/mprj_io_vtrip_sel[19] gpio_control_in_2\[5\]/resetn
+ gpio_control_in_2\[4\]/resetn gpio_control_in_2\[5\]/serial_clock gpio_control_in_2\[4\]/serial_clock
+ gpio_control_in_2\[5\]/serial_data_in gpio_control_in_2\[4\]/serial_data_in gpio_control_in_2\[5\]/serial_load
+ gpio_control_in_2\[4\]/serial_load mprj/io_in[19] mprj/io_oeb[19] mprj/io_out[19]
+ vccd_core vccd1_core VSUBS vssd1_core gpio_control_in_2\[5\]/zero gpio_control_block
Xgpio_defaults_block_0 VSUBS vccd_core gpio_defaults_block_0/gpio_defaults[0] gpio_defaults_block_0/gpio_defaults[10]
+ gpio_defaults_block_0/gpio_defaults[11] gpio_defaults_block_0/gpio_defaults[12]
+ gpio_defaults_block_0/gpio_defaults[1] gpio_defaults_block_0/gpio_defaults[2] gpio_defaults_block_0/gpio_defaults[3]
+ gpio_defaults_block_0/gpio_defaults[4] gpio_defaults_block_0/gpio_defaults[5] gpio_defaults_block_0/gpio_defaults[6]
+ gpio_defaults_block_0/gpio_defaults[7] gpio_defaults_block_0/gpio_defaults[8] gpio_defaults_block_0/gpio_defaults[9]
+ gpio_defaults_block_1803
Xgpio_defaults_block_1 VSUBS vccd_core gpio_defaults_block_1/gpio_defaults[0] gpio_defaults_block_1/gpio_defaults[10]
+ gpio_defaults_block_1/gpio_defaults[11] gpio_defaults_block_1/gpio_defaults[12]
+ gpio_defaults_block_1/gpio_defaults[1] gpio_defaults_block_1/gpio_defaults[2] gpio_defaults_block_1/gpio_defaults[3]
+ gpio_defaults_block_1/gpio_defaults[4] gpio_defaults_block_1/gpio_defaults[5] gpio_defaults_block_1/gpio_defaults[6]
+ gpio_defaults_block_1/gpio_defaults[7] gpio_defaults_block_1/gpio_defaults[8] gpio_defaults_block_1/gpio_defaults[9]
+ gpio_defaults_block_1803
Xuser_id_value user_id_value/mask_rev[0] user_id_value/mask_rev[10] user_id_value/mask_rev[11]
+ user_id_value/mask_rev[12] user_id_value/mask_rev[13] user_id_value/mask_rev[14]
+ user_id_value/mask_rev[15] user_id_value/mask_rev[16] user_id_value/mask_rev[17]
+ user_id_value/mask_rev[18] user_id_value/mask_rev[19] user_id_value/mask_rev[1]
+ user_id_value/mask_rev[20] user_id_value/mask_rev[21] user_id_value/mask_rev[22]
+ user_id_value/mask_rev[23] user_id_value/mask_rev[24] user_id_value/mask_rev[25]
+ user_id_value/mask_rev[26] user_id_value/mask_rev[27] user_id_value/mask_rev[28]
+ user_id_value/mask_rev[29] user_id_value/mask_rev[2] user_id_value/mask_rev[30]
+ user_id_value/mask_rev[31] user_id_value/mask_rev[3] user_id_value/mask_rev[4] user_id_value/mask_rev[5]
+ user_id_value/mask_rev[6] user_id_value/mask_rev[7] user_id_value/mask_rev[8] user_id_value/mask_rev[9]
+ vccd_core VSUBS user_id_programming
Xgpio_control_in_2\[3\] gpio_defaults_block_28/gpio_defaults[0] gpio_defaults_block_28/gpio_defaults[10]
+ gpio_defaults_block_28/gpio_defaults[11] gpio_defaults_block_28/gpio_defaults[12]
+ gpio_defaults_block_28/gpio_defaults[1] gpio_defaults_block_28/gpio_defaults[2]
+ gpio_defaults_block_28/gpio_defaults[3] gpio_defaults_block_28/gpio_defaults[4]
+ gpio_defaults_block_28/gpio_defaults[5] gpio_defaults_block_28/gpio_defaults[6]
+ gpio_defaults_block_28/gpio_defaults[7] gpio_defaults_block_28/gpio_defaults[8]
+ gpio_defaults_block_28/gpio_defaults[9] housekeeping/mgmt_gpio_in[28] gpio_control_in_2\[3\]/one
+ housekeeping/mgmt_gpio_in[28] gpio_control_in_2\[3\]/one padframe/mprj_io_analog_en[17]
+ padframe/mprj_io_analog_pol[17] padframe/mprj_io_analog_sel[17] padframe/mprj_io_dm[51]
+ padframe/mprj_io_dm[52] padframe/mprj_io_dm[53] padframe/mprj_io_holdover[17] padframe/mprj_io_ib_mode_sel[17]
+ padframe/mprj_io_in[17] padframe/mprj_io_inp_dis[17] padframe/mprj_io_out[17] padframe/mprj_io_oeb[17]
+ padframe/mprj_io_slow_sel[17] padframe/mprj_io_vtrip_sel[17] gpio_control_in_2\[3\]/resetn
+ gpio_control_in_2\[2\]/resetn gpio_control_in_2\[3\]/serial_clock gpio_control_in_2\[2\]/serial_clock
+ gpio_control_in_2\[3\]/serial_data_in gpio_control_in_2\[2\]/serial_data_in gpio_control_in_2\[3\]/serial_load
+ gpio_control_in_2\[2\]/serial_load mprj/io_in[17] mprj/io_oeb[17] mprj/io_out[17]
+ vccd_core vccd1_core VSUBS vssd1_core gpio_control_in_2\[3\]/zero gpio_control_block
Xgpio_defaults_block_2 VSUBS vccd_core gpio_defaults_block_2/gpio_defaults[0] gpio_defaults_block_2/gpio_defaults[10]
+ gpio_defaults_block_2/gpio_defaults[11] gpio_defaults_block_2/gpio_defaults[12]
+ gpio_defaults_block_2/gpio_defaults[1] gpio_defaults_block_2/gpio_defaults[2] gpio_defaults_block_2/gpio_defaults[3]
+ gpio_defaults_block_2/gpio_defaults[4] gpio_defaults_block_2/gpio_defaults[5] gpio_defaults_block_2/gpio_defaults[6]
+ gpio_defaults_block_2/gpio_defaults[7] gpio_defaults_block_2/gpio_defaults[8] gpio_defaults_block_2/gpio_defaults[9]
+ gpio_defaults_block_0403
Xgpio_defaults_block_3 VSUBS vccd_core gpio_defaults_block_3/gpio_defaults[0] gpio_defaults_block_3/gpio_defaults[10]
+ gpio_defaults_block_3/gpio_defaults[11] gpio_defaults_block_3/gpio_defaults[12]
+ gpio_defaults_block_3/gpio_defaults[1] gpio_defaults_block_3/gpio_defaults[2] gpio_defaults_block_3/gpio_defaults[3]
+ gpio_defaults_block_3/gpio_defaults[4] gpio_defaults_block_3/gpio_defaults[5] gpio_defaults_block_3/gpio_defaults[6]
+ gpio_defaults_block_3/gpio_defaults[7] gpio_defaults_block_3/gpio_defaults[8] gpio_defaults_block_3/gpio_defaults[9]
+ gpio_defaults_block_0403
Xgpio_control_bidir_1\[0\] gpio_defaults_block_0/gpio_defaults[0] gpio_defaults_block_0/gpio_defaults[10]
+ gpio_defaults_block_0/gpio_defaults[11] gpio_defaults_block_0/gpio_defaults[12]
+ gpio_defaults_block_0/gpio_defaults[1] gpio_defaults_block_0/gpio_defaults[2] gpio_defaults_block_0/gpio_defaults[3]
+ gpio_defaults_block_0/gpio_defaults[4] gpio_defaults_block_0/gpio_defaults[5] gpio_defaults_block_0/gpio_defaults[6]
+ gpio_defaults_block_0/gpio_defaults[7] gpio_defaults_block_0/gpio_defaults[8] gpio_defaults_block_0/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[0] gpio_control_bidir_1\[0\]/mgmt_gpio_oeb gpio_control_bidir_1\[0\]/mgmt_gpio_out
+ gpio_control_bidir_1\[0\]/one padframe/mprj_io_analog_en[0] padframe/mprj_io_analog_pol[0]
+ padframe/mprj_io_analog_sel[0] padframe/mprj_io_dm[0] padframe/mprj_io_dm[1] padframe/mprj_io_dm[2]
+ padframe/mprj_io_holdover[0] padframe/mprj_io_ib_mode_sel[0] padframe/mprj_io_in[0]
+ padframe/mprj_io_inp_dis[0] padframe/mprj_io_out[0] padframe/mprj_io_oeb[0] padframe/mprj_io_slow_sel[0]
+ padframe/mprj_io_vtrip_sel[0] housekeeping/serial_resetn gpio_control_bidir_1\[1\]/resetn
+ housekeeping/serial_clock gpio_control_bidir_1\[1\]/serial_clock housekeeping/serial_data_1
+ gpio_control_bidir_1\[1\]/serial_data_in housekeeping/serial_load gpio_control_bidir_1\[1\]/serial_load
+ mprj/io_in[0] mprj/io_oeb[0] mprj/io_out[0] vccd_core vccd1_core VSUBS vssd1_core
+ gpio_control_bidir_1\[0\]/zero gpio_control_block
Xgpio_defaults_block_5 VSUBS vccd_core gpio_defaults_block_5/gpio_defaults[0] gpio_defaults_block_5/gpio_defaults[10]
+ gpio_defaults_block_5/gpio_defaults[11] gpio_defaults_block_5/gpio_defaults[12]
+ gpio_defaults_block_5/gpio_defaults[1] gpio_defaults_block_5/gpio_defaults[2] gpio_defaults_block_5/gpio_defaults[3]
+ gpio_defaults_block_5/gpio_defaults[4] gpio_defaults_block_5/gpio_defaults[5] gpio_defaults_block_5/gpio_defaults[6]
+ gpio_defaults_block_5/gpio_defaults[7] gpio_defaults_block_5/gpio_defaults[8] gpio_defaults_block_5/gpio_defaults[9]
+ gpio_defaults_block
Xgpio_defaults_block_4 VSUBS vccd_core gpio_defaults_block_4/gpio_defaults[0] gpio_defaults_block_4/gpio_defaults[10]
+ gpio_defaults_block_4/gpio_defaults[11] gpio_defaults_block_4/gpio_defaults[12]
+ gpio_defaults_block_4/gpio_defaults[1] gpio_defaults_block_4/gpio_defaults[2] gpio_defaults_block_4/gpio_defaults[3]
+ gpio_defaults_block_4/gpio_defaults[4] gpio_defaults_block_4/gpio_defaults[5] gpio_defaults_block_4/gpio_defaults[6]
+ gpio_defaults_block_4/gpio_defaults[7] gpio_defaults_block_4/gpio_defaults[8] gpio_defaults_block_4/gpio_defaults[9]
+ gpio_defaults_block_0403
Xgpio_control_in_2\[1\] gpio_defaults_block_26/gpio_defaults[0] gpio_defaults_block_26/gpio_defaults[10]
+ gpio_defaults_block_26/gpio_defaults[11] gpio_defaults_block_26/gpio_defaults[12]
+ gpio_defaults_block_26/gpio_defaults[1] gpio_defaults_block_26/gpio_defaults[2]
+ gpio_defaults_block_26/gpio_defaults[3] gpio_defaults_block_26/gpio_defaults[4]
+ gpio_defaults_block_26/gpio_defaults[5] gpio_defaults_block_26/gpio_defaults[6]
+ gpio_defaults_block_26/gpio_defaults[7] gpio_defaults_block_26/gpio_defaults[8]
+ gpio_defaults_block_26/gpio_defaults[9] housekeeping/mgmt_gpio_in[26] gpio_control_in_2\[1\]/one
+ housekeeping/mgmt_gpio_in[26] gpio_control_in_2\[1\]/one padframe/mprj_io_analog_en[15]
+ padframe/mprj_io_analog_pol[15] padframe/mprj_io_analog_sel[15] padframe/mprj_io_dm[45]
+ padframe/mprj_io_dm[46] padframe/mprj_io_dm[47] padframe/mprj_io_holdover[15] padframe/mprj_io_ib_mode_sel[15]
+ padframe/mprj_io_in[15] padframe/mprj_io_inp_dis[15] padframe/mprj_io_out[15] padframe/mprj_io_oeb[15]
+ padframe/mprj_io_slow_sel[15] padframe/mprj_io_vtrip_sel[15] gpio_control_in_2\[1\]/resetn
+ gpio_control_in_2\[0\]/resetn gpio_control_in_2\[1\]/serial_clock gpio_control_in_2\[0\]/serial_clock
+ gpio_control_in_2\[1\]/serial_data_in gpio_control_in_2\[0\]/serial_data_in gpio_control_in_2\[1\]/serial_load
+ gpio_control_in_2\[0\]/serial_load mprj/io_in[15] mprj/io_oeb[15] mprj/io_out[15]
+ vccd_core vccd1_core VSUBS vssd1_core gpio_control_in_2\[1\]/zero gpio_control_block
Xgpio_defaults_block_6 VSUBS vccd_core gpio_defaults_block_6/gpio_defaults[0] gpio_defaults_block_6/gpio_defaults[10]
+ gpio_defaults_block_6/gpio_defaults[11] gpio_defaults_block_6/gpio_defaults[12]
+ gpio_defaults_block_6/gpio_defaults[1] gpio_defaults_block_6/gpio_defaults[2] gpio_defaults_block_6/gpio_defaults[3]
+ gpio_defaults_block_6/gpio_defaults[4] gpio_defaults_block_6/gpio_defaults[5] gpio_defaults_block_6/gpio_defaults[6]
+ gpio_defaults_block_6/gpio_defaults[7] gpio_defaults_block_6/gpio_defaults[8] gpio_defaults_block_6/gpio_defaults[9]
+ gpio_defaults_block
Xgpio_defaults_block_7 VSUBS vccd_core gpio_defaults_block_7/gpio_defaults[0] gpio_defaults_block_7/gpio_defaults[10]
+ gpio_defaults_block_7/gpio_defaults[11] gpio_defaults_block_7/gpio_defaults[12]
+ gpio_defaults_block_7/gpio_defaults[1] gpio_defaults_block_7/gpio_defaults[2] gpio_defaults_block_7/gpio_defaults[3]
+ gpio_defaults_block_7/gpio_defaults[4] gpio_defaults_block_7/gpio_defaults[5] gpio_defaults_block_7/gpio_defaults[6]
+ gpio_defaults_block_7/gpio_defaults[7] gpio_defaults_block_7/gpio_defaults[8] gpio_defaults_block_7/gpio_defaults[9]
+ gpio_defaults_block
Xgpio_defaults_block_8 VSUBS vccd_core gpio_defaults_block_8/gpio_defaults[0] gpio_defaults_block_8/gpio_defaults[10]
+ gpio_defaults_block_8/gpio_defaults[11] gpio_defaults_block_8/gpio_defaults[12]
+ gpio_defaults_block_8/gpio_defaults[1] gpio_defaults_block_8/gpio_defaults[2] gpio_defaults_block_8/gpio_defaults[3]
+ gpio_defaults_block_8/gpio_defaults[4] gpio_defaults_block_8/gpio_defaults[5] gpio_defaults_block_8/gpio_defaults[6]
+ gpio_defaults_block_8/gpio_defaults[7] gpio_defaults_block_8/gpio_defaults[8] gpio_defaults_block_8/gpio_defaults[9]
+ gpio_defaults_block
Xgpio_control_in_1a\[4\] gpio_defaults_block_6/gpio_defaults[0] gpio_defaults_block_6/gpio_defaults[10]
+ gpio_defaults_block_6/gpio_defaults[11] gpio_defaults_block_6/gpio_defaults[12]
+ gpio_defaults_block_6/gpio_defaults[1] gpio_defaults_block_6/gpio_defaults[2] gpio_defaults_block_6/gpio_defaults[3]
+ gpio_defaults_block_6/gpio_defaults[4] gpio_defaults_block_6/gpio_defaults[5] gpio_defaults_block_6/gpio_defaults[6]
+ gpio_defaults_block_6/gpio_defaults[7] gpio_defaults_block_6/gpio_defaults[8] gpio_defaults_block_6/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[6] gpio_control_in_1a\[4\]/one housekeeping/mgmt_gpio_in[6]
+ gpio_control_in_1a\[4\]/one padframe/mprj_io_analog_en[6] padframe/mprj_io_analog_pol[6]
+ padframe/mprj_io_analog_sel[6] padframe/mprj_io_dm[18] padframe/mprj_io_dm[19] padframe/mprj_io_dm[20]
+ padframe/mprj_io_holdover[6] padframe/mprj_io_ib_mode_sel[6] padframe/mprj_io_in[6]
+ padframe/mprj_io_inp_dis[6] padframe/mprj_io_out[6] padframe/mprj_io_oeb[6] padframe/mprj_io_slow_sel[6]
+ padframe/mprj_io_vtrip_sel[6] gpio_control_in_1a\[4\]/resetn gpio_control_in_1a\[5\]/resetn
+ gpio_control_in_1a\[4\]/serial_clock gpio_control_in_1a\[5\]/serial_clock gpio_control_in_1a\[4\]/serial_data_in
+ gpio_control_in_1a\[5\]/serial_data_in gpio_control_in_1a\[4\]/serial_load gpio_control_in_1a\[5\]/serial_load
+ mprj/io_in[6] mprj/io_oeb[6] mprj/io_out[6] vccd_core vccd1_core VSUBS vssd1_core
+ gpio_control_in_1a\[4\]/zero gpio_control_block
Xmgmt_buffers soc/core_clk clocking/user_clk soc/core_rstn mprj/la_data_in[0] mprj/la_data_in[100]
+ mprj/la_data_in[101] mprj/la_data_in[102] mprj/la_data_in[103] mprj/la_data_in[104]
+ mprj/la_data_in[105] mprj/la_data_in[106] mprj/la_data_in[107] mprj/la_data_in[108]
+ mprj/la_data_in[109] mprj/la_data_in[10] mprj/la_data_in[110] mprj/la_data_in[111]
+ mprj/la_data_in[112] mprj/la_data_in[113] mprj/la_data_in[114] mprj/la_data_in[115]
+ mprj/la_data_in[116] mprj/la_data_in[117] mprj/la_data_in[118] mprj/la_data_in[119]
+ mprj/la_data_in[11] mprj/la_data_in[120] mprj/la_data_in[121] mprj/la_data_in[122]
+ mprj/la_data_in[123] mprj/la_data_in[124] mprj/la_data_in[125] mprj/la_data_in[126]
+ mprj/la_data_in[127] mprj/la_data_in[12] mprj/la_data_in[13] mprj/la_data_in[14]
+ mprj/la_data_in[15] mprj/la_data_in[16] mprj/la_data_in[17] mprj/la_data_in[18]
+ mprj/la_data_in[19] mprj/la_data_in[1] mprj/la_data_in[20] mprj/la_data_in[21] mprj/la_data_in[22]
+ mprj/la_data_in[23] mprj/la_data_in[24] mprj/la_data_in[25] mprj/la_data_in[26]
+ mprj/la_data_in[27] mprj/la_data_in[28] mprj/la_data_in[29] mprj/la_data_in[2] mprj/la_data_in[30]
+ mprj/la_data_in[31] mprj/la_data_in[32] mprj/la_data_in[33] mprj/la_data_in[34]
+ mprj/la_data_in[35] mprj/la_data_in[36] mprj/la_data_in[37] mprj/la_data_in[38]
+ mprj/la_data_in[39] mprj/la_data_in[3] mprj/la_data_in[40] mprj/la_data_in[41] mprj/la_data_in[42]
+ mprj/la_data_in[43] mprj/la_data_in[44] mprj/la_data_in[45] mprj/la_data_in[46]
+ mprj/la_data_in[47] mprj/la_data_in[48] mprj/la_data_in[49] mprj/la_data_in[4] mprj/la_data_in[50]
+ mprj/la_data_in[51] mprj/la_data_in[52] mprj/la_data_in[53] mprj/la_data_in[54]
+ mprj/la_data_in[55] mprj/la_data_in[56] mprj/la_data_in[57] mprj/la_data_in[58]
+ mprj/la_data_in[59] mprj/la_data_in[5] mprj/la_data_in[60] mprj/la_data_in[61] mprj/la_data_in[62]
+ mprj/la_data_in[63] mprj/la_data_in[64] mprj/la_data_in[65] mprj/la_data_in[66]
+ mprj/la_data_in[67] mprj/la_data_in[68] mprj/la_data_in[69] mprj/la_data_in[6] mprj/la_data_in[70]
+ mprj/la_data_in[71] mprj/la_data_in[72] mprj/la_data_in[73] mprj/la_data_in[74]
+ mprj/la_data_in[75] mprj/la_data_in[76] mprj/la_data_in[77] mprj/la_data_in[78]
+ mprj/la_data_in[79] mprj/la_data_in[7] mprj/la_data_in[80] mprj/la_data_in[81] mprj/la_data_in[82]
+ mprj/la_data_in[83] mprj/la_data_in[84] mprj/la_data_in[85] mprj/la_data_in[86]
+ mprj/la_data_in[87] mprj/la_data_in[88] mprj/la_data_in[89] mprj/la_data_in[8] mprj/la_data_in[90]
+ mprj/la_data_in[91] mprj/la_data_in[92] mprj/la_data_in[93] mprj/la_data_in[94]
+ mprj/la_data_in[95] mprj/la_data_in[96] mprj/la_data_in[97] mprj/la_data_in[98]
+ mprj/la_data_in[99] mprj/la_data_in[9] soc/la_input[0] soc/la_input[100] soc/la_input[101]
+ soc/la_input[102] soc/la_input[103] soc/la_input[104] soc/la_input[105] soc/la_input[106]
+ soc/la_input[107] soc/la_input[108] soc/la_input[109] soc/la_input[10] soc/la_input[110]
+ soc/la_input[111] soc/la_input[112] soc/la_input[113] soc/la_input[114] soc/la_input[115]
+ soc/la_input[116] soc/la_input[117] soc/la_input[118] soc/la_input[119] soc/la_input[11]
+ soc/la_input[120] soc/la_input[121] soc/la_input[122] soc/la_input[123] soc/la_input[124]
+ soc/la_input[125] soc/la_input[126] soc/la_input[127] soc/la_input[12] soc/la_input[13]
+ soc/la_input[14] soc/la_input[15] soc/la_input[16] soc/la_input[17] soc/la_input[18]
+ soc/la_input[19] soc/la_input[1] soc/la_input[20] soc/la_input[21] soc/la_input[22]
+ soc/la_input[23] soc/la_input[24] soc/la_input[25] soc/la_input[26] soc/la_input[27]
+ soc/la_input[28] soc/la_input[29] soc/la_input[2] soc/la_input[30] soc/la_input[31]
+ soc/la_input[32] soc/la_input[33] soc/la_input[34] soc/la_input[35] soc/la_input[36]
+ soc/la_input[37] soc/la_input[38] soc/la_input[39] soc/la_input[3] soc/la_input[40]
+ soc/la_input[41] soc/la_input[42] soc/la_input[43] soc/la_input[44] soc/la_input[45]
+ soc/la_input[46] soc/la_input[47] soc/la_input[48] soc/la_input[49] soc/la_input[4]
+ soc/la_input[50] soc/la_input[51] soc/la_input[52] soc/la_input[53] soc/la_input[54]
+ soc/la_input[55] soc/la_input[56] soc/la_input[57] soc/la_input[58] soc/la_input[59]
+ soc/la_input[5] soc/la_input[60] soc/la_input[61] soc/la_input[62] soc/la_input[63]
+ soc/la_input[64] soc/la_input[65] soc/la_input[66] soc/la_input[67] soc/la_input[68]
+ soc/la_input[69] soc/la_input[6] soc/la_input[70] soc/la_input[71] soc/la_input[72]
+ soc/la_input[73] soc/la_input[74] soc/la_input[75] soc/la_input[76] soc/la_input[77]
+ soc/la_input[78] soc/la_input[79] soc/la_input[7] soc/la_input[80] soc/la_input[81]
+ soc/la_input[82] soc/la_input[83] soc/la_input[84] soc/la_input[85] soc/la_input[86]
+ soc/la_input[87] soc/la_input[88] soc/la_input[89] soc/la_input[8] soc/la_input[90]
+ soc/la_input[91] soc/la_input[92] soc/la_input[93] soc/la_input[94] soc/la_input[95]
+ soc/la_input[96] soc/la_input[97] soc/la_input[98] soc/la_input[99] soc/la_input[9]
+ mprj/la_data_out[0] mprj/la_data_out[100] mprj/la_data_out[101] mprj/la_data_out[102]
+ mprj/la_data_out[103] mprj/la_data_out[104] mprj/la_data_out[105] mprj/la_data_out[106]
+ mprj/la_data_out[107] mprj/la_data_out[108] mprj/la_data_out[109] mprj/la_data_out[10]
+ mprj/la_data_out[110] mprj/la_data_out[111] mprj/la_data_out[112] mprj/la_data_out[113]
+ mprj/la_data_out[114] mprj/la_data_out[115] mprj/la_data_out[116] mprj/la_data_out[117]
+ mprj/la_data_out[118] mprj/la_data_out[119] mprj/la_data_out[11] mprj/la_data_out[120]
+ mprj/la_data_out[121] mprj/la_data_out[122] mprj/la_data_out[123] mprj/la_data_out[124]
+ mprj/la_data_out[125] mprj/la_data_out[126] mprj/la_data_out[127] mprj/la_data_out[12]
+ mprj/la_data_out[13] mprj/la_data_out[14] mprj/la_data_out[15] mprj/la_data_out[16]
+ mprj/la_data_out[17] mprj/la_data_out[18] mprj/la_data_out[19] mprj/la_data_out[1]
+ mprj/la_data_out[20] mprj/la_data_out[21] mprj/la_data_out[22] mprj/la_data_out[23]
+ mprj/la_data_out[24] mprj/la_data_out[25] mprj/la_data_out[26] mprj/la_data_out[27]
+ mprj/la_data_out[28] mprj/la_data_out[29] mprj/la_data_out[2] mprj/la_data_out[30]
+ mprj/la_data_out[31] mprj/la_data_out[32] mprj/la_data_out[33] mprj/la_data_out[34]
+ mprj/la_data_out[35] mprj/la_data_out[36] mprj/la_data_out[37] mprj/la_data_out[38]
+ mprj/la_data_out[39] mprj/la_data_out[3] mprj/la_data_out[40] mprj/la_data_out[41]
+ mprj/la_data_out[42] mprj/la_data_out[43] mprj/la_data_out[44] mprj/la_data_out[45]
+ mprj/la_data_out[46] mprj/la_data_out[47] mprj/la_data_out[48] mprj/la_data_out[49]
+ mprj/la_data_out[4] mprj/la_data_out[50] mprj/la_data_out[51] mprj/la_data_out[52]
+ mprj/la_data_out[53] mprj/la_data_out[54] mprj/la_data_out[55] mprj/la_data_out[56]
+ mprj/la_data_out[57] mprj/la_data_out[58] mprj/la_data_out[59] mprj/la_data_out[5]
+ mprj/la_data_out[60] mprj/la_data_out[61] mprj/la_data_out[62] mprj/la_data_out[63]
+ mprj/la_data_out[64] mprj/la_data_out[65] mprj/la_data_out[66] mprj/la_data_out[67]
+ mprj/la_data_out[68] mprj/la_data_out[69] mprj/la_data_out[6] mprj/la_data_out[70]
+ mprj/la_data_out[71] mprj/la_data_out[72] mprj/la_data_out[73] mprj/la_data_out[74]
+ mprj/la_data_out[75] mprj/la_data_out[76] mprj/la_data_out[77] mprj/la_data_out[78]
+ mprj/la_data_out[79] mprj/la_data_out[7] mprj/la_data_out[80] mprj/la_data_out[81]
+ mprj/la_data_out[82] mprj/la_data_out[83] mprj/la_data_out[84] mprj/la_data_out[85]
+ mprj/la_data_out[86] mprj/la_data_out[87] mprj/la_data_out[88] mprj/la_data_out[89]
+ mprj/la_data_out[8] mprj/la_data_out[90] mprj/la_data_out[91] mprj/la_data_out[92]
+ mprj/la_data_out[93] mprj/la_data_out[94] mprj/la_data_out[95] mprj/la_data_out[96]
+ mprj/la_data_out[97] mprj/la_data_out[98] mprj/la_data_out[99] mprj/la_data_out[9]
+ soc/la_output[0] soc/la_output[100] soc/la_output[101] soc/la_output[102] soc/la_output[103]
+ soc/la_output[104] soc/la_output[105] soc/la_output[106] soc/la_output[107] soc/la_output[108]
+ soc/la_output[109] soc/la_output[10] soc/la_output[110] soc/la_output[111] soc/la_output[112]
+ soc/la_output[113] soc/la_output[114] soc/la_output[115] soc/la_output[116] soc/la_output[117]
+ soc/la_output[118] soc/la_output[119] soc/la_output[11] soc/la_output[120] soc/la_output[121]
+ soc/la_output[122] soc/la_output[123] soc/la_output[124] soc/la_output[125] soc/la_output[126]
+ soc/la_output[127] soc/la_output[12] soc/la_output[13] soc/la_output[14] soc/la_output[15]
+ soc/la_output[16] soc/la_output[17] soc/la_output[18] soc/la_output[19] soc/la_output[1]
+ soc/la_output[20] soc/la_output[21] soc/la_output[22] soc/la_output[23] soc/la_output[24]
+ soc/la_output[25] soc/la_output[26] soc/la_output[27] soc/la_output[28] soc/la_output[29]
+ soc/la_output[2] soc/la_output[30] soc/la_output[31] soc/la_output[32] soc/la_output[33]
+ soc/la_output[34] soc/la_output[35] soc/la_output[36] soc/la_output[37] soc/la_output[38]
+ soc/la_output[39] soc/la_output[3] soc/la_output[40] soc/la_output[41] soc/la_output[42]
+ soc/la_output[43] soc/la_output[44] soc/la_output[45] soc/la_output[46] soc/la_output[47]
+ soc/la_output[48] soc/la_output[49] soc/la_output[4] soc/la_output[50] soc/la_output[51]
+ soc/la_output[52] soc/la_output[53] soc/la_output[54] soc/la_output[55] soc/la_output[56]
+ soc/la_output[57] soc/la_output[58] soc/la_output[59] soc/la_output[5] soc/la_output[60]
+ soc/la_output[61] soc/la_output[62] soc/la_output[63] soc/la_output[64] soc/la_output[65]
+ soc/la_output[66] soc/la_output[67] soc/la_output[68] soc/la_output[69] soc/la_output[6]
+ soc/la_output[70] soc/la_output[71] soc/la_output[72] soc/la_output[73] soc/la_output[74]
+ soc/la_output[75] soc/la_output[76] soc/la_output[77] soc/la_output[78] soc/la_output[79]
+ soc/la_output[7] soc/la_output[80] soc/la_output[81] soc/la_output[82] soc/la_output[83]
+ soc/la_output[84] soc/la_output[85] soc/la_output[86] soc/la_output[87] soc/la_output[88]
+ soc/la_output[89] soc/la_output[8] soc/la_output[90] soc/la_output[91] soc/la_output[92]
+ soc/la_output[93] soc/la_output[94] soc/la_output[95] soc/la_output[96] soc/la_output[97]
+ soc/la_output[98] soc/la_output[99] soc/la_output[9] soc/la_iena[0] soc/la_iena[100]
+ soc/la_iena[101] soc/la_iena[102] soc/la_iena[103] soc/la_iena[104] soc/la_iena[105]
+ soc/la_iena[106] soc/la_iena[107] soc/la_iena[108] soc/la_iena[109] soc/la_iena[10]
+ soc/la_iena[110] soc/la_iena[111] soc/la_iena[112] soc/la_iena[113] soc/la_iena[114]
+ soc/la_iena[115] soc/la_iena[116] soc/la_iena[117] soc/la_iena[118] soc/la_iena[119]
+ soc/la_iena[11] soc/la_iena[120] soc/la_iena[121] soc/la_iena[122] soc/la_iena[123]
+ soc/la_iena[124] soc/la_iena[125] soc/la_iena[126] soc/la_iena[127] soc/la_iena[12]
+ soc/la_iena[13] soc/la_iena[14] soc/la_iena[15] soc/la_iena[16] soc/la_iena[17]
+ soc/la_iena[18] soc/la_iena[19] soc/la_iena[1] soc/la_iena[20] soc/la_iena[21] soc/la_iena[22]
+ soc/la_iena[23] soc/la_iena[24] soc/la_iena[25] soc/la_iena[26] soc/la_iena[27]
+ soc/la_iena[28] soc/la_iena[29] soc/la_iena[2] soc/la_iena[30] soc/la_iena[31] soc/la_iena[32]
+ soc/la_iena[33] soc/la_iena[34] soc/la_iena[35] soc/la_iena[36] soc/la_iena[37]
+ soc/la_iena[38] soc/la_iena[39] soc/la_iena[3] soc/la_iena[40] soc/la_iena[41] soc/la_iena[42]
+ soc/la_iena[43] soc/la_iena[44] soc/la_iena[45] soc/la_iena[46] soc/la_iena[47]
+ soc/la_iena[48] soc/la_iena[49] soc/la_iena[4] soc/la_iena[50] soc/la_iena[51] soc/la_iena[52]
+ soc/la_iena[53] soc/la_iena[54] soc/la_iena[55] soc/la_iena[56] soc/la_iena[57]
+ soc/la_iena[58] soc/la_iena[59] soc/la_iena[5] soc/la_iena[60] soc/la_iena[61] soc/la_iena[62]
+ soc/la_iena[63] soc/la_iena[64] soc/la_iena[65] soc/la_iena[66] soc/la_iena[67]
+ soc/la_iena[68] soc/la_iena[69] soc/la_iena[6] soc/la_iena[70] soc/la_iena[71] soc/la_iena[72]
+ soc/la_iena[73] soc/la_iena[74] soc/la_iena[75] soc/la_iena[76] soc/la_iena[77]
+ soc/la_iena[78] soc/la_iena[79] soc/la_iena[7] soc/la_iena[80] soc/la_iena[81] soc/la_iena[82]
+ soc/la_iena[83] soc/la_iena[84] soc/la_iena[85] soc/la_iena[86] soc/la_iena[87]
+ soc/la_iena[88] soc/la_iena[89] soc/la_iena[8] soc/la_iena[90] soc/la_iena[91] soc/la_iena[92]
+ soc/la_iena[93] soc/la_iena[94] soc/la_iena[95] soc/la_iena[96] soc/la_iena[97]
+ soc/la_iena[98] soc/la_iena[99] soc/la_iena[9] mprj/la_oenb[0] mprj/la_oenb[100]
+ mprj/la_oenb[101] mprj/la_oenb[102] mprj/la_oenb[103] mprj/la_oenb[104] mprj/la_oenb[105]
+ mprj/la_oenb[106] mprj/la_oenb[107] mprj/la_oenb[108] mprj/la_oenb[109] mprj/la_oenb[10]
+ mprj/la_oenb[110] mprj/la_oenb[111] mprj/la_oenb[112] mprj/la_oenb[113] mprj/la_oenb[114]
+ mprj/la_oenb[115] mprj/la_oenb[116] mprj/la_oenb[117] mprj/la_oenb[118] mprj/la_oenb[119]
+ mprj/la_oenb[11] mprj/la_oenb[120] mprj/la_oenb[121] mprj/la_oenb[122] mprj/la_oenb[123]
+ mprj/la_oenb[124] mprj/la_oenb[125] mprj/la_oenb[126] mprj/la_oenb[127] mprj/la_oenb[12]
+ mprj/la_oenb[13] mprj/la_oenb[14] mprj/la_oenb[15] mprj/la_oenb[16] mprj/la_oenb[17]
+ mprj/la_oenb[18] mprj/la_oenb[19] mprj/la_oenb[1] mprj/la_oenb[20] mprj/la_oenb[21]
+ mprj/la_oenb[22] mprj/la_oenb[23] mprj/la_oenb[24] mprj/la_oenb[25] mprj/la_oenb[26]
+ mprj/la_oenb[27] mprj/la_oenb[28] mprj/la_oenb[29] mprj/la_oenb[2] mprj/la_oenb[30]
+ mprj/la_oenb[31] mprj/la_oenb[32] mprj/la_oenb[33] mprj/la_oenb[34] mprj/la_oenb[35]
+ mprj/la_oenb[36] mprj/la_oenb[37] mprj/la_oenb[38] mprj/la_oenb[39] mprj/la_oenb[3]
+ mprj/la_oenb[40] mprj/la_oenb[41] mprj/la_oenb[42] mprj/la_oenb[43] mprj/la_oenb[44]
+ mprj/la_oenb[45] mprj/la_oenb[46] mprj/la_oenb[47] mprj/la_oenb[48] mprj/la_oenb[49]
+ mprj/la_oenb[4] mprj/la_oenb[50] mprj/la_oenb[51] mprj/la_oenb[52] mprj/la_oenb[53]
+ mprj/la_oenb[54] mprj/la_oenb[55] mprj/la_oenb[56] mprj/la_oenb[57] mprj/la_oenb[58]
+ mprj/la_oenb[59] mprj/la_oenb[5] mprj/la_oenb[60] mprj/la_oenb[61] mprj/la_oenb[62]
+ mprj/la_oenb[63] mprj/la_oenb[64] mprj/la_oenb[65] mprj/la_oenb[66] mprj/la_oenb[67]
+ mprj/la_oenb[68] mprj/la_oenb[69] mprj/la_oenb[6] mprj/la_oenb[70] mprj/la_oenb[71]
+ mprj/la_oenb[72] mprj/la_oenb[73] mprj/la_oenb[74] mprj/la_oenb[75] mprj/la_oenb[76]
+ mprj/la_oenb[77] mprj/la_oenb[78] mprj/la_oenb[79] mprj/la_oenb[7] mprj/la_oenb[80]
+ mprj/la_oenb[81] mprj/la_oenb[82] mprj/la_oenb[83] mprj/la_oenb[84] mprj/la_oenb[85]
+ mprj/la_oenb[86] mprj/la_oenb[87] mprj/la_oenb[88] mprj/la_oenb[89] mprj/la_oenb[8]
+ mprj/la_oenb[90] mprj/la_oenb[91] mprj/la_oenb[92] mprj/la_oenb[93] mprj/la_oenb[94]
+ mprj/la_oenb[95] mprj/la_oenb[96] mprj/la_oenb[97] mprj/la_oenb[98] mprj/la_oenb[99]
+ mprj/la_oenb[9] soc/la_oenb[0] soc/la_oenb[100] soc/la_oenb[101] soc/la_oenb[102]
+ soc/la_oenb[103] soc/la_oenb[104] soc/la_oenb[105] soc/la_oenb[106] soc/la_oenb[107]
+ soc/la_oenb[108] soc/la_oenb[109] soc/la_oenb[10] soc/la_oenb[110] soc/la_oenb[111]
+ soc/la_oenb[112] soc/la_oenb[113] soc/la_oenb[114] soc/la_oenb[115] soc/la_oenb[116]
+ soc/la_oenb[117] soc/la_oenb[118] soc/la_oenb[119] soc/la_oenb[11] soc/la_oenb[120]
+ soc/la_oenb[121] soc/la_oenb[122] soc/la_oenb[123] soc/la_oenb[124] soc/la_oenb[125]
+ soc/la_oenb[126] soc/la_oenb[127] soc/la_oenb[12] soc/la_oenb[13] soc/la_oenb[14]
+ soc/la_oenb[15] soc/la_oenb[16] soc/la_oenb[17] soc/la_oenb[18] soc/la_oenb[19]
+ soc/la_oenb[1] soc/la_oenb[20] soc/la_oenb[21] soc/la_oenb[22] soc/la_oenb[23] soc/la_oenb[24]
+ soc/la_oenb[25] soc/la_oenb[26] soc/la_oenb[27] soc/la_oenb[28] soc/la_oenb[29]
+ soc/la_oenb[2] soc/la_oenb[30] soc/la_oenb[31] soc/la_oenb[32] soc/la_oenb[33] soc/la_oenb[34]
+ soc/la_oenb[35] soc/la_oenb[36] soc/la_oenb[37] soc/la_oenb[38] soc/la_oenb[39]
+ soc/la_oenb[3] soc/la_oenb[40] soc/la_oenb[41] soc/la_oenb[42] soc/la_oenb[43] soc/la_oenb[44]
+ soc/la_oenb[45] soc/la_oenb[46] soc/la_oenb[47] soc/la_oenb[48] soc/la_oenb[49]
+ soc/la_oenb[4] soc/la_oenb[50] soc/la_oenb[51] soc/la_oenb[52] soc/la_oenb[53] soc/la_oenb[54]
+ soc/la_oenb[55] soc/la_oenb[56] soc/la_oenb[57] soc/la_oenb[58] soc/la_oenb[59]
+ soc/la_oenb[5] soc/la_oenb[60] soc/la_oenb[61] soc/la_oenb[62] soc/la_oenb[63] soc/la_oenb[64]
+ soc/la_oenb[65] soc/la_oenb[66] soc/la_oenb[67] soc/la_oenb[68] soc/la_oenb[69]
+ soc/la_oenb[6] soc/la_oenb[70] soc/la_oenb[71] soc/la_oenb[72] soc/la_oenb[73] soc/la_oenb[74]
+ soc/la_oenb[75] soc/la_oenb[76] soc/la_oenb[77] soc/la_oenb[78] soc/la_oenb[79]
+ soc/la_oenb[7] soc/la_oenb[80] soc/la_oenb[81] soc/la_oenb[82] soc/la_oenb[83] soc/la_oenb[84]
+ soc/la_oenb[85] soc/la_oenb[86] soc/la_oenb[87] soc/la_oenb[88] soc/la_oenb[89]
+ soc/la_oenb[8] soc/la_oenb[90] soc/la_oenb[91] soc/la_oenb[92] soc/la_oenb[93] soc/la_oenb[94]
+ soc/la_oenb[95] soc/la_oenb[96] soc/la_oenb[97] soc/la_oenb[98] soc/la_oenb[99]
+ soc/la_oenb[9] soc/mprj_ack_i mprj/wbs_ack_o soc/mprj_adr_o[0] soc/mprj_adr_o[10]
+ soc/mprj_adr_o[11] soc/mprj_adr_o[12] soc/mprj_adr_o[13] soc/mprj_adr_o[14] soc/mprj_adr_o[15]
+ soc/mprj_adr_o[16] soc/mprj_adr_o[17] soc/mprj_adr_o[18] soc/mprj_adr_o[19] soc/mprj_adr_o[1]
+ soc/mprj_adr_o[20] soc/mprj_adr_o[21] soc/mprj_adr_o[22] soc/mprj_adr_o[23] soc/mprj_adr_o[24]
+ soc/mprj_adr_o[25] soc/mprj_adr_o[26] soc/mprj_adr_o[27] soc/mprj_adr_o[28] soc/mprj_adr_o[29]
+ soc/mprj_adr_o[2] soc/mprj_adr_o[30] soc/mprj_adr_o[31] soc/mprj_adr_o[3] soc/mprj_adr_o[4]
+ soc/mprj_adr_o[5] soc/mprj_adr_o[6] soc/mprj_adr_o[7] soc/mprj_adr_o[8] soc/mprj_adr_o[9]
+ mprj/wbs_adr_i[0] mprj/wbs_adr_i[10] mprj/wbs_adr_i[11] mprj/wbs_adr_i[12] mprj/wbs_adr_i[13]
+ mprj/wbs_adr_i[14] mprj/wbs_adr_i[15] mprj/wbs_adr_i[16] mprj/wbs_adr_i[17] mprj/wbs_adr_i[18]
+ mprj/wbs_adr_i[19] mprj/wbs_adr_i[1] mprj/wbs_adr_i[20] mprj/wbs_adr_i[21] mprj/wbs_adr_i[22]
+ mprj/wbs_adr_i[23] mprj/wbs_adr_i[24] mprj/wbs_adr_i[25] mprj/wbs_adr_i[26] mprj/wbs_adr_i[27]
+ mprj/wbs_adr_i[28] mprj/wbs_adr_i[29] mprj/wbs_adr_i[2] mprj/wbs_adr_i[30] mprj/wbs_adr_i[31]
+ mprj/wbs_adr_i[3] mprj/wbs_adr_i[4] mprj/wbs_adr_i[5] mprj/wbs_adr_i[6] mprj/wbs_adr_i[7]
+ mprj/wbs_adr_i[8] mprj/wbs_adr_i[9] soc/mprj_cyc_o mprj/wbs_cyc_i soc/mprj_dat_i[0]
+ soc/mprj_dat_i[10] soc/mprj_dat_i[11] soc/mprj_dat_i[12] soc/mprj_dat_i[13] soc/mprj_dat_i[14]
+ soc/mprj_dat_i[15] soc/mprj_dat_i[16] soc/mprj_dat_i[17] soc/mprj_dat_i[18] soc/mprj_dat_i[19]
+ soc/mprj_dat_i[1] soc/mprj_dat_i[20] soc/mprj_dat_i[21] soc/mprj_dat_i[22] soc/mprj_dat_i[23]
+ soc/mprj_dat_i[24] soc/mprj_dat_i[25] soc/mprj_dat_i[26] soc/mprj_dat_i[27] soc/mprj_dat_i[28]
+ soc/mprj_dat_i[29] soc/mprj_dat_i[2] soc/mprj_dat_i[30] soc/mprj_dat_i[31] soc/mprj_dat_i[3]
+ soc/mprj_dat_i[4] soc/mprj_dat_i[5] soc/mprj_dat_i[6] soc/mprj_dat_i[7] soc/mprj_dat_i[8]
+ soc/mprj_dat_i[9] mprj/wbs_dat_o[0] mprj/wbs_dat_o[10] mprj/wbs_dat_o[11] mprj/wbs_dat_o[12]
+ mprj/wbs_dat_o[13] mprj/wbs_dat_o[14] mprj/wbs_dat_o[15] mprj/wbs_dat_o[16] mprj/wbs_dat_o[17]
+ mprj/wbs_dat_o[18] mprj/wbs_dat_o[19] mprj/wbs_dat_o[1] mprj/wbs_dat_o[20] mprj/wbs_dat_o[21]
+ mprj/wbs_dat_o[22] mprj/wbs_dat_o[23] mprj/wbs_dat_o[24] mprj/wbs_dat_o[25] mprj/wbs_dat_o[26]
+ mprj/wbs_dat_o[27] mprj/wbs_dat_o[28] mprj/wbs_dat_o[29] mprj/wbs_dat_o[2] mprj/wbs_dat_o[30]
+ mprj/wbs_dat_o[31] mprj/wbs_dat_o[3] mprj/wbs_dat_o[4] mprj/wbs_dat_o[5] mprj/wbs_dat_o[6]
+ mprj/wbs_dat_o[7] mprj/wbs_dat_o[8] mprj/wbs_dat_o[9] soc/mprj_dat_o[0] soc/mprj_dat_o[10]
+ soc/mprj_dat_o[11] soc/mprj_dat_o[12] soc/mprj_dat_o[13] soc/mprj_dat_o[14] soc/mprj_dat_o[15]
+ soc/mprj_dat_o[16] soc/mprj_dat_o[17] soc/mprj_dat_o[18] soc/mprj_dat_o[19] soc/mprj_dat_o[1]
+ soc/mprj_dat_o[20] soc/mprj_dat_o[21] soc/mprj_dat_o[22] soc/mprj_dat_o[23] soc/mprj_dat_o[24]
+ soc/mprj_dat_o[25] soc/mprj_dat_o[26] soc/mprj_dat_o[27] soc/mprj_dat_o[28] soc/mprj_dat_o[29]
+ soc/mprj_dat_o[2] soc/mprj_dat_o[30] soc/mprj_dat_o[31] soc/mprj_dat_o[3] soc/mprj_dat_o[4]
+ soc/mprj_dat_o[5] soc/mprj_dat_o[6] soc/mprj_dat_o[7] soc/mprj_dat_o[8] soc/mprj_dat_o[9]
+ mprj/wbs_dat_i[0] mprj/wbs_dat_i[10] mprj/wbs_dat_i[11] mprj/wbs_dat_i[12] mprj/wbs_dat_i[13]
+ mprj/wbs_dat_i[14] mprj/wbs_dat_i[15] mprj/wbs_dat_i[16] mprj/wbs_dat_i[17] mprj/wbs_dat_i[18]
+ mprj/wbs_dat_i[19] mprj/wbs_dat_i[1] mprj/wbs_dat_i[20] mprj/wbs_dat_i[21] mprj/wbs_dat_i[22]
+ mprj/wbs_dat_i[23] mprj/wbs_dat_i[24] mprj/wbs_dat_i[25] mprj/wbs_dat_i[26] mprj/wbs_dat_i[27]
+ mprj/wbs_dat_i[28] mprj/wbs_dat_i[29] mprj/wbs_dat_i[2] mprj/wbs_dat_i[30] mprj/wbs_dat_i[31]
+ mprj/wbs_dat_i[3] mprj/wbs_dat_i[4] mprj/wbs_dat_i[5] mprj/wbs_dat_i[6] mprj/wbs_dat_i[7]
+ mprj/wbs_dat_i[8] mprj/wbs_dat_i[9] mgmt_buffers/mprj_iena_wb soc/mprj_sel_o[0]
+ soc/mprj_sel_o[1] soc/mprj_sel_o[2] soc/mprj_sel_o[3] mprj/wbs_sel_i[0] mprj/wbs_sel_i[1]
+ mprj/wbs_sel_i[2] mprj/wbs_sel_i[3] soc/mprj_stb_o mprj/wbs_stb_i soc/mprj_we_o
+ mprj/wbs_we_i housekeeping/usr1_vcc_pwrgood housekeeping/usr1_vdd_pwrgood housekeeping/usr2_vcc_pwrgood
+ housekeeping/usr2_vdd_pwrgood mprj/wb_clk_i mprj/user_clock2 soc/irq[0] soc/irq[1]
+ soc/irq[2] mprj/user_irq[0] mprj/user_irq[1] mprj/user_irq[2] mgmt_buffers/user_irq_ena[0]
+ mgmt_buffers/user_irq_ena[1] mgmt_buffers/user_irq_ena[2] mprj/wb_rst_i vccd_core
+ vccd1_core vccd2_core vdda1_core vdda2_core vssa1_core vssa2_core VSUBS vssd1_core
+ vssd2_core mgmt_protect
Xrstb_level rstb_level/A pll/resetb por/vdd3v3 por/vss3v3 vccd_core VSUBS xres_buf
Xgpio_defaults_block_9 VSUBS vccd_core gpio_defaults_block_9/gpio_defaults[0] gpio_defaults_block_9/gpio_defaults[10]
+ gpio_defaults_block_9/gpio_defaults[11] gpio_defaults_block_9/gpio_defaults[12]
+ gpio_defaults_block_9/gpio_defaults[1] gpio_defaults_block_9/gpio_defaults[2] gpio_defaults_block_9/gpio_defaults[3]
+ gpio_defaults_block_9/gpio_defaults[4] gpio_defaults_block_9/gpio_defaults[5] gpio_defaults_block_9/gpio_defaults[6]
+ gpio_defaults_block_9/gpio_defaults[7] gpio_defaults_block_9/gpio_defaults[8] gpio_defaults_block_9/gpio_defaults[9]
+ gpio_defaults_block
Xgpio_control_bidir_2\[1\] gpio_defaults_block_36/gpio_defaults[0] gpio_defaults_block_36/gpio_defaults[10]
+ gpio_defaults_block_36/gpio_defaults[11] gpio_defaults_block_36/gpio_defaults[12]
+ gpio_defaults_block_36/gpio_defaults[1] gpio_defaults_block_36/gpio_defaults[2]
+ gpio_defaults_block_36/gpio_defaults[3] gpio_defaults_block_36/gpio_defaults[4]
+ gpio_defaults_block_36/gpio_defaults[5] gpio_defaults_block_36/gpio_defaults[6]
+ gpio_defaults_block_36/gpio_defaults[7] gpio_defaults_block_36/gpio_defaults[8]
+ gpio_defaults_block_36/gpio_defaults[9] housekeeping/mgmt_gpio_in[36] housekeeping/mgmt_gpio_oeb[36]
+ housekeeping/mgmt_gpio_out[36] gpio_control_bidir_2\[1\]/one padframe/mprj_io_analog_en[25]
+ padframe/mprj_io_analog_pol[25] padframe/mprj_io_analog_sel[25] padframe/mprj_io_dm[75]
+ padframe/mprj_io_dm[76] padframe/mprj_io_dm[77] padframe/mprj_io_holdover[25] padframe/mprj_io_ib_mode_sel[25]
+ padframe/mprj_io_in[25] padframe/mprj_io_inp_dis[25] padframe/mprj_io_out[25] padframe/mprj_io_oeb[25]
+ padframe/mprj_io_slow_sel[25] padframe/mprj_io_vtrip_sel[25] gpio_control_bidir_2\[1\]/resetn
+ gpio_control_bidir_2\[0\]/resetn gpio_control_bidir_2\[1\]/serial_clock gpio_control_bidir_2\[0\]/serial_clock
+ gpio_control_bidir_2\[1\]/serial_data_in gpio_control_bidir_2\[0\]/serial_data_in
+ gpio_control_bidir_2\[1\]/serial_load gpio_control_bidir_2\[0\]/serial_load mprj/io_in[25]
+ mprj/io_oeb[25] mprj/io_out[25] vccd_core vccd1_core VSUBS vssd1_core gpio_control_bidir_2\[1\]/zero
+ gpio_control_block
Xgpio_control_in_1\[5\] gpio_defaults_block_13/gpio_defaults[0] gpio_defaults_block_13/gpio_defaults[10]
+ gpio_defaults_block_13/gpio_defaults[11] gpio_defaults_block_13/gpio_defaults[12]
+ gpio_defaults_block_13/gpio_defaults[1] gpio_defaults_block_13/gpio_defaults[2]
+ gpio_defaults_block_13/gpio_defaults[3] gpio_defaults_block_13/gpio_defaults[4]
+ gpio_defaults_block_13/gpio_defaults[5] gpio_defaults_block_13/gpio_defaults[6]
+ gpio_defaults_block_13/gpio_defaults[7] gpio_defaults_block_13/gpio_defaults[8]
+ gpio_defaults_block_13/gpio_defaults[9] housekeeping/mgmt_gpio_in[13] gpio_control_in_1\[5\]/one
+ housekeeping/mgmt_gpio_in[13] gpio_control_in_1\[5\]/one padframe/mprj_io_analog_en[13]
+ padframe/mprj_io_analog_pol[13] padframe/mprj_io_analog_sel[13] padframe/mprj_io_dm[39]
+ padframe/mprj_io_dm[40] padframe/mprj_io_dm[41] padframe/mprj_io_holdover[13] padframe/mprj_io_ib_mode_sel[13]
+ padframe/mprj_io_in[13] padframe/mprj_io_inp_dis[13] padframe/mprj_io_out[13] padframe/mprj_io_oeb[13]
+ padframe/mprj_io_slow_sel[13] padframe/mprj_io_vtrip_sel[13] gpio_control_in_1\[5\]/resetn
+ gpio_control_in_1\[5\]/resetn_out gpio_control_in_1\[5\]/serial_clock gpio_control_in_1\[5\]/serial_clock_out
+ gpio_control_in_1\[5\]/serial_data_in gpio_control_in_1\[5\]/serial_data_out gpio_control_in_1\[5\]/serial_load
+ gpio_control_in_1\[5\]/serial_load_out mprj/io_in[13] mprj/io_oeb[13] mprj/io_out[13]
+ vccd_core vccd1_core VSUBS vssd1_core gpio_control_in_1\[5\]/zero gpio_control_block
Xgpio_control_in_1a\[2\] gpio_defaults_block_4/gpio_defaults[0] gpio_defaults_block_4/gpio_defaults[10]
+ gpio_defaults_block_4/gpio_defaults[11] gpio_defaults_block_4/gpio_defaults[12]
+ gpio_defaults_block_4/gpio_defaults[1] gpio_defaults_block_4/gpio_defaults[2] gpio_defaults_block_4/gpio_defaults[3]
+ gpio_defaults_block_4/gpio_defaults[4] gpio_defaults_block_4/gpio_defaults[5] gpio_defaults_block_4/gpio_defaults[6]
+ gpio_defaults_block_4/gpio_defaults[7] gpio_defaults_block_4/gpio_defaults[8] gpio_defaults_block_4/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[4] gpio_control_in_1a\[2\]/one housekeeping/mgmt_gpio_in[4]
+ gpio_control_in_1a\[2\]/one padframe/mprj_io_analog_en[4] padframe/mprj_io_analog_pol[4]
+ padframe/mprj_io_analog_sel[4] padframe/mprj_io_dm[12] padframe/mprj_io_dm[13] padframe/mprj_io_dm[14]
+ padframe/mprj_io_holdover[4] padframe/mprj_io_ib_mode_sel[4] padframe/mprj_io_in[4]
+ padframe/mprj_io_inp_dis[4] padframe/mprj_io_out[4] padframe/mprj_io_oeb[4] padframe/mprj_io_slow_sel[4]
+ padframe/mprj_io_vtrip_sel[4] gpio_control_in_1a\[2\]/resetn gpio_control_in_1a\[3\]/resetn
+ gpio_control_in_1a\[2\]/serial_clock gpio_control_in_1a\[3\]/serial_clock gpio_control_in_1a\[2\]/serial_data_in
+ gpio_control_in_1a\[3\]/serial_data_in gpio_control_in_1a\[2\]/serial_load gpio_control_in_1a\[3\]/serial_load
+ mprj/io_in[4] mprj/io_oeb[4] mprj/io_out[4] vccd_core vccd1_core VSUBS vssd1_core
+ gpio_control_in_1a\[2\]/zero gpio_control_block
Xgpio_control_in_2\[8\] gpio_defaults_block_33/gpio_defaults[0] gpio_defaults_block_33/gpio_defaults[10]
+ gpio_defaults_block_33/gpio_defaults[11] gpio_defaults_block_33/gpio_defaults[12]
+ gpio_defaults_block_33/gpio_defaults[1] gpio_defaults_block_33/gpio_defaults[2]
+ gpio_defaults_block_33/gpio_defaults[3] gpio_defaults_block_33/gpio_defaults[4]
+ gpio_defaults_block_33/gpio_defaults[5] gpio_defaults_block_33/gpio_defaults[6]
+ gpio_defaults_block_33/gpio_defaults[7] gpio_defaults_block_33/gpio_defaults[8]
+ gpio_defaults_block_33/gpio_defaults[9] housekeeping/mgmt_gpio_in[33] gpio_control_in_2\[8\]/one
+ housekeeping/mgmt_gpio_in[33] gpio_control_in_2\[8\]/one padframe/mprj_io_analog_en[22]
+ padframe/mprj_io_analog_pol[22] padframe/mprj_io_analog_sel[22] padframe/mprj_io_dm[66]
+ padframe/mprj_io_dm[67] padframe/mprj_io_dm[68] padframe/mprj_io_holdover[22] padframe/mprj_io_ib_mode_sel[22]
+ padframe/mprj_io_in[22] padframe/mprj_io_inp_dis[22] padframe/mprj_io_out[22] padframe/mprj_io_oeb[22]
+ padframe/mprj_io_slow_sel[22] padframe/mprj_io_vtrip_sel[22] gpio_control_in_2\[8\]/resetn
+ gpio_control_in_2\[7\]/resetn gpio_control_in_2\[8\]/serial_clock gpio_control_in_2\[7\]/serial_clock
+ gpio_control_in_2\[8\]/serial_data_in gpio_control_in_2\[7\]/serial_data_in gpio_control_in_2\[8\]/serial_load
+ gpio_control_in_2\[7\]/serial_load mprj/io_in[22] mprj/io_oeb[22] mprj/io_out[22]
+ vccd_core vccd1_core VSUBS vssd1_core gpio_control_in_2\[8\]/zero gpio_control_block
Xgpio_control_in_1\[3\] gpio_defaults_block_11/gpio_defaults[0] gpio_defaults_block_11/gpio_defaults[10]
+ gpio_defaults_block_11/gpio_defaults[11] gpio_defaults_block_11/gpio_defaults[12]
+ gpio_defaults_block_11/gpio_defaults[1] gpio_defaults_block_11/gpio_defaults[2]
+ gpio_defaults_block_11/gpio_defaults[3] gpio_defaults_block_11/gpio_defaults[4]
+ gpio_defaults_block_11/gpio_defaults[5] gpio_defaults_block_11/gpio_defaults[6]
+ gpio_defaults_block_11/gpio_defaults[7] gpio_defaults_block_11/gpio_defaults[8]
+ gpio_defaults_block_11/gpio_defaults[9] housekeeping/mgmt_gpio_in[11] gpio_control_in_1\[3\]/one
+ housekeeping/mgmt_gpio_in[11] gpio_control_in_1\[3\]/one padframe/mprj_io_analog_en[11]
+ padframe/mprj_io_analog_pol[11] padframe/mprj_io_analog_sel[11] padframe/mprj_io_dm[33]
+ padframe/mprj_io_dm[34] padframe/mprj_io_dm[35] padframe/mprj_io_holdover[11] padframe/mprj_io_ib_mode_sel[11]
+ padframe/mprj_io_in[11] padframe/mprj_io_inp_dis[11] padframe/mprj_io_out[11] padframe/mprj_io_oeb[11]
+ padframe/mprj_io_slow_sel[11] padframe/mprj_io_vtrip_sel[11] gpio_control_in_1\[3\]/resetn
+ gpio_control_in_1\[4\]/resetn gpio_control_in_1\[3\]/serial_clock gpio_control_in_1\[4\]/serial_clock
+ gpio_control_in_1\[3\]/serial_data_in gpio_control_in_1\[4\]/serial_data_in gpio_control_in_1\[3\]/serial_load
+ gpio_control_in_1\[4\]/serial_load mprj/io_in[11] mprj/io_oeb[11] mprj/io_out[11]
+ vccd_core vccd1_core VSUBS vssd1_core gpio_control_in_1\[3\]/zero gpio_control_block
Xgpio_control_in_1a\[0\] gpio_defaults_block_2/gpio_defaults[0] gpio_defaults_block_2/gpio_defaults[10]
+ gpio_defaults_block_2/gpio_defaults[11] gpio_defaults_block_2/gpio_defaults[12]
+ gpio_defaults_block_2/gpio_defaults[1] gpio_defaults_block_2/gpio_defaults[2] gpio_defaults_block_2/gpio_defaults[3]
+ gpio_defaults_block_2/gpio_defaults[4] gpio_defaults_block_2/gpio_defaults[5] gpio_defaults_block_2/gpio_defaults[6]
+ gpio_defaults_block_2/gpio_defaults[7] gpio_defaults_block_2/gpio_defaults[8] gpio_defaults_block_2/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[2] gpio_control_in_1a\[0\]/one housekeeping/mgmt_gpio_in[2]
+ gpio_control_in_1a\[0\]/one padframe/mprj_io_analog_en[2] padframe/mprj_io_analog_pol[2]
+ padframe/mprj_io_analog_sel[2] padframe/mprj_io_dm[6] padframe/mprj_io_dm[7] padframe/mprj_io_dm[8]
+ padframe/mprj_io_holdover[2] padframe/mprj_io_ib_mode_sel[2] padframe/mprj_io_in[2]
+ padframe/mprj_io_inp_dis[2] padframe/mprj_io_out[2] padframe/mprj_io_oeb[2] padframe/mprj_io_slow_sel[2]
+ padframe/mprj_io_vtrip_sel[2] gpio_control_in_1a\[0\]/resetn gpio_control_in_1a\[1\]/resetn
+ gpio_control_in_1a\[0\]/serial_clock gpio_control_in_1a\[1\]/serial_clock gpio_control_in_1a\[0\]/serial_data_in
+ gpio_control_in_1a\[1\]/serial_data_in gpio_control_in_1a\[0\]/serial_load gpio_control_in_1a\[1\]/serial_load
+ mprj/io_in[2] mprj/io_oeb[2] mprj/io_out[2] vccd_core vccd1_core VSUBS vssd1_core
+ gpio_control_in_1a\[0\]/zero gpio_control_block
Xgpio_control_in_2\[6\] gpio_defaults_block_31/gpio_defaults[0] gpio_defaults_block_31/gpio_defaults[10]
+ gpio_defaults_block_31/gpio_defaults[11] gpio_defaults_block_31/gpio_defaults[12]
+ gpio_defaults_block_31/gpio_defaults[1] gpio_defaults_block_31/gpio_defaults[2]
+ gpio_defaults_block_31/gpio_defaults[3] gpio_defaults_block_31/gpio_defaults[4]
+ gpio_defaults_block_31/gpio_defaults[5] gpio_defaults_block_31/gpio_defaults[6]
+ gpio_defaults_block_31/gpio_defaults[7] gpio_defaults_block_31/gpio_defaults[8]
+ gpio_defaults_block_31/gpio_defaults[9] housekeeping/mgmt_gpio_in[31] gpio_control_in_2\[6\]/one
+ housekeeping/mgmt_gpio_in[31] gpio_control_in_2\[6\]/one padframe/mprj_io_analog_en[20]
+ padframe/mprj_io_analog_pol[20] padframe/mprj_io_analog_sel[20] padframe/mprj_io_dm[60]
+ padframe/mprj_io_dm[61] padframe/mprj_io_dm[62] padframe/mprj_io_holdover[20] padframe/mprj_io_ib_mode_sel[20]
+ padframe/mprj_io_in[20] padframe/mprj_io_inp_dis[20] padframe/mprj_io_out[20] padframe/mprj_io_oeb[20]
+ padframe/mprj_io_slow_sel[20] padframe/mprj_io_vtrip_sel[20] gpio_control_in_2\[6\]/resetn
+ gpio_control_in_2\[5\]/resetn gpio_control_in_2\[6\]/serial_clock gpio_control_in_2\[5\]/serial_clock
+ gpio_control_in_2\[6\]/serial_data_in gpio_control_in_2\[5\]/serial_data_in gpio_control_in_2\[6\]/serial_load
+ gpio_control_in_2\[5\]/serial_load mprj/io_in[20] mprj/io_oeb[20] mprj/io_out[20]
+ vccd_core vccd1_core VSUBS vssd1_core gpio_control_in_2\[6\]/zero gpio_control_block
Xgpio_control_in_1\[1\] gpio_defaults_block_9/gpio_defaults[0] gpio_defaults_block_9/gpio_defaults[10]
+ gpio_defaults_block_9/gpio_defaults[11] gpio_defaults_block_9/gpio_defaults[12]
+ gpio_defaults_block_9/gpio_defaults[1] gpio_defaults_block_9/gpio_defaults[2] gpio_defaults_block_9/gpio_defaults[3]
+ gpio_defaults_block_9/gpio_defaults[4] gpio_defaults_block_9/gpio_defaults[5] gpio_defaults_block_9/gpio_defaults[6]
+ gpio_defaults_block_9/gpio_defaults[7] gpio_defaults_block_9/gpio_defaults[8] gpio_defaults_block_9/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[9] gpio_control_in_1\[1\]/one housekeeping/mgmt_gpio_in[9]
+ gpio_control_in_1\[1\]/one padframe/mprj_io_analog_en[9] padframe/mprj_io_analog_pol[9]
+ padframe/mprj_io_analog_sel[9] padframe/mprj_io_dm[27] padframe/mprj_io_dm[28] padframe/mprj_io_dm[29]
+ padframe/mprj_io_holdover[9] padframe/mprj_io_ib_mode_sel[9] padframe/mprj_io_in[9]
+ padframe/mprj_io_inp_dis[9] padframe/mprj_io_out[9] padframe/mprj_io_oeb[9] padframe/mprj_io_slow_sel[9]
+ padframe/mprj_io_vtrip_sel[9] gpio_control_in_1\[1\]/resetn gpio_control_in_1\[2\]/resetn
+ gpio_control_in_1\[1\]/serial_clock gpio_control_in_1\[2\]/serial_clock gpio_control_in_1\[1\]/serial_data_in
+ gpio_control_in_1\[2\]/serial_data_in gpio_control_in_1\[1\]/serial_load gpio_control_in_1\[2\]/serial_load
+ mprj/io_in[9] mprj/io_oeb[9] mprj/io_out[9] vccd_core vccd1_core VSUBS vssd1_core
+ gpio_control_in_1\[1\]/zero gpio_control_block
Xmprj mprj/gpio_analog[0] mprj/gpio_analog[10] mprj/gpio_analog[11] mprj/gpio_analog[12]
+ mprj/gpio_analog[13] mprj/gpio_analog[14] mprj/gpio_analog[15] mprj/gpio_analog[16]
+ mprj/gpio_analog[17] mprj/gpio_analog[1] mprj/gpio_analog[2] mprj/gpio_analog[3]
+ mprj/gpio_analog[4] mprj/gpio_analog[5] mprj/gpio_analog[6] mprj/gpio_analog[7]
+ mprj/gpio_analog[8] mprj/gpio_analog[9] mprj/gpio_noesd[0] mprj/gpio_noesd[10] mprj/gpio_noesd[11]
+ mprj/gpio_noesd[12] mprj/gpio_noesd[13] mprj/gpio_noesd[14] mprj/gpio_noesd[15]
+ mprj/gpio_noesd[16] mprj/gpio_noesd[17] mprj/gpio_noesd[1] mprj/gpio_noesd[2] mprj/gpio_noesd[3]
+ mprj/gpio_noesd[4] mprj/gpio_noesd[5] mprj/gpio_noesd[6] mprj/gpio_noesd[7] mprj/gpio_noesd[8]
+ mprj/gpio_noesd[9] mprj/io_analog[0] mprj/io_analog[10] mprj/io_analog[1] mprj/io_analog[2]
+ mprj/io_analog[3] mprj/io_analog[7] mprj/io_analog[8] mprj/io_analog[9] mprj/io_analog[4]
+ mprj/io_analog[5] mprj/io_analog[6] mprj/io_clamp_high[0] mprj/io_clamp_high[1]
+ mprj/io_clamp_high[2] mprj/io_clamp_low[0] mprj/io_clamp_low[1] mprj/io_clamp_low[2]
+ mprj/io_in[0] mprj/io_in[10] mprj/io_in[11] mprj/io_in[12] mprj/io_in[13] mprj/io_in[14]
+ mprj/io_in[15] mprj/io_in[16] mprj/io_in[17] mprj/io_in[18] mprj/io_in[19] mprj/io_in[1]
+ mprj/io_in[20] mprj/io_in[21] mprj/io_in[22] mprj/io_in[23] mprj/io_in[24] mprj/io_in[25]
+ mprj/io_in[26] mprj/io_in[2] mprj/io_in[3] mprj/io_in[4] mprj/io_in[5] mprj/io_in[6]
+ mprj/io_in[7] mprj/io_in[8] mprj/io_in[9] mprj/io_in_3v3[0] mprj/io_in_3v3[10] mprj/io_in_3v3[11]
+ mprj/io_in_3v3[12] mprj/io_in_3v3[13] mprj/io_in_3v3[14] mprj/io_in_3v3[15] mprj/io_in_3v3[16]
+ mprj/io_in_3v3[17] mprj/io_in_3v3[18] mprj/io_in_3v3[19] mprj/io_in_3v3[1] mprj/io_in_3v3[20]
+ mprj/io_in_3v3[21] mprj/io_in_3v3[22] mprj/io_in_3v3[23] mprj/io_in_3v3[24] mprj/io_in_3v3[25]
+ mprj/io_in_3v3[26] mprj/io_in_3v3[2] mprj/io_in_3v3[3] mprj/io_in_3v3[4] mprj/io_in_3v3[5]
+ mprj/io_in_3v3[6] mprj/io_in_3v3[7] mprj/io_in_3v3[8] mprj/io_in_3v3[9] mprj/io_oeb[0]
+ mprj/io_oeb[10] mprj/io_oeb[11] mprj/io_oeb[12] mprj/io_oeb[13] mprj/io_oeb[14]
+ mprj/io_oeb[15] mprj/io_oeb[16] mprj/io_oeb[17] mprj/io_oeb[18] mprj/io_oeb[19]
+ mprj/io_oeb[1] mprj/io_oeb[20] mprj/io_oeb[21] mprj/io_oeb[22] mprj/io_oeb[23] mprj/io_oeb[24]
+ mprj/io_oeb[25] mprj/io_oeb[26] mprj/io_oeb[2] mprj/io_oeb[3] mprj/io_oeb[4] mprj/io_oeb[5]
+ mprj/io_oeb[6] mprj/io_oeb[7] mprj/io_oeb[8] mprj/io_oeb[9] mprj/io_out[0] mprj/io_out[10]
+ mprj/io_out[11] mprj/io_out[12] mprj/io_out[13] mprj/io_out[14] mprj/io_out[15]
+ mprj/io_out[16] mprj/io_out[17] mprj/io_out[18] mprj/io_out[19] mprj/io_out[1] mprj/io_out[20]
+ mprj/io_out[21] mprj/io_out[22] mprj/io_out[23] mprj/io_out[24] mprj/io_out[25]
+ mprj/io_out[26] mprj/io_out[2] mprj/io_out[3] mprj/io_out[4] mprj/io_out[5] mprj/io_out[6]
+ mprj/io_out[7] mprj/io_out[8] mprj/io_out[9] mprj/la_data_in[0] mprj/la_data_in[100]
+ mprj/la_data_in[101] mprj/la_data_in[102] mprj/la_data_in[103] mprj/la_data_in[104]
+ mprj/la_data_in[105] mprj/la_data_in[106] mprj/la_data_in[107] mprj/la_data_in[108]
+ mprj/la_data_in[109] mprj/la_data_in[10] mprj/la_data_in[110] mprj/la_data_in[111]
+ mprj/la_data_in[112] mprj/la_data_in[113] mprj/la_data_in[114] mprj/la_data_in[115]
+ mprj/la_data_in[116] mprj/la_data_in[117] mprj/la_data_in[118] mprj/la_data_in[119]
+ mprj/la_data_in[11] mprj/la_data_in[120] mprj/la_data_in[121] mprj/la_data_in[122]
+ mprj/la_data_in[123] mprj/la_data_in[124] mprj/la_data_in[125] mprj/la_data_in[126]
+ mprj/la_data_in[127] mprj/la_data_in[12] mprj/la_data_in[13] mprj/la_data_in[14]
+ mprj/la_data_in[15] mprj/la_data_in[16] mprj/la_data_in[17] mprj/la_data_in[18]
+ mprj/la_data_in[19] mprj/la_data_in[1] mprj/la_data_in[20] mprj/la_data_in[21] mprj/la_data_in[22]
+ mprj/la_data_in[23] mprj/la_data_in[24] mprj/la_data_in[25] mprj/la_data_in[26]
+ mprj/la_data_in[27] mprj/la_data_in[28] mprj/la_data_in[29] mprj/la_data_in[2] mprj/la_data_in[30]
+ mprj/la_data_in[31] mprj/la_data_in[32] mprj/la_data_in[33] mprj/la_data_in[34]
+ mprj/la_data_in[35] mprj/la_data_in[36] mprj/la_data_in[37] mprj/la_data_in[38]
+ mprj/la_data_in[39] mprj/la_data_in[3] mprj/la_data_in[40] mprj/la_data_in[41] mprj/la_data_in[42]
+ mprj/la_data_in[43] mprj/la_data_in[44] mprj/la_data_in[45] mprj/la_data_in[46]
+ mprj/la_data_in[47] mprj/la_data_in[48] mprj/la_data_in[49] mprj/la_data_in[4] mprj/la_data_in[50]
+ mprj/la_data_in[51] mprj/la_data_in[52] mprj/la_data_in[53] mprj/la_data_in[54]
+ mprj/la_data_in[55] mprj/la_data_in[56] mprj/la_data_in[57] mprj/la_data_in[58]
+ mprj/la_data_in[59] mprj/la_data_in[5] mprj/la_data_in[60] mprj/la_data_in[61] mprj/la_data_in[62]
+ mprj/la_data_in[63] mprj/la_data_in[64] mprj/la_data_in[65] mprj/la_data_in[66]
+ mprj/la_data_in[67] mprj/la_data_in[68] mprj/la_data_in[69] mprj/la_data_in[6] mprj/la_data_in[70]
+ mprj/la_data_in[71] mprj/la_data_in[72] mprj/la_data_in[73] mprj/la_data_in[74]
+ mprj/la_data_in[75] mprj/la_data_in[76] mprj/la_data_in[77] mprj/la_data_in[78]
+ mprj/la_data_in[79] mprj/la_data_in[7] mprj/la_data_in[80] mprj/la_data_in[81] mprj/la_data_in[82]
+ mprj/la_data_in[83] mprj/la_data_in[84] mprj/la_data_in[85] mprj/la_data_in[86]
+ mprj/la_data_in[87] mprj/la_data_in[88] mprj/la_data_in[89] mprj/la_data_in[8] mprj/la_data_in[90]
+ mprj/la_data_in[91] mprj/la_data_in[92] mprj/la_data_in[93] mprj/la_data_in[94]
+ mprj/la_data_in[95] mprj/la_data_in[96] mprj/la_data_in[97] mprj/la_data_in[98]
+ mprj/la_data_in[99] mprj/la_data_in[9] mprj/la_data_out[0] mprj/la_data_out[100]
+ mprj/la_data_out[101] mprj/la_data_out[102] mprj/la_data_out[103] mprj/la_data_out[104]
+ mprj/la_data_out[105] mprj/la_data_out[106] mprj/la_data_out[107] mprj/la_data_out[108]
+ mprj/la_data_out[109] mprj/la_data_out[10] mprj/la_data_out[110] mprj/la_data_out[111]
+ mprj/la_data_out[112] mprj/la_data_out[113] mprj/la_data_out[114] mprj/la_data_out[115]
+ mprj/la_data_out[116] mprj/la_data_out[117] mprj/la_data_out[118] mprj/la_data_out[119]
+ mprj/la_data_out[11] mprj/la_data_out[120] mprj/la_data_out[121] mprj/la_data_out[122]
+ mprj/la_data_out[123] mprj/la_data_out[124] mprj/la_data_out[125] mprj/la_data_out[126]
+ mprj/la_data_out[127] mprj/la_data_out[12] mprj/la_data_out[13] mprj/la_data_out[14]
+ mprj/la_data_out[15] mprj/la_data_out[16] mprj/la_data_out[17] mprj/la_data_out[18]
+ mprj/la_data_out[19] mprj/la_data_out[1] mprj/la_data_out[20] mprj/la_data_out[21]
+ mprj/la_data_out[22] mprj/la_data_out[23] mprj/la_data_out[24] mprj/la_data_out[25]
+ mprj/la_data_out[26] mprj/la_data_out[27] mprj/la_data_out[28] mprj/la_data_out[29]
+ mprj/la_data_out[2] mprj/la_data_out[30] mprj/la_data_out[31] mprj/la_data_out[32]
+ mprj/la_data_out[33] mprj/la_data_out[34] mprj/la_data_out[35] mprj/la_data_out[36]
+ mprj/la_data_out[37] mprj/la_data_out[38] mprj/la_data_out[39] mprj/la_data_out[3]
+ mprj/la_data_out[40] mprj/la_data_out[41] mprj/la_data_out[42] mprj/la_data_out[43]
+ mprj/la_data_out[44] mprj/la_data_out[45] mprj/la_data_out[46] mprj/la_data_out[47]
+ mprj/la_data_out[48] mprj/la_data_out[49] mprj/la_data_out[4] mprj/la_data_out[50]
+ mprj/la_data_out[51] mprj/la_data_out[52] mprj/la_data_out[53] mprj/la_data_out[54]
+ mprj/la_data_out[55] mprj/la_data_out[56] mprj/la_data_out[57] mprj/la_data_out[58]
+ mprj/la_data_out[59] mprj/la_data_out[5] mprj/la_data_out[60] mprj/la_data_out[61]
+ mprj/la_data_out[62] mprj/la_data_out[63] mprj/la_data_out[64] mprj/la_data_out[65]
+ mprj/la_data_out[66] mprj/la_data_out[67] mprj/la_data_out[68] mprj/la_data_out[69]
+ mprj/la_data_out[6] mprj/la_data_out[70] mprj/la_data_out[71] mprj/la_data_out[72]
+ mprj/la_data_out[73] mprj/la_data_out[74] mprj/la_data_out[75] mprj/la_data_out[76]
+ mprj/la_data_out[77] mprj/la_data_out[78] mprj/la_data_out[79] mprj/la_data_out[7]
+ mprj/la_data_out[80] mprj/la_data_out[81] mprj/la_data_out[82] mprj/la_data_out[83]
+ mprj/la_data_out[84] mprj/la_data_out[85] mprj/la_data_out[86] mprj/la_data_out[87]
+ mprj/la_data_out[88] mprj/la_data_out[89] mprj/la_data_out[8] mprj/la_data_out[90]
+ mprj/la_data_out[91] mprj/la_data_out[92] mprj/la_data_out[93] mprj/la_data_out[94]
+ mprj/la_data_out[95] mprj/la_data_out[96] mprj/la_data_out[97] mprj/la_data_out[98]
+ mprj/la_data_out[99] mprj/la_data_out[9] mprj/la_oenb[0] mprj/la_oenb[100] mprj/la_oenb[101]
+ mprj/la_oenb[102] mprj/la_oenb[103] mprj/la_oenb[104] mprj/la_oenb[105] mprj/la_oenb[106]
+ mprj/la_oenb[107] mprj/la_oenb[108] mprj/la_oenb[109] mprj/la_oenb[10] mprj/la_oenb[110]
+ mprj/la_oenb[111] mprj/la_oenb[112] mprj/la_oenb[113] mprj/la_oenb[114] mprj/la_oenb[115]
+ mprj/la_oenb[116] mprj/la_oenb[117] mprj/la_oenb[118] mprj/la_oenb[119] mprj/la_oenb[11]
+ mprj/la_oenb[120] mprj/la_oenb[121] mprj/la_oenb[122] mprj/la_oenb[123] mprj/la_oenb[124]
+ mprj/la_oenb[125] mprj/la_oenb[126] mprj/la_oenb[127] mprj/la_oenb[12] mprj/la_oenb[13]
+ mprj/la_oenb[14] mprj/la_oenb[15] mprj/la_oenb[16] mprj/la_oenb[17] mprj/la_oenb[18]
+ mprj/la_oenb[19] mprj/la_oenb[1] mprj/la_oenb[20] mprj/la_oenb[21] mprj/la_oenb[22]
+ mprj/la_oenb[23] mprj/la_oenb[24] mprj/la_oenb[25] mprj/la_oenb[26] mprj/la_oenb[27]
+ mprj/la_oenb[28] mprj/la_oenb[29] mprj/la_oenb[2] mprj/la_oenb[30] mprj/la_oenb[31]
+ mprj/la_oenb[32] mprj/la_oenb[33] mprj/la_oenb[34] mprj/la_oenb[35] mprj/la_oenb[36]
+ mprj/la_oenb[37] mprj/la_oenb[38] mprj/la_oenb[39] mprj/la_oenb[3] mprj/la_oenb[40]
+ mprj/la_oenb[41] mprj/la_oenb[42] mprj/la_oenb[43] mprj/la_oenb[44] mprj/la_oenb[45]
+ mprj/la_oenb[46] mprj/la_oenb[47] mprj/la_oenb[48] mprj/la_oenb[49] mprj/la_oenb[4]
+ mprj/la_oenb[50] mprj/la_oenb[51] mprj/la_oenb[52] mprj/la_oenb[53] mprj/la_oenb[54]
+ mprj/la_oenb[55] mprj/la_oenb[56] mprj/la_oenb[57] mprj/la_oenb[58] mprj/la_oenb[59]
+ mprj/la_oenb[5] mprj/la_oenb[60] mprj/la_oenb[61] mprj/la_oenb[62] mprj/la_oenb[63]
+ mprj/la_oenb[64] mprj/la_oenb[65] mprj/la_oenb[66] mprj/la_oenb[67] mprj/la_oenb[68]
+ mprj/la_oenb[69] mprj/la_oenb[6] mprj/la_oenb[70] mprj/la_oenb[71] mprj/la_oenb[72]
+ mprj/la_oenb[73] mprj/la_oenb[74] mprj/la_oenb[75] mprj/la_oenb[76] mprj/la_oenb[77]
+ mprj/la_oenb[78] mprj/la_oenb[79] mprj/la_oenb[7] mprj/la_oenb[80] mprj/la_oenb[81]
+ mprj/la_oenb[82] mprj/la_oenb[83] mprj/la_oenb[84] mprj/la_oenb[85] mprj/la_oenb[86]
+ mprj/la_oenb[87] mprj/la_oenb[88] mprj/la_oenb[89] mprj/la_oenb[8] mprj/la_oenb[90]
+ mprj/la_oenb[91] mprj/la_oenb[92] mprj/la_oenb[93] mprj/la_oenb[94] mprj/la_oenb[95]
+ mprj/la_oenb[96] mprj/la_oenb[97] mprj/la_oenb[98] mprj/la_oenb[99] mprj/la_oenb[9]
+ mprj/user_clock2 mprj/user_irq[0] mprj/user_irq[1] mprj/user_irq[2] vccd1_core vccd2_core
+ vdda1_core vdda2_core vssa1_core vssa2_core vssd1_core vssd2_core mprj/wb_clk_i
+ mprj/wb_rst_i mprj/wbs_ack_o mprj/wbs_adr_i[0] mprj/wbs_adr_i[10] mprj/wbs_adr_i[11]
+ mprj/wbs_adr_i[12] mprj/wbs_adr_i[13] mprj/wbs_adr_i[14] mprj/wbs_adr_i[15] mprj/wbs_adr_i[16]
+ mprj/wbs_adr_i[17] mprj/wbs_adr_i[18] mprj/wbs_adr_i[19] mprj/wbs_adr_i[1] mprj/wbs_adr_i[20]
+ mprj/wbs_adr_i[21] mprj/wbs_adr_i[22] mprj/wbs_adr_i[23] mprj/wbs_adr_i[24] mprj/wbs_adr_i[25]
+ mprj/wbs_adr_i[26] mprj/wbs_adr_i[27] mprj/wbs_adr_i[28] mprj/wbs_adr_i[29] mprj/wbs_adr_i[2]
+ mprj/wbs_adr_i[30] mprj/wbs_adr_i[31] mprj/wbs_adr_i[3] mprj/wbs_adr_i[4] mprj/wbs_adr_i[5]
+ mprj/wbs_adr_i[6] mprj/wbs_adr_i[7] mprj/wbs_adr_i[8] mprj/wbs_adr_i[9] mprj/wbs_cyc_i
+ mprj/wbs_dat_i[0] mprj/wbs_dat_i[10] mprj/wbs_dat_i[11] mprj/wbs_dat_i[12] mprj/wbs_dat_i[13]
+ mprj/wbs_dat_i[14] mprj/wbs_dat_i[15] mprj/wbs_dat_i[16] mprj/wbs_dat_i[17] mprj/wbs_dat_i[18]
+ mprj/wbs_dat_i[19] mprj/wbs_dat_i[1] mprj/wbs_dat_i[20] mprj/wbs_dat_i[21] mprj/wbs_dat_i[22]
+ mprj/wbs_dat_i[23] mprj/wbs_dat_i[24] mprj/wbs_dat_i[25] mprj/wbs_dat_i[26] mprj/wbs_dat_i[27]
+ mprj/wbs_dat_i[28] mprj/wbs_dat_i[29] mprj/wbs_dat_i[2] mprj/wbs_dat_i[30] mprj/wbs_dat_i[31]
+ mprj/wbs_dat_i[3] mprj/wbs_dat_i[4] mprj/wbs_dat_i[5] mprj/wbs_dat_i[6] mprj/wbs_dat_i[7]
+ mprj/wbs_dat_i[8] mprj/wbs_dat_i[9] mprj/wbs_dat_o[0] mprj/wbs_dat_o[10] mprj/wbs_dat_o[11]
+ mprj/wbs_dat_o[12] mprj/wbs_dat_o[13] mprj/wbs_dat_o[14] mprj/wbs_dat_o[15] mprj/wbs_dat_o[16]
+ mprj/wbs_dat_o[17] mprj/wbs_dat_o[18] mprj/wbs_dat_o[19] mprj/wbs_dat_o[1] mprj/wbs_dat_o[20]
+ mprj/wbs_dat_o[21] mprj/wbs_dat_o[22] mprj/wbs_dat_o[23] mprj/wbs_dat_o[24] mprj/wbs_dat_o[25]
+ mprj/wbs_dat_o[26] mprj/wbs_dat_o[27] mprj/wbs_dat_o[28] mprj/wbs_dat_o[29] mprj/wbs_dat_o[2]
+ mprj/wbs_dat_o[30] mprj/wbs_dat_o[31] mprj/wbs_dat_o[3] mprj/wbs_dat_o[4] mprj/wbs_dat_o[5]
+ mprj/wbs_dat_o[6] mprj/wbs_dat_o[7] mprj/wbs_dat_o[8] mprj/wbs_dat_o[9] mprj/wbs_sel_i[0]
+ mprj/wbs_sel_i[1] mprj/wbs_sel_i[2] mprj/wbs_sel_i[3] mprj/wbs_stb_i mprj/wbs_we_i
+ user_analog_project_wrapper
Xgpio_control_in_2\[4\] gpio_defaults_block_29/gpio_defaults[0] gpio_defaults_block_29/gpio_defaults[10]
+ gpio_defaults_block_29/gpio_defaults[11] gpio_defaults_block_29/gpio_defaults[12]
+ gpio_defaults_block_29/gpio_defaults[1] gpio_defaults_block_29/gpio_defaults[2]
+ gpio_defaults_block_29/gpio_defaults[3] gpio_defaults_block_29/gpio_defaults[4]
+ gpio_defaults_block_29/gpio_defaults[5] gpio_defaults_block_29/gpio_defaults[6]
+ gpio_defaults_block_29/gpio_defaults[7] gpio_defaults_block_29/gpio_defaults[8]
+ gpio_defaults_block_29/gpio_defaults[9] housekeeping/mgmt_gpio_in[29] gpio_control_in_2\[4\]/one
+ housekeeping/mgmt_gpio_in[29] gpio_control_in_2\[4\]/one padframe/mprj_io_analog_en[18]
+ padframe/mprj_io_analog_pol[18] padframe/mprj_io_analog_sel[18] padframe/mprj_io_dm[54]
+ padframe/mprj_io_dm[55] padframe/mprj_io_dm[56] padframe/mprj_io_holdover[18] padframe/mprj_io_ib_mode_sel[18]
+ padframe/mprj_io_in[18] padframe/mprj_io_inp_dis[18] padframe/mprj_io_out[18] padframe/mprj_io_oeb[18]
+ padframe/mprj_io_slow_sel[18] padframe/mprj_io_vtrip_sel[18] gpio_control_in_2\[4\]/resetn
+ gpio_control_in_2\[3\]/resetn gpio_control_in_2\[4\]/serial_clock gpio_control_in_2\[3\]/serial_clock
+ gpio_control_in_2\[4\]/serial_data_in gpio_control_in_2\[3\]/serial_data_in gpio_control_in_2\[4\]/serial_load
+ gpio_control_in_2\[3\]/serial_load mprj/io_in[18] mprj/io_oeb[18] mprj/io_out[18]
+ vccd_core vccd1_core VSUBS vssd1_core gpio_control_in_2\[4\]/zero gpio_control_block
Xgpio_control_bidir_1\[1\] gpio_defaults_block_1/gpio_defaults[0] gpio_defaults_block_1/gpio_defaults[10]
+ gpio_defaults_block_1/gpio_defaults[11] gpio_defaults_block_1/gpio_defaults[12]
+ gpio_defaults_block_1/gpio_defaults[1] gpio_defaults_block_1/gpio_defaults[2] gpio_defaults_block_1/gpio_defaults[3]
+ gpio_defaults_block_1/gpio_defaults[4] gpio_defaults_block_1/gpio_defaults[5] gpio_defaults_block_1/gpio_defaults[6]
+ gpio_defaults_block_1/gpio_defaults[7] gpio_defaults_block_1/gpio_defaults[8] gpio_defaults_block_1/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[1] gpio_control_bidir_1\[1\]/mgmt_gpio_oeb gpio_control_bidir_1\[1\]/mgmt_gpio_out
+ gpio_control_bidir_1\[1\]/one padframe/mprj_io_analog_en[1] padframe/mprj_io_analog_pol[1]
+ padframe/mprj_io_analog_sel[1] padframe/mprj_io_dm[3] padframe/mprj_io_dm[4] padframe/mprj_io_dm[5]
+ padframe/mprj_io_holdover[1] padframe/mprj_io_ib_mode_sel[1] padframe/mprj_io_in[1]
+ padframe/mprj_io_inp_dis[1] padframe/mprj_io_out[1] padframe/mprj_io_oeb[1] padframe/mprj_io_slow_sel[1]
+ padframe/mprj_io_vtrip_sel[1] gpio_control_bidir_1\[1\]/resetn gpio_control_in_1a\[0\]/resetn
+ gpio_control_bidir_1\[1\]/serial_clock gpio_control_in_1a\[0\]/serial_clock gpio_control_bidir_1\[1\]/serial_data_in
+ gpio_control_in_1a\[0\]/serial_data_in gpio_control_bidir_1\[1\]/serial_load gpio_control_in_1a\[0\]/serial_load
+ mprj/io_in[1] mprj/io_oeb[1] mprj/io_out[1] vccd_core vccd1_core VSUBS vssd1_core
+ gpio_control_bidir_1\[1\]/zero gpio_control_block
Xhousekeeping VSUBS vccd_core soc/debug_in soc/debug_mode soc/debug_oeb soc/debug_out
+ soc/irq[3] soc/irq[4] soc/irq[5] user_id_value/mask_rev[0] user_id_value/mask_rev[10]
+ user_id_value/mask_rev[11] user_id_value/mask_rev[12] user_id_value/mask_rev[13]
+ user_id_value/mask_rev[14] user_id_value/mask_rev[15] user_id_value/mask_rev[16]
+ user_id_value/mask_rev[17] user_id_value/mask_rev[18] user_id_value/mask_rev[19]
+ user_id_value/mask_rev[1] user_id_value/mask_rev[20] user_id_value/mask_rev[21]
+ user_id_value/mask_rev[22] user_id_value/mask_rev[23] user_id_value/mask_rev[24]
+ user_id_value/mask_rev[25] user_id_value/mask_rev[26] user_id_value/mask_rev[27]
+ user_id_value/mask_rev[28] user_id_value/mask_rev[29] user_id_value/mask_rev[2]
+ user_id_value/mask_rev[30] user_id_value/mask_rev[31] user_id_value/mask_rev[3]
+ user_id_value/mask_rev[4] user_id_value/mask_rev[5] user_id_value/mask_rev[6] user_id_value/mask_rev[7]
+ user_id_value/mask_rev[8] user_id_value/mask_rev[9] housekeeping/mgmt_gpio_in[0]
+ housekeeping/mgmt_gpio_in[10] housekeeping/mgmt_gpio_in[11] housekeeping/mgmt_gpio_in[12]
+ housekeeping/mgmt_gpio_in[13] housekeeping/mgmt_gpio_in[14] housekeeping/mgmt_gpio_in[15]
+ housekeeping/mgmt_gpio_in[16] housekeeping/mgmt_gpio_in[17] housekeeping/mgmt_gpio_in[18]
+ housekeeping/mgmt_gpio_in[19] housekeeping/mgmt_gpio_in[1] housekeeping/mgmt_gpio_in[20]
+ housekeeping/mgmt_gpio_in[21] housekeeping/mgmt_gpio_in[22] housekeeping/mgmt_gpio_in[23]
+ housekeeping/mgmt_gpio_in[24] housekeeping/mgmt_gpio_in[25] housekeeping/mgmt_gpio_in[26]
+ housekeeping/mgmt_gpio_in[27] housekeeping/mgmt_gpio_in[28] housekeeping/mgmt_gpio_in[29]
+ housekeeping/mgmt_gpio_in[2] housekeeping/mgmt_gpio_in[30] housekeeping/mgmt_gpio_in[31]
+ housekeeping/mgmt_gpio_in[32] housekeeping/mgmt_gpio_in[33] housekeeping/mgmt_gpio_in[34]
+ housekeeping/mgmt_gpio_in[35] housekeeping/mgmt_gpio_in[36] housekeeping/mgmt_gpio_in[37]
+ housekeeping/mgmt_gpio_in[3] housekeeping/mgmt_gpio_in[4] housekeeping/mgmt_gpio_in[5]
+ housekeeping/mgmt_gpio_in[6] housekeeping/mgmt_gpio_in[7] housekeeping/mgmt_gpio_in[8]
+ housekeeping/mgmt_gpio_in[9] housekeeping/mgmt_gpio_oeb[0] housekeeping/mgmt_gpio_oeb[10]
+ housekeeping/mgmt_gpio_oeb[11] housekeeping/mgmt_gpio_oeb[12] housekeeping/mgmt_gpio_oeb[13]
+ housekeeping/mgmt_gpio_oeb[14] housekeeping/mgmt_gpio_oeb[15] housekeeping/mgmt_gpio_oeb[16]
+ housekeeping/mgmt_gpio_oeb[17] housekeeping/mgmt_gpio_oeb[18] housekeeping/mgmt_gpio_oeb[19]
+ housekeeping/mgmt_gpio_oeb[1] housekeeping/mgmt_gpio_oeb[20] housekeeping/mgmt_gpio_oeb[21]
+ housekeeping/mgmt_gpio_oeb[22] housekeeping/mgmt_gpio_oeb[23] housekeeping/mgmt_gpio_oeb[24]
+ housekeeping/mgmt_gpio_oeb[25] housekeeping/mgmt_gpio_oeb[26] housekeeping/mgmt_gpio_oeb[27]
+ housekeeping/mgmt_gpio_oeb[28] housekeeping/mgmt_gpio_oeb[29] housekeeping/mgmt_gpio_oeb[2]
+ housekeeping/mgmt_gpio_oeb[30] housekeeping/mgmt_gpio_oeb[31] housekeeping/mgmt_gpio_oeb[32]
+ housekeeping/mgmt_gpio_oeb[33] housekeeping/mgmt_gpio_oeb[34] housekeeping/mgmt_gpio_oeb[35]
+ housekeeping/mgmt_gpio_oeb[36] housekeeping/mgmt_gpio_oeb[37] housekeeping/mgmt_gpio_oeb[3]
+ housekeeping/mgmt_gpio_oeb[4] housekeeping/mgmt_gpio_oeb[5] housekeeping/mgmt_gpio_oeb[6]
+ housekeeping/mgmt_gpio_oeb[7] housekeeping/mgmt_gpio_oeb[8] housekeeping/mgmt_gpio_oeb[9]
+ housekeeping/mgmt_gpio_out[0] housekeeping/mgmt_gpio_in[10] housekeeping/mgmt_gpio_in[11]
+ housekeeping/mgmt_gpio_in[12] housekeeping/mgmt_gpio_in[13] housekeeping/mgmt_gpio_in[14]
+ housekeeping/mgmt_gpio_in[15] housekeeping/mgmt_gpio_in[16] housekeeping/mgmt_gpio_in[17]
+ housekeeping/mgmt_gpio_in[18] housekeeping/mgmt_gpio_in[19] housekeeping/mgmt_gpio_out[1]
+ housekeeping/mgmt_gpio_in[20] housekeeping/mgmt_gpio_in[21] housekeeping/mgmt_gpio_in[22]
+ housekeeping/mgmt_gpio_in[23] housekeeping/mgmt_gpio_in[24] housekeeping/mgmt_gpio_in[25]
+ housekeeping/mgmt_gpio_in[26] housekeeping/mgmt_gpio_in[27] housekeeping/mgmt_gpio_in[28]
+ housekeeping/mgmt_gpio_in[29] housekeeping/mgmt_gpio_in[2] housekeeping/mgmt_gpio_in[30]
+ housekeeping/mgmt_gpio_in[31] housekeeping/mgmt_gpio_in[32] housekeeping/mgmt_gpio_in[33]
+ housekeeping/mgmt_gpio_in[34] housekeeping/mgmt_gpio_out[35] housekeeping/mgmt_gpio_out[36]
+ housekeeping/mgmt_gpio_out[37] housekeeping/mgmt_gpio_in[3] housekeeping/mgmt_gpio_in[4]
+ housekeeping/mgmt_gpio_in[5] housekeeping/mgmt_gpio_in[6] housekeeping/mgmt_gpio_in[7]
+ housekeeping/mgmt_gpio_in[8] housekeeping/mgmt_gpio_in[9] padframe/flash_clk_core
+ padframe/flash_clk_oeb_core padframe/flash_csb_core padframe/flash_csb_oeb_core
+ padframe/flash_io0_di_core padframe/flash_io0_do_core padframe/flash_io0_ieb_core
+ padframe/flash_io0_oeb_core padframe/flash_io1_di_core padframe/flash_io1_do_core
+ padframe/flash_io1_ieb_core padframe/flash_io1_oeb_core clocking/sel2[0] clocking/sel2[1]
+ clocking/sel2[2] clocking/ext_clk_sel pll/dco pll/div[0] pll/div[1] pll/div[2] pll/div[3]
+ pll/div[4] pll/enable clocking/sel[0] clocking/sel[1] clocking/sel[2] pll/ext_trim[0]
+ pll/ext_trim[10] pll/ext_trim[11] pll/ext_trim[12] pll/ext_trim[13] pll/ext_trim[14]
+ pll/ext_trim[15] pll/ext_trim[16] pll/ext_trim[17] pll/ext_trim[18] pll/ext_trim[19]
+ pll/ext_trim[1] pll/ext_trim[20] pll/ext_trim[21] pll/ext_trim[22] pll/ext_trim[23]
+ pll/ext_trim[24] pll/ext_trim[25] pll/ext_trim[2] pll/ext_trim[3] pll/ext_trim[4]
+ pll/ext_trim[5] pll/ext_trim[6] pll/ext_trim[7] pll/ext_trim[8] pll/ext_trim[9]
+ por/porb_l housekeeping/pwr_ctrl_out[0] housekeeping/pwr_ctrl_out[1] housekeeping/pwr_ctrl_out[2]
+ housekeeping/pwr_ctrl_out[3] soc/qspi_enabled housekeeping/reset soc/ser_rx soc/ser_tx
+ housekeeping/serial_clock housekeeping/serial_data_1 housekeeping/serial_data_2
+ housekeeping/serial_load housekeeping/serial_resetn soc/spi_csb soc/spi_enabled
+ soc/spi_sck soc/spi_sdi soc/spi_sdo soc/spi_sdoenb soc/flash_clk soc/flash_csb soc/flash_io0_di
+ soc/flash_io0_do soc/flash_io0_oeb soc/flash_io1_di soc/flash_io1_do soc/flash_io1_oeb
+ soc/flash_io2_di soc/flash_io2_do soc/flash_io2_oeb soc/flash_io3_di soc/flash_io3_do
+ soc/flash_io3_oeb soc/sram_ro_addr[0] soc/sram_ro_addr[1] soc/sram_ro_addr[2] soc/sram_ro_addr[3]
+ soc/sram_ro_addr[4] soc/sram_ro_addr[5] soc/sram_ro_addr[6] soc/sram_ro_addr[7]
+ soc/sram_ro_clk soc/sram_ro_csb soc/sram_ro_data[0] soc/sram_ro_data[10] soc/sram_ro_data[11]
+ soc/sram_ro_data[12] soc/sram_ro_data[13] soc/sram_ro_data[14] soc/sram_ro_data[15]
+ soc/sram_ro_data[16] soc/sram_ro_data[17] soc/sram_ro_data[18] soc/sram_ro_data[19]
+ soc/sram_ro_data[1] soc/sram_ro_data[20] soc/sram_ro_data[21] soc/sram_ro_data[22]
+ soc/sram_ro_data[23] soc/sram_ro_data[24] soc/sram_ro_data[25] soc/sram_ro_data[26]
+ soc/sram_ro_data[27] soc/sram_ro_data[28] soc/sram_ro_data[29] soc/sram_ro_data[2]
+ soc/sram_ro_data[30] soc/sram_ro_data[31] soc/sram_ro_data[3] soc/sram_ro_data[4]
+ soc/sram_ro_data[5] soc/sram_ro_data[6] soc/sram_ro_data[7] soc/sram_ro_data[8]
+ soc/sram_ro_data[9] soc/trap soc/uart_enabled clocking/user_clk housekeeping/usr1_vcc_pwrgood
+ housekeeping/usr1_vdd_pwrgood housekeeping/usr2_vcc_pwrgood housekeeping/usr2_vdd_pwrgood
+ soc/hk_ack_i soc/mprj_adr_o[0] soc/mprj_adr_o[10] soc/mprj_adr_o[11] soc/mprj_adr_o[12]
+ soc/mprj_adr_o[13] soc/mprj_adr_o[14] soc/mprj_adr_o[15] soc/mprj_adr_o[16] soc/mprj_adr_o[17]
+ soc/mprj_adr_o[18] soc/mprj_adr_o[19] soc/mprj_adr_o[1] soc/mprj_adr_o[20] soc/mprj_adr_o[21]
+ soc/mprj_adr_o[22] soc/mprj_adr_o[23] soc/mprj_adr_o[24] soc/mprj_adr_o[25] soc/mprj_adr_o[26]
+ soc/mprj_adr_o[27] soc/mprj_adr_o[28] soc/mprj_adr_o[29] soc/mprj_adr_o[2] soc/mprj_adr_o[30]
+ soc/mprj_adr_o[31] soc/mprj_adr_o[3] soc/mprj_adr_o[4] soc/mprj_adr_o[5] soc/mprj_adr_o[6]
+ soc/mprj_adr_o[7] soc/mprj_adr_o[8] soc/mprj_adr_o[9] soc/core_clk soc/hk_cyc_o
+ soc/mprj_dat_o[0] soc/mprj_dat_o[10] soc/mprj_dat_o[11] soc/mprj_dat_o[12] soc/mprj_dat_o[13]
+ soc/mprj_dat_o[14] soc/mprj_dat_o[15] soc/mprj_dat_o[16] soc/mprj_dat_o[17] soc/mprj_dat_o[18]
+ soc/mprj_dat_o[19] soc/mprj_dat_o[1] soc/mprj_dat_o[20] soc/mprj_dat_o[21] soc/mprj_dat_o[22]
+ soc/mprj_dat_o[23] soc/mprj_dat_o[24] soc/mprj_dat_o[25] soc/mprj_dat_o[26] soc/mprj_dat_o[27]
+ soc/mprj_dat_o[28] soc/mprj_dat_o[29] soc/mprj_dat_o[2] soc/mprj_dat_o[30] soc/mprj_dat_o[31]
+ soc/mprj_dat_o[3] soc/mprj_dat_o[4] soc/mprj_dat_o[5] soc/mprj_dat_o[6] soc/mprj_dat_o[7]
+ soc/mprj_dat_o[8] soc/mprj_dat_o[9] soc/hk_dat_i[0] soc/hk_dat_i[10] soc/hk_dat_i[11]
+ soc/hk_dat_i[12] soc/hk_dat_i[13] soc/hk_dat_i[14] soc/hk_dat_i[15] soc/hk_dat_i[16]
+ soc/hk_dat_i[17] soc/hk_dat_i[18] soc/hk_dat_i[19] soc/hk_dat_i[1] soc/hk_dat_i[20]
+ soc/hk_dat_i[21] soc/hk_dat_i[22] soc/hk_dat_i[23] soc/hk_dat_i[24] soc/hk_dat_i[25]
+ soc/hk_dat_i[26] soc/hk_dat_i[27] soc/hk_dat_i[28] soc/hk_dat_i[29] soc/hk_dat_i[2]
+ soc/hk_dat_i[30] soc/hk_dat_i[31] soc/hk_dat_i[3] soc/hk_dat_i[4] soc/hk_dat_i[5]
+ soc/hk_dat_i[6] soc/hk_dat_i[7] soc/hk_dat_i[8] soc/hk_dat_i[9] soc/core_rstn soc/mprj_sel_o[0]
+ soc/mprj_sel_o[1] soc/mprj_sel_o[2] soc/mprj_sel_o[3] soc/hk_stb_o soc/mprj_we_o
+ housekeeping
Xgpio_control_in_2\[2\] gpio_defaults_block_27/gpio_defaults[0] gpio_defaults_block_27/gpio_defaults[10]
+ gpio_defaults_block_27/gpio_defaults[11] gpio_defaults_block_27/gpio_defaults[12]
+ gpio_defaults_block_27/gpio_defaults[1] gpio_defaults_block_27/gpio_defaults[2]
+ gpio_defaults_block_27/gpio_defaults[3] gpio_defaults_block_27/gpio_defaults[4]
+ gpio_defaults_block_27/gpio_defaults[5] gpio_defaults_block_27/gpio_defaults[6]
+ gpio_defaults_block_27/gpio_defaults[7] gpio_defaults_block_27/gpio_defaults[8]
+ gpio_defaults_block_27/gpio_defaults[9] housekeeping/mgmt_gpio_in[27] gpio_control_in_2\[2\]/one
+ housekeeping/mgmt_gpio_in[27] gpio_control_in_2\[2\]/one padframe/mprj_io_analog_en[16]
+ padframe/mprj_io_analog_pol[16] padframe/mprj_io_analog_sel[16] padframe/mprj_io_dm[48]
+ padframe/mprj_io_dm[49] padframe/mprj_io_dm[50] padframe/mprj_io_holdover[16] padframe/mprj_io_ib_mode_sel[16]
+ padframe/mprj_io_in[16] padframe/mprj_io_inp_dis[16] padframe/mprj_io_out[16] padframe/mprj_io_oeb[16]
+ padframe/mprj_io_slow_sel[16] padframe/mprj_io_vtrip_sel[16] gpio_control_in_2\[2\]/resetn
+ gpio_control_in_2\[1\]/resetn gpio_control_in_2\[2\]/serial_clock gpio_control_in_2\[1\]/serial_clock
+ gpio_control_in_2\[2\]/serial_data_in gpio_control_in_2\[1\]/serial_data_in gpio_control_in_2\[2\]/serial_load
+ gpio_control_in_2\[1\]/serial_load mprj/io_in[16] mprj/io_oeb[16] mprj/io_out[16]
+ vccd_core vccd1_core VSUBS vssd1_core gpio_control_in_2\[2\]/zero gpio_control_block
Xgpio_defaults_block_30 VSUBS vccd_core gpio_defaults_block_30/gpio_defaults[0] gpio_defaults_block_30/gpio_defaults[10]
+ gpio_defaults_block_30/gpio_defaults[11] gpio_defaults_block_30/gpio_defaults[12]
+ gpio_defaults_block_30/gpio_defaults[1] gpio_defaults_block_30/gpio_defaults[2]
+ gpio_defaults_block_30/gpio_defaults[3] gpio_defaults_block_30/gpio_defaults[4]
+ gpio_defaults_block_30/gpio_defaults[5] gpio_defaults_block_30/gpio_defaults[6]
+ gpio_defaults_block_30/gpio_defaults[7] gpio_defaults_block_30/gpio_defaults[8]
+ gpio_defaults_block_30/gpio_defaults[9] gpio_defaults_block
Xgpio_defaults_block_10 VSUBS vccd_core gpio_defaults_block_10/gpio_defaults[0] gpio_defaults_block_10/gpio_defaults[10]
+ gpio_defaults_block_10/gpio_defaults[11] gpio_defaults_block_10/gpio_defaults[12]
+ gpio_defaults_block_10/gpio_defaults[1] gpio_defaults_block_10/gpio_defaults[2]
+ gpio_defaults_block_10/gpio_defaults[3] gpio_defaults_block_10/gpio_defaults[4]
+ gpio_defaults_block_10/gpio_defaults[5] gpio_defaults_block_10/gpio_defaults[6]
+ gpio_defaults_block_10/gpio_defaults[7] gpio_defaults_block_10/gpio_defaults[8]
+ gpio_defaults_block_10/gpio_defaults[9] gpio_defaults_block
Xgpio_defaults_block_31 VSUBS vccd_core gpio_defaults_block_31/gpio_defaults[0] gpio_defaults_block_31/gpio_defaults[10]
+ gpio_defaults_block_31/gpio_defaults[11] gpio_defaults_block_31/gpio_defaults[12]
+ gpio_defaults_block_31/gpio_defaults[1] gpio_defaults_block_31/gpio_defaults[2]
+ gpio_defaults_block_31/gpio_defaults[3] gpio_defaults_block_31/gpio_defaults[4]
+ gpio_defaults_block_31/gpio_defaults[5] gpio_defaults_block_31/gpio_defaults[6]
+ gpio_defaults_block_31/gpio_defaults[7] gpio_defaults_block_31/gpio_defaults[8]
+ gpio_defaults_block_31/gpio_defaults[9] gpio_defaults_block
Xgpio_control_in_1a\[5\] gpio_defaults_block_7/gpio_defaults[0] gpio_defaults_block_7/gpio_defaults[10]
+ gpio_defaults_block_7/gpio_defaults[11] gpio_defaults_block_7/gpio_defaults[12]
+ gpio_defaults_block_7/gpio_defaults[1] gpio_defaults_block_7/gpio_defaults[2] gpio_defaults_block_7/gpio_defaults[3]
+ gpio_defaults_block_7/gpio_defaults[4] gpio_defaults_block_7/gpio_defaults[5] gpio_defaults_block_7/gpio_defaults[6]
+ gpio_defaults_block_7/gpio_defaults[7] gpio_defaults_block_7/gpio_defaults[8] gpio_defaults_block_7/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[7] gpio_control_in_1a\[5\]/one housekeeping/mgmt_gpio_in[7]
+ gpio_control_in_1a\[5\]/one padframe/mprj_io_analog_en[7] padframe/mprj_io_analog_pol[7]
+ padframe/mprj_io_analog_sel[7] padframe/mprj_io_dm[21] padframe/mprj_io_dm[22] padframe/mprj_io_dm[23]
+ padframe/mprj_io_holdover[7] padframe/mprj_io_ib_mode_sel[7] padframe/mprj_io_in[7]
+ padframe/mprj_io_inp_dis[7] padframe/mprj_io_out[7] padframe/mprj_io_oeb[7] padframe/mprj_io_slow_sel[7]
+ padframe/mprj_io_vtrip_sel[7] gpio_control_in_1a\[5\]/resetn gpio_control_in_1\[0\]/resetn
+ gpio_control_in_1a\[5\]/serial_clock gpio_control_in_1\[0\]/serial_clock gpio_control_in_1a\[5\]/serial_data_in
+ gpio_control_in_1\[0\]/serial_data_in gpio_control_in_1a\[5\]/serial_load gpio_control_in_1\[0\]/serial_load
+ mprj/io_in[7] mprj/io_oeb[7] mprj/io_out[7] vccd_core vccd1_core VSUBS vssd1_core
+ gpio_control_in_1a\[5\]/zero gpio_control_block
Xgpio_defaults_block_32 VSUBS vccd_core gpio_defaults_block_32/gpio_defaults[0] gpio_defaults_block_32/gpio_defaults[10]
+ gpio_defaults_block_32/gpio_defaults[11] gpio_defaults_block_32/gpio_defaults[12]
+ gpio_defaults_block_32/gpio_defaults[1] gpio_defaults_block_32/gpio_defaults[2]
+ gpio_defaults_block_32/gpio_defaults[3] gpio_defaults_block_32/gpio_defaults[4]
+ gpio_defaults_block_32/gpio_defaults[5] gpio_defaults_block_32/gpio_defaults[6]
+ gpio_defaults_block_32/gpio_defaults[7] gpio_defaults_block_32/gpio_defaults[8]
+ gpio_defaults_block_32/gpio_defaults[9] gpio_defaults_block
Xgpio_control_bidir_2\[2\] gpio_defaults_block_37/gpio_defaults[0] gpio_defaults_block_37/gpio_defaults[10]
+ gpio_defaults_block_37/gpio_defaults[11] gpio_defaults_block_37/gpio_defaults[12]
+ gpio_defaults_block_37/gpio_defaults[1] gpio_defaults_block_37/gpio_defaults[2]
+ gpio_defaults_block_37/gpio_defaults[3] gpio_defaults_block_37/gpio_defaults[4]
+ gpio_defaults_block_37/gpio_defaults[5] gpio_defaults_block_37/gpio_defaults[6]
+ gpio_defaults_block_37/gpio_defaults[7] gpio_defaults_block_37/gpio_defaults[8]
+ gpio_defaults_block_37/gpio_defaults[9] housekeeping/mgmt_gpio_in[37] housekeeping/mgmt_gpio_oeb[37]
+ housekeeping/mgmt_gpio_out[37] gpio_control_bidir_2\[2\]/one padframe/mprj_io_analog_en[26]
+ padframe/mprj_io_analog_pol[26] padframe/mprj_io_analog_sel[26] padframe/mprj_io_dm[78]
+ padframe/mprj_io_dm[79] padframe/mprj_io_dm[80] padframe/mprj_io_holdover[26] padframe/mprj_io_ib_mode_sel[26]
+ padframe/mprj_io_in[26] padframe/mprj_io_inp_dis[26] padframe/mprj_io_out[26] padframe/mprj_io_oeb[26]
+ padframe/mprj_io_slow_sel[26] padframe/mprj_io_vtrip_sel[26] housekeeping/serial_resetn
+ gpio_control_bidir_2\[1\]/resetn housekeeping/serial_clock gpio_control_bidir_2\[1\]/serial_clock
+ housekeeping/serial_data_2 gpio_control_bidir_2\[1\]/serial_data_in housekeeping/serial_load
+ gpio_control_bidir_2\[1\]/serial_load mprj/io_in[26] mprj/io_oeb[26] mprj/io_out[26]
+ vccd_core vccd1_core VSUBS vssd1_core gpio_control_bidir_2\[2\]/zero gpio_control_block
.ends

