* NGSPICE file created from caravel_clocking.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd1_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd1_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_4 abstract view
.subckt sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtn_1 abstract view
.subckt sky130_fd_sc_hd__dfrtn_1 CLK_N D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

.subckt caravel_clocking VGND VPWR core_clk ext_clk ext_clk_sel ext_reset pll_clk
+ pll_clk90 resetb resetb_sync sel2[0] sel2[1] sel2[2] sel[0] sel[1] sel[2] user_clk
X_294_ _302_/B VGND VGND VPWR VPWR _294_/Y sky130_fd_sc_hd__inv_2
Xrebuffer7 _431_/Q VGND VGND VPWR VPWR _314_/A2 sky130_fd_sc_hd__dlygate4sd1_1
X_363_ _445_/Q _444_/Q VGND VGND VPWR VPWR _363_/Y sky130_fd_sc_hd__xnor2_1
X_432_ _351_/Y _432_/D _343_/S VGND VGND VPWR VPWR _432_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_9_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_346_ _346_/A VGND VGND VPWR VPWR _410_/S sky130_fd_sc_hd__inv_2
XFILLER_12_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_415_ _411_/A1 _415_/D VGND VGND VPWR VPWR _415_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_277_ _454_/Q VGND VGND VPWR VPWR _279_/B sky130_fd_sc_hd__inv_2
XFILLER_5_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_329_ _325_/Y _328_/Y _286_/Y VGND VGND VPWR VPWR _443_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0_pll_clk clkbuf_0_pll_clk/X VGND VGND VPWR VPWR _411_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrebuffer8 _314_/A2 VGND VGND VPWR VPWR _381_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
X_293_ _449_/Q _448_/Q VGND VGND VPWR VPWR _293_/Y sky130_fd_sc_hd__nor2_1
X_362_ _444_/Q VGND VGND VPWR VPWR _362_/Y sky130_fd_sc_hd__clkinv_2
X_431_ _351_/Y _431_/D _343_/S VGND VGND VPWR VPWR _431_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_12_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_276_ _276_/A _276_/B _451_/Q VGND VGND VPWR VPWR _345_/A sky130_fd_sc_hd__nand3_1
X_345_ _345_/A VGND VGND VPWR VPWR _404_/S sky130_fd_sc_hd__inv_2
X_414_ _411_/A1 _430_/Q VGND VGND VPWR VPWR _414_/Q sky130_fd_sc_hd__dfxtp_1
X_259_ _266_/A VGND VGND VPWR VPWR _263_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_328_ _326_/Y _327_/X _279_/C VGND VGND VPWR VPWR _328_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_18_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput10 _393_/X VGND VGND VPWR VPWR core_clk sky130_fd_sc_hd__clkbuf_1
XTAP_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrebuffer9 _381_/A1 VGND VGND VPWR VPWR _382_/A1 sky130_fd_sc_hd__dlygate4sd1_1
X_292_ _405_/X _286_/Y _291_/Y VGND VGND VPWR VPWR _451_/D sky130_fd_sc_hd__a21bo_1
X_334__6 _453_/CLK VGND VGND VPWR VPWR _441_/CLK sky130_fd_sc_hd__inv_2
X_361_ _453_/Q _361_/B VGND VGND VPWR VPWR _361_/X sky130_fd_sc_hd__xor2_1
X_430_ _351_/Y _430_/D _343_/S VGND VGND VPWR VPWR _430_/Q sky130_fd_sc_hd__dfrtp_4
X_344_ _344_/A VGND VGND VPWR VPWR _420_/D sky130_fd_sc_hd__buf_1
X_413_ _455_/Q _413_/A1 _413_/S VGND VGND VPWR VPWR _413_/X sky130_fd_sc_hd__mux2_1
X_275_ _452_/Q VGND VGND VPWR VPWR _276_/B sky130_fd_sc_hd__inv_2
XFILLER_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_258_ _258_/A _258_/B VGND VGND VPWR VPWR _266_/A sky130_fd_sc_hd__nand2_1
X_327_ _416_/D _416_/Q VGND VGND VPWR VPWR _327_/X sky130_fd_sc_hd__and2_1
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput11 _375_/Y VGND VGND VPWR VPWR resetb_sync sky130_fd_sc_hd__buf_2
XFILLER_15_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_291_ _291_/A _451_/Q _316_/C VGND VGND VPWR VPWR _291_/Y sky130_fd_sc_hd__nand3_1
X_360_ _452_/Q _451_/Q VGND VGND VPWR VPWR _361_/B sky130_fd_sc_hd__nor2_1
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_343_ hold1/A _343_/A1 _343_/S VGND VGND VPWR VPWR _344_/A sky130_fd_sc_hd__mux2_2
X_412_ _412_/A0 _426_/Q _425_/D VGND VGND VPWR VPWR _412_/X sky130_fd_sc_hd__mux2_1
X_274_ _453_/Q VGND VGND VPWR VPWR _276_/A sky130_fd_sc_hd__inv_2
X_257_ _257_/A _257_/B _257_/C VGND VGND VPWR VPWR _459_/D sky130_fd_sc_hd__nand3_1
X_326_ _416_/D _416_/Q VGND VGND VPWR VPWR _326_/Y sky130_fd_sc_hd__nor2_1
XFILLER_18_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_309_ _309_/A _309_/B _406_/S VGND VGND VPWR VPWR _316_/A sky130_fd_sc_hd__nand3_1
XFILLER_6_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput12 _394_/X VGND VGND VPWR VPWR user_clk sky130_fd_sc_hd__clkbuf_1
XTAP_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_290_ _402_/X _286_/Y _289_/Y VGND VGND VPWR VPWR _452_/D sky130_fd_sc_hd__a21bo_1
XFILLER_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_0_pll_clk pll_clk VGND VGND VPWR VPWR clkbuf_0_pll_clk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_10_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_273_ _273_/A _273_/B VGND VGND VPWR VPWR _455_/D sky130_fd_sc_hd__nand2_1
XFILLER_5_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_411_ _439_/Q _411_/A1 _411_/S VGND VGND VPWR VPWR _411_/X sky130_fd_sc_hd__mux2_1
X_342_ _439_/Q _342_/B VGND VGND VPWR VPWR _439_/D sky130_fd_sc_hd__xnor2_1
XFILLER_2_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_256_ _253_/Y _258_/A _250_/B VGND VGND VPWR VPWR _257_/B sky130_fd_sc_hd__o21bai_1
XFILLER_13_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_325_ _325_/A _325_/B _414_/Q VGND VGND VPWR VPWR _325_/Y sky130_fd_sc_hd__nand3_1
XFILLER_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_239_ _461_/Q VGND VGND VPWR VPWR _240_/B sky130_fd_sc_hd__inv_2
X_308_ _442_/Q _441_/Q _440_/Q VGND VGND VPWR VPWR _406_/S sky130_fd_sc_hd__nor3b_2
XFILLER_19_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_272_ _346_/A _272_/B _272_/C VGND VGND VPWR VPWR _273_/B sky130_fd_sc_hd__nand3_1
X_410_ _438_/Q _373_/Y _410_/S VGND VGND VPWR VPWR _410_/X sky130_fd_sc_hd__mux2_1
X_341_ _430_/Q _364_/A _444_/Q VGND VGND VPWR VPWR _342_/B sky130_fd_sc_hd__nand3b_1
XFILLER_5_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_255_ _437_/Q _438_/Q _436_/Q _254_/Y VGND VGND VPWR VPWR _258_/A sky130_fd_sc_hd__o211ai_1
X_324_ _415_/Q _324_/B_N VGND VGND VPWR VPWR _325_/B sky130_fd_sc_hd__or2b_1
XFILLER_9_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_238_ _462_/Q VGND VGND VPWR VPWR _240_/A sky130_fd_sc_hd__inv_2
X_307_ _447_/Q VGND VGND VPWR VPWR _309_/B sky130_fd_sc_hd__inv_2
XFILLER_19_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_271_ _346_/A _272_/B _272_/C VGND VGND VPWR VPWR _273_/A sky130_fd_sc_hd__a21o_1
X_340_ _446_/Q _445_/Q VGND VGND VPWR VPWR _364_/A sky130_fd_sc_hd__nor2_1
X_469_ _413_/A1 _469_/D _343_/S VGND VGND VPWR VPWR _469_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_14_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_254_ _462_/Q _461_/Q VGND VGND VPWR VPWR _254_/Y sky130_fd_sc_hd__nor2_1
X_323_ _415_/D _415_/Q VGND VGND VPWR VPWR _325_/A sky130_fd_sc_hd__or2b_1
XFILLER_2_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_237_ _460_/Q _258_/B _390_/X VGND VGND VPWR VPWR _237_/Y sky130_fd_sc_hd__nand3b_1
X_306_ _306_/A _306_/B VGND VGND VPWR VPWR _397_/S sky130_fd_sc_hd__nor2_2
XFILLER_16_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_270_ _455_/Q VGND VGND VPWR VPWR _272_/C sky130_fd_sc_hd__inv_2
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_468_ _413_/A1 _468_/D _343_/S VGND VGND VPWR VPWR _468_/Q sky130_fd_sc_hd__dfstp_1
X_399_ _398_/X _416_/D _443_/Q VGND VGND VPWR VPWR _399_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_322_ _322_/A VGND VGND VPWR VPWR _444_/D sky130_fd_sc_hd__clkbuf_1
X_253_ _253_/A _253_/B _456_/Q VGND VGND VPWR VPWR _253_/Y sky130_fd_sc_hd__nand3_1
XFILLER_13_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_236_ _467_/Q _234_/Y _235_/Y VGND VGND VPWR VPWR _236_/Y sky130_fd_sc_hd__o21bai_1
Xclkbuf_1_1_0_pll_clk90 clkbuf_0_pll_clk90/X VGND VGND VPWR VPWR _413_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_1_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_219_ _465_/Q VGND VGND VPWR VPWR _221_/A sky130_fd_sc_hd__inv_2
XFILLER_18_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_467_ _413_/A1 _467_/D _343_/S VGND VGND VPWR VPWR _467_/Q sky130_fd_sc_hd__dfrtp_4
X_398_ _361_/X _432_/Q _404_/S VGND VGND VPWR VPWR _398_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_252_ _457_/Q VGND VGND VPWR VPWR _253_/B sky130_fd_sc_hd__inv_2
X_321_ _400_/X _444_/Q _430_/Q VGND VGND VPWR VPWR _322_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0_0_pll_clk90 clkbuf_0_pll_clk90/X VGND VGND VPWR VPWR _465_/CLK sky130_fd_sc_hd__clkbuf_2
X_235_ _243_/B VGND VGND VPWR VPWR _235_/Y sky130_fd_sc_hd__inv_2
X_304_ _294_/Y _448_/Q _296_/Y VGND VGND VPWR VPWR _448_/D sky130_fd_sc_hd__a21bo_1
XFILLER_1_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_242__1 _465_/CLK VGND VGND VPWR VPWR _461_/CLK sky130_fd_sc_hd__inv_2
XFILLER_10_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_218_ _210_/Y _214_/Y _217_/Y VGND VGND VPWR VPWR _467_/D sky130_fd_sc_hd__o21a_1
Xclkbuf_1_1_0_ext_clk clkbuf_0_ext_clk/X VGND VGND VPWR VPWR _412_/A0 sky130_fd_sc_hd__clkbuf_2
XTAP_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_0_pll_clk clkbuf_0_pll_clk/X VGND VGND VPWR VPWR _453_/CLK sky130_fd_sc_hd__clkbuf_2
X_466_ _413_/A1 _466_/D _343_/S VGND VGND VPWR VPWR _466_/Q sky130_fd_sc_hd__dfstp_1
X_397_ _286_/Y _443_/Q _397_/S VGND VGND VPWR VPWR _397_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_251_ _458_/Q VGND VGND VPWR VPWR _253_/A sky130_fd_sc_hd__inv_2
X_320_ _320_/A VGND VGND VPWR VPWR _445_/D sky130_fd_sc_hd__clkbuf_1
X_449_ _449_/CLK _449_/D _343_/S VGND VGND VPWR VPWR _449_/Q sky130_fd_sc_hd__dfstp_1
X_234_ _461_/Q _460_/Q VGND VGND VPWR VPWR _234_/Y sky130_fd_sc_hd__nor2_1
XFILLER_1_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_303_ _299_/B _302_/X _295_/Y VGND VGND VPWR VPWR _449_/D sky130_fd_sc_hd__o21ai_1
XFILLER_19_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_217_ _247_/A _258_/B VGND VGND VPWR VPWR _217_/Y sky130_fd_sc_hd__nand2_2
XFILLER_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_396_ _395_/X _438_/Q _467_/Q VGND VGND VPWR VPWR _396_/X sky130_fd_sc_hd__mux2_1
X_465_ _465_/CLK _465_/D _343_/S VGND VGND VPWR VPWR _465_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_4_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_250_ _250_/A _250_/B _408_/S VGND VGND VPWR VPWR _257_/A sky130_fd_sc_hd__nand3_1
XFILLER_13_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_305__5 _453_/CLK VGND VGND VPWR VPWR _447_/CLK sky130_fd_sc_hd__inv_2
X_379_ _368_/Y _436_/Q _391_/S VGND VGND VPWR VPWR _379_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_448_ _453_/CLK _448_/D _343_/S VGND VGND VPWR VPWR _448_/Q sky130_fd_sc_hd__dfrtn_1
X_233_ _380_/X _217_/Y _232_/Y VGND VGND VPWR VPWR _463_/D sky130_fd_sc_hd__a21bo_1
X_302_ _448_/Q _302_/B VGND VGND VPWR VPWR _302_/X sky130_fd_sc_hd__and2b_1
XFILLER_6_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_216_ _467_/Q VGND VGND VPWR VPWR _258_/B sky130_fd_sc_hd__inv_2
XFILLER_15_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_464_ _465_/CLK _464_/D _343_/S VGND VGND VPWR VPWR _464_/Q sky130_fd_sc_hd__dfstp_1
X_395_ _367_/X _438_/Q _408_/S VGND VGND VPWR VPWR _395_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_447_ _447_/CLK _447_/D _343_/S VGND VGND VPWR VPWR _447_/Q sky130_fd_sc_hd__dfstp_1
X_232_ _232_/A _257_/C _463_/Q VGND VGND VPWR VPWR _232_/Y sky130_fd_sc_hd__nand3_1
XFILLER_19_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_215_ _437_/Q _438_/Q _436_/Q VGND VGND VPWR VPWR _247_/A sky130_fd_sc_hd__o21ai_2
XFILLER_15_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_394_ _412_/X _354_/Y _425_/Q VGND VGND VPWR VPWR _394_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_463_ _413_/A1 _463_/D _343_/S VGND VGND VPWR VPWR _463_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_13_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_446_ _411_/A1 _446_/D _343_/S VGND VGND VPWR VPWR _446_/Q sky130_fd_sc_hd__dfrtp_1
X_377_ _470_/Q _377_/B VGND VGND VPWR VPWR _470_/D sky130_fd_sc_hd__xor2_1
Xclkbuf_0_ext_clk ext_clk VGND VGND VPWR VPWR clkbuf_0_ext_clk/X sky130_fd_sc_hd__clkbuf_16
X_231_ _392_/X _217_/Y _230_/Y VGND VGND VPWR VPWR _464_/D sky130_fd_sc_hd__a21bo_1
X_300_ _450_/Q _295_/Y _296_/Y _306_/B VGND VGND VPWR VPWR _450_/D sky130_fd_sc_hd__o2bb2ai_1
XFILLER_1_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_429_ _351_/Y _429_/D _343_/S VGND VGND VPWR VPWR _432_/D sky130_fd_sc_hd__dfrtp_1
XFILLER_19_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput1 ext_clk_sel VGND VGND VPWR VPWR _374_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_18_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_214_ _211_/Y _212_/X _223_/C VGND VGND VPWR VPWR _214_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_15_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_393_ _412_/X _351_/Y _425_/Q VGND VGND VPWR VPWR _393_/X sky130_fd_sc_hd__mux2_1
X_462_ _465_/CLK _462_/D _343_/S VGND VGND VPWR VPWR _462_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_4_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_376_ _469_/Q _436_/Q _468_/Q VGND VGND VPWR VPWR _377_/B sky130_fd_sc_hd__nor3_1
X_445_ _411_/A1 _445_/D _343_/S VGND VGND VPWR VPWR _445_/Q sky130_fd_sc_hd__dfrtp_1
X_230_ _232_/A _257_/C _464_/Q VGND VGND VPWR VPWR _230_/Y sky130_fd_sc_hd__nand3_1
X_359_ _452_/Q _451_/Q VGND VGND VPWR VPWR _359_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_1_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_428_ _351_/Y _428_/D _343_/S VGND VGND VPWR VPWR _431_/D sky130_fd_sc_hd__dfstp_1
Xinput2 ext_reset VGND VGND VPWR VPWR _375_/A sky130_fd_sc_hd__clkbuf_1
XTAP_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_213_ _437_/Q _438_/Q _436_/Q VGND VGND VPWR VPWR _223_/C sky130_fd_sc_hd__o21a_1
XFILLER_15_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_392_ _391_/X _418_/D _467_/Q VGND VGND VPWR VPWR _392_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_461_ _461_/CLK _461_/D _343_/S VGND VGND VPWR VPWR _461_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_1_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_375_ _375_/A _421_/Q VGND VGND VPWR VPWR _375_/Y sky130_fd_sc_hd__nor2_1
X_444_ _453_/CLK _444_/D _343_/S VGND VGND VPWR VPWR _444_/Q sky130_fd_sc_hd__dfstp_2
X_358_ _451_/Q VGND VGND VPWR VPWR _358_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_427_ _351_/Y _427_/D _343_/S VGND VGND VPWR VPWR _430_/D sky130_fd_sc_hd__dfrtp_1
Xinput3 resetb VGND VGND VPWR VPWR _343_/S sky130_fd_sc_hd__buf_12
XTAP_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_289_ _291_/A _452_/Q _316_/C VGND VGND VPWR VPWR _289_/Y sky130_fd_sc_hd__nand3_1
XTAP_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_212_ _419_/Q _438_/Q VGND VGND VPWR VPWR _212_/X sky130_fd_sc_hd__and2_1
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_391_ _369_/Y _418_/D _391_/S VGND VGND VPWR VPWR _391_/X sky130_fd_sc_hd__mux2_1
X_460_ _465_/CLK _460_/D _343_/S VGND VGND VPWR VPWR _460_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_4_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_443_ _411_/A1 _443_/D _343_/S VGND VGND VPWR VPWR _443_/Q sky130_fd_sc_hd__dfrtp_4
X_374_ _374_/A VGND VGND VPWR VPWR _424_/D sky130_fd_sc_hd__inv_2
XFILLER_0_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_426_ _411_/A1 hold1/X _343_/S VGND VGND VPWR VPWR _426_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput4 sel2[0] VGND VGND VPWR VPWR _433_/D sky130_fd_sc_hd__clkbuf_1
XTAP_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_288_ _399_/X _286_/Y _287_/Y VGND VGND VPWR VPWR _453_/D sky130_fd_sc_hd__a21bo_1
X_357_ _442_/Q _357_/B VGND VGND VPWR VPWR _357_/X sky130_fd_sc_hd__xor2_1
XTAP_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_211_ _419_/Q _438_/Q VGND VGND VPWR VPWR _211_/Y sky130_fd_sc_hd__nor2_1
X_409_ _408_/X _437_/Q _467_/Q VGND VGND VPWR VPWR _409_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_390_ _217_/Y _467_/Q _390_/S VGND VGND VPWR VPWR _390_/X sky130_fd_sc_hd__mux2_4
XFILLER_8_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_373_ _469_/Q _468_/Q VGND VGND VPWR VPWR _373_/Y sky130_fd_sc_hd__xnor2_1
X_442_ _453_/CLK _442_/D _343_/S VGND VGND VPWR VPWR _442_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_1_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_425_ _411_/A1 _425_/D _343_/S VGND VGND VPWR VPWR _425_/Q sky130_fd_sc_hd__dfrtp_1
Xinput5 sel2[1] VGND VGND VPWR VPWR _434_/D sky130_fd_sc_hd__clkbuf_1
X_356_ _441_/Q _440_/Q VGND VGND VPWR VPWR _357_/B sky130_fd_sc_hd__nor2_1
X_287_ _291_/A _453_/Q _316_/C VGND VGND VPWR VPWR _287_/Y sky130_fd_sc_hd__nand3_1
XTAP_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_408_ _365_/Y _437_/Q _408_/S VGND VGND VPWR VPWR _408_/X sky130_fd_sc_hd__mux2_1
X_210_ _210_/A _210_/B _417_/Q VGND VGND VPWR VPWR _210_/Y sky130_fd_sc_hd__nand3_1
X_339_ _337_/Y _335_/A _338_/Y VGND VGND VPWR VPWR _440_/D sky130_fd_sc_hd__o21ai_1
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_372_ _468_/Q VGND VGND VPWR VPWR _372_/Y sky130_fd_sc_hd__clkinv_2
X_441_ _441_/CLK _441_/D _343_/S VGND VGND VPWR VPWR _441_/Q sky130_fd_sc_hd__dfstp_1
Xclkbuf_1_0_0_ext_clk clkbuf_0_ext_clk/X VGND VGND VPWR VPWR _343_/A1 sky130_fd_sc_hd__clkbuf_2
X_355_ _441_/Q _440_/Q VGND VGND VPWR VPWR _355_/Y sky130_fd_sc_hd__xnor2_1
X_286_ _306_/A _330_/B VGND VGND VPWR VPWR _286_/Y sky130_fd_sc_hd__nand2_2
X_424_ _411_/A1 _424_/D _343_/S VGND VGND VPWR VPWR _425_/D sky130_fd_sc_hd__dfrtp_1
Xinput6 sel2[2] VGND VGND VPWR VPWR _435_/D sky130_fd_sc_hd__clkbuf_1
XTAP_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_269_ _436_/Q VGND VGND VPWR VPWR _272_/B sky130_fd_sc_hd__inv_2
XFILLER_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_407_ _406_/X _432_/Q _443_/Q VGND VGND VPWR VPWR _407_/X sky130_fd_sc_hd__mux2_1
X_338_ _338_/A _386_/X VGND VGND VPWR VPWR _338_/Y sky130_fd_sc_hd__nand2_1
XFILLER_15_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_440_ _453_/CLK _440_/D _343_/S VGND VGND VPWR VPWR _440_/Q sky130_fd_sc_hd__dfrtn_1
X_371_ _465_/Q _371_/B VGND VGND VPWR VPWR _371_/X sky130_fd_sc_hd__xor2_1
X_423_ _393_/X _423_/D _343_/S VGND VGND VPWR VPWR _423_/Q sky130_fd_sc_hd__dfstp_1
X_354_ _272_/B _413_/X _232_/A _353_/Y VGND VGND VPWR VPWR _354_/Y sky130_fd_sc_hd__o2bb2ai_2
XFILLER_14_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_285_ _285_/A _316_/C _285_/C VGND VGND VPWR VPWR _454_/D sky130_fd_sc_hd__nand3_1
XTAP_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput7 sel[0] VGND VGND VPWR VPWR _427_/D sky130_fd_sc_hd__clkbuf_1
XTAP_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_268_ _469_/Q _470_/Q _468_/Q VGND VGND VPWR VPWR _346_/A sky130_fd_sc_hd__nor3b_1
X_337_ _440_/Q VGND VGND VPWR VPWR _337_/Y sky130_fd_sc_hd__inv_2
X_406_ _357_/X _432_/Q _406_/S VGND VGND VPWR VPWR _406_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_370_ _464_/Q _463_/Q VGND VGND VPWR VPWR _371_/B sky130_fd_sc_hd__nor2_1
X_422_ _393_/X _423_/Q _343_/S VGND VGND VPWR VPWR _422_/Q sky130_fd_sc_hd__dfstp_1
X_353_ _466_/Q _459_/Q VGND VGND VPWR VPWR _353_/Y sky130_fd_sc_hd__xnor2_1
X_284_ _291_/A _345_/A _279_/B VGND VGND VPWR VPWR _285_/C sky130_fd_sc_hd__o21bai_1
XFILLER_6_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput8 sel[1] VGND VGND VPWR VPWR _428_/D sky130_fd_sc_hd__clkbuf_1
XTAP_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_267_ _265_/Y _263_/A _266_/Y VGND VGND VPWR VPWR _456_/D sky130_fd_sc_hd__o21ai_1
X_405_ _404_/X _430_/Q _443_/Q VGND VGND VPWR VPWR _405_/X sky130_fd_sc_hd__mux2_1
X_336_ _312_/B _335_/A _335_/Y VGND VGND VPWR VPWR _441_/D sky130_fd_sc_hd__o21ai_1
XFILLER_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_319_ _403_/X _445_/Q _430_/Q VGND VGND VPWR VPWR _320_/A sky130_fd_sc_hd__mux2_1
XFILLER_11_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_421_ _393_/X _422_/Q _343_/S VGND VGND VPWR VPWR _421_/Q sky130_fd_sc_hd__dfstp_1
X_352_ _418_/D _438_/Q VGND VGND VPWR VPWR _413_/S sky130_fd_sc_hd__nor2_1
XTAP_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput9 sel[2] VGND VGND VPWR VPWR _429_/D sky130_fd_sc_hd__clkbuf_1
XTAP_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_283_ _306_/A VGND VGND VPWR VPWR _291_/A sky130_fd_sc_hd__clkbuf_2
XTAP_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_266_ _266_/A _384_/X VGND VGND VPWR VPWR _266_/Y sky130_fd_sc_hd__nand2_1
X_335_ _335_/A _382_/X VGND VGND VPWR VPWR _335_/Y sky130_fd_sc_hd__nand2_1
X_404_ _358_/Y _430_/Q _404_/S VGND VGND VPWR VPWR _404_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_249_ _458_/Q _457_/Q _456_/Q VGND VGND VPWR VPWR _408_/S sky130_fd_sc_hd__nor3b_2
X_318_ _446_/Q _318_/B VGND VGND VPWR VPWR _446_/D sky130_fd_sc_hd__xor2_1
XFILLER_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1 hold1/A VGND VGND VPWR VPWR hold1/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_378__13 VGND VGND VPWR VPWR _378__13/HI _423_/D sky130_fd_sc_hd__conb_1
XFILLER_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_420_ _453_/CLK _420_/D VGND VGND VPWR VPWR hold1/A sky130_fd_sc_hd__dfxtp_1
X_351_ _291_/A _349_/Y _350_/X VGND VGND VPWR VPWR _351_/Y sky130_fd_sc_hd__o21bai_2
XFILLER_5_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_282_ _432_/Q _431_/Q _430_/Q VGND VGND VPWR VPWR _306_/A sky130_fd_sc_hd__o21ai_2
XTAP_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_403_ _432_/Q _363_/Y _403_/S VGND VGND VPWR VPWR _403_/X sky130_fd_sc_hd__mux2_1
X_265_ _456_/Q VGND VGND VPWR VPWR _265_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_248_ _459_/Q VGND VGND VPWR VPWR _250_/B sky130_fd_sc_hd__inv_2
XFILLER_11_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_317_ _430_/Q _445_/Q _444_/Q VGND VGND VPWR VPWR _318_/B sky130_fd_sc_hd__nor3_1
XFILLER_19_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_246__2 _465_/CLK VGND VGND VPWR VPWR _459_/CLK sky130_fd_sc_hd__inv_2
XFILLER_5_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_281_ _330_/B VGND VGND VPWR VPWR _316_/C sky130_fd_sc_hd__clkbuf_2
X_350_ _430_/Q _411_/X VGND VGND VPWR VPWR _350_/X sky130_fd_sc_hd__and2b_2
XTAP_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_264_ _253_/B _263_/A _263_/Y VGND VGND VPWR VPWR _457_/D sky130_fd_sc_hd__o21ai_1
XFILLER_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_333_ _312_/A _335_/A _332_/Y VGND VGND VPWR VPWR _442_/D sky130_fd_sc_hd__o21ai_1
X_402_ _401_/X _415_/D _443_/Q VGND VGND VPWR VPWR _402_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_247_ _247_/A _247_/B VGND VGND VPWR VPWR _390_/S sky130_fd_sc_hd__nor2_1
X_316_ _316_/A _316_/B _316_/C VGND VGND VPWR VPWR _447_/D sky130_fd_sc_hd__nand3_1
XFILLER_6_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_280_ _443_/Q VGND VGND VPWR VPWR _330_/B sky130_fd_sc_hd__inv_2
XTAP_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_263_ _263_/A _409_/X VGND VGND VPWR VPWR _263_/Y sky130_fd_sc_hd__nand2_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_332_ _335_/A _407_/X VGND VGND VPWR VPWR _332_/Y sky130_fd_sc_hd__nand2_1
XFILLER_2_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_401_ _359_/Y _415_/D _404_/S VGND VGND VPWR VPWR _401_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_315_ _312_/Y _330_/A _309_/B VGND VGND VPWR VPWR _316_/B sky130_fd_sc_hd__o21bai_1
X_229_ _389_/X _217_/Y _228_/Y VGND VGND VPWR VPWR _465_/D sky130_fd_sc_hd__a21bo_1
XFILLER_17_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_262__3 _465_/CLK VGND VGND VPWR VPWR _457_/CLK sky130_fd_sc_hd__inv_2
XFILLER_14_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_331_ _338_/A VGND VGND VPWR VPWR _335_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_400_ _415_/D _362_/Y _403_/S VGND VGND VPWR VPWR _400_/X sky130_fd_sc_hd__mux2_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_245_ _235_/Y _460_/Q _237_/Y VGND VGND VPWR VPWR _460_/D sky130_fd_sc_hd__a21bo_1
X_314_ _432_/Q _314_/A2 _430_/Q _313_/Y VGND VGND VPWR VPWR _330_/A sky130_fd_sc_hd__o211ai_1
XFILLER_9_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_228_ _232_/A _257_/C _465_/Q VGND VGND VPWR VPWR _228_/Y sky130_fd_sc_hd__nand3_1
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_261_ _253_/A _263_/A _260_/Y VGND VGND VPWR VPWR _458_/D sky130_fd_sc_hd__o21ai_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_330_ _330_/A _330_/B VGND VGND VPWR VPWR _338_/A sky130_fd_sc_hd__nand2_1
XFILLER_17_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_459_ _459_/CLK _459_/D _343_/S VGND VGND VPWR VPWR _459_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_11_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_244_ _240_/B _243_/X _236_/Y VGND VGND VPWR VPWR _461_/D sky130_fd_sc_hd__o21ai_1
X_313_ _450_/Q _449_/Q VGND VGND VPWR VPWR _313_/Y sky130_fd_sc_hd__nor2_1
X_227_ _227_/A _257_/C _227_/C VGND VGND VPWR VPWR _466_/D sky130_fd_sc_hd__nand3_1
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_260_ _263_/A _396_/X VGND VGND VPWR VPWR _260_/Y sky130_fd_sc_hd__nand2_1
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_458_ _465_/CLK _458_/D _343_/S VGND VGND VPWR VPWR _458_/Q sky130_fd_sc_hd__dfrtn_1
X_389_ _388_/X _438_/Q _467_/Q VGND VGND VPWR VPWR _389_/X sky130_fd_sc_hd__mux2_1
X_243_ _460_/Q _243_/B VGND VGND VPWR VPWR _243_/X sky130_fd_sc_hd__and2b_1
X_312_ _312_/A _312_/B _440_/Q VGND VGND VPWR VPWR _312_/Y sky130_fd_sc_hd__nand3_1
XFILLER_7_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_226_ _232_/A _347_/A _223_/B VGND VGND VPWR VPWR _227_/C sky130_fd_sc_hd__o21bai_1
XFILLER_10_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_209_ _418_/D _418_/Q VGND VGND VPWR VPWR _210_/B sky130_fd_sc_hd__or2b_1
XFILLER_0_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xsplit12 _432_/Q VGND VGND VPWR VPWR _416_/D sky130_fd_sc_hd__clkbuf_2
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_457_ _457_/CLK _457_/D _343_/S VGND VGND VPWR VPWR _457_/Q sky130_fd_sc_hd__dfstp_1
X_388_ _371_/X _438_/Q _391_/S VGND VGND VPWR VPWR _388_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_311_ _441_/Q VGND VGND VPWR VPWR _312_/B sky130_fd_sc_hd__inv_2
X_225_ _247_/A VGND VGND VPWR VPWR _232_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_6_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_208_ _418_/Q _437_/Q VGND VGND VPWR VPWR _210_/A sky130_fd_sc_hd__or2b_1
XFILLER_0_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_456_ _465_/CLK _456_/D _343_/S VGND VGND VPWR VPWR _456_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_15_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_387_ _418_/D _372_/Y _410_/S VGND VGND VPWR VPWR _387_/X sky130_fd_sc_hd__mux2_1
X_310_ _442_/Q VGND VGND VPWR VPWR _312_/A sky130_fd_sc_hd__inv_2
X_241_ _462_/Q _236_/Y _237_/Y _247_/B VGND VGND VPWR VPWR _462_/D sky130_fd_sc_hd__o2bb2ai_1
X_439_ _411_/A1 _439_/D _343_/S VGND VGND VPWR VPWR _439_/Q sky130_fd_sc_hd__dfstp_1
X_224_ _258_/B VGND VGND VPWR VPWR _257_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_207_ _207_/A VGND VGND VPWR VPWR _468_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsplit1 _437_/Q VGND VGND VPWR VPWR _418_/D sky130_fd_sc_hd__buf_2
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer10 _390_/X VGND VGND VPWR VPWR _243_/B sky130_fd_sc_hd__clkbuf_1
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_455_ _413_/A1 _455_/D _343_/S VGND VGND VPWR VPWR _455_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_386_ _385_/X _430_/Q _443_/Q VGND VGND VPWR VPWR _386_/X sky130_fd_sc_hd__mux2_1
X_240_ _240_/A _240_/B VGND VGND VPWR VPWR _247_/B sky130_fd_sc_hd__nand2_1
X_438_ _354_/Y _438_/D _343_/S VGND VGND VPWR VPWR _438_/Q sky130_fd_sc_hd__dfrtp_4
X_369_ _464_/Q _463_/Q VGND VGND VPWR VPWR _369_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_9_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_223_ _347_/A _223_/B _223_/C VGND VGND VPWR VPWR _227_/A sky130_fd_sc_hd__nand3b_1
XFILLER_10_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_206_ _387_/X _468_/Q _436_/Q VGND VGND VPWR VPWR _207_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsplit2 split2/A VGND VGND VPWR VPWR _415_/D sky130_fd_sc_hd__clkbuf_2
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer11 _397_/S VGND VGND VPWR VPWR _309_/A sky130_fd_sc_hd__dlygate4sd1_1
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_385_ _337_/Y _430_/Q _406_/S VGND VGND VPWR VPWR _385_/X sky130_fd_sc_hd__mux2_1
X_454_ _411_/A1 _454_/D _343_/S VGND VGND VPWR VPWR _454_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_437_ _354_/Y _437_/D _343_/S VGND VGND VPWR VPWR _437_/Q sky130_fd_sc_hd__dfstp_4
Xrebuffer2 _390_/S VGND VGND VPWR VPWR _250_/A sky130_fd_sc_hd__dlygate4sd1_1
X_368_ _463_/Q VGND VGND VPWR VPWR _368_/Y sky130_fd_sc_hd__clkinv_2
X_299_ _299_/A _299_/B VGND VGND VPWR VPWR _306_/B sky130_fd_sc_hd__nand2_1
X_222_ _466_/Q VGND VGND VPWR VPWR _223_/B sky130_fd_sc_hd__inv_2
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_205_ _205_/A VGND VGND VPWR VPWR _469_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0_pll_clk90 pll_clk90 VGND VGND VPWR VPWR clkbuf_0_pll_clk90/X sky130_fd_sc_hd__clkbuf_16
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_470_ _413_/A1 _470_/D _343_/S VGND VGND VPWR VPWR _470_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_384_ _383_/X _436_/Q _467_/Q VGND VGND VPWR VPWR _384_/X sky130_fd_sc_hd__mux2_1
X_453_ _453_/CLK _453_/D _343_/S VGND VGND VPWR VPWR _453_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_11_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_367_ _458_/Q _367_/B VGND VGND VPWR VPWR _367_/X sky130_fd_sc_hd__xor2_1
X_436_ _354_/Y _436_/D _343_/S VGND VGND VPWR VPWR _436_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_13_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrebuffer3 _397_/X VGND VGND VPWR VPWR _302_/B sky130_fd_sc_hd__buf_2
X_298_ _449_/Q VGND VGND VPWR VPWR _299_/B sky130_fd_sc_hd__inv_2
X_221_ _221_/A _221_/B _463_/Q VGND VGND VPWR VPWR _347_/A sky130_fd_sc_hd__nand3_1
X_419_ _413_/A1 _438_/Q VGND VGND VPWR VPWR _419_/Q sky130_fd_sc_hd__dfxtp_1
X_204_ _410_/X _469_/Q _436_/Q VGND VGND VPWR VPWR _205_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_301__4 _453_/CLK VGND VGND VPWR VPWR _449_/CLK sky130_fd_sc_hd__inv_2
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_383_ _265_/Y _436_/Q _408_/S VGND VGND VPWR VPWR _383_/X sky130_fd_sc_hd__mux2_1
X_452_ _453_/CLK _452_/D _343_/S VGND VGND VPWR VPWR _452_/Q sky130_fd_sc_hd__dfstp_1
X_366_ _457_/Q _456_/Q VGND VGND VPWR VPWR _367_/B sky130_fd_sc_hd__nor2_1
X_435_ _354_/Y _435_/D _343_/S VGND VGND VPWR VPWR _438_/D sky130_fd_sc_hd__dfrtp_1
Xrebuffer4 _431_/Q VGND VGND VPWR VPWR split2/A sky130_fd_sc_hd__dlygate4sd1_1
X_297_ _450_/Q VGND VGND VPWR VPWR _299_/A sky130_fd_sc_hd__inv_2
XFILLER_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_220_ _464_/Q VGND VGND VPWR VPWR _221_/B sky130_fd_sc_hd__inv_2
XFILLER_10_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_418_ _465_/CLK _418_/D VGND VGND VPWR VPWR _418_/Q sky130_fd_sc_hd__dfxtp_1
X_349_ _454_/Q _447_/Q VGND VGND VPWR VPWR _349_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_18_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_451_ _411_/A1 _451_/D _343_/S VGND VGND VPWR VPWR _451_/Q sky130_fd_sc_hd__dfrtp_2
X_382_ _381_/X _382_/A1 _443_/Q VGND VGND VPWR VPWR _382_/X sky130_fd_sc_hd__mux2_1
X_365_ _457_/Q _456_/Q VGND VGND VPWR VPWR _365_/Y sky130_fd_sc_hd__xnor2_1
X_434_ _354_/Y _434_/D _343_/S VGND VGND VPWR VPWR _437_/D sky130_fd_sc_hd__dfstp_1
X_296_ _448_/Q _330_/B _397_/X VGND VGND VPWR VPWR _296_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer5 split2/A VGND VGND VPWR VPWR _324_/B_N sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_12_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_417_ _413_/A1 _436_/Q VGND VGND VPWR VPWR _417_/Q sky130_fd_sc_hd__dfxtp_1
X_279_ _345_/A _279_/B _279_/C VGND VGND VPWR VPWR _285_/A sky130_fd_sc_hd__nand3b_1
X_348_ _416_/D _415_/D VGND VGND VPWR VPWR _411_/S sky130_fd_sc_hd__nor2_1
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_381_ _355_/Y _381_/A1 _406_/S VGND VGND VPWR VPWR _381_/X sky130_fd_sc_hd__mux2_1
X_450_ _453_/CLK _450_/D _343_/S VGND VGND VPWR VPWR _450_/Q sky130_fd_sc_hd__dfrtn_1
XTAP_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_433_ _354_/Y _433_/D _343_/S VGND VGND VPWR VPWR _436_/D sky130_fd_sc_hd__dfrtp_1
XFILLER_13_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_295_ _443_/Q _293_/Y _294_/Y VGND VGND VPWR VPWR _295_/Y sky130_fd_sc_hd__o21bai_1
X_364_ _364_/A _444_/Q VGND VGND VPWR VPWR _403_/S sky130_fd_sc_hd__nand2_1
Xrebuffer6 _431_/Q VGND VGND VPWR VPWR _278_/A2 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_9_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_347_ _347_/A VGND VGND VPWR VPWR _391_/S sky130_fd_sc_hd__inv_2
XFILLER_12_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_278_ _416_/D _278_/A2 _430_/Q VGND VGND VPWR VPWR _279_/C sky130_fd_sc_hd__o21a_1
X_416_ _411_/A1 _416_/D VGND VGND VPWR VPWR _416_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_380_ _379_/X _436_/Q _467_/Q VGND VGND VPWR VPWR _380_/X sky130_fd_sc_hd__mux2_1
XTAP_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

