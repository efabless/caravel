* NGSPICE file created from caravel_clocking.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_1 abstract view
.subckt sky130_fd_sc_hd__a41oi_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtn_1 abstract view
.subckt sky130_fd_sc_hd__dfrtn_1 CLK_N D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_1 abstract view
.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

.subckt caravel_clocking VGND VPWR core_clk ext_clk ext_clk_sel ext_reset pll_clk
+ pll_clk90 resetb resetb_sync sel2[0] sel2[1] sel2[2] sel[0] sel[1] sel[2] user_clk
XTAP_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_294_ _287_/Y _301_/B _292_/Y _251_/Y _227_/S VGND VGND VPWR VPWR _294_/Y sky130_fd_sc_hd__a41oi_1
X_363_ _301_/A _365_/B _429_/Q VGND VGND VPWR VPWR _363_/Y sky130_fd_sc_hd__nand3b_1
X_432_ _432_/CLK _432_/D _380_/S VGND VGND VPWR VPWR _432_/Q sky130_fd_sc_hd__dfstp_1
X_346_ _462_/Q _461_/Q _463_/Q VGND VGND VPWR VPWR _347_/B sky130_fd_sc_hd__o21ai_1
XFILLER_12_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_277_ _335_/A _450_/D _408_/A _259_/Y _247_/Y VGND VGND VPWR VPWR _393_/B sky130_fd_sc_hd__o2111ai_4
X_329_ _436_/Q _437_/Q _438_/Q VGND VGND VPWR VPWR _331_/A sky130_fd_sc_hd__or3_1
XFILLER_18_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__037_ clkbuf_0__037_/X VGND VGND VPWR VPWR _212_/A0 sky130_fd_sc_hd__clkbuf_16
XTAP_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__283__A1 _388_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_431_ _208_/A1 _431_/D fanout27/X VGND VGND VPWR VPWR _431_/Q sky130_fd_sc_hd__dfrtn_1
X_293_ _426_/D _425_/D _377_/A _287_/Y _292_/Y VGND VGND VPWR VPWR _293_/X sky130_fd_sc_hd__o2111a_1
X_362_ _428_/Q _301_/B _358_/Y _361_/Y VGND VGND VPWR VPWR _428_/D sky130_fd_sc_hd__o22a_1
XFILLER_10_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__468__RESET_B fanout29/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_276_ _335_/A _472_/Q _408_/A VGND VGND VPWR VPWR _388_/A sky130_fd_sc_hd__o21a_4
X_345_ _462_/Q _461_/Q _463_/Q VGND VGND VPWR VPWR _347_/A sky130_fd_sc_hd__or3_1
XANTENNA__238__A1 _335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_328_ _436_/Q _437_/Q VGND VGND VPWR VPWR _328_/Y sky130_fd_sc_hd__xnor2_1
X_259_ _460_/Q VGND VGND VPWR VPWR _259_/Y sky130_fd_sc_hd__clkinv_4
XANTENNA__408__A _408_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_292_ _430_/Q _431_/Q _429_/Q VGND VGND VPWR VPWR _292_/Y sky130_fd_sc_hd__nor3b_2
X_430_ _430_/CLK _430_/D _380_/S VGND VGND VPWR VPWR _430_/Q sky130_fd_sc_hd__dfstp_1
X_361_ _359_/Y _360_/X _301_/B VGND VGND VPWR VPWR _361_/Y sky130_fd_sc_hd__o21ai_1
X_275_ _335_/A _450_/D VGND VGND VPWR VPWR _275_/Y sky130_fd_sc_hd__nor2_1
X_344_ _462_/Q _461_/Q VGND VGND VPWR VPWR _344_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_5_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__401__A2 _388_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_258_ _465_/Q VGND VGND VPWR VPWR _258_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_9_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_327_ _327_/A _327_/B VGND VGND VPWR VPWR _327_/Y sky130_fd_sc_hd__nand2_1
XFILLER_18_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__277__B1 _408_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput11 _349_/Y VGND VGND VPWR VPWR resetb_sync sky130_fd_sc_hd__buf_12
XANTENNA__422__SET_B fanout28/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_291_ _365_/B VGND VGND VPWR VPWR _291_/Y sky130_fd_sc_hd__inv_2
X_360_ _426_/D _426_/Q VGND VGND VPWR VPWR _360_/X sky130_fd_sc_hd__and2_1
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_343_ _343_/A _343_/B VGND VGND VPWR VPWR _343_/Y sky130_fd_sc_hd__nand2_1
X_274_ _459_/Q _460_/Q VGND VGND VPWR VPWR _274_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_326_ _430_/Q _429_/Q _431_/Q VGND VGND VPWR VPWR _327_/B sky130_fd_sc_hd__o21ai_1
X_257_ _436_/Q VGND VGND VPWR VPWR _303_/C sky130_fd_sc_hd__clkinv_4
XFILLER_9_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_309_ _424_/D _309_/B VGND VGND VPWR VPWR _309_/X sky130_fd_sc_hd__and2b_2
XANTENNA__421__RESET_B fanout28/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_0_divider.out _312_/X VGND VGND VPWR VPWR clkbuf_0_divider.out/X sky130_fd_sc_hd__clkbuf_16
XANTENNA__277__A1 _335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input8_A sel[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_290_ _426_/D _425_/D _377_/A _255_/Y _250_/Y VGND VGND VPWR VPWR _365_/B sky130_fd_sc_hd__o2111ai_4
Xclkbuf_0_pll_clk pll_clk VGND VGND VPWR VPWR clkbuf_0_pll_clk/X sky130_fd_sc_hd__clkbuf_16
X_342_ _455_/Q _454_/Q _456_/Q VGND VGND VPWR VPWR _343_/B sky130_fd_sc_hd__o21ai_1
X_273_ _459_/Q _231_/X _396_/S VGND VGND VPWR VPWR _459_/D sky130_fd_sc_hd__mux2_1
XFILLER_4_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_325_ _430_/Q _429_/Q _431_/Q VGND VGND VPWR VPWR _327_/A sky130_fd_sc_hd__or3_1
X_256_ _429_/Q VGND VGND VPWR VPWR _256_/Y sky130_fd_sc_hd__clkinv_2
X_239_ _308_/C _449_/D _308_/Y VGND VGND VPWR VPWR _239_/X sky130_fd_sc_hd__mux2_1
X_308_ _462_/Q _463_/Q _308_/C VGND VGND VPWR VPWR _308_/Y sky130_fd_sc_hd__nor3_2
XANTENNA__461__RESET_B fanout28/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__277__A2 _450_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f_pll_clk90 clkbuf_0_pll_clk90/X VGND VGND VPWR VPWR _463_/CLK sky130_fd_sc_hd__clkbuf_16
X_272_ _272_/A VGND VGND VPWR VPWR _272_/Y sky130_fd_sc_hd__inv_2
X_341_ _455_/Q _454_/Q _456_/Q VGND VGND VPWR VPWR _343_/A sky130_fd_sc_hd__or3_1
X_410_ _410_/A _410_/B VGND VGND VPWR VPWR _467_/D sky130_fd_sc_hd__or2_1
XANTENNA__398__A1 _242_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_324_ _430_/Q _429_/Q VGND VGND VPWR VPWR _324_/Y sky130_fd_sc_hd__xnor2_1
X_255_ _435_/Q VGND VGND VPWR VPWR _255_/Y sky130_fd_sc_hd__clkinv_4
X_266__7 _411__8/A VGND VGND VPWR VPWR _417_/CLK sky130_fd_sc_hd__inv_4
XFILLER_1_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_238_ _237_/X _335_/A _306_/A VGND VGND VPWR VPWR _272_/A sky130_fd_sc_hd__mux2_1
X_307_ _462_/Q _463_/Q VGND VGND VPWR VPWR _307_/Y sky130_fd_sc_hd__nor2_1
XFILLER_1_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_340_ _455_/Q _454_/Q VGND VGND VPWR VPWR _340_/Y sky130_fd_sc_hd__xnor2_1
X_469_ _212_/A1 _469_/D fanout28/X VGND VGND VPWR VPWR _472_/D sky130_fd_sc_hd__dfstp_1
X_323_ _254_/Y _287_/Y _322_/X VGND VGND VPWR VPWR _323_/X sky130_fd_sc_hd__a21o_1
X_254_ _433_/Q VGND VGND VPWR VPWR _254_/Y sky130_fd_sc_hd__inv_2
X_237_ _343_/Y _335_/A _279_/Y VGND VGND VPWR VPWR _237_/X sky130_fd_sc_hd__mux2_1
X_306_ _306_/A _388_/A VGND VGND VPWR VPWR _306_/X sky130_fd_sc_hd__or2_1
XANTENNA__313__A_N _408_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__470__RESET_B fanout29/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input6_A sel2[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_270_ _270_/A VGND VGND VPWR VPWR _270_/Y sky130_fd_sc_hd__inv_2
X_468_ _473_/CLK _468_/D fanout29/X VGND VGND VPWR VPWR _471_/D sky130_fd_sc_hd__dfrtp_1
XANTENNA__398__A3 _388_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_399_ _242_/S _388_/A _242_/X VGND VGND VPWR VPWR _399_/Y sky130_fd_sc_hd__o21bai_1
XANTENNA__457__SET_B fanout28/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_322_ _434_/Q _433_/Q _435_/Q VGND VGND VPWR VPWR _322_/X sky130_fd_sc_hd__o21a_1
XFILLER_9_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f_net10 clkbuf_0_net10/X VGND VGND VPWR VPWR core_clk sky130_fd_sc_hd__clkbuf_16
X_253_ _439_/Q VGND VGND VPWR VPWR _253_/Y sky130_fd_sc_hd__clkinv_2
X_305_ _465_/Q _382_/C VGND VGND VPWR VPWR _305_/Y sky130_fd_sc_hd__nand2_1
X_236_ _235_/X _450_/D _242_/S VGND VGND VPWR VPWR _249_/A sky130_fd_sc_hd__mux2_1
XANTENNA_fanout27_A fanout29/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_219_ _218_/X _425_/D _301_/A VGND VGND VPWR VPWR _252_/A sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_0_pll_clk_A pll_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__240__S _242_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__417__SET_B fanout28/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_467_ _211_/A1 _467_/D fanout29/X VGND VGND VPWR VPWR _467_/Q sky130_fd_sc_hd__dfrtp_1
X_398_ _242_/S _308_/C _388_/A _397_/Y VGND VGND VPWR VPWR _461_/D sky130_fd_sc_hd__o31ai_1
X_252_ _252_/A VGND VGND VPWR VPWR _252_/Y sky130_fd_sc_hd__inv_2
X_321_ _321_/A _321_/B VGND VGND VPWR VPWR _321_/Y sky130_fd_sc_hd__nor2_1
X_235_ _340_/Y _450_/D _279_/Y VGND VGND VPWR VPWR _235_/X sky130_fd_sc_hd__mux2_1
X_304_ _466_/Q _467_/Q VGND VGND VPWR VPWR _382_/C sky130_fd_sc_hd__nor2_1
X_218_ _324_/Y _425_/D _292_/Y VGND VGND VPWR VPWR _218_/X sky130_fd_sc_hd__mux2_1
XTAP_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xuser_clk_out_buffer _212_/X VGND VGND VPWR VPWR user_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_8_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_397_ _242_/S _388_/A _240_/X VGND VGND VPWR VPWR _397_/Y sky130_fd_sc_hd__o21ai_1
X_466_ _211_/A1 _466_/D fanout28/X VGND VGND VPWR VPWR _466_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__316__A2 _388_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_251_ _432_/Q VGND VGND VPWR VPWR _251_/Y sky130_fd_sc_hd__clkinv_4
X_320_ _425_/D _377_/A _426_/D VGND VGND VPWR VPWR _321_/B sky130_fd_sc_hd__o21a_1
XANTENNA__243__A1 _335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__234__A1 _408_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_449_ _211_/A1 _449_/D VGND VGND VPWR VPWR _449_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f_divider.out clkbuf_0_divider.out/X VGND VGND VPWR VPWR _210_/A1 sky130_fd_sc_hd__clkbuf_16
X_234_ _233_/X _408_/A _242_/S VGND VGND VPWR VPWR _270_/A sky130_fd_sc_hd__mux2_1
X_303_ _437_/Q _438_/Q _303_/C VGND VGND VPWR VPWR _303_/Y sky130_fd_sc_hd__nor3_2
X_217_ _216_/X _377_/A _301_/A VGND VGND VPWR VPWR _267_/A sky130_fd_sc_hd__mux2_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_465_ _211_/A1 _465_/D fanout28/X VGND VGND VPWR VPWR _465_/Q sky130_fd_sc_hd__dfstp_2
X_396_ _460_/Q _232_/X _396_/S VGND VGND VPWR VPWR _460_/D sky130_fd_sc_hd__mux2_1
XANTENNA__473__RESET_B fanout29/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_250_ _434_/Q VGND VGND VPWR VPWR _250_/Y sky130_fd_sc_hd__clkinv_4
XANTENNA_input4_A sel2[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout20 _445_/Q VGND VGND VPWR VPWR _424_/D sky130_fd_sc_hd__clkbuf_2
X_448_ _448_/CLK _448_/D VGND VGND VPWR VPWR _448_/Q sky130_fd_sc_hd__dfxtp_1
X_379_ _379_/A _379_/B VGND VGND VPWR VPWR _441_/D sky130_fd_sc_hd__or2_1
X_233_ _261_/Y _408_/A _279_/Y VGND VGND VPWR VPWR _233_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_302_ _437_/Q _438_/Q VGND VGND VPWR VPWR _302_/Y sky130_fd_sc_hd__nor2_1
X_216_ _256_/Y _424_/D _292_/Y VGND VGND VPWR VPWR _216_/X sky130_fd_sc_hd__mux2_1
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__469__SET_B fanout28/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__246__A0 _335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_464_ _208_/A1 _464_/D fanout27/X VGND VGND VPWR VPWR _464_/Q sky130_fd_sc_hd__dfstp_1
X_395_ _458_/Q _230_/X _396_/S VGND VGND VPWR VPWR _458_/D sky130_fd_sc_hd__mux2_1
XANTENNA__452__SET_B fanout28/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout21 _242_/S VGND VGND VPWR VPWR _306_/A sky130_fd_sc_hd__clkbuf_4
X_378_ _377_/A _440_/Q _439_/Q _441_/Q VGND VGND VPWR VPWR _379_/B sky130_fd_sc_hd__o31a_1
X_447_ _447_/CLK _447_/D fanout27/X VGND VGND VPWR VPWR _447_/Q sky130_fd_sc_hd__dfrtp_1
X_232_ _339_/X _337_/B _306_/A VGND VGND VPWR VPWR _232_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_301_ _301_/A _301_/B VGND VGND VPWR VPWR _301_/X sky130_fd_sc_hd__or2_1
Xclkbuf_1_0__f__037_ clkbuf_0__037_/X VGND VGND VPWR VPWR _210_/A0 sky130_fd_sc_hd__clkbuf_16
XFILLER_1_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_215_ _323_/X _321_/B _301_/A VGND VGND VPWR VPWR _215_/X sky130_fd_sc_hd__mux2_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__467__RESET_B fanout29/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_394_ _272_/Y _283_/Y _393_/Y VGND VGND VPWR VPWR _456_/D sky130_fd_sc_hd__o21ai_1
X_463_ _463_/CLK _463_/D fanout28/X VGND VGND VPWR VPWR _463_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__237__A1 _335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout22 _453_/Q VGND VGND VPWR VPWR _242_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__400__A1 _242_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_1_1__f_pll_clk90 clkbuf_0_pll_clk90/X VGND VGND VPWR VPWR _211_/A1 sky130_fd_sc_hd__clkbuf_16
X_377_ _377_/A _440_/Q _439_/Q _441_/Q VGND VGND VPWR VPWR _379_/A sky130_fd_sc_hd__nor4_1
X_446_ _447_/CLK _446_/D fanout27/X VGND VGND VPWR VPWR _446_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_0_ext_clk ext_clk VGND VGND VPWR VPWR clkbuf_0_ext_clk/X sky130_fd_sc_hd__clkbuf_16
X_231_ _334_/Y _337_/Y _306_/A VGND VGND VPWR VPWR _231_/X sky130_fd_sc_hd__mux2_1
X_300_ _439_/Q _354_/C VGND VGND VPWR VPWR _300_/Y sky130_fd_sc_hd__nand2_1
X_429_ _448_/CLK _429_/D _380_/S VGND VGND VPWR VPWR _429_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_10_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput1 ext_clk_sel VGND VGND VPWR VPWR _263_/A sky130_fd_sc_hd__clkbuf_1
XTAP_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_214_ _318_/Y _321_/Y _301_/A VGND VGND VPWR VPWR _214_/X sky130_fd_sc_hd__mux2_1
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_414__6 _448_/CLK VGND VGND VPWR VPWR _434_/CLK sky130_fd_sc_hd__inv_4
XFILLER_7_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_462_ _463_/CLK _462_/D fanout26/X VGND VGND VPWR VPWR _462_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_4_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_393_ _306_/A _393_/B _456_/Q VGND VGND VPWR VPWR _393_/Y sky130_fd_sc_hd__nand3b_1
Xfanout23 _227_/S VGND VGND VPWR VPWR _301_/A sky130_fd_sc_hd__clkbuf_4
X_376_ _229_/X _440_/Q _377_/A VGND VGND VPWR VPWR _440_/D sky130_fd_sc_hd__mux2_1
X_445_ _447_/CLK _445_/D fanout27/X VGND VGND VPWR VPWR _445_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_input2_A ext_reset VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_230_ _260_/Y _333_/Y _306_/A VGND VGND VPWR VPWR _230_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_359_ _447_/Q _426_/Q VGND VGND VPWR VPWR _359_/Y sky130_fd_sc_hd__nor2_1
X_428_ _208_/A1 _428_/D fanout27/X VGND VGND VPWR VPWR _428_/Q sky130_fd_sc_hd__dfrtp_1
Xinput2 ext_reset VGND VGND VPWR VPWR _349_/A sky130_fd_sc_hd__clkbuf_1
XTAP_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_213_ _254_/Y _317_/Y _301_/A VGND VGND VPWR VPWR _213_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__276__B1 _408_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0_net10 _210_/X VGND VGND VPWR VPWR clkbuf_0_net10/X sky130_fd_sc_hd__clkbuf_16
X_392_ _270_/Y _283_/Y _391_/Y VGND VGND VPWR VPWR _454_/D sky130_fd_sc_hd__o21ai_1
X_461_ _211_/A1 _461_/D fanout28/X VGND VGND VPWR VPWR _461_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_4_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_411__8 _411__8/A VGND VGND VPWR VPWR _418_/CLK sky130_fd_sc_hd__inv_4
XFILLER_1_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout24 _428_/Q VGND VGND VPWR VPWR _227_/S sky130_fd_sc_hd__clkbuf_4
Xfanout13 _473_/Q VGND VGND VPWR VPWR _335_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__400__A3 _388_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_375_ _228_/X _439_/Q _377_/A VGND VGND VPWR VPWR _439_/D sky130_fd_sc_hd__mux2_1
X_444_ _210_/A1 _444_/D fanout27/X VGND VGND VPWR VPWR _447_/D sky130_fd_sc_hd__dfrtp_1
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_427_ _208_/A1 _427_/D fanout27/X VGND VGND VPWR VPWR _427_/Q sky130_fd_sc_hd__dfstp_1
X_358_ _358_/A _358_/B _424_/Q VGND VGND VPWR VPWR _358_/Y sky130_fd_sc_hd__nand3_1
Xinput3 resetb VGND VGND VPWR VPWR input3/X sky130_fd_sc_hd__clkbuf_1
XTAP_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_289_ _426_/D _446_/Q _424_/D VGND VGND VPWR VPWR _301_/B sky130_fd_sc_hd__o21a_4
XTAP_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_212_ _212_/A0 _212_/A1 _421_/Q VGND VGND VPWR VPWR _212_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__276__A1 _335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__335__A _335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_391_ _306_/A _393_/B _454_/Q VGND VGND VPWR VPWR _391_/Y sky130_fd_sc_hd__nand3b_1
X_460_ _463_/CLK _460_/D fanout26/X VGND VGND VPWR VPWR _460_/Q sky130_fd_sc_hd__dfrtn_1
Xfanout25 input3/X VGND VGND VPWR VPWR _380_/S sky130_fd_sc_hd__buf_4
XFILLER_13_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout14 _472_/Q VGND VGND VPWR VPWR _450_/D sky130_fd_sc_hd__clkbuf_4
X_443_ _447_/CLK _443_/D fanout27/X VGND VGND VPWR VPWR _446_/D sky130_fd_sc_hd__dfstp_1
X_374_ _227_/S _438_/Q _301_/B _373_/Y VGND VGND VPWR VPWR _438_/D sky130_fd_sc_hd__o31a_1
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput4 sel2[0] VGND VGND VPWR VPWR _468_/D sky130_fd_sc_hd__clkbuf_1
X_357_ _425_/D _425_/Q VGND VGND VPWR VPWR _358_/B sky130_fd_sc_hd__nand2b_1
XTAP_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_426_ _208_/A1 _426_/D VGND VGND VPWR VPWR _426_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_288_ _426_/D _446_/Q VGND VGND VPWR VPWR _288_/Y sky130_fd_sc_hd__nor2_1
X_211_ _452_/Q _211_/A1 _275_/Y VGND VGND VPWR VPWR _313_/B sky130_fd_sc_hd__mux2_1
X_409_ _408_/A _466_/Q _465_/Q _467_/Q VGND VGND VPWR VPWR _410_/B sky130_fd_sc_hd__o31a_1
XFILLER_2_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_390_ _242_/S _388_/A _388_/Y _389_/Y VGND VGND VPWR VPWR _453_/D sky130_fd_sc_hd__o22a_1
XANTENNA__335__B _450_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout26 input3/X VGND VGND VPWR VPWR fanout26/X sky130_fd_sc_hd__buf_2
XANTENNA__397__A1 _242_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout15 _471_/Q VGND VGND VPWR VPWR _408_/A sky130_fd_sc_hd__clkbuf_4
Xclkbuf_1_1__f_pll_clk clkbuf_0_pll_clk/X VGND VGND VPWR VPWR _208_/A1 sky130_fd_sc_hd__clkbuf_16
X_442_ _447_/CLK _442_/D fanout27/X VGND VGND VPWR VPWR _445_/D sky130_fd_sc_hd__dfrtp_1
X_373_ _227_/S _301_/B _227_/X VGND VGND VPWR VPWR _373_/Y sky130_fd_sc_hd__o21bai_1
Xinput5 sel2[1] VGND VGND VPWR VPWR _469_/D sky130_fd_sc_hd__clkbuf_1
X_425_ _208_/A1 _425_/D VGND VGND VPWR VPWR _425_/Q sky130_fd_sc_hd__dfxtp_1
X_287_ _434_/Q _435_/Q VGND VGND VPWR VPWR _287_/Y sky130_fd_sc_hd__nor2_1
X_356_ _425_/Q _425_/D VGND VGND VPWR VPWR _358_/A sky130_fd_sc_hd__nand2b_1
XTAP_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_210_ _210_/A0 _210_/A1 _421_/Q VGND VGND VPWR VPWR _210_/X sky130_fd_sc_hd__mux2_1
X_408_ _408_/A _466_/Q _465_/Q _467_/Q VGND VGND VPWR VPWR _410_/A sky130_fd_sc_hd__nor4_1
Xclkbuf_1_0__f_divider2.out clkbuf_0_divider2.out/X VGND VGND VPWR VPWR _212_/A1 sky130_fd_sc_hd__clkbuf_16
X_339_ _260_/Y _274_/Y _338_/X VGND VGND VPWR VPWR _339_/X sky130_fd_sc_hd__a21o_1
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__335__C _408_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout21_A _242_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout16 _471_/Q VGND VGND VPWR VPWR _449_/D sky130_fd_sc_hd__clkbuf_2
XANTENNA__397__A2 _388_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout27 fanout29/X VGND VGND VPWR VPWR fanout27/X sky130_fd_sc_hd__buf_4
X_441_ _448_/CLK _441_/D _380_/S VGND VGND VPWR VPWR _441_/Q sky130_fd_sc_hd__dfrtp_1
X_372_ _227_/S _437_/Q _301_/B _371_/Y VGND VGND VPWR VPWR _437_/D sky130_fd_sc_hd__o31a_1
X_355_ _355_/A _355_/B VGND VGND VPWR VPWR _427_/D sky130_fd_sc_hd__nand2_1
X_286_ _434_/Q _214_/X _368_/S VGND VGND VPWR VPWR _434_/D sky130_fd_sc_hd__mux2_1
X_424_ _208_/A1 _424_/D VGND VGND VPWR VPWR _424_/Q sky130_fd_sc_hd__dfxtp_1
Xinput6 sel2[2] VGND VGND VPWR VPWR _470_/D sky130_fd_sc_hd__clkbuf_1
XTAP_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_338_ _459_/Q _458_/Q _460_/Q VGND VGND VPWR VPWR _338_/X sky130_fd_sc_hd__o21a_1
X_269_ _269_/A VGND VGND VPWR VPWR _269_/Y sky130_fd_sc_hd__inv_2
X_407_ _246_/X _466_/Q _449_/D VGND VGND VPWR VPWR _466_/D sky130_fd_sc_hd__mux2_1
XANTENNA__351__B1 _242_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__275__A _335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_0__037_ _209_/X VGND VGND VPWR VPWR clkbuf_0__037_/X sky130_fd_sc_hd__clkbuf_16
Xfanout28 fanout29/X VGND VGND VPWR VPWR fanout28/X sky130_fd_sc_hd__buf_4
Xfanout17 _447_/Q VGND VGND VPWR VPWR _426_/D sky130_fd_sc_hd__clkbuf_4
X_371_ _227_/S _301_/B _225_/X VGND VGND VPWR VPWR _371_/Y sky130_fd_sc_hd__o21bai_1
X_440_ _448_/CLK _440_/D _380_/S VGND VGND VPWR VPWR _440_/Q sky130_fd_sc_hd__dfrtp_1
X_423_ _448_/CLK _448_/Q fanout26/X VGND VGND VPWR VPWR _423_/Q sky130_fd_sc_hd__dfrtp_1
X_285_ _249_/Y _283_/Y _284_/Y VGND VGND VPWR VPWR _455_/D sky130_fd_sc_hd__o21ai_1
X_354_ _377_/A _439_/Q _354_/C _354_/D VGND VGND VPWR VPWR _355_/B sky130_fd_sc_hd__nand4b_1
XTAP_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput7 sel[0] VGND VGND VPWR VPWR _442_/D sky130_fd_sc_hd__clkbuf_1
XTAP_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_406_ _245_/X _465_/Q _449_/D VGND VGND VPWR VPWR _465_/D sky130_fd_sc_hd__mux2_1
XFILLER_2_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_337_ _337_/A _337_/B VGND VGND VPWR VPWR _337_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_0_pll_clk90_A pll_clk90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__463__RESET_B fanout28/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__275__B _450_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_1_0__f_divider.out clkbuf_0_divider.out/X VGND VGND VPWR VPWR _447_/CLK sky130_fd_sc_hd__clkbuf_16
Xfanout29 input3/X VGND VGND VPWR VPWR fanout29/X sky130_fd_sc_hd__clkbuf_4
Xfanout18 _446_/Q VGND VGND VPWR VPWR _425_/D sky130_fd_sc_hd__clkbuf_4
X_370_ _227_/S _303_/C _301_/B _369_/Y VGND VGND VPWR VPWR _436_/D sky130_fd_sc_hd__o31ai_1
X_284_ _306_/A _393_/B _455_/Q VGND VGND VPWR VPWR _284_/Y sky130_fd_sc_hd__nand3b_1
X_422_ _211_/A1 _422_/D fanout28/X VGND VGND VPWR VPWR _422_/Q sky130_fd_sc_hd__dfstp_1
X_353_ _377_/A _300_/Y _427_/Q VGND VGND VPWR VPWR _355_/A sky130_fd_sc_hd__o21ai_1
Xclkbuf_1_0__f_pll_clk clkbuf_0_pll_clk/X VGND VGND VPWR VPWR _448_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput8 sel[1] VGND VGND VPWR VPWR _443_/D sky130_fd_sc_hd__clkbuf_1
XTAP_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_336_ _450_/D _408_/A _335_/A VGND VGND VPWR VPWR _337_/B sky130_fd_sc_hd__o21a_1
X_267_ _267_/A VGND VGND VPWR VPWR _267_/Y sky130_fd_sc_hd__inv_2
X_405_ _464_/Q _403_/Y _404_/Y VGND VGND VPWR VPWR _464_/D sky130_fd_sc_hd__o21ai_1
X_319_ _426_/D _425_/D _377_/A VGND VGND VPWR VPWR _321_/A sky130_fd_sc_hd__nor3_1
Xfanout19 _424_/D VGND VGND VPWR VPWR _377_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input9_A sel[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__242__A1 _450_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__233__A1 _408_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__236__S _242_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_421_ _448_/CLK _421_/D fanout28/X VGND VGND VPWR VPWR _421_/Q sky130_fd_sc_hd__dfrtp_1
X_352_ _422_/Q _350_/Y _351_/Y VGND VGND VPWR VPWR _422_/D sky130_fd_sc_hd__o21ai_1
X_283_ _388_/A _259_/Y _247_/Y _306_/A VGND VGND VPWR VPWR _283_/Y sky130_fd_sc_hd__a31oi_2
XTAP_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput9 sel[2] VGND VGND VPWR VPWR _444_/D sky130_fd_sc_hd__clkbuf_1
XTAP_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_335_ _335_/A _450_/D _408_/A VGND VGND VPWR VPWR _337_/A sky130_fd_sc_hd__nor3_1
X_404_ _403_/Y _464_/Q _227_/S VGND VGND VPWR VPWR _404_/Y sky130_fd_sc_hd__a21oi_1
X_249_ _249_/A VGND VGND VPWR VPWR _249_/Y sky130_fd_sc_hd__inv_2
XANTENNA__409__A1 _408_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_318_ _434_/Q _433_/Q VGND VGND VPWR VPWR _318_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__336__B1 _335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_415__2 _211_/A1 VGND VGND VPWR VPWR _457_/CLK sky130_fd_sc_hd__inv_4
XANTENNA__465__SET_B fanout28/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_0_divider2.out _316_/X VGND VGND VPWR VPWR clkbuf_0_divider2.out/X sky130_fd_sc_hd__clkbuf_16
XFILLER_5_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_282_ _248_/Y _280_/X _281_/Y VGND VGND VPWR VPWR _457_/D sky130_fd_sc_hd__o21ai_1
X_351_ _350_/Y _422_/Q _242_/S VGND VGND VPWR VPWR _351_/Y sky130_fd_sc_hd__a21oi_1
X_420_ _208_/A1 _420_/D fanout27/X VGND VGND VPWR VPWR _421_/D sky130_fd_sc_hd__dfrtp_1
XANTENNA__390__A1 _242_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__381__A1 _408_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_403_ _447_/Q _446_/Q _424_/D _436_/Q _302_/Y VGND VGND VPWR VPWR _403_/Y sky130_fd_sc_hd__o2111ai_1
X_334_ _459_/Q _458_/Q VGND VGND VPWR VPWR _334_/Y sky130_fd_sc_hd__xnor2_1
X_265_ _452_/Q VGND VGND VPWR VPWR _382_/D sky130_fd_sc_hd__inv_2
X_248_ _457_/Q VGND VGND VPWR VPWR _248_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_317_ _425_/D _377_/A VGND VGND VPWR VPWR _317_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__336__A1 _450_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__245__A0 _450_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_281_ _274_/Y _388_/A _279_/Y _248_/Y _453_/Q VGND VGND VPWR VPWR _281_/Y sky130_fd_sc_hd__a41oi_1
X_350_ _473_/Q _472_/Q _449_/D _461_/Q _307_/Y VGND VGND VPWR VPWR _350_/Y sky130_fd_sc_hd__o2111ai_1
XTAP_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__390__A2 _388_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__466__RESET_B fanout28/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_402_ _242_/S _463_/Q _388_/A _401_/Y VGND VGND VPWR VPWR _463_/D sky130_fd_sc_hd__o31a_1
XFILLER_2_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_333_ _450_/D _408_/A VGND VGND VPWR VPWR _333_/Y sky130_fd_sc_hd__xnor2_1
X_264_ _427_/Q VGND VGND VPWR VPWR _354_/D sky130_fd_sc_hd__inv_2
X_316_ _315_/X _388_/A _314_/Y _313_/X VGND VGND VPWR VPWR _316_/X sky130_fd_sc_hd__a31o_2
X_247_ _459_/Q VGND VGND VPWR VPWR _247_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_14_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__336__A2 _408_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__236__A1 _450_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_280_ _335_/A _450_/D _408_/A _274_/Y _279_/Y VGND VGND VPWR VPWR _280_/X sky130_fd_sc_hd__o2111a_1
XANTENNA_input7_A sel[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_1_1__f_divider2.out clkbuf_0_divider2.out/X VGND VGND VPWR VPWR _473_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_401_ _306_/A _388_/A _244_/X VGND VGND VPWR VPWR _401_/Y sky130_fd_sc_hd__o21bai_1
X_332_ _440_/Q _439_/Q VGND VGND VPWR VPWR _332_/Y sky130_fd_sc_hd__xnor2_1
X_263_ _263_/A VGND VGND VPWR VPWR _420_/D sky130_fd_sc_hd__inv_2
XANTENNA__281__A2 _388_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_315_ _457_/Q _422_/Q VGND VGND VPWR VPWR _315_/X sky130_fd_sc_hd__or2_1
X_246_ _335_/A _348_/Y _305_/Y VGND VGND VPWR VPWR _246_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout28_A fanout29/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_229_ _426_/D _332_/Y _300_/Y VGND VGND VPWR VPWR _229_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f_ext_clk clkbuf_0_ext_clk/X VGND VGND VPWR VPWR _209_/A0 sky130_fd_sc_hd__clkbuf_16
X_262_ _461_/Q VGND VGND VPWR VPWR _308_/C sky130_fd_sc_hd__clkinv_4
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_331_ _331_/A _331_/B VGND VGND VPWR VPWR _331_/Y sky130_fd_sc_hd__nand2_1
X_400_ _242_/S _462_/Q _388_/A _399_/Y VGND VGND VPWR VPWR _462_/D sky130_fd_sc_hd__o31a_1
XFILLER_2_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_245_ _450_/D _258_/Y _305_/Y VGND VGND VPWR VPWR _245_/X sky130_fd_sc_hd__mux2_1
X_314_ _457_/Q _422_/Q VGND VGND VPWR VPWR _314_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__387__A_N _335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_228_ _425_/D _253_/Y _300_/Y VGND VGND VPWR VPWR _228_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__306__B _388_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_261_ _454_/Q VGND VGND VPWR VPWR _261_/Y sky130_fd_sc_hd__clkinv_2
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_330_ _436_/Q _437_/Q _438_/Q VGND VGND VPWR VPWR _331_/B sky130_fd_sc_hd__o21ai_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__437__SET_B fanout29/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_459_ _459_/CLK _459_/D fanout26/X VGND VGND VPWR VPWR _459_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_2_14 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_313_ _408_/A _313_/B VGND VGND VPWR VPWR _313_/X sky130_fd_sc_hd__and2b_2
X_244_ _243_/X _335_/A _306_/A VGND VGND VPWR VPWR _244_/X sky130_fd_sc_hd__mux2_1
X_227_ _226_/X _426_/D _227_/S VGND VGND VPWR VPWR _227_/X sky130_fd_sc_hd__mux2_1
XANTENNA__402__A1 _242_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_260_ _458_/Q VGND VGND VPWR VPWR _260_/Y sky130_fd_sc_hd__inv_2
XANTENNA_input5_A sel2[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__333__A _450_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_389_ _389_/A _389_/B _449_/Q VGND VGND VPWR VPWR _389_/Y sky130_fd_sc_hd__nand3_1
XFILLER_2_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_458_ _463_/CLK _458_/D fanout26/X VGND VGND VPWR VPWR _458_/Q sky130_fd_sc_hd__dfrtn_1
X_268__4 _448_/CLK VGND VGND VPWR VPWR _430_/CLK sky130_fd_sc_hd__inv_4
XTAP_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_243_ _347_/Y _335_/A _308_/Y VGND VGND VPWR VPWR _243_/X sky130_fd_sc_hd__mux2_1
X_312_ _311_/X _301_/B _310_/Y _309_/X VGND VGND VPWR VPWR _312_/X sky130_fd_sc_hd__a31o_2
X_226_ _331_/Y _447_/Q _303_/Y VGND VGND VPWR VPWR _226_/X sky130_fd_sc_hd__mux2_1
X_209_ _209_/A0 _423_/Q _421_/D VGND VGND VPWR VPWR _209_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__438__RESET_B fanout29/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_412__9 core_clk VGND VGND VPWR VPWR _419_/CLK sky130_fd_sc_hd__inv_4
XTAP_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__333__B _408_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__453__RESET_B fanout28/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_457_ _457_/CLK _457_/D fanout28/X VGND VGND VPWR VPWR _457_/Q sky130_fd_sc_hd__dfstp_1
X_388_ _388_/A _388_/B _388_/C VGND VGND VPWR VPWR _388_/Y sky130_fd_sc_hd__nand3_1
XTAP_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_311_ _432_/Q _464_/Q VGND VGND VPWR VPWR _311_/X sky130_fd_sc_hd__or2_1
X_242_ _241_/X _450_/D _242_/S VGND VGND VPWR VPWR _242_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0__f_ext_clk clkbuf_0_ext_clk/X VGND VGND VPWR VPWR _380_/A1 sky130_fd_sc_hd__clkbuf_16
X_225_ _224_/X _425_/D _227_/S VGND VGND VPWR VPWR _225_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__402__A3 _388_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_208_ _427_/Q _208_/A1 _288_/Y VGND VGND VPWR VPWR _309_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_473_ _473_/CLK _473_/D fanout29/X VGND VGND VPWR VPWR _473_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__472__SET_B fanout28/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_456_ _463_/CLK _456_/D fanout26/X VGND VGND VPWR VPWR _456_/Q sky130_fd_sc_hd__dfrtn_1
X_387_ _335_/A _451_/Q VGND VGND VPWR VPWR _388_/C sky130_fd_sc_hd__nand2b_1
XTAP_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_310_ _432_/Q _464_/Q VGND VGND VPWR VPWR _310_/Y sky130_fd_sc_hd__nand2_1
X_241_ _344_/Y _450_/D _308_/Y VGND VGND VPWR VPWR _241_/X sky130_fd_sc_hd__mux2_1
X_439_ _448_/CLK _439_/D _380_/S VGND VGND VPWR VPWR _439_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_11_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_224_ _328_/Y _446_/Q _303_/Y VGND VGND VPWR VPWR _224_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_207_ _306_/X _306_/A _278_/Y VGND VGND VPWR VPWR _396_/S sky130_fd_sc_hd__mux2_1
X_472_ _212_/A1 _472_/D fanout28/X VGND VGND VPWR VPWR _472_/Q sky130_fd_sc_hd__dfstp_1
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_455_ _455_/CLK _455_/D fanout26/X VGND VGND VPWR VPWR _455_/Q sky130_fd_sc_hd__dfstp_1
X_386_ _450_/Q _472_/Q VGND VGND VPWR VPWR _389_/B sky130_fd_sc_hd__nand2b_1
XTAP_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input3_A resetb VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_240_ _239_/X _449_/D _242_/S VGND VGND VPWR VPWR _240_/X sky130_fd_sc_hd__mux2_1
X_369_ _227_/S _301_/B _223_/X VGND VGND VPWR VPWR _369_/Y sky130_fd_sc_hd__o21ai_1
X_438_ _208_/A1 _438_/D fanout29/X VGND VGND VPWR VPWR _438_/Q sky130_fd_sc_hd__dfrtp_1
X_223_ _222_/X _424_/D _227_/S VGND VGND VPWR VPWR _223_/X sky130_fd_sc_hd__mux2_1
XANTENNA__399__A1 _242_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_206_ _301_/X _301_/A _291_/Y VGND VGND VPWR VPWR _368_/S sky130_fd_sc_hd__mux2_1
XFILLER_0_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_471_ _473_/CLK _471_/D fanout29/X VGND VGND VPWR VPWR _471_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_454_ _463_/CLK _454_/D fanout26/X VGND VGND VPWR VPWR _454_/Q sky130_fd_sc_hd__dfrtn_1
X_385_ _451_/Q _473_/Q VGND VGND VPWR VPWR _388_/B sky130_fd_sc_hd__nand2b_1
XTAP_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_299_ _440_/Q _441_/Q VGND VGND VPWR VPWR _354_/C sky130_fd_sc_hd__nor2_1
X_368_ _435_/Q _215_/X _368_/S VGND VGND VPWR VPWR _435_/D sky130_fd_sc_hd__mux2_1
X_437_ _208_/A1 _437_/D fanout29/X VGND VGND VPWR VPWR _437_/Q sky130_fd_sc_hd__dfstp_1
X_222_ _303_/C _424_/D _303_/Y VGND VGND VPWR VPWR _222_/X sky130_fd_sc_hd__mux2_1
XANTENNA__399__A2 _388_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_0_pll_clk90 pll_clk90 VGND VGND VPWR VPWR clkbuf_0_pll_clk90/X sky130_fd_sc_hd__clkbuf_16
XFILLER_0_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__241__A1 _450_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_470_ _473_/CLK _470_/D fanout29/X VGND VGND VPWR VPWR _473_/D sky130_fd_sc_hd__dfrtp_1
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_384_ _472_/Q _450_/Q VGND VGND VPWR VPWR _389_/A sky130_fd_sc_hd__nand2b_1
X_453_ _211_/A1 _453_/D fanout28/X VGND VGND VPWR VPWR _453_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__471__RESET_B fanout29/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__450__D _450_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_0_ext_clk_A ext_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__234__S _242_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_298_ _252_/Y _296_/Y _297_/Y VGND VGND VPWR VPWR _430_/D sky130_fd_sc_hd__o21ai_1
X_436_ _208_/A1 _436_/D fanout27/X VGND VGND VPWR VPWR _436_/Q sky130_fd_sc_hd__dfrtp_2
X_367_ _433_/Q _213_/X _368_/S VGND VGND VPWR VPWR _433_/D sky130_fd_sc_hd__mux2_1
X_221_ _220_/X _426_/D _301_/A VGND VGND VPWR VPWR _269_/A sky130_fd_sc_hd__mux2_1
X_419_ _419_/CLK _419_/D _380_/S VGND VGND VPWR VPWR _419_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__242__S _242_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_1_1__f_net10 clkbuf_0_net10/X VGND VGND VPWR VPWR _411__8/A sky130_fd_sc_hd__clkbuf_16
XANTENNA__388__A _388_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_383_ _383_/A _383_/B VGND VGND VPWR VPWR _452_/D sky130_fd_sc_hd__nand2_1
X_452_ _211_/A1 _452_/D fanout28/X VGND VGND VPWR VPWR _452_/Q sky130_fd_sc_hd__dfstp_1
XTAP_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_297_ _301_/A _365_/B _430_/Q VGND VGND VPWR VPWR _297_/Y sky130_fd_sc_hd__nand3b_1
X_366_ _269_/Y _296_/Y _365_/Y VGND VGND VPWR VPWR _431_/D sky130_fd_sc_hd__o21ai_1
X_435_ _448_/CLK _435_/D _380_/S VGND VGND VPWR VPWR _435_/Q sky130_fd_sc_hd__dfrtn_1
XANTENNA__280__B1 _408_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input1_A ext_clk_sel VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_220_ _327_/Y _426_/D _292_/Y VGND VGND VPWR VPWR _220_/X sky130_fd_sc_hd__mux2_1
X_349_ _349_/A _417_/Q VGND VGND VPWR VPWR _349_/Y sky130_fd_sc_hd__nor2_1
X_418_ _418_/CLK _419_/Q _380_/S VGND VGND VPWR VPWR _418_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_382_ _449_/D _465_/Q _382_/C _382_/D VGND VGND VPWR VPWR _383_/B sky130_fd_sc_hd__nand4b_1
X_451_ _211_/A1 _473_/Q VGND VGND VPWR VPWR _451_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_296_ _301_/B _255_/Y _250_/Y _301_/A VGND VGND VPWR VPWR _296_/Y sky130_fd_sc_hd__a31oi_2
X_365_ _301_/A _365_/B _431_/Q VGND VGND VPWR VPWR _365_/Y sky130_fd_sc_hd__nand3b_1
X_434_ _434_/CLK _434_/D _380_/S VGND VGND VPWR VPWR _434_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA__280__A1 _335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_417_ _417_/CLK _418_/Q fanout28/X VGND VGND VPWR VPWR _417_/Q sky130_fd_sc_hd__dfstp_1
X_279_ _455_/Q _456_/Q _454_/Q VGND VGND VPWR VPWR _279_/Y sky130_fd_sc_hd__nor3b_2
X_348_ _466_/Q _465_/Q VGND VGND VPWR VPWR _348_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__244__A1 _335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__235__A1 _450_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_416__3 _463_/CLK VGND VGND VPWR VPWR _459_/CLK sky130_fd_sc_hd__inv_4
XFILLER_18_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_419__30 VGND VGND VPWR VPWR _419__30/HI _419_/D sky130_fd_sc_hd__conb_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_381_ _408_/A _305_/Y _452_/Q VGND VGND VPWR VPWR _383_/A sky130_fd_sc_hd__o21ai_1
X_450_ _211_/A1 _450_/D VGND VGND VPWR VPWR _450_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_433_ _448_/CLK _433_/D _380_/S VGND VGND VPWR VPWR _433_/Q sky130_fd_sc_hd__dfrtn_1
XANTENNA__280__A2 _450_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_364_ _267_/Y _296_/Y _363_/Y VGND VGND VPWR VPWR _429_/D sky130_fd_sc_hd__o21ai_1
X_295_ _251_/Y _293_/X _294_/Y VGND VGND VPWR VPWR _432_/D sky130_fd_sc_hd__o21ai_1
X_347_ _347_/A _347_/B VGND VGND VPWR VPWR _347_/Y sky130_fd_sc_hd__nand2_1
X_278_ _393_/B VGND VGND VPWR VPWR _278_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_271__1 _463_/CLK VGND VGND VPWR VPWR _455_/CLK sky130_fd_sc_hd__inv_4
X_413__5 _208_/A1 VGND VGND VPWR VPWR _432_/CLK sky130_fd_sc_hd__inv_4
XFILLER_6_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_380_ _448_/Q _380_/A1 _380_/S VGND VGND VPWR VPWR _448_/D sky130_fd_sc_hd__mux2_1
XFILLER_15_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

