magic
tech sky130A
magscale 1 2
timestamp 1637778834
<< obsli1 >>
rect 1104 85 7975 8211
<< obsm1 >>
rect 14 76 8450 8220
<< metal2 >>
rect 18 8200 74 9000
rect 662 8200 718 9000
rect 1950 8200 2006 9000
rect 2594 8200 2650 9000
rect 3238 8200 3294 9000
rect 4526 8200 4582 9000
rect 5170 8200 5226 9000
rect 5814 8200 5870 9000
rect 7102 8200 7158 9000
rect 7746 8200 7802 9000
rect 8390 8200 8446 9000
rect 18 0 74 800
rect 662 0 718 800
rect 1306 0 1362 800
rect 2594 0 2650 800
rect 3238 0 3294 800
rect 3882 0 3938 800
rect 5170 0 5226 800
rect 5814 0 5870 800
rect 6458 0 6514 800
rect 7746 0 7802 800
rect 8390 0 8446 800
<< obsm2 >>
rect 130 8144 606 8945
rect 774 8144 1894 8945
rect 2062 8144 2538 8945
rect 2706 8144 3182 8945
rect 3350 8144 4470 8945
rect 4638 8144 5114 8945
rect 5282 8144 5758 8945
rect 5926 8144 7046 8945
rect 7214 8144 7690 8945
rect 7858 8144 8334 8945
rect 20 856 8444 8144
rect 130 31 606 856
rect 774 31 1250 856
rect 1418 31 2538 856
rect 2706 31 3182 856
rect 3350 31 3826 856
rect 3994 31 5114 856
rect 5282 31 5758 856
rect 5926 31 6402 856
rect 6570 31 7690 856
rect 7858 31 8334 856
<< metal3 >>
rect 0 8848 800 8968
rect 8200 8168 9000 8288
rect 0 7488 800 7608
rect 8200 7488 9000 7608
rect 0 6808 800 6928
rect 8200 6808 9000 6928
rect 0 6128 800 6248
rect 8200 5448 9000 5568
rect 0 4768 800 4888
rect 8200 4768 9000 4888
rect 0 4088 800 4208
rect 8200 4088 9000 4208
rect 0 3408 800 3528
rect 8200 2728 9000 2848
rect 0 2048 800 2168
rect 8200 2048 9000 2168
rect 0 1368 800 1488
rect 8200 1368 9000 1488
rect 0 688 800 808
rect 8200 8 9000 128
<< obsm3 >>
rect 880 8768 8200 8941
rect 800 8368 8200 8768
rect 800 8088 8120 8368
rect 800 7688 8200 8088
rect 880 7408 8120 7688
rect 800 7008 8200 7408
rect 880 6728 8120 7008
rect 800 6328 8200 6728
rect 880 6048 8200 6328
rect 800 5648 8200 6048
rect 800 5368 8120 5648
rect 800 4968 8200 5368
rect 880 4688 8120 4968
rect 800 4288 8200 4688
rect 880 4008 8120 4288
rect 800 3608 8200 4008
rect 880 3328 8200 3608
rect 800 2928 8200 3328
rect 800 2648 8120 2928
rect 800 2248 8200 2648
rect 880 1968 8120 2248
rect 800 1568 8200 1968
rect 880 1288 8120 1568
rect 800 888 8200 1288
rect 880 608 8200 888
rect 800 208 8200 608
rect 800 35 8120 208
<< metal4 >>
rect 1144 1040 1464 7664
rect 3144 1040 3464 7664
rect 5144 1040 5464 7664
rect 7144 1040 7464 7664
<< metal5 >>
rect 1104 5280 7820 5600
rect 1104 3280 7820 3600
rect 1104 1280 7820 1600
<< labels >>
rlabel metal3 s 0 2048 800 2168 6 spare_xfq[0]
port 1 nsew signal output
rlabel metal2 s 6458 0 6514 800 6 spare_xfq[1]
port 2 nsew signal output
rlabel metal2 s 4526 8200 4582 9000 6 spare_xfqn[0]
port 3 nsew signal output
rlabel metal3 s 0 6808 800 6928 6 spare_xfqn[1]
port 4 nsew signal output
rlabel metal2 s 8390 0 8446 800 6 spare_xi[0]
port 5 nsew signal output
rlabel metal3 s 8200 8 9000 128 6 spare_xi[1]
port 6 nsew signal output
rlabel metal3 s 8200 5448 9000 5568 6 spare_xi[2]
port 7 nsew signal output
rlabel metal2 s 18 8200 74 9000 6 spare_xi[3]
port 8 nsew signal output
rlabel metal3 s 0 7488 800 7608 6 spare_xib
port 9 nsew signal output
rlabel metal2 s 7102 8200 7158 9000 6 spare_xmx[0]
port 10 nsew signal output
rlabel metal2 s 5170 0 5226 800 6 spare_xmx[1]
port 11 nsew signal output
rlabel metal3 s 8200 6808 9000 6928 6 spare_xna[0]
port 12 nsew signal output
rlabel metal3 s 8200 1368 9000 1488 6 spare_xna[1]
port 13 nsew signal output
rlabel metal2 s 1306 0 1362 800 6 spare_xno[0]
port 14 nsew signal output
rlabel metal3 s 0 6128 800 6248 6 spare_xno[1]
port 15 nsew signal output
rlabel metal3 s 0 4088 800 4208 6 spare_xz[0]
port 16 nsew signal output
rlabel metal2 s 5170 8200 5226 9000 6 spare_xz[10]
port 17 nsew signal output
rlabel metal2 s 7746 8200 7802 9000 6 spare_xz[11]
port 18 nsew signal output
rlabel metal3 s 0 4768 800 4888 6 spare_xz[12]
port 19 nsew signal output
rlabel metal3 s 8200 7488 9000 7608 6 spare_xz[13]
port 20 nsew signal output
rlabel metal2 s 1950 8200 2006 9000 6 spare_xz[14]
port 21 nsew signal output
rlabel metal2 s 18 0 74 800 6 spare_xz[15]
port 22 nsew signal output
rlabel metal3 s 0 1368 800 1488 6 spare_xz[16]
port 23 nsew signal output
rlabel metal3 s 8200 4768 9000 4888 6 spare_xz[17]
port 24 nsew signal output
rlabel metal2 s 662 8200 718 9000 6 spare_xz[18]
port 25 nsew signal output
rlabel metal3 s 0 688 800 808 6 spare_xz[19]
port 26 nsew signal output
rlabel metal2 s 7746 0 7802 800 6 spare_xz[1]
port 27 nsew signal output
rlabel metal2 s 5814 8200 5870 9000 6 spare_xz[20]
port 28 nsew signal output
rlabel metal3 s 8200 2048 9000 2168 6 spare_xz[21]
port 29 nsew signal output
rlabel metal2 s 662 0 718 800 6 spare_xz[22]
port 30 nsew signal output
rlabel metal2 s 2594 0 2650 800 6 spare_xz[23]
port 31 nsew signal output
rlabel metal2 s 3238 0 3294 800 6 spare_xz[24]
port 32 nsew signal output
rlabel metal3 s 8200 2728 9000 2848 6 spare_xz[25]
port 33 nsew signal output
rlabel metal2 s 3882 0 3938 800 6 spare_xz[26]
port 34 nsew signal output
rlabel metal3 s 8200 8168 9000 8288 6 spare_xz[2]
port 35 nsew signal output
rlabel metal2 s 8390 8200 8446 9000 6 spare_xz[3]
port 36 nsew signal output
rlabel metal2 s 2594 8200 2650 9000 6 spare_xz[4]
port 37 nsew signal output
rlabel metal2 s 3238 8200 3294 9000 6 spare_xz[5]
port 38 nsew signal output
rlabel metal2 s 5814 0 5870 800 6 spare_xz[6]
port 39 nsew signal output
rlabel metal3 s 0 3408 800 3528 6 spare_xz[7]
port 40 nsew signal output
rlabel metal3 s 0 8848 800 8968 6 spare_xz[8]
port 41 nsew signal output
rlabel metal3 s 8200 4088 9000 4208 6 spare_xz[9]
port 42 nsew signal output
rlabel metal5 s 1104 1280 7820 1600 6 vccd
port 43 nsew power input
rlabel metal5 s 1104 5280 7820 5600 6 vccd
port 43 nsew power input
rlabel metal4 s 1144 1040 1464 7664 6 vccd
port 43 nsew power input
rlabel metal4 s 5144 1040 5464 7664 6 vccd
port 43 nsew power input
rlabel metal5 s 1104 3280 7820 3600 6 vssd
port 44 nsew ground input
rlabel metal4 s 3144 1040 3464 7664 6 vssd
port 44 nsew ground input
rlabel metal4 s 7144 1040 7464 7664 6 vssd
port 44 nsew ground input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 9000 9000
string LEFview TRUE
string GDS_FILE /home/ma/ef/caravel_openframe/openlane/spare_logic_block/runs/spare_logic_block/results/magic/spare_logic_block.gds
string GDS_END 175312
string GDS_START 71630
<< end >>

