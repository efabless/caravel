magic
tech sky130A
magscale 1 2
timestamp 1666350041
<< checkpaint >>
rect -1260 996747 718860 1038860
rect -1260 996340 42060 996747
rect 75940 996340 93460 996747
rect 127340 996340 144860 996747
rect 178740 996340 196260 996747
rect 219740 996340 256060 996747
rect 272340 996340 308660 996747
rect 332140 996340 349660 996747
rect 374140 996340 410460 996747
rect 472540 996340 490060 996747
rect 523940 996340 541460 996747
rect 574340 996340 591860 996747
rect 625740 996340 643260 996747
rect -1260 971460 40853 996340
rect 676340 995540 718860 996747
rect -1260 953940 41260 971460
rect 676747 967860 718860 995540
rect -1260 930447 40853 953940
rect 676340 950340 718860 967860
rect -1260 910740 43030 930447
rect 676747 923860 718860 950340
rect -1260 886060 40853 910740
rect 674570 904930 718860 923860
rect -1260 868540 41260 886060
rect 670350 884688 718860 904930
rect 676747 879692 718860 884688
rect -1260 843860 40853 868540
rect 674147 861108 718860 879692
rect -1260 826340 41260 843860
rect 676747 834660 718860 861108
rect -1260 825530 40853 826340
rect -1260 805288 56720 825530
rect 676340 817140 718860 834660
rect -1260 801692 40853 805288
rect -1260 783108 43453 801692
rect 676747 790492 718860 817140
rect -1260 782330 40853 783108
rect -1260 762088 56720 782330
rect 674147 771908 718860 790492
rect -1260 758492 40853 762088
rect -1260 739908 43453 758492
rect 676747 745492 718860 771908
rect -1260 739130 40853 739908
rect -1260 718888 56720 739130
rect 674147 726908 718860 745492
rect 676747 724330 718860 726908
rect -1260 715292 40853 718888
rect -1260 696708 43453 715292
rect 670360 704088 718860 724330
rect 676747 700492 718860 704088
rect -1260 695930 40853 696708
rect -1260 675688 56720 695930
rect 674147 681908 718860 700492
rect 676747 679130 718860 681908
rect -1260 672092 40853 675688
rect -1260 653508 43453 672092
rect 670360 658888 718860 679130
rect 676747 655292 718860 658888
rect -1260 652730 40853 653508
rect -1260 632488 56720 652730
rect 674147 636708 718860 655292
rect 676747 634130 718860 636708
rect -1260 628892 40853 632488
rect -1260 610308 43453 628892
rect 670360 613888 718860 634130
rect -1260 609530 40853 610308
rect 676747 610292 718860 613888
rect -1260 589288 56720 609530
rect 674147 591708 718860 610292
rect -1260 585692 40853 589288
rect 676747 588930 718860 591708
rect -1260 567108 43453 585692
rect 670360 568688 718860 588930
rect -1260 566330 40853 567108
rect -1260 546088 56720 566330
rect 676747 565092 718860 568688
rect 674147 546508 718860 565092
rect -1260 542492 40853 546088
rect 676747 543930 718860 546508
rect -1260 523908 43453 542492
rect -1260 499260 40853 523908
rect 670360 523688 718860 543930
rect 676747 520060 718860 523688
rect 676340 502540 718860 520060
rect 676747 499930 718860 502540
rect -1260 481740 41260 499260
rect -1260 459247 40853 481740
rect 670360 479688 718860 499930
rect 676747 476060 718860 479688
rect -1260 439540 43030 459247
rect 674570 456353 718860 476060
rect 676747 448974 718860 456353
rect -1260 438730 40853 439540
rect -1260 418488 56720 438730
rect 674265 437914 718860 448974
rect 676747 431860 718860 437914
rect -1260 414892 40853 418488
rect -1260 396308 43453 414892
rect 676340 414340 718860 431860
rect 676747 411730 718860 414340
rect -1260 395530 40853 396308
rect -1260 375288 56720 395530
rect 670360 391488 718860 411730
rect 676747 387892 718860 391488
rect -1260 371692 40853 375288
rect -1260 353108 43453 371692
rect 674147 369308 718860 387892
rect 676747 366530 718860 369308
rect -1260 352330 40853 353108
rect -1260 332088 56720 352330
rect 670360 346288 718860 366530
rect 676747 342692 718860 346288
rect -1260 328492 40853 332088
rect -1260 309908 43453 328492
rect 674147 324108 718860 342692
rect 676747 321530 718860 324108
rect -1260 309130 40853 309908
rect -1260 288888 56720 309130
rect 670360 301288 718860 321530
rect 676747 297692 718860 301288
rect -1260 285292 40853 288888
rect -1260 266708 43453 285292
rect 674147 279108 718860 297692
rect 676747 276530 718860 279108
rect -1260 265930 40853 266708
rect -1260 245688 56720 265930
rect 127986 247048 552310 263808
rect 670360 256288 718860 276530
rect 676747 252692 718860 256288
rect -1260 242092 40853 245688
rect 127986 242152 263154 247048
rect -1260 223508 43453 242092
rect 127986 241936 193510 242152
rect 215018 241936 263154 242152
rect 88438 232308 97750 241452
rect 108438 232308 117750 241452
rect 127986 240960 263154 241936
rect 263870 241536 333994 246328
rect 334618 244872 552310 247048
rect 334618 240960 379718 244872
rect 411254 244283 552310 244872
rect 387974 243509 392258 244283
rect 127986 238784 379718 240960
rect 385478 240049 392258 243509
rect 393062 240049 396194 243509
rect 407270 240049 552310 244283
rect 411254 238784 552310 240049
rect 127986 231816 552310 238784
rect 578438 232308 587750 241452
rect 674147 234108 718860 252692
rect 676747 231330 718860 234108
rect -1260 222730 40853 223508
rect -1260 202488 56720 222730
rect 640680 220372 649992 229516
rect 670360 211088 718860 231330
rect -1260 198892 40853 202488
rect -1260 180308 43453 198892
rect -1260 126460 40853 180308
rect -1260 108940 41260 126460
rect -1260 86499 40853 108940
rect 592240 100870 666596 209022
rect 676747 207492 718860 211088
rect 674147 188908 718860 207492
rect 676747 186330 718860 188908
rect 670360 166088 718860 186330
rect 676747 162492 718860 166088
rect 674147 143908 718860 162492
rect 676747 141130 718860 143908
rect 670360 120888 718860 141130
rect 676747 117292 718860 120888
rect 674147 98708 718860 117292
rect -1260 66740 42960 86499
rect 627952 80724 648304 95852
rect 656430 87906 663902 95418
rect -1260 42060 40853 66740
rect 625650 54520 646922 75088
rect 140928 45929 146556 51017
rect 457470 47380 467242 52716
rect 656287 49147 662299 50181
rect 656287 46721 662309 49147
rect 656297 45687 662309 46721
rect -1260 40853 41260 42060
rect 132502 41260 147150 45277
rect 77540 40853 95060 41260
rect 131216 40853 148963 41260
rect 150442 41029 160306 45277
rect 185108 40853 203692 43453
rect 237701 40853 257460 42960
rect 293708 40853 312292 43453
rect 348508 40853 367092 43453
rect 403308 40853 421892 43453
rect 427902 41029 442550 45277
rect 445842 41029 455706 45277
rect 458108 40853 476692 43453
rect 512908 40853 531492 43453
rect 676747 41260 718860 98708
rect 567740 40853 585260 41260
rect 621540 40853 639060 41260
rect 675540 40853 718860 41260
rect -1260 -1260 718860 40853
<< metal1 >>
rect 676030 897104 676036 897116
rect 663766 897076 676036 897104
rect 652018 896996 652024 897048
rect 652076 897036 652082 897048
rect 663766 897036 663794 897076
rect 676030 897064 676036 897076
rect 676088 897064 676094 897116
rect 652076 897008 663794 897036
rect 652076 896996 652082 897008
rect 654778 895772 654784 895824
rect 654836 895812 654842 895824
rect 675846 895812 675852 895824
rect 654836 895784 675852 895812
rect 654836 895772 654842 895784
rect 675846 895772 675852 895784
rect 675904 895772 675910 895824
rect 672718 895636 672724 895688
rect 672776 895676 672782 895688
rect 676030 895676 676036 895688
rect 672776 895648 676036 895676
rect 672776 895636 672782 895648
rect 676030 895636 676036 895648
rect 676088 895636 676094 895688
rect 672166 894412 672172 894464
rect 672224 894452 672230 894464
rect 675846 894452 675852 894464
rect 672224 894424 675852 894452
rect 672224 894412 672230 894424
rect 675846 894412 675852 894424
rect 675904 894412 675910 894464
rect 673362 894276 673368 894328
rect 673420 894316 673426 894328
rect 676030 894316 676036 894328
rect 673420 894288 676036 894316
rect 673420 894276 673426 894288
rect 676030 894276 676036 894288
rect 676088 894276 676094 894328
rect 671982 892984 671988 893036
rect 672040 893024 672046 893036
rect 676030 893024 676036 893036
rect 672040 892996 676036 893024
rect 672040 892984 672046 892996
rect 676030 892984 676036 892996
rect 676088 892984 676094 893036
rect 670970 892848 670976 892900
rect 671028 892888 671034 892900
rect 675846 892888 675852 892900
rect 671028 892860 675852 892888
rect 671028 892848 671034 892860
rect 675846 892848 675852 892860
rect 675904 892848 675910 892900
rect 676214 891488 676220 891540
rect 676272 891528 676278 891540
rect 676858 891528 676864 891540
rect 676272 891500 676864 891528
rect 676272 891488 676278 891500
rect 676858 891488 676864 891500
rect 676916 891488 676922 891540
rect 674834 890740 674840 890792
rect 674892 890780 674898 890792
rect 676030 890780 676036 890792
rect 674892 890752 676036 890780
rect 674892 890740 674898 890752
rect 676030 890740 676036 890752
rect 676088 890740 676094 890792
rect 676030 889992 676036 890044
rect 676088 890032 676094 890044
rect 677042 890032 677048 890044
rect 676088 890004 677048 890032
rect 676088 889992 676094 890004
rect 677042 889992 677048 890004
rect 677100 889992 677106 890044
rect 674650 888904 674656 888956
rect 674708 888944 674714 888956
rect 676030 888944 676036 888956
rect 674708 888916 676036 888944
rect 674708 888904 674714 888916
rect 676030 888904 676036 888916
rect 676088 888904 676094 888956
rect 675018 888768 675024 888820
rect 675076 888808 675082 888820
rect 675846 888808 675852 888820
rect 675076 888780 675852 888808
rect 675076 888768 675082 888780
rect 675846 888768 675852 888780
rect 675904 888768 675910 888820
rect 674282 888496 674288 888548
rect 674340 888536 674346 888548
rect 676030 888536 676036 888548
rect 674340 888508 676036 888536
rect 674340 888496 674346 888508
rect 676030 888496 676036 888508
rect 676088 888496 676094 888548
rect 673178 886864 673184 886916
rect 673236 886904 673242 886916
rect 676030 886904 676036 886916
rect 673236 886876 676036 886904
rect 673236 886864 673242 886876
rect 676030 886864 676036 886876
rect 676088 886864 676094 886916
rect 671798 885640 671804 885692
rect 671856 885680 671862 885692
rect 676030 885680 676036 885692
rect 671856 885652 676036 885680
rect 671856 885640 671862 885652
rect 676030 885640 676036 885652
rect 676088 885640 676094 885692
rect 675202 881016 675208 881068
rect 675260 881056 675266 881068
rect 683298 881056 683304 881068
rect 675260 881028 683304 881056
rect 675260 881016 675266 881028
rect 683298 881016 683304 881028
rect 683356 881016 683362 881068
rect 675570 880580 675576 880592
rect 663766 880552 675576 880580
rect 653398 880472 653404 880524
rect 653456 880512 653462 880524
rect 663766 880512 663794 880552
rect 675570 880540 675576 880552
rect 675628 880540 675634 880592
rect 653456 880484 663794 880512
rect 653456 880472 653462 880484
rect 675754 880404 675760 880456
rect 675812 880444 675818 880456
rect 679618 880444 679624 880456
rect 675812 880416 679624 880444
rect 675812 880404 675818 880416
rect 679618 880404 679624 880416
rect 679676 880404 679682 880456
rect 675386 879316 675392 879368
rect 675444 879356 675450 879368
rect 677042 879356 677048 879368
rect 675444 879328 677048 879356
rect 675444 879316 675450 879328
rect 677042 879316 677048 879328
rect 677100 879316 677106 879368
rect 674834 879180 674840 879232
rect 674892 879220 674898 879232
rect 675294 879220 675300 879232
rect 674892 879192 675300 879220
rect 674892 879180 674898 879192
rect 675294 879180 675300 879192
rect 675352 879180 675358 879232
rect 674834 879044 674840 879096
rect 674892 879084 674898 879096
rect 678238 879084 678244 879096
rect 674892 879056 678244 879084
rect 674892 879044 674898 879056
rect 678238 879044 678244 879056
rect 678296 879044 678302 879096
rect 676858 878540 676864 878552
rect 675588 878512 676864 878540
rect 675588 877724 675616 878512
rect 676858 878500 676864 878512
rect 676916 878500 676922 878552
rect 675496 877696 675616 877724
rect 675496 876580 675524 877696
rect 675478 876528 675484 876580
rect 675536 876528 675542 876580
rect 674466 876188 674472 876240
rect 674524 876228 674530 876240
rect 674834 876228 674840 876240
rect 674524 876200 674840 876228
rect 674524 876188 674530 876200
rect 674834 876188 674840 876200
rect 674892 876188 674898 876240
rect 674834 872856 674840 872908
rect 674892 872896 674898 872908
rect 675386 872896 675392 872908
rect 674892 872868 675392 872896
rect 674892 872856 674898 872868
rect 675386 872856 675392 872868
rect 675444 872856 675450 872908
rect 674282 870272 674288 870324
rect 674340 870312 674346 870324
rect 674926 870312 674932 870324
rect 674340 870284 674932 870312
rect 674340 870272 674346 870284
rect 674926 870272 674932 870284
rect 674984 870272 674990 870324
rect 657538 869388 657544 869440
rect 657596 869428 657602 869440
rect 657596 869400 675064 869428
rect 657596 869388 657602 869400
rect 675036 869032 675064 869400
rect 675202 869320 675208 869372
rect 675260 869320 675266 869372
rect 675220 869168 675248 869320
rect 675202 869116 675208 869168
rect 675260 869116 675266 869168
rect 675018 868980 675024 869032
rect 675076 868980 675082 869032
rect 651466 868844 651472 868896
rect 651524 868884 651530 868896
rect 654778 868884 654784 868896
rect 651524 868856 654784 868884
rect 651524 868844 651530 868856
rect 654778 868844 654784 868856
rect 654836 868844 654842 868896
rect 654134 868028 654140 868080
rect 654192 868068 654198 868080
rect 674834 868068 674840 868080
rect 654192 868040 674840 868068
rect 654192 868028 654198 868040
rect 674834 868028 674840 868040
rect 674892 868028 674898 868080
rect 651466 866600 651472 866652
rect 651524 866640 651530 866652
rect 672718 866640 672724 866652
rect 651524 866612 672724 866640
rect 651524 866600 651530 866612
rect 672718 866600 672724 866612
rect 672776 866600 672782 866652
rect 651374 865172 651380 865224
rect 651432 865212 651438 865224
rect 653398 865212 653404 865224
rect 651432 865184 653404 865212
rect 651432 865172 651438 865184
rect 653398 865172 653404 865184
rect 653456 865172 653462 865224
rect 651466 863812 651472 863864
rect 651524 863852 651530 863864
rect 657538 863852 657544 863864
rect 651524 863824 657544 863852
rect 651524 863812 651530 863824
rect 657538 863812 657544 863824
rect 657596 863812 657602 863864
rect 651466 862452 651472 862504
rect 651524 862492 651530 862504
rect 654134 862492 654140 862504
rect 651524 862464 654140 862492
rect 651524 862452 651530 862464
rect 654134 862452 654140 862464
rect 654192 862452 654198 862504
rect 35618 817096 35624 817148
rect 35676 817096 35682 817148
rect 35802 817096 35808 817148
rect 35860 817136 35866 817148
rect 44818 817136 44824 817148
rect 35860 817108 44824 817136
rect 35860 817096 35866 817108
rect 44818 817096 44824 817108
rect 44876 817096 44882 817148
rect 35636 817000 35664 817096
rect 61378 817000 61384 817012
rect 35636 816972 61384 817000
rect 61378 816960 61384 816972
rect 61436 816960 61442 817012
rect 35618 815736 35624 815788
rect 35676 815776 35682 815788
rect 43438 815776 43444 815788
rect 35676 815748 43444 815776
rect 35676 815736 35682 815748
rect 43438 815736 43444 815748
rect 43496 815736 43502 815788
rect 35802 815600 35808 815652
rect 35860 815640 35866 815652
rect 44174 815640 44180 815652
rect 35860 815612 44180 815640
rect 35860 815600 35866 815612
rect 44174 815600 44180 815612
rect 44232 815600 44238 815652
rect 35802 814376 35808 814428
rect 35860 814416 35866 814428
rect 44358 814416 44364 814428
rect 35860 814388 44364 814416
rect 35860 814376 35866 814388
rect 44358 814376 44364 814388
rect 44416 814376 44422 814428
rect 35618 814240 35624 814292
rect 35676 814280 35682 814292
rect 44542 814280 44548 814292
rect 35676 814252 44548 814280
rect 35676 814240 35682 814252
rect 44542 814240 44548 814252
rect 44600 814240 44606 814292
rect 41322 812812 41328 812864
rect 41380 812852 41386 812864
rect 43254 812852 43260 812864
rect 41380 812824 43260 812852
rect 41380 812812 41386 812824
rect 43254 812812 43260 812824
rect 43312 812812 43318 812864
rect 41322 811452 41328 811504
rect 41380 811492 41386 811504
rect 41782 811492 41788 811504
rect 41380 811464 41788 811492
rect 41380 811452 41386 811464
rect 41782 811452 41788 811464
rect 41840 811452 41846 811504
rect 31662 809344 31668 809396
rect 31720 809384 31726 809396
rect 42426 809384 42432 809396
rect 31720 809356 42432 809384
rect 31720 809344 31726 809356
rect 42426 809344 42432 809356
rect 42484 809344 42490 809396
rect 41322 808664 41328 808716
rect 41380 808704 41386 808716
rect 43070 808704 43076 808716
rect 41380 808676 43076 808704
rect 41380 808664 41386 808676
rect 43070 808664 43076 808676
rect 43128 808664 43134 808716
rect 43438 807916 43444 807968
rect 43496 807956 43502 807968
rect 62758 807956 62764 807968
rect 43496 807928 62764 807956
rect 43496 807916 43502 807928
rect 62758 807916 62764 807928
rect 62816 807916 62822 807968
rect 41322 807440 41328 807492
rect 41380 807480 41386 807492
rect 42886 807480 42892 807492
rect 41380 807452 42892 807480
rect 41380 807440 41386 807452
rect 42886 807440 42892 807452
rect 42944 807440 42950 807492
rect 41138 807304 41144 807356
rect 41196 807344 41202 807356
rect 43438 807344 43444 807356
rect 41196 807316 43444 807344
rect 41196 807304 41202 807316
rect 43438 807304 43444 807316
rect 43496 807304 43502 807356
rect 41322 806080 41328 806132
rect 41380 806120 41386 806132
rect 43806 806120 43812 806132
rect 41380 806092 43812 806120
rect 41380 806080 41386 806092
rect 43806 806080 43812 806092
rect 43864 806080 43870 806132
rect 41138 805944 41144 805996
rect 41196 805984 41202 805996
rect 64138 805984 64144 805996
rect 41196 805956 64144 805984
rect 41196 805944 41202 805956
rect 64138 805944 64144 805956
rect 64196 805944 64202 805996
rect 30282 805196 30288 805248
rect 30340 805236 30346 805248
rect 42702 805236 42708 805248
rect 30340 805208 42708 805236
rect 30340 805196 30346 805208
rect 42702 805196 42708 805208
rect 42760 805196 42766 805248
rect 32214 802408 32220 802460
rect 32272 802448 32278 802460
rect 41782 802448 41788 802460
rect 32272 802420 41788 802448
rect 32272 802408 32278 802420
rect 41782 802408 41788 802420
rect 41840 802408 41846 802460
rect 33778 801184 33784 801236
rect 33836 801224 33842 801236
rect 42610 801224 42616 801236
rect 33836 801196 42616 801224
rect 33836 801184 33842 801196
rect 42610 801184 42616 801196
rect 42668 801184 42674 801236
rect 31018 801048 31024 801100
rect 31076 801088 31082 801100
rect 40494 801088 40500 801100
rect 31076 801060 40500 801088
rect 31076 801048 31082 801060
rect 40494 801048 40500 801060
rect 40552 801048 40558 801100
rect 43622 799076 43628 799128
rect 43680 799116 43686 799128
rect 53098 799116 53104 799128
rect 43680 799088 53104 799116
rect 43680 799076 43686 799088
rect 53098 799076 53104 799088
rect 53156 799076 53162 799128
rect 45002 797648 45008 797700
rect 45060 797688 45066 797700
rect 57238 797688 57244 797700
rect 45060 797660 57244 797688
rect 45060 797648 45066 797660
rect 57238 797648 57244 797660
rect 57296 797648 57302 797700
rect 42242 796832 42248 796884
rect 42300 796872 42306 796884
rect 42610 796872 42616 796884
rect 42300 796844 42616 796872
rect 42300 796832 42306 796844
rect 42610 796832 42616 796844
rect 42668 796832 42674 796884
rect 42702 794724 42708 794776
rect 42760 794764 42766 794776
rect 43438 794764 43444 794776
rect 42760 794736 43444 794764
rect 42760 794724 42766 794736
rect 43438 794724 43444 794736
rect 43496 794724 43502 794776
rect 653398 790780 653404 790832
rect 653456 790820 653462 790832
rect 675386 790820 675392 790832
rect 653456 790792 675392 790820
rect 653456 790780 653462 790792
rect 675386 790780 675392 790792
rect 675444 790780 675450 790832
rect 53098 790712 53104 790764
rect 53156 790752 53162 790764
rect 62206 790752 62212 790764
rect 53156 790724 62212 790752
rect 53156 790712 53162 790724
rect 62206 790712 62212 790724
rect 62264 790712 62270 790764
rect 42242 789692 42248 789744
rect 42300 789692 42306 789744
rect 42260 789540 42288 789692
rect 42242 789488 42248 789540
rect 42300 789488 42306 789540
rect 670602 789352 670608 789404
rect 670660 789392 670666 789404
rect 675110 789392 675116 789404
rect 670660 789364 675116 789392
rect 670660 789352 670666 789364
rect 675110 789352 675116 789364
rect 675168 789352 675174 789404
rect 57238 789148 57244 789200
rect 57296 789188 57302 789200
rect 62114 789188 62120 789200
rect 57296 789160 62120 789188
rect 57296 789148 57302 789160
rect 62114 789148 62120 789160
rect 62172 789148 62178 789200
rect 42610 786632 42616 786684
rect 42668 786672 42674 786684
rect 62114 786672 62120 786684
rect 42668 786644 62120 786672
rect 42668 786632 42674 786644
rect 62114 786632 62120 786644
rect 62172 786632 62178 786684
rect 44818 785136 44824 785188
rect 44876 785176 44882 785188
rect 62114 785176 62120 785188
rect 44876 785148 62120 785176
rect 44876 785136 44882 785148
rect 62114 785136 62120 785148
rect 62172 785136 62178 785188
rect 674466 783844 674472 783896
rect 674524 783884 674530 783896
rect 675110 783884 675116 783896
rect 674524 783856 675116 783884
rect 674524 783844 674530 783856
rect 675110 783844 675116 783856
rect 675168 783844 675174 783896
rect 674742 782620 674748 782672
rect 674800 782660 674806 782672
rect 675202 782660 675208 782672
rect 674800 782632 675208 782660
rect 674800 782620 674806 782632
rect 675202 782620 675208 782632
rect 675260 782620 675266 782672
rect 655514 781056 655520 781108
rect 655572 781096 655578 781108
rect 675202 781096 675208 781108
rect 655572 781068 675208 781096
rect 655572 781056 655578 781068
rect 675202 781056 675208 781068
rect 675260 781056 675266 781108
rect 655054 778336 655060 778388
rect 655112 778376 655118 778388
rect 675202 778376 675208 778388
rect 655112 778348 675208 778376
rect 655112 778336 655118 778348
rect 675202 778336 675208 778348
rect 675260 778336 675266 778388
rect 651466 777588 651472 777640
rect 651524 777628 651530 777640
rect 660298 777628 660304 777640
rect 651524 777600 660304 777628
rect 651524 777588 651530 777600
rect 660298 777588 660304 777600
rect 660356 777588 660362 777640
rect 674282 776976 674288 777028
rect 674340 777016 674346 777028
rect 675294 777016 675300 777028
rect 674340 776988 675300 777016
rect 674340 776976 674346 776988
rect 675294 776976 675300 776988
rect 675352 776976 675358 777028
rect 651466 775548 651472 775600
rect 651524 775588 651530 775600
rect 669958 775588 669964 775600
rect 651524 775560 669964 775588
rect 651524 775548 651530 775560
rect 669958 775548 669964 775560
rect 670016 775548 670022 775600
rect 670786 775548 670792 775600
rect 670844 775588 670850 775600
rect 674834 775588 674840 775600
rect 670844 775560 674840 775588
rect 670844 775548 670850 775560
rect 674834 775548 674840 775560
rect 674892 775548 674898 775600
rect 651374 775276 651380 775328
rect 651432 775316 651438 775328
rect 653398 775316 653404 775328
rect 651432 775288 653404 775316
rect 651432 775276 651438 775288
rect 653398 775276 653404 775288
rect 653456 775276 653462 775328
rect 35802 774188 35808 774240
rect 35860 774228 35866 774240
rect 41690 774228 41696 774240
rect 35860 774200 41696 774228
rect 35860 774188 35866 774200
rect 41690 774188 41696 774200
rect 41748 774188 41754 774240
rect 42058 774188 42064 774240
rect 42116 774228 42122 774240
rect 59998 774228 60004 774240
rect 42116 774200 60004 774228
rect 42116 774188 42122 774200
rect 59998 774188 60004 774200
rect 60056 774188 60062 774240
rect 651466 774120 651472 774172
rect 651524 774160 651530 774172
rect 655514 774160 655520 774172
rect 651524 774132 655520 774160
rect 651524 774120 651530 774132
rect 655514 774120 655520 774132
rect 655572 774120 655578 774172
rect 651466 773780 651472 773832
rect 651524 773820 651530 773832
rect 655054 773820 655060 773832
rect 651524 773792 655060 773820
rect 651524 773780 651530 773792
rect 655054 773780 655060 773792
rect 655112 773780 655118 773832
rect 35434 773372 35440 773424
rect 35492 773412 35498 773424
rect 41506 773412 41512 773424
rect 35492 773384 41512 773412
rect 35492 773372 35498 773384
rect 41506 773372 41512 773384
rect 41564 773372 41570 773424
rect 41690 773208 41696 773220
rect 41386 773180 41696 773208
rect 35802 773100 35808 773152
rect 35860 773140 35866 773152
rect 41386 773140 41414 773180
rect 41690 773168 41696 773180
rect 41748 773168 41754 773220
rect 42058 773168 42064 773220
rect 42116 773208 42122 773220
rect 44174 773208 44180 773220
rect 42116 773180 44180 773208
rect 42116 773168 42122 773180
rect 44174 773168 44180 773180
rect 44232 773168 44238 773220
rect 35860 773112 41414 773140
rect 35860 773100 35866 773112
rect 41690 773072 41696 773084
rect 41524 773044 41696 773072
rect 35618 772964 35624 773016
rect 35676 773004 35682 773016
rect 41524 773004 41552 773044
rect 41690 773032 41696 773044
rect 41748 773032 41754 773084
rect 42058 773032 42064 773084
rect 42116 773072 42122 773084
rect 46198 773072 46204 773084
rect 42116 773044 46204 773072
rect 42116 773032 42122 773044
rect 46198 773032 46204 773044
rect 46256 773032 46262 773084
rect 35676 772976 41552 773004
rect 35676 772964 35682 772976
rect 35250 772828 35256 772880
rect 35308 772868 35314 772880
rect 41690 772868 41696 772880
rect 35308 772840 41696 772868
rect 35308 772828 35314 772840
rect 41690 772828 41696 772840
rect 41748 772828 41754 772880
rect 42058 772828 42064 772880
rect 42116 772868 42122 772880
rect 61378 772868 61384 772880
rect 42116 772840 61384 772868
rect 42116 772828 42122 772840
rect 61378 772828 61384 772840
rect 61436 772828 61442 772880
rect 35802 771808 35808 771860
rect 35860 771848 35866 771860
rect 39482 771848 39488 771860
rect 35860 771820 39488 771848
rect 35860 771808 35866 771820
rect 39482 771808 39488 771820
rect 39540 771808 39546 771860
rect 42058 771604 42064 771656
rect 42116 771644 42122 771656
rect 44542 771644 44548 771656
rect 42116 771616 44548 771644
rect 42116 771604 42122 771616
rect 44542 771604 44548 771616
rect 44600 771604 44606 771656
rect 35618 771536 35624 771588
rect 35676 771576 35682 771588
rect 41690 771576 41696 771588
rect 35676 771548 41696 771576
rect 35676 771536 35682 771548
rect 41690 771536 41696 771548
rect 41748 771536 41754 771588
rect 35802 771400 35808 771452
rect 35860 771440 35866 771452
rect 41690 771440 41696 771452
rect 35860 771412 41696 771440
rect 35860 771400 35866 771412
rect 41690 771400 41696 771412
rect 41748 771400 41754 771452
rect 42058 771400 42064 771452
rect 42116 771440 42122 771452
rect 44358 771440 44364 771452
rect 42116 771412 44364 771440
rect 42116 771400 42122 771412
rect 44358 771400 44364 771412
rect 44416 771400 44422 771452
rect 35802 770448 35808 770500
rect 35860 770488 35866 770500
rect 39114 770488 39120 770500
rect 35860 770460 39120 770488
rect 35860 770448 35866 770460
rect 39114 770448 39120 770460
rect 39172 770448 39178 770500
rect 35802 770176 35808 770228
rect 35860 770216 35866 770228
rect 39850 770216 39856 770228
rect 35860 770188 39856 770216
rect 35860 770176 35866 770188
rect 39850 770176 39856 770188
rect 39908 770176 39914 770228
rect 35618 770040 35624 770092
rect 35676 770080 35682 770092
rect 41690 770080 41696 770092
rect 35676 770052 41696 770080
rect 35676 770040 35682 770052
rect 41690 770040 41696 770052
rect 41748 770040 41754 770092
rect 42058 770040 42064 770092
rect 42116 770080 42122 770092
rect 45370 770080 45376 770092
rect 42116 770052 45376 770080
rect 42116 770040 42122 770052
rect 45370 770040 45376 770052
rect 45428 770040 45434 770092
rect 35802 768952 35808 769004
rect 35860 768992 35866 769004
rect 41690 768992 41696 769004
rect 35860 768964 41696 768992
rect 35860 768952 35866 768964
rect 41690 768952 41696 768964
rect 41748 768952 41754 769004
rect 35802 768816 35808 768868
rect 35860 768856 35866 768868
rect 39758 768856 39764 768868
rect 35860 768828 39764 768856
rect 35860 768816 35866 768828
rect 39758 768816 39764 768828
rect 39816 768816 39822 768868
rect 35618 768680 35624 768732
rect 35676 768720 35682 768732
rect 40034 768720 40040 768732
rect 35676 768692 40040 768720
rect 35676 768680 35682 768692
rect 40034 768680 40040 768692
rect 40092 768680 40098 768732
rect 35802 767320 35808 767372
rect 35860 767360 35866 767372
rect 36538 767360 36544 767372
rect 35860 767332 36544 767360
rect 35860 767320 35866 767332
rect 36538 767320 36544 767332
rect 36596 767320 36602 767372
rect 35802 766096 35808 766148
rect 35860 766136 35866 766148
rect 39574 766136 39580 766148
rect 35860 766108 39580 766136
rect 35860 766096 35866 766108
rect 39574 766096 39580 766108
rect 39632 766096 39638 766148
rect 35802 764804 35808 764856
rect 35860 764844 35866 764856
rect 40126 764844 40132 764856
rect 35860 764816 40132 764844
rect 35860 764804 35866 764816
rect 40126 764804 40132 764816
rect 40184 764804 40190 764856
rect 35802 764532 35808 764584
rect 35860 764572 35866 764584
rect 41690 764572 41696 764584
rect 35860 764544 41696 764572
rect 35860 764532 35866 764544
rect 41690 764532 41696 764544
rect 41748 764532 41754 764584
rect 42058 764532 42064 764584
rect 42116 764572 42122 764584
rect 44174 764572 44180 764584
rect 42116 764544 44180 764572
rect 42116 764532 42122 764544
rect 44174 764532 44180 764544
rect 44232 764532 44238 764584
rect 35618 763376 35624 763428
rect 35676 763416 35682 763428
rect 35676 763388 38654 763416
rect 35676 763376 35682 763388
rect 38626 763348 38654 763388
rect 40494 763348 40500 763360
rect 38626 763320 40500 763348
rect 40494 763308 40500 763320
rect 40552 763308 40558 763360
rect 42058 763308 42064 763360
rect 42116 763348 42122 763360
rect 42116 763320 51074 763348
rect 42116 763308 42122 763320
rect 35802 763172 35808 763224
rect 35860 763212 35866 763224
rect 41690 763212 41696 763224
rect 35860 763184 41696 763212
rect 35860 763172 35866 763184
rect 41690 763172 41696 763184
rect 41748 763172 41754 763224
rect 51046 763212 51074 763320
rect 58618 763212 58624 763224
rect 51046 763184 58624 763212
rect 58618 763172 58624 763184
rect 58676 763172 58682 763224
rect 35802 761880 35808 761932
rect 35860 761920 35866 761932
rect 39942 761920 39948 761932
rect 35860 761892 39948 761920
rect 35860 761880 35866 761892
rect 39942 761880 39948 761892
rect 40000 761880 40006 761932
rect 35158 759772 35164 759824
rect 35216 759812 35222 759824
rect 41690 759812 41696 759824
rect 35216 759784 41696 759812
rect 35216 759772 35222 759784
rect 41690 759772 41696 759784
rect 41748 759772 41754 759824
rect 32398 759636 32404 759688
rect 32456 759676 32462 759688
rect 41598 759676 41604 759688
rect 32456 759648 41604 759676
rect 32456 759636 32462 759648
rect 41598 759636 41604 759648
rect 41656 759636 41662 759688
rect 33778 758276 33784 758328
rect 33836 758316 33842 758328
rect 39850 758316 39856 758328
rect 33836 758288 39856 758316
rect 33836 758276 33842 758288
rect 39850 758276 39856 758288
rect 39908 758276 39914 758328
rect 44726 755488 44732 755540
rect 44784 755528 44790 755540
rect 62758 755528 62764 755540
rect 44784 755500 62764 755528
rect 44784 755488 44790 755500
rect 62758 755488 62764 755500
rect 62816 755488 62822 755540
rect 42242 754264 42248 754316
rect 42300 754304 42306 754316
rect 44726 754304 44732 754316
rect 42300 754276 44732 754304
rect 42300 754264 42306 754276
rect 44726 754264 44732 754276
rect 44784 754264 44790 754316
rect 42426 754128 42432 754180
rect 42484 754168 42490 754180
rect 42794 754168 42800 754180
rect 42484 754140 42800 754168
rect 42484 754128 42490 754140
rect 42794 754128 42800 754140
rect 42852 754128 42858 754180
rect 42242 751476 42248 751528
rect 42300 751476 42306 751528
rect 42260 751188 42288 751476
rect 42242 751136 42248 751188
rect 42300 751136 42306 751188
rect 61378 747124 61384 747176
rect 61436 747164 61442 747176
rect 63034 747164 63040 747176
rect 61436 747136 63040 747164
rect 61436 747124 61442 747136
rect 63034 747124 63040 747136
rect 63092 747124 63098 747176
rect 45094 746512 45100 746564
rect 45152 746552 45158 746564
rect 62114 746552 62120 746564
rect 45152 746524 62120 746552
rect 45152 746512 45158 746524
rect 62114 746512 62120 746524
rect 62172 746512 62178 746564
rect 671338 743996 671344 744048
rect 671396 744036 671402 744048
rect 675386 744036 675392 744048
rect 671396 744008 675392 744036
rect 671396 743996 671402 744008
rect 675386 743996 675392 744008
rect 675444 743996 675450 744048
rect 42518 743860 42524 743912
rect 42576 743900 42582 743912
rect 62114 743900 62120 743912
rect 42576 743872 62120 743900
rect 42576 743860 42582 743872
rect 62114 743860 62120 743872
rect 62172 743860 62178 743912
rect 46198 743724 46204 743776
rect 46256 743764 46262 743776
rect 62114 743764 62120 743776
rect 46256 743736 62120 743764
rect 46256 743724 46262 743736
rect 62114 743724 62120 743736
rect 62172 743724 62178 743776
rect 671154 743180 671160 743232
rect 671212 743220 671218 743232
rect 675294 743220 675300 743232
rect 671212 743192 675300 743220
rect 671212 743180 671218 743192
rect 675294 743180 675300 743192
rect 675352 743180 675358 743232
rect 672350 742772 672356 742824
rect 672408 742812 672414 742824
rect 675478 742812 675484 742824
rect 672408 742784 675484 742812
rect 672408 742772 672414 742784
rect 675478 742772 675484 742784
rect 675536 742772 675542 742824
rect 59998 742364 60004 742416
rect 60056 742404 60062 742416
rect 62114 742404 62120 742416
rect 60056 742376 62120 742404
rect 60056 742364 60062 742376
rect 62114 742364 62120 742376
rect 62172 742364 62178 742416
rect 669222 741072 669228 741124
rect 669280 741112 669286 741124
rect 674834 741112 674840 741124
rect 669280 741084 674840 741112
rect 669280 741072 669286 741084
rect 674834 741072 674840 741084
rect 674892 741072 674898 741124
rect 674834 740596 674840 740648
rect 674892 740636 674898 740648
rect 675386 740636 675392 740648
rect 674892 740608 675392 740636
rect 674892 740596 674898 740608
rect 675386 740596 675392 740608
rect 675444 740596 675450 740648
rect 652018 736176 652024 736228
rect 652076 736216 652082 736228
rect 653398 736216 653404 736228
rect 652076 736188 653404 736216
rect 652076 736176 652082 736188
rect 653398 736176 653404 736188
rect 653456 736176 653462 736228
rect 675202 735740 675208 735752
rect 663766 735712 675208 735740
rect 657538 735564 657544 735616
rect 657596 735604 657602 735616
rect 663766 735604 663794 735712
rect 675202 735700 675208 735712
rect 675260 735700 675266 735752
rect 657596 735576 663794 735604
rect 657596 735564 657602 735576
rect 675110 734244 675116 734256
rect 663766 734216 675116 734244
rect 654778 734136 654784 734188
rect 654836 734176 654842 734188
rect 663766 734176 663794 734216
rect 675110 734204 675116 734216
rect 675168 734204 675174 734256
rect 654836 734148 663794 734176
rect 654836 734136 654842 734148
rect 668670 733864 668676 733916
rect 668728 733904 668734 733916
rect 668728 733876 675340 733904
rect 668728 733864 668734 733876
rect 651466 733388 651472 733440
rect 651524 733428 651530 733440
rect 668026 733428 668032 733440
rect 651524 733400 668032 733428
rect 651524 733388 651530 733400
rect 668026 733388 668032 733400
rect 668084 733388 668090 733440
rect 675312 733372 675340 733876
rect 675294 733320 675300 733372
rect 675352 733320 675358 733372
rect 651466 732776 651472 732828
rect 651524 732816 651530 732828
rect 661678 732816 661684 732828
rect 651524 732788 661684 732816
rect 651524 732776 651530 732788
rect 661678 732776 661684 732788
rect 661736 732776 661742 732828
rect 651466 731416 651472 731468
rect 651524 731456 651530 731468
rect 658918 731456 658924 731468
rect 651524 731428 658924 731456
rect 651524 731416 651530 731428
rect 658918 731416 658924 731428
rect 658976 731416 658982 731468
rect 651466 731280 651472 731332
rect 651524 731320 651530 731332
rect 671338 731320 671344 731332
rect 651524 731292 671344 731320
rect 651524 731280 651530 731292
rect 671338 731280 671344 731292
rect 671396 731280 671402 731332
rect 41690 730300 41696 730312
rect 41386 730272 41696 730300
rect 41138 730192 41144 730244
rect 41196 730232 41202 730244
rect 41386 730232 41414 730272
rect 41690 730260 41696 730272
rect 41748 730260 41754 730312
rect 42058 730260 42064 730312
rect 42116 730300 42122 730312
rect 46198 730300 46204 730312
rect 42116 730272 46204 730300
rect 42116 730260 42122 730272
rect 46198 730260 46204 730272
rect 46256 730260 46262 730312
rect 41196 730204 41414 730232
rect 41196 730192 41202 730204
rect 43438 730124 43444 730176
rect 43496 730164 43502 730176
rect 43496 730136 51074 730164
rect 43496 730124 43502 730136
rect 51046 730096 51074 730136
rect 61378 730096 61384 730108
rect 51046 730068 61384 730096
rect 61378 730056 61384 730068
rect 61436 730056 61442 730108
rect 651466 729988 651472 730040
rect 651524 730028 651530 730040
rect 657538 730028 657544 730040
rect 651524 730000 657544 730028
rect 651524 729988 651530 730000
rect 657538 729988 657544 730000
rect 657596 729988 657602 730040
rect 43622 729308 43628 729360
rect 43680 729348 43686 729360
rect 62758 729348 62764 729360
rect 43680 729320 62764 729348
rect 43680 729308 43686 729320
rect 62758 729308 62764 729320
rect 62816 729308 62822 729360
rect 41322 729036 41328 729088
rect 41380 729076 41386 729088
rect 41690 729076 41696 729088
rect 41380 729048 41696 729076
rect 41380 729036 41386 729048
rect 41690 729036 41696 729048
rect 41748 729036 41754 729088
rect 42058 728628 42064 728680
rect 42116 728668 42122 728680
rect 43070 728668 43076 728680
rect 42116 728640 43076 728668
rect 42116 728628 42122 728640
rect 43070 728628 43076 728640
rect 43128 728628 43134 728680
rect 651466 728492 651472 728544
rect 651524 728532 651530 728544
rect 654778 728532 654784 728544
rect 651524 728504 654784 728532
rect 651524 728492 651530 728504
rect 654778 728492 654784 728504
rect 654836 728492 654842 728544
rect 671798 728288 671804 728340
rect 671856 728328 671862 728340
rect 671856 728300 674176 728328
rect 671856 728288 671862 728300
rect 673178 728084 673184 728136
rect 673236 728124 673242 728136
rect 673236 728096 674058 728124
rect 673236 728084 673242 728096
rect 674466 727880 674472 727932
rect 674524 727920 674530 727932
rect 683482 727920 683488 727932
rect 674524 727892 683488 727920
rect 674524 727880 674530 727892
rect 683482 727880 683488 727892
rect 683540 727880 683546 727932
rect 674834 727472 674840 727524
rect 674892 727472 674898 727524
rect 675110 727472 675116 727524
rect 675168 727512 675174 727524
rect 675478 727512 675484 727524
rect 675168 727484 675484 727512
rect 675168 727472 675174 727484
rect 675478 727472 675484 727484
rect 675536 727472 675542 727524
rect 41046 727404 41052 727456
rect 41104 727444 41110 727456
rect 41690 727444 41696 727456
rect 41104 727416 41696 727444
rect 41104 727404 41110 727416
rect 41690 727404 41696 727416
rect 41748 727404 41754 727456
rect 42058 727404 42064 727456
rect 42116 727444 42122 727456
rect 45002 727444 45008 727456
rect 42116 727416 45008 727444
rect 42116 727404 42122 727416
rect 45002 727404 45008 727416
rect 45060 727404 45066 727456
rect 40770 727268 40776 727320
rect 40828 727308 40834 727320
rect 41690 727308 41696 727320
rect 40828 727280 41696 727308
rect 40828 727268 40834 727280
rect 41690 727268 41696 727280
rect 41748 727268 41754 727320
rect 42058 727268 42064 727320
rect 42116 727308 42122 727320
rect 45370 727308 45376 727320
rect 42116 727280 45376 727308
rect 42116 727268 42122 727280
rect 45370 727268 45376 727280
rect 45428 727268 45434 727320
rect 674852 727274 674880 727472
rect 674852 727246 674972 727274
rect 674944 727240 674972 727246
rect 678238 727240 678244 727252
rect 674944 727212 678244 727240
rect 678238 727200 678244 727212
rect 678296 727200 678302 727252
rect 674650 726656 674656 726708
rect 674708 726696 674714 726708
rect 683298 726696 683304 726708
rect 674708 726668 683304 726696
rect 674708 726656 674714 726668
rect 683298 726656 683304 726668
rect 683356 726656 683362 726708
rect 674282 726520 674288 726572
rect 674340 726560 674346 726572
rect 684126 726560 684132 726572
rect 674340 726532 684132 726560
rect 674340 726520 674346 726532
rect 684126 726520 684132 726532
rect 684184 726520 684190 726572
rect 41322 726180 41328 726232
rect 41380 726220 41386 726232
rect 41690 726220 41696 726232
rect 41380 726192 41696 726220
rect 41380 726180 41386 726192
rect 41690 726180 41696 726192
rect 41748 726180 41754 726232
rect 41138 725908 41144 725960
rect 41196 725948 41202 725960
rect 41598 725948 41604 725960
rect 41196 725920 41604 725948
rect 41196 725908 41202 725920
rect 41598 725908 41604 725920
rect 41656 725908 41662 725960
rect 42058 725908 42064 725960
rect 42116 725948 42122 725960
rect 42702 725948 42708 725960
rect 42116 725920 42708 725948
rect 42116 725908 42122 725920
rect 42702 725908 42708 725920
rect 42760 725908 42766 725960
rect 673730 722168 673736 722220
rect 673788 722208 673794 722220
rect 673914 722208 673920 722220
rect 673788 722180 673920 722208
rect 673788 722168 673794 722180
rect 673914 722168 673920 722180
rect 673972 722168 673978 722220
rect 675110 721692 675116 721744
rect 675168 721692 675174 721744
rect 675294 721692 675300 721744
rect 675352 721692 675358 721744
rect 675128 721268 675156 721692
rect 675312 721268 675340 721692
rect 675110 721216 675116 721268
rect 675168 721216 675174 721268
rect 675294 721216 675300 721268
rect 675352 721216 675358 721268
rect 675110 720808 675116 720860
rect 675168 720808 675174 720860
rect 675294 720808 675300 720860
rect 675352 720808 675358 720860
rect 675128 720520 675156 720808
rect 675312 720520 675340 720808
rect 675110 720468 675116 720520
rect 675168 720468 675174 720520
rect 675294 720468 675300 720520
rect 675352 720468 675358 720520
rect 42058 718972 42064 719024
rect 42116 719012 42122 719024
rect 57238 719012 57244 719024
rect 42116 718984 57244 719012
rect 42116 718972 42122 718984
rect 57238 718972 57244 718984
rect 57296 718972 57302 719024
rect 42242 717204 42248 717256
rect 42300 717244 42306 717256
rect 42702 717244 42708 717256
rect 42300 717216 42708 717244
rect 42300 717204 42306 717216
rect 42702 717204 42708 717216
rect 42760 717204 42766 717256
rect 653398 716252 653404 716304
rect 653456 716292 653462 716304
rect 673822 716292 673828 716304
rect 653456 716264 673828 716292
rect 653456 716252 653462 716264
rect 673822 716252 673828 716264
rect 673880 716252 673886 716304
rect 672166 716116 672172 716168
rect 672224 716156 672230 716168
rect 673362 716156 673368 716168
rect 672224 716128 673368 716156
rect 672224 716116 672230 716128
rect 673362 716116 673368 716128
rect 673420 716116 673426 716168
rect 669958 715708 669964 715760
rect 670016 715748 670022 715760
rect 672810 715748 672816 715760
rect 670016 715720 672816 715748
rect 670016 715708 670022 715720
rect 672810 715708 672816 715720
rect 672868 715708 672874 715760
rect 35158 715640 35164 715692
rect 35216 715680 35222 715692
rect 35216 715652 41552 715680
rect 35216 715640 35222 715652
rect 33778 715504 33784 715556
rect 33836 715544 33842 715556
rect 40770 715544 40776 715556
rect 33836 715516 40776 715544
rect 33836 715504 33842 715516
rect 40770 715504 40776 715516
rect 40828 715504 40834 715556
rect 41524 715216 41552 715652
rect 41506 715164 41512 715216
rect 41564 715164 41570 715216
rect 660298 714960 660304 715012
rect 660356 715000 660362 715012
rect 673822 715000 673828 715012
rect 660356 714972 673828 715000
rect 660356 714960 660362 714972
rect 673822 714960 673828 714972
rect 673880 714960 673886 715012
rect 670142 714824 670148 714876
rect 670200 714864 670206 714876
rect 673362 714864 673368 714876
rect 670200 714836 673368 714864
rect 670200 714824 670206 714836
rect 673362 714824 673368 714836
rect 673420 714824 673426 714876
rect 671798 714008 671804 714060
rect 671856 714048 671862 714060
rect 673822 714048 673828 714060
rect 671856 714020 673828 714048
rect 671856 714008 671862 714020
rect 673822 714008 673828 714020
rect 673880 714008 673886 714060
rect 670970 713668 670976 713720
rect 671028 713708 671034 713720
rect 673822 713708 673828 713720
rect 671028 713680 673828 713708
rect 671028 713668 671034 713680
rect 673822 713668 673828 713680
rect 673880 713668 673886 713720
rect 671338 713192 671344 713244
rect 671396 713232 671402 713244
rect 673822 713232 673828 713244
rect 671396 713204 673828 713232
rect 671396 713192 671402 713204
rect 673822 713192 673828 713204
rect 673880 713192 673886 713244
rect 671982 712852 671988 712904
rect 672040 712892 672046 712904
rect 673822 712892 673828 712904
rect 672040 712864 673828 712892
rect 672040 712852 672046 712864
rect 673822 712852 673828 712864
rect 673880 712852 673886 712904
rect 671982 712376 671988 712428
rect 672040 712416 672046 712428
rect 673822 712416 673828 712428
rect 672040 712388 673828 712416
rect 672040 712376 672046 712388
rect 673822 712376 673828 712388
rect 673880 712376 673886 712428
rect 43622 712104 43628 712156
rect 43680 712144 43686 712156
rect 50338 712144 50344 712156
rect 43680 712116 50344 712144
rect 43680 712104 43686 712116
rect 50338 712104 50344 712116
rect 50396 712104 50402 712156
rect 669774 711628 669780 711680
rect 669832 711668 669838 711680
rect 673822 711668 673828 711680
rect 669832 711640 673828 711668
rect 669832 711628 669838 711640
rect 673822 711628 673828 711640
rect 673880 711628 673886 711680
rect 670786 709996 670792 710048
rect 670844 710036 670850 710048
rect 673822 710036 673828 710048
rect 670844 710008 673828 710036
rect 670844 709996 670850 710008
rect 673822 709996 673828 710008
rect 673880 709996 673886 710048
rect 670602 709588 670608 709640
rect 670660 709628 670666 709640
rect 673822 709628 673828 709640
rect 670660 709600 673828 709628
rect 670660 709588 670666 709600
rect 673822 709588 673828 709600
rect 673880 709588 673886 709640
rect 43622 709316 43628 709368
rect 43680 709356 43686 709368
rect 44450 709356 44456 709368
rect 43680 709328 44456 709356
rect 43680 709316 43686 709328
rect 44450 709316 44456 709328
rect 44508 709316 44514 709368
rect 674282 707956 674288 708008
rect 674340 707996 674346 708008
rect 676030 707996 676036 708008
rect 674340 707968 676036 707996
rect 674340 707956 674346 707968
rect 676030 707956 676036 707968
rect 676088 707956 676094 708008
rect 674466 705576 674472 705628
rect 674524 705616 674530 705628
rect 676030 705616 676036 705628
rect 674524 705588 676036 705616
rect 674524 705576 674530 705588
rect 676030 705576 676036 705588
rect 676088 705576 676094 705628
rect 42242 705508 42248 705560
rect 42300 705548 42306 705560
rect 43438 705548 43444 705560
rect 42300 705520 43444 705548
rect 42300 705508 42306 705520
rect 43438 705508 43444 705520
rect 43496 705508 43502 705560
rect 668394 705508 668400 705560
rect 668452 705548 668458 705560
rect 673362 705548 673368 705560
rect 668452 705520 673368 705548
rect 668452 705508 668458 705520
rect 673362 705508 673368 705520
rect 673420 705508 673426 705560
rect 674282 705304 674288 705356
rect 674340 705344 674346 705356
rect 683114 705344 683120 705356
rect 674340 705316 683120 705344
rect 674340 705304 674346 705316
rect 683114 705304 683120 705316
rect 683172 705304 683178 705356
rect 50338 705100 50344 705152
rect 50396 705140 50402 705152
rect 62114 705140 62120 705152
rect 50396 705112 62120 705140
rect 50396 705100 50402 705112
rect 62114 705100 62120 705112
rect 62172 705100 62178 705152
rect 674282 703876 674288 703928
rect 674340 703916 674346 703928
rect 676030 703916 676036 703928
rect 674340 703888 676036 703916
rect 674340 703876 674346 703888
rect 676030 703876 676036 703888
rect 676088 703876 676094 703928
rect 667842 703808 667848 703860
rect 667900 703848 667906 703860
rect 673178 703848 673184 703860
rect 667900 703820 673184 703848
rect 667900 703808 667906 703820
rect 673178 703808 673184 703820
rect 673236 703808 673242 703860
rect 44450 703740 44456 703792
rect 44508 703780 44514 703792
rect 62114 703780 62120 703792
rect 44508 703752 62120 703780
rect 44508 703740 44514 703752
rect 62114 703740 62120 703752
rect 62172 703740 62178 703792
rect 42242 702176 42248 702228
rect 42300 702176 42306 702228
rect 42260 701956 42288 702176
rect 42242 701904 42248 701956
rect 42300 701904 42306 701956
rect 654778 701156 654784 701208
rect 654836 701196 654842 701208
rect 673178 701196 673184 701208
rect 654836 701168 673184 701196
rect 654836 701156 654842 701168
rect 673178 701156 673184 701168
rect 673236 701156 673242 701208
rect 42702 701088 42708 701140
rect 42760 701128 42766 701140
rect 42760 701100 51074 701128
rect 42760 701088 42766 701100
rect 51046 701060 51074 701100
rect 62206 701060 62212 701072
rect 51046 701032 62212 701060
rect 62206 701020 62212 701032
rect 62264 701020 62270 701072
rect 666462 701020 666468 701072
rect 666520 701060 666526 701072
rect 672994 701060 673000 701072
rect 666520 701032 673000 701060
rect 666520 701020 666526 701032
rect 672994 701020 673000 701032
rect 673052 701020 673058 701072
rect 46198 698164 46204 698216
rect 46256 698204 46262 698216
rect 62114 698204 62120 698216
rect 46256 698176 62120 698204
rect 46256 698164 46262 698176
rect 62114 698164 62120 698176
rect 62172 698164 62178 698216
rect 656802 690004 656808 690056
rect 656860 690044 656866 690056
rect 673178 690044 673184 690056
rect 656860 690016 673184 690044
rect 656860 690004 656866 690016
rect 673178 690004 673184 690016
rect 673236 690004 673242 690056
rect 652754 688780 652760 688832
rect 652812 688820 652818 688832
rect 673178 688820 673184 688832
rect 652812 688792 673184 688820
rect 652812 688780 652818 688792
rect 673178 688780 673184 688792
rect 673236 688780 673242 688832
rect 651466 688644 651472 688696
rect 651524 688684 651530 688696
rect 657538 688684 657544 688696
rect 651524 688656 657544 688684
rect 651524 688644 651530 688656
rect 657538 688644 657544 688656
rect 657596 688644 657602 688696
rect 42702 687284 42708 687336
rect 42760 687324 42766 687336
rect 42760 687296 51074 687324
rect 42760 687284 42766 687296
rect 51046 687256 51074 687296
rect 61378 687256 61384 687268
rect 51046 687228 61384 687256
rect 61378 687216 61384 687228
rect 61436 687216 61442 687268
rect 651466 687216 651472 687268
rect 651524 687256 651530 687268
rect 669958 687256 669964 687268
rect 651524 687228 669964 687256
rect 651524 687216 651530 687228
rect 669958 687216 669964 687228
rect 670016 687216 670022 687268
rect 675110 687256 675116 687268
rect 674484 687228 675116 687256
rect 674484 687132 674512 687228
rect 675110 687216 675116 687228
rect 675168 687216 675174 687268
rect 674466 687080 674472 687132
rect 674524 687080 674530 687132
rect 651466 687012 651472 687064
rect 651524 687052 651530 687064
rect 654778 687052 654784 687064
rect 651524 687024 654784 687052
rect 651524 687012 651530 687024
rect 654778 687012 654784 687024
rect 654836 687012 654842 687064
rect 43438 686468 43444 686520
rect 43496 686508 43502 686520
rect 62758 686508 62764 686520
rect 43496 686480 62764 686508
rect 43496 686468 43502 686480
rect 62758 686468 62764 686480
rect 62816 686468 62822 686520
rect 651650 686468 651656 686520
rect 651708 686508 651714 686520
rect 667198 686508 667204 686520
rect 651708 686480 667204 686508
rect 651708 686468 651714 686480
rect 667198 686468 667204 686480
rect 667256 686468 667262 686520
rect 41138 685992 41144 686044
rect 41196 686032 41202 686044
rect 41690 686032 41696 686044
rect 41196 686004 41696 686032
rect 41196 685992 41202 686004
rect 41690 685992 41696 686004
rect 41748 685992 41754 686044
rect 42058 685992 42064 686044
rect 42116 686032 42122 686044
rect 45370 686032 45376 686044
rect 42116 686004 45376 686032
rect 42116 685992 42122 686004
rect 45370 685992 45376 686004
rect 45428 685992 45434 686044
rect 668210 685924 668216 685976
rect 668268 685964 668274 685976
rect 673638 685964 673644 685976
rect 668268 685936 673644 685964
rect 668268 685924 668274 685936
rect 673638 685924 673644 685936
rect 673696 685924 673702 685976
rect 40862 685856 40868 685908
rect 40920 685896 40926 685908
rect 41690 685896 41696 685908
rect 40920 685868 41696 685896
rect 40920 685856 40926 685868
rect 41690 685856 41696 685868
rect 41748 685856 41754 685908
rect 42058 685856 42064 685908
rect 42116 685896 42122 685908
rect 45186 685896 45192 685908
rect 42116 685868 45192 685896
rect 42116 685856 42122 685868
rect 45186 685856 45192 685868
rect 45244 685856 45250 685908
rect 651466 685516 651472 685568
rect 651524 685556 651530 685568
rect 656802 685556 656808 685568
rect 651524 685528 656808 685556
rect 651524 685516 651530 685528
rect 656802 685516 656808 685528
rect 656860 685516 656866 685568
rect 41322 683408 41328 683460
rect 41380 683448 41386 683460
rect 41690 683448 41696 683460
rect 41380 683420 41696 683448
rect 41380 683408 41386 683420
rect 41690 683408 41696 683420
rect 41748 683408 41754 683460
rect 41046 682932 41052 682984
rect 41104 682972 41110 682984
rect 41690 682972 41696 682984
rect 41104 682944 41696 682972
rect 41104 682932 41110 682944
rect 41690 682932 41696 682944
rect 41748 682932 41754 682984
rect 674650 682388 674656 682440
rect 674708 682428 674714 682440
rect 683206 682428 683212 682440
rect 674708 682400 683212 682428
rect 674708 682388 674714 682400
rect 683206 682388 683212 682400
rect 683264 682388 683270 682440
rect 41138 676200 41144 676252
rect 41196 676240 41202 676252
rect 41690 676240 41696 676252
rect 41196 676212 41696 676240
rect 41196 676200 41202 676212
rect 41690 676200 41696 676212
rect 41748 676200 41754 676252
rect 42058 676200 42064 676252
rect 42116 676240 42122 676252
rect 55858 676240 55864 676252
rect 42116 676212 55864 676240
rect 42116 676200 42122 676212
rect 55858 676200 55864 676212
rect 55916 676200 55922 676252
rect 31662 674092 31668 674144
rect 31720 674132 31726 674144
rect 41506 674132 41512 674144
rect 31720 674104 41512 674132
rect 31720 674092 31726 674104
rect 41506 674092 41512 674104
rect 41564 674092 41570 674144
rect 35158 672732 35164 672784
rect 35216 672772 35222 672784
rect 41690 672772 41696 672784
rect 35216 672744 41696 672772
rect 35216 672732 35222 672744
rect 41690 672732 41696 672744
rect 41748 672732 41754 672784
rect 42058 672664 42064 672716
rect 42116 672704 42122 672716
rect 42518 672704 42524 672716
rect 42116 672676 42524 672704
rect 42116 672664 42122 672676
rect 42518 672664 42524 672676
rect 42576 672664 42582 672716
rect 33778 671304 33784 671356
rect 33836 671344 33842 671356
rect 41690 671344 41696 671356
rect 33836 671316 41696 671344
rect 33836 671304 33842 671316
rect 41690 671304 41696 671316
rect 41748 671304 41754 671356
rect 673730 671304 673736 671356
rect 673788 671344 673794 671356
rect 673788 671316 673960 671344
rect 673788 671304 673794 671316
rect 668026 671100 668032 671152
rect 668084 671140 668090 671152
rect 673730 671140 673736 671152
rect 668084 671112 673736 671140
rect 668084 671100 668090 671112
rect 673730 671100 673736 671112
rect 673788 671100 673794 671152
rect 661678 670692 661684 670744
rect 661736 670732 661742 670744
rect 673932 670732 673960 671316
rect 661736 670704 673960 670732
rect 661736 670692 661742 670704
rect 670142 670148 670148 670200
rect 670200 670188 670206 670200
rect 672166 670188 672172 670200
rect 670200 670160 672172 670188
rect 670200 670148 670206 670160
rect 672166 670148 672172 670160
rect 672224 670148 672230 670200
rect 670142 669672 670148 669724
rect 670200 669712 670206 669724
rect 672166 669712 672172 669724
rect 670200 669684 672172 669712
rect 670200 669672 670206 669684
rect 672166 669672 672172 669684
rect 672224 669672 672230 669724
rect 673546 669576 673552 669588
rect 663766 669548 673552 669576
rect 658918 669468 658924 669520
rect 658976 669508 658982 669520
rect 663766 669508 663794 669548
rect 673546 669536 673552 669548
rect 673604 669536 673610 669588
rect 658976 669480 663794 669508
rect 658976 669468 658982 669480
rect 42334 669332 42340 669384
rect 42392 669372 42398 669384
rect 53098 669372 53104 669384
rect 42392 669344 53104 669372
rect 42392 669332 42398 669344
rect 53098 669332 53104 669344
rect 53156 669332 53162 669384
rect 671798 669332 671804 669384
rect 671856 669372 671862 669384
rect 671856 669344 673776 669372
rect 671856 669332 671862 669344
rect 673546 669196 673552 669248
rect 673604 669236 673610 669248
rect 673748 669236 673776 669344
rect 673604 669208 673776 669236
rect 673604 669196 673610 669208
rect 669774 668652 669780 668704
rect 669832 668692 669838 668704
rect 673546 668692 673552 668704
rect 669832 668664 673552 668692
rect 669832 668652 669838 668664
rect 673546 668652 673552 668664
rect 673604 668652 673610 668704
rect 671338 668244 671344 668296
rect 671396 668284 671402 668296
rect 673546 668284 673552 668296
rect 671396 668256 673552 668284
rect 671396 668244 671402 668256
rect 673546 668244 673552 668256
rect 673604 668244 673610 668296
rect 59998 667944 60004 667956
rect 42260 667916 60004 667944
rect 42260 667276 42288 667916
rect 59998 667904 60004 667916
rect 60056 667904 60062 667956
rect 671430 667904 671436 667956
rect 671488 667944 671494 667956
rect 673546 667944 673552 667956
rect 671488 667916 673552 667944
rect 671488 667904 671494 667916
rect 673546 667904 673552 667916
rect 673604 667904 673610 667956
rect 675202 667836 675208 667888
rect 675260 667876 675266 667888
rect 676030 667876 676036 667888
rect 675260 667848 676036 667876
rect 675260 667836 675266 667848
rect 676030 667836 676036 667848
rect 676088 667836 676094 667888
rect 42242 667224 42248 667276
rect 42300 667224 42306 667276
rect 671982 666884 671988 666936
rect 672040 666924 672046 666936
rect 673546 666924 673552 666936
rect 672040 666896 673552 666924
rect 672040 666884 672046 666896
rect 673546 666884 673552 666896
rect 673604 666884 673610 666936
rect 671798 666680 671804 666732
rect 671856 666720 671862 666732
rect 673546 666720 673552 666732
rect 671856 666692 673552 666720
rect 671856 666680 671862 666692
rect 673546 666680 673552 666692
rect 673604 666680 673610 666732
rect 671154 665660 671160 665712
rect 671212 665700 671218 665712
rect 673546 665700 673552 665712
rect 671212 665672 673552 665700
rect 671212 665660 671218 665672
rect 673546 665660 673552 665672
rect 673604 665660 673610 665712
rect 42334 665388 42340 665440
rect 42392 665428 42398 665440
rect 43622 665428 43628 665440
rect 42392 665400 43628 665428
rect 42392 665388 42398 665400
rect 43622 665388 43628 665400
rect 43680 665388 43686 665440
rect 671246 665320 671252 665372
rect 671304 665360 671310 665372
rect 671798 665360 671804 665372
rect 671304 665332 671804 665360
rect 671304 665320 671310 665332
rect 671798 665320 671804 665332
rect 671856 665320 671862 665372
rect 669590 665184 669596 665236
rect 669648 665224 669654 665236
rect 673546 665224 673552 665236
rect 669648 665196 673552 665224
rect 669648 665184 669654 665196
rect 673546 665184 673552 665196
rect 673604 665184 673610 665236
rect 670326 664300 670332 664352
rect 670384 664340 670390 664352
rect 673546 664340 673552 664352
rect 670384 664312 673552 664340
rect 670384 664300 670390 664312
rect 673546 664300 673552 664312
rect 673604 664300 673610 664352
rect 674834 663892 674840 663944
rect 674892 663932 674898 663944
rect 676214 663932 676220 663944
rect 674892 663904 676220 663932
rect 674892 663892 674898 663904
rect 676214 663892 676220 663904
rect 676272 663892 676278 663944
rect 42426 663824 42432 663876
rect 42484 663824 42490 663876
rect 42444 663060 42472 663824
rect 669222 663756 669228 663808
rect 669280 663796 669286 663808
rect 673546 663796 673552 663808
rect 669280 663768 673552 663796
rect 669280 663756 669286 663768
rect 673546 663756 673552 663768
rect 673604 663756 673610 663808
rect 673546 663348 673552 663400
rect 673604 663388 673610 663400
rect 673914 663388 673920 663400
rect 673604 663360 673920 663388
rect 673604 663348 673610 663360
rect 673914 663348 673920 663360
rect 673972 663348 673978 663400
rect 42426 663008 42432 663060
rect 42484 663008 42490 663060
rect 674650 662940 674656 662992
rect 674708 662980 674714 662992
rect 676214 662980 676220 662992
rect 674708 662952 676220 662980
rect 674708 662940 674714 662952
rect 676214 662940 676220 662952
rect 676272 662940 676278 662992
rect 668670 662736 668676 662788
rect 668728 662776 668734 662788
rect 673914 662776 673920 662788
rect 668728 662748 673920 662776
rect 668728 662736 668734 662748
rect 673914 662736 673920 662748
rect 673972 662736 673978 662788
rect 671614 661512 671620 661564
rect 671672 661552 671678 661564
rect 673914 661552 673920 661564
rect 671672 661524 673920 661552
rect 671672 661512 671678 661524
rect 673914 661512 673920 661524
rect 673972 661512 673978 661564
rect 669222 661104 669228 661156
rect 669280 661144 669286 661156
rect 673914 661144 673920 661156
rect 669280 661116 673920 661144
rect 669280 661104 669286 661116
rect 673914 661104 673920 661116
rect 673972 661104 673978 661156
rect 53098 660900 53104 660952
rect 53156 660940 53162 660952
rect 62114 660940 62120 660952
rect 53156 660912 62120 660940
rect 53156 660900 53162 660912
rect 62114 660900 62120 660912
rect 62172 660900 62178 660952
rect 42150 660492 42156 660544
rect 42208 660532 42214 660544
rect 43070 660532 43076 660544
rect 42208 660504 43076 660532
rect 42208 660492 42214 660504
rect 43070 660492 43076 660504
rect 43128 660492 43134 660544
rect 668946 660084 668952 660136
rect 669004 660124 669010 660136
rect 673914 660124 673920 660136
rect 669004 660096 673920 660124
rect 669004 660084 669010 660096
rect 673914 660084 673920 660096
rect 673972 660084 673978 660136
rect 674650 659812 674656 659864
rect 674708 659852 674714 659864
rect 683114 659852 683120 659864
rect 674708 659824 683120 659852
rect 674708 659812 674714 659824
rect 683114 659812 683120 659824
rect 683172 659812 683178 659864
rect 59998 659540 60004 659592
rect 60056 659580 60062 659592
rect 62114 659580 62120 659592
rect 60056 659552 62120 659580
rect 60056 659540 60062 659552
rect 62114 659540 62120 659552
rect 62172 659540 62178 659592
rect 62114 657540 62120 657552
rect 45526 657512 62120 657540
rect 42518 657364 42524 657416
rect 42576 657404 42582 657416
rect 45526 657404 45554 657512
rect 62114 657500 62120 657512
rect 62172 657500 62178 657552
rect 42576 657376 45554 657404
rect 42576 657364 42582 657376
rect 653398 655528 653404 655580
rect 653456 655568 653462 655580
rect 673914 655568 673920 655580
rect 653456 655540 673920 655568
rect 653456 655528 653462 655540
rect 673914 655528 673920 655540
rect 673972 655528 673978 655580
rect 44818 655460 44824 655512
rect 44876 655500 44882 655512
rect 62114 655500 62120 655512
rect 44876 655472 62120 655500
rect 44876 655460 44882 655472
rect 62114 655460 62120 655472
rect 62172 655460 62178 655512
rect 667014 647300 667020 647352
rect 667072 647340 667078 647352
rect 674006 647340 674012 647352
rect 667072 647312 674012 647340
rect 667072 647300 667078 647312
rect 674006 647300 674012 647312
rect 674064 647300 674070 647352
rect 655514 645872 655520 645924
rect 655572 645912 655578 645924
rect 674006 645912 674012 645924
rect 655572 645884 674012 645912
rect 655572 645872 655578 645884
rect 674006 645872 674012 645884
rect 674064 645872 674070 645924
rect 35802 644444 35808 644496
rect 35860 644484 35866 644496
rect 41690 644484 41696 644496
rect 35860 644456 41696 644484
rect 35860 644444 35866 644456
rect 41690 644444 41696 644456
rect 41748 644444 41754 644496
rect 42058 644444 42064 644496
rect 42116 644484 42122 644496
rect 54478 644484 54484 644496
rect 42116 644456 54484 644484
rect 42116 644444 42122 644456
rect 54478 644444 54484 644456
rect 54536 644444 54542 644496
rect 35802 643492 35808 643544
rect 35860 643532 35866 643544
rect 40494 643532 40500 643544
rect 35860 643504 40500 643532
rect 35860 643492 35866 643504
rect 40494 643492 40500 643504
rect 40552 643492 40558 643544
rect 41690 643328 41696 643340
rect 41386 643300 41696 643328
rect 35526 643220 35532 643272
rect 35584 643260 35590 643272
rect 41386 643260 41414 643300
rect 41690 643288 41696 643300
rect 41748 643288 41754 643340
rect 42058 643288 42064 643340
rect 42116 643328 42122 643340
rect 45370 643328 45376 643340
rect 42116 643300 45376 643328
rect 42116 643288 42122 643300
rect 45370 643288 45376 643300
rect 45428 643288 45434 643340
rect 35584 643232 41414 643260
rect 35584 643220 35590 643232
rect 35342 643084 35348 643136
rect 35400 643124 35406 643136
rect 41690 643124 41696 643136
rect 35400 643096 41696 643124
rect 35400 643084 35406 643096
rect 41690 643084 41696 643096
rect 41748 643084 41754 643136
rect 42058 643084 42064 643136
rect 42116 643124 42122 643136
rect 61378 643124 61384 643136
rect 42116 643096 61384 643124
rect 42116 643084 42122 643096
rect 61378 643084 61384 643096
rect 61436 643084 61442 643136
rect 655330 643084 655336 643136
rect 655388 643124 655394 643136
rect 674006 643124 674012 643136
rect 655388 643096 674012 643124
rect 655388 643084 655394 643096
rect 674006 643084 674012 643096
rect 674064 643084 674070 643136
rect 38562 642472 38568 642524
rect 38620 642512 38626 642524
rect 41690 642512 41696 642524
rect 38620 642484 41696 642512
rect 38620 642472 38626 642484
rect 41690 642472 41696 642484
rect 41748 642472 41754 642524
rect 42058 642336 42064 642388
rect 42116 642376 42122 642388
rect 62942 642376 62948 642388
rect 42116 642348 62948 642376
rect 42116 642336 42122 642348
rect 62942 642336 62948 642348
rect 63000 642336 63006 642388
rect 651466 642336 651472 642388
rect 651524 642376 651530 642388
rect 660298 642376 660304 642388
rect 651524 642348 660304 642376
rect 651524 642336 651530 642348
rect 660298 642336 660304 642348
rect 660356 642336 660362 642388
rect 35618 641996 35624 642048
rect 35676 642036 35682 642048
rect 39482 642036 39488 642048
rect 35676 642008 39488 642036
rect 35676 641996 35682 642008
rect 39482 641996 39488 642008
rect 39540 641996 39546 642048
rect 35802 641724 35808 641776
rect 35860 641764 35866 641776
rect 41690 641764 41696 641776
rect 35860 641736 41696 641764
rect 35860 641724 35866 641736
rect 41690 641724 41696 641736
rect 41748 641724 41754 641776
rect 42058 641724 42064 641776
rect 42116 641764 42122 641776
rect 44634 641764 44640 641776
rect 42116 641736 44640 641764
rect 42116 641724 42122 641736
rect 44634 641724 44640 641736
rect 44692 641724 44698 641776
rect 35802 640772 35808 640824
rect 35860 640812 35866 640824
rect 35860 640772 35894 640812
rect 35866 640744 35894 640772
rect 39574 640744 39580 640756
rect 35866 640716 39580 640744
rect 39574 640704 39580 640716
rect 39632 640704 39638 640756
rect 35802 640432 35808 640484
rect 35860 640472 35866 640484
rect 39942 640472 39948 640484
rect 35860 640444 39948 640472
rect 35860 640432 35866 640444
rect 39942 640432 39948 640444
rect 40000 640432 40006 640484
rect 35618 640296 35624 640348
rect 35676 640336 35682 640348
rect 41690 640336 41696 640348
rect 35676 640308 41696 640336
rect 35676 640296 35682 640308
rect 41690 640296 41696 640308
rect 41748 640296 41754 640348
rect 42058 640296 42064 640348
rect 42116 640336 42122 640348
rect 45370 640336 45376 640348
rect 42116 640308 45376 640336
rect 42116 640296 42122 640308
rect 45370 640296 45376 640308
rect 45428 640296 45434 640348
rect 651466 640296 651472 640348
rect 651524 640336 651530 640348
rect 668578 640336 668584 640348
rect 651524 640308 668584 640336
rect 651524 640296 651530 640308
rect 668578 640296 668584 640308
rect 668636 640296 668642 640348
rect 651374 640092 651380 640144
rect 651432 640132 651438 640144
rect 653398 640132 653404 640144
rect 651432 640104 653404 640132
rect 651432 640092 651438 640104
rect 653398 640092 653404 640104
rect 653456 640092 653462 640144
rect 35802 639072 35808 639124
rect 35860 639112 35866 639124
rect 41690 639112 41696 639124
rect 35860 639084 41696 639112
rect 35860 639072 35866 639084
rect 41690 639072 41696 639084
rect 41748 639072 41754 639124
rect 35526 638936 35532 638988
rect 35584 638976 35590 638988
rect 37918 638976 37924 638988
rect 35584 638948 37924 638976
rect 35584 638936 35590 638948
rect 37918 638936 37924 638948
rect 37976 638936 37982 638988
rect 651650 638868 651656 638920
rect 651708 638908 651714 638920
rect 655330 638908 655336 638920
rect 651708 638880 655336 638908
rect 651708 638868 651714 638880
rect 655330 638868 655336 638880
rect 655388 638868 655394 638920
rect 651466 638732 651472 638784
rect 651524 638772 651530 638784
rect 655514 638772 655520 638784
rect 651524 638744 655520 638772
rect 651524 638732 651530 638744
rect 655514 638732 655520 638744
rect 655572 638732 655578 638784
rect 35342 638188 35348 638240
rect 35400 638228 35406 638240
rect 41690 638228 41696 638240
rect 35400 638200 41696 638228
rect 35400 638188 35406 638200
rect 41690 638188 41696 638200
rect 41748 638188 41754 638240
rect 35802 637576 35808 637628
rect 35860 637616 35866 637628
rect 36538 637616 36544 637628
rect 35860 637588 36544 637616
rect 35860 637576 35866 637588
rect 36538 637576 36544 637588
rect 36596 637576 36602 637628
rect 672350 637372 672356 637424
rect 672408 637412 672414 637424
rect 672810 637412 672816 637424
rect 672408 637384 672816 637412
rect 672408 637372 672414 637384
rect 672810 637372 672816 637384
rect 672868 637372 672874 637424
rect 35618 637168 35624 637220
rect 35676 637208 35682 637220
rect 35676 637180 35894 637208
rect 35676 637168 35682 637180
rect 35866 636936 35894 637180
rect 675478 636964 675484 637016
rect 675536 637004 675542 637016
rect 683298 637004 683304 637016
rect 675536 636976 683304 637004
rect 675536 636964 675542 636976
rect 683298 636964 683304 636976
rect 683356 636964 683362 637016
rect 40402 636936 40408 636948
rect 35866 636908 40408 636936
rect 40402 636896 40408 636908
rect 40460 636896 40466 636948
rect 674374 636828 674380 636880
rect 674432 636868 674438 636880
rect 683942 636868 683948 636880
rect 674432 636840 683948 636868
rect 674432 636828 674438 636840
rect 683942 636828 683948 636840
rect 684000 636828 684006 636880
rect 674282 636692 674288 636744
rect 674340 636732 674346 636744
rect 675478 636732 675484 636744
rect 674340 636704 675484 636732
rect 674340 636692 674346 636704
rect 675478 636692 675484 636704
rect 675536 636692 675542 636744
rect 35618 636488 35624 636540
rect 35676 636528 35682 636540
rect 39850 636528 39856 636540
rect 35676 636500 39856 636528
rect 35676 636488 35682 636500
rect 39850 636488 39856 636500
rect 39908 636488 39914 636540
rect 35802 636216 35808 636268
rect 35860 636256 35866 636268
rect 35860 636228 38654 636256
rect 35860 636216 35866 636228
rect 38626 636188 38654 636228
rect 39022 636188 39028 636200
rect 38626 636160 39028 636188
rect 39022 636148 39028 636160
rect 39080 636148 39086 636200
rect 675110 635468 675116 635520
rect 675168 635508 675174 635520
rect 675478 635508 675484 635520
rect 675168 635480 675484 635508
rect 675168 635468 675174 635480
rect 675478 635468 675484 635480
rect 675536 635468 675542 635520
rect 35802 634924 35808 634976
rect 35860 634964 35866 634976
rect 39482 634964 39488 634976
rect 35860 634936 39488 634964
rect 35860 634924 35866 634936
rect 39482 634924 39488 634936
rect 39540 634924 39546 634976
rect 35802 633836 35808 633888
rect 35860 633876 35866 633888
rect 40126 633876 40132 633888
rect 35860 633848 40132 633876
rect 35860 633836 35866 633848
rect 40126 633836 40132 633848
rect 40184 633836 40190 633888
rect 39758 633672 39764 633684
rect 36004 633644 39764 633672
rect 35802 633564 35808 633616
rect 35860 633604 35866 633616
rect 36004 633604 36032 633644
rect 39758 633632 39764 633644
rect 39816 633632 39822 633684
rect 35860 633576 36032 633604
rect 35860 633564 35866 633576
rect 35618 633428 35624 633480
rect 35676 633468 35682 633480
rect 41598 633468 41604 633480
rect 35676 633440 41604 633468
rect 35676 633428 35682 633440
rect 41598 633428 41604 633440
rect 41656 633428 41662 633480
rect 42058 633428 42064 633480
rect 42116 633468 42122 633480
rect 63402 633468 63408 633480
rect 42116 633440 63408 633468
rect 42116 633428 42122 633440
rect 63402 633428 63408 633440
rect 63460 633428 63466 633480
rect 672350 632680 672356 632732
rect 672408 632720 672414 632732
rect 672718 632720 672724 632732
rect 672408 632692 672724 632720
rect 672408 632680 672414 632692
rect 672718 632680 672724 632692
rect 672776 632680 672782 632732
rect 36538 630572 36544 630624
rect 36596 630612 36602 630624
rect 41598 630612 41604 630624
rect 36596 630584 41604 630612
rect 36596 630572 36602 630584
rect 41598 630572 41604 630584
rect 41656 630572 41662 630624
rect 35158 628668 35164 628720
rect 35216 628708 35222 628720
rect 40494 628708 40500 628720
rect 35216 628680 40500 628708
rect 35216 628668 35222 628680
rect 40494 628668 40500 628680
rect 40552 628668 40558 628720
rect 673546 627648 673552 627700
rect 673604 627688 673610 627700
rect 673914 627688 673920 627700
rect 673604 627660 673920 627688
rect 673604 627648 673610 627660
rect 673914 627648 673920 627660
rect 673972 627648 673978 627700
rect 674282 626220 674288 626272
rect 674340 626260 674346 626272
rect 674834 626260 674840 626272
rect 674340 626232 674840 626260
rect 674340 626220 674346 626232
rect 674834 626220 674840 626232
rect 674892 626220 674898 626272
rect 674282 626016 674288 626068
rect 674340 626056 674346 626068
rect 676214 626056 676220 626068
rect 674340 626028 676220 626056
rect 674340 626016 674346 626028
rect 676214 626016 676220 626028
rect 676272 626016 676278 626068
rect 44450 625812 44456 625864
rect 44508 625852 44514 625864
rect 63126 625852 63132 625864
rect 44508 625824 63132 625852
rect 44508 625812 44514 625824
rect 63126 625812 63132 625824
rect 63184 625812 63190 625864
rect 667198 625608 667204 625660
rect 667256 625648 667262 625660
rect 674006 625648 674012 625660
rect 667256 625620 674012 625648
rect 667256 625608 667262 625620
rect 674006 625608 674012 625620
rect 674064 625608 674070 625660
rect 674282 625608 674288 625660
rect 674340 625648 674346 625660
rect 676214 625648 676220 625660
rect 674340 625620 676220 625648
rect 674340 625608 674346 625620
rect 676214 625608 676220 625620
rect 676272 625608 676278 625660
rect 674006 625376 674012 625388
rect 663766 625348 674012 625376
rect 657538 625268 657544 625320
rect 657596 625308 657602 625320
rect 663766 625308 663794 625348
rect 674006 625336 674012 625348
rect 674064 625336 674070 625388
rect 657596 625280 663794 625308
rect 657596 625268 657602 625280
rect 669958 625200 669964 625252
rect 670016 625240 670022 625252
rect 674006 625240 674012 625252
rect 670016 625212 674012 625240
rect 670016 625200 670022 625212
rect 674006 625200 674012 625212
rect 674064 625200 674070 625252
rect 674282 625200 674288 625252
rect 674340 625240 674346 625252
rect 676214 625240 676220 625252
rect 674340 625212 676220 625240
rect 674340 625200 674346 625212
rect 676214 625200 676220 625212
rect 676272 625200 676278 625252
rect 670234 625064 670240 625116
rect 670292 625104 670298 625116
rect 674006 625104 674012 625116
rect 670292 625076 674012 625104
rect 670292 625064 670298 625076
rect 674006 625064 674012 625076
rect 674064 625064 674070 625116
rect 674282 625064 674288 625116
rect 674340 625104 674346 625116
rect 676490 625104 676496 625116
rect 674340 625076 676496 625104
rect 674340 625064 674346 625076
rect 676490 625064 676496 625076
rect 676548 625064 676554 625116
rect 669774 624588 669780 624640
rect 669832 624628 669838 624640
rect 674006 624628 674012 624640
rect 669832 624600 674012 624628
rect 669832 624588 669838 624600
rect 674006 624588 674012 624600
rect 674064 624588 674070 624640
rect 674282 624452 674288 624504
rect 674340 624492 674346 624504
rect 676214 624492 676220 624504
rect 674340 624464 676220 624492
rect 674340 624452 674346 624464
rect 676214 624452 676220 624464
rect 676272 624452 676278 624504
rect 674282 624316 674288 624368
rect 674340 624356 674346 624368
rect 676030 624356 676036 624368
rect 674340 624328 676036 624356
rect 674340 624316 674346 624328
rect 676030 624316 676036 624328
rect 676088 624316 676094 624368
rect 669866 624248 669872 624300
rect 669924 624288 669930 624300
rect 674006 624288 674012 624300
rect 669924 624260 674012 624288
rect 669924 624248 669930 624260
rect 674006 624248 674012 624260
rect 674064 624248 674070 624300
rect 670234 623840 670240 623892
rect 670292 623880 670298 623892
rect 674006 623880 674012 623892
rect 670292 623852 674012 623880
rect 670292 623840 670298 623852
rect 674006 623840 674012 623852
rect 674064 623840 674070 623892
rect 671430 623636 671436 623688
rect 671488 623676 671494 623688
rect 674006 623676 674012 623688
rect 671488 623648 674012 623676
rect 671488 623636 671494 623648
rect 674006 623636 674012 623648
rect 674064 623636 674070 623688
rect 674282 623568 674288 623620
rect 674340 623608 674346 623620
rect 676214 623608 676220 623620
rect 674340 623580 676220 623608
rect 674340 623568 674346 623580
rect 676214 623568 676220 623580
rect 676272 623568 676278 623620
rect 670050 623024 670056 623076
rect 670108 623064 670114 623076
rect 674006 623064 674012 623076
rect 670108 623036 674012 623064
rect 670108 623024 670114 623036
rect 674006 623024 674012 623036
rect 674064 623024 674070 623076
rect 671246 622820 671252 622872
rect 671304 622860 671310 622872
rect 674006 622860 674012 622872
rect 671304 622832 674012 622860
rect 671304 622820 671310 622832
rect 674006 622820 674012 622832
rect 674064 622820 674070 622872
rect 674282 622820 674288 622872
rect 674340 622860 674346 622872
rect 676214 622860 676220 622872
rect 674340 622832 676220 622860
rect 674340 622820 674346 622832
rect 676214 622820 676220 622832
rect 676272 622820 676278 622872
rect 671430 622208 671436 622260
rect 671488 622248 671494 622260
rect 674006 622248 674012 622260
rect 671488 622220 674012 622248
rect 671488 622208 671494 622220
rect 674006 622208 674012 622220
rect 674064 622208 674070 622260
rect 42242 621664 42248 621716
rect 42300 621704 42306 621716
rect 44542 621704 44548 621716
rect 42300 621676 44548 621704
rect 42300 621664 42306 621676
rect 44542 621664 44548 621676
rect 44600 621664 44606 621716
rect 674282 621188 674288 621240
rect 674340 621228 674346 621240
rect 676214 621228 676220 621240
rect 674340 621200 676220 621228
rect 674340 621188 674346 621200
rect 676214 621188 676220 621200
rect 676272 621188 676278 621240
rect 666462 621120 666468 621172
rect 666520 621160 666526 621172
rect 674006 621160 674012 621172
rect 666520 621132 674012 621160
rect 666520 621120 666526 621132
rect 674006 621120 674012 621132
rect 674064 621120 674070 621172
rect 670602 620780 670608 620832
rect 670660 620820 670666 620832
rect 674006 620820 674012 620832
rect 670660 620792 674012 620820
rect 670660 620780 670666 620792
rect 674006 620780 674012 620792
rect 674064 620780 674070 620832
rect 674282 620780 674288 620832
rect 674340 620820 674346 620832
rect 676214 620820 676220 620832
rect 674340 620792 676220 620820
rect 674340 620780 674346 620792
rect 676214 620780 676220 620792
rect 676272 620780 676278 620832
rect 42242 620372 42248 620424
rect 42300 620412 42306 620424
rect 42702 620412 42708 620424
rect 42300 620384 42708 620412
rect 42300 620372 42306 620384
rect 42702 620372 42708 620384
rect 42760 620372 42766 620424
rect 674834 620168 674840 620220
rect 674892 620208 674898 620220
rect 683114 620208 683120 620220
rect 674892 620180 683120 620208
rect 674892 620168 674898 620180
rect 683114 620168 683120 620180
rect 683172 620168 683178 620220
rect 674282 619760 674288 619812
rect 674340 619800 674346 619812
rect 676030 619800 676036 619812
rect 674340 619772 676036 619800
rect 674340 619760 674346 619772
rect 676030 619760 676036 619772
rect 676088 619760 676094 619812
rect 668210 619692 668216 619744
rect 668268 619732 668274 619744
rect 674006 619732 674012 619744
rect 668268 619704 674012 619732
rect 668268 619692 668274 619704
rect 674006 619692 674012 619704
rect 674064 619692 674070 619744
rect 42242 619624 42248 619676
rect 42300 619664 42306 619676
rect 44266 619664 44272 619676
rect 42300 619636 44272 619664
rect 42300 619624 42306 619636
rect 44266 619624 44272 619636
rect 44324 619624 44330 619676
rect 673178 619284 673184 619336
rect 673236 619324 673242 619336
rect 674006 619324 674012 619336
rect 673236 619296 674012 619324
rect 673236 619284 673242 619296
rect 674006 619284 674012 619296
rect 674064 619284 674070 619336
rect 674282 619148 674288 619200
rect 674340 619188 674346 619200
rect 676490 619188 676496 619200
rect 674340 619160 676496 619188
rect 674340 619148 674346 619160
rect 676490 619148 676496 619160
rect 676548 619148 676554 619200
rect 674282 618332 674288 618384
rect 674340 618372 674346 618384
rect 676214 618372 676220 618384
rect 674340 618344 676220 618372
rect 674340 618332 674346 618344
rect 676214 618332 676220 618344
rect 676272 618332 676278 618384
rect 668394 618264 668400 618316
rect 668452 618304 668458 618316
rect 674006 618304 674012 618316
rect 668452 618276 674012 618304
rect 668452 618264 668458 618276
rect 674006 618264 674012 618276
rect 674064 618264 674070 618316
rect 674466 618196 674472 618248
rect 674524 618236 674530 618248
rect 676030 618236 676036 618248
rect 674524 618208 676036 618236
rect 674524 618196 674530 618208
rect 676030 618196 676036 618208
rect 676088 618196 676094 618248
rect 670970 618060 670976 618112
rect 671028 618100 671034 618112
rect 674006 618100 674012 618112
rect 671028 618072 674012 618100
rect 671028 618060 671034 618072
rect 674006 618060 674012 618072
rect 674064 618060 674070 618112
rect 674282 617924 674288 617976
rect 674340 617964 674346 617976
rect 676214 617964 676220 617976
rect 674340 617936 676220 617964
rect 674340 617924 674346 617936
rect 676214 617924 676220 617936
rect 676272 617924 676278 617976
rect 42242 617312 42248 617364
rect 42300 617352 42306 617364
rect 43070 617352 43076 617364
rect 42300 617324 43076 617352
rect 42300 617312 42306 617324
rect 43070 617312 43076 617324
rect 43128 617312 43134 617364
rect 44726 616768 44732 616820
rect 44784 616808 44790 616820
rect 62114 616808 62120 616820
rect 44784 616780 62120 616808
rect 44784 616768 44790 616780
rect 62114 616768 62120 616780
rect 62172 616768 62178 616820
rect 669406 616700 669412 616752
rect 669464 616740 669470 616752
rect 674006 616740 674012 616752
rect 669464 616712 674012 616740
rect 669464 616700 669470 616712
rect 674006 616700 674012 616712
rect 674064 616700 674070 616752
rect 674282 616632 674288 616684
rect 674340 616672 674346 616684
rect 676214 616672 676220 616684
rect 674340 616644 676220 616672
rect 674340 616632 674346 616644
rect 676214 616632 676220 616644
rect 676272 616632 676278 616684
rect 43070 616496 43076 616548
rect 43128 616536 43134 616548
rect 43806 616536 43812 616548
rect 43128 616508 43812 616536
rect 43128 616496 43134 616508
rect 43806 616496 43812 616508
rect 43864 616496 43870 616548
rect 672810 615612 672816 615664
rect 672868 615652 672874 615664
rect 674006 615652 674012 615664
rect 672868 615624 674012 615652
rect 672868 615612 672874 615624
rect 674006 615612 674012 615624
rect 674064 615612 674070 615664
rect 674282 615476 674288 615528
rect 674340 615516 674346 615528
rect 683114 615516 683120 615528
rect 674340 615488 683120 615516
rect 674340 615476 674346 615488
rect 683114 615476 683120 615488
rect 683172 615476 683178 615528
rect 670602 614864 670608 614916
rect 670660 614904 670666 614916
rect 674006 614904 674012 614916
rect 670660 614876 674012 614904
rect 670660 614864 670666 614876
rect 674006 614864 674012 614876
rect 674064 614864 674070 614916
rect 43530 614660 43536 614712
rect 43588 614700 43594 614712
rect 44358 614700 44364 614712
rect 43588 614672 44364 614700
rect 43588 614660 43594 614672
rect 44358 614660 44364 614672
rect 44416 614660 44422 614712
rect 42702 614116 42708 614168
rect 42760 614156 42766 614168
rect 62114 614156 62120 614168
rect 42760 614128 62120 614156
rect 42760 614116 42766 614128
rect 62114 614116 62120 614128
rect 62172 614116 62178 614168
rect 673546 613504 673552 613556
rect 673604 613544 673610 613556
rect 673604 613516 673776 613544
rect 673604 613504 673610 613516
rect 673748 613352 673776 613516
rect 673730 613300 673736 613352
rect 673788 613300 673794 613352
rect 42886 612756 42892 612808
rect 42944 612756 42950 612808
rect 42904 612660 42932 612756
rect 42904 612632 43668 612660
rect 43640 612592 43668 612632
rect 54478 612620 54484 612672
rect 54536 612660 54542 612672
rect 62114 612660 62120 612672
rect 54536 612632 62120 612660
rect 54536 612620 54542 612632
rect 62114 612620 62120 612632
rect 62172 612620 62178 612672
rect 43640 612564 43691 612592
rect 43070 612484 43076 612536
rect 43128 612524 43134 612536
rect 43128 612496 43562 612524
rect 43128 612484 43134 612496
rect 43663 612306 43691 612564
rect 43898 612212 43904 612264
rect 43956 612252 43962 612264
rect 44542 612252 44548 612264
rect 43956 612224 44548 612252
rect 43956 612212 43962 612224
rect 44542 612212 44548 612224
rect 44600 612212 44606 612264
rect 43766 612196 43818 612202
rect 43766 612138 43818 612144
rect 47026 612048 47032 612060
rect 44008 612020 47032 612048
rect 43875 611924 43927 611930
rect 43875 611866 43927 611872
rect 44008 611762 44036 612020
rect 47026 612008 47032 612020
rect 47084 612008 47090 612060
rect 47210 611912 47216 611924
rect 44100 611884 47216 611912
rect 44100 611558 44128 611884
rect 47210 611872 47216 611884
rect 47268 611872 47274 611924
rect 44358 611640 44364 611652
rect 44223 611612 44364 611640
rect 44223 611354 44251 611612
rect 44358 611600 44364 611612
rect 44416 611600 44422 611652
rect 653398 611328 653404 611380
rect 653456 611368 653462 611380
rect 674006 611368 674012 611380
rect 653456 611340 674012 611368
rect 653456 611328 653462 611340
rect 674006 611328 674012 611340
rect 674064 611328 674070 611380
rect 674282 611328 674288 611380
rect 674340 611368 674346 611380
rect 675386 611368 675392 611380
rect 674340 611340 675392 611368
rect 674340 611328 674346 611340
rect 675386 611328 675392 611340
rect 675444 611328 675450 611380
rect 44818 611232 44824 611244
rect 44447 611204 44824 611232
rect 44312 611124 44318 611176
rect 44370 611124 44376 611176
rect 44447 610946 44475 611204
rect 44818 611192 44824 611204
rect 44876 611192 44882 611244
rect 44542 611056 44548 611108
rect 44600 611056 44606 611108
rect 44560 610742 44588 611056
rect 657538 600312 657544 600364
rect 657596 600352 657602 600364
rect 670878 600352 670884 600364
rect 657596 600324 670884 600352
rect 657596 600312 657602 600324
rect 670878 600312 670884 600324
rect 670936 600312 670942 600364
rect 670786 599128 670792 599140
rect 666526 599100 670792 599128
rect 666526 599060 666554 599100
rect 670786 599088 670792 599100
rect 670844 599088 670850 599140
rect 663766 599032 666554 599060
rect 654778 598952 654784 599004
rect 654836 598992 654842 599004
rect 663766 598992 663794 599032
rect 654836 598964 663794 598992
rect 654836 598952 654842 598964
rect 674650 598884 674656 598936
rect 674708 598884 674714 598936
rect 674668 598664 674696 598884
rect 674650 598612 674656 598664
rect 674708 598612 674714 598664
rect 651466 597524 651472 597576
rect 651524 597564 651530 597576
rect 667382 597564 667388 597576
rect 651524 597536 667388 597564
rect 651524 597524 651530 597536
rect 667382 597524 667388 597536
rect 667440 597524 667446 597576
rect 42886 597388 42892 597440
rect 42944 597388 42950 597440
rect 42904 597032 42932 597388
rect 42886 596980 42892 597032
rect 42944 596980 42950 597032
rect 672350 596232 672356 596284
rect 672408 596272 672414 596284
rect 672718 596272 672724 596284
rect 672408 596244 672724 596272
rect 672408 596232 672414 596244
rect 672718 596232 672724 596244
rect 672776 596232 672782 596284
rect 651466 596164 651472 596216
rect 651524 596204 651530 596216
rect 661678 596204 661684 596216
rect 651524 596176 661684 596204
rect 651524 596164 651530 596176
rect 661678 596164 661684 596176
rect 661736 596164 661742 596216
rect 39942 595756 39948 595808
rect 40000 595796 40006 595808
rect 41690 595796 41696 595808
rect 40000 595768 41696 595796
rect 40000 595756 40006 595768
rect 41690 595756 41696 595768
rect 41748 595756 41754 595808
rect 651650 595484 651656 595536
rect 651708 595524 651714 595536
rect 653398 595524 653404 595536
rect 651708 595496 653404 595524
rect 651708 595484 651714 595496
rect 653398 595484 653404 595496
rect 653456 595484 653462 595536
rect 651466 594804 651472 594856
rect 651524 594844 651530 594856
rect 658918 594844 658924 594856
rect 651524 594816 658924 594844
rect 651524 594804 651530 594816
rect 658918 594804 658924 594816
rect 658976 594804 658982 594856
rect 651466 594668 651472 594720
rect 651524 594708 651530 594720
rect 657538 594708 657544 594720
rect 651524 594680 657544 594708
rect 651524 594668 651530 594680
rect 657538 594668 657544 594680
rect 657596 594668 657602 594720
rect 38562 594124 38568 594176
rect 38620 594164 38626 594176
rect 41690 594164 41696 594176
rect 38620 594136 41696 594164
rect 38620 594124 38626 594136
rect 41690 594124 41696 594136
rect 41748 594124 41754 594176
rect 651466 593036 651472 593088
rect 651524 593076 651530 593088
rect 654778 593076 654784 593088
rect 651524 593048 654784 593076
rect 651524 593036 651530 593048
rect 654778 593036 654784 593048
rect 654836 593036 654842 593088
rect 674834 592492 674840 592544
rect 674892 592532 674898 592544
rect 683390 592532 683396 592544
rect 674892 592504 683396 592532
rect 674892 592492 674898 592504
rect 683390 592492 683396 592504
rect 683448 592492 683454 592544
rect 675570 588548 675576 588600
rect 675628 588588 675634 588600
rect 684034 588588 684040 588600
rect 675628 588560 684040 588588
rect 675628 588548 675634 588560
rect 684034 588548 684040 588560
rect 684092 588548 684098 588600
rect 35434 587120 35440 587172
rect 35492 587160 35498 587172
rect 41506 587160 41512 587172
rect 35492 587132 41512 587160
rect 35492 587120 35498 587132
rect 41506 587120 41512 587132
rect 41564 587120 41570 587172
rect 36538 586100 36544 586152
rect 36596 586140 36602 586152
rect 39666 586140 39672 586152
rect 36596 586112 39672 586140
rect 36596 586100 36602 586112
rect 39666 586100 39672 586112
rect 39724 586100 39730 586152
rect 32398 585896 32404 585948
rect 32456 585936 32462 585948
rect 41690 585936 41696 585948
rect 32456 585908 41696 585936
rect 32456 585896 32462 585908
rect 41690 585896 41696 585908
rect 41748 585896 41754 585948
rect 31018 585760 31024 585812
rect 31076 585800 31082 585812
rect 39758 585800 39764 585812
rect 31076 585772 39764 585800
rect 31076 585760 31082 585772
rect 39758 585760 39764 585772
rect 39816 585760 39822 585812
rect 652018 581000 652024 581052
rect 652076 581040 652082 581052
rect 673914 581040 673920 581052
rect 652076 581012 673920 581040
rect 652076 581000 652082 581012
rect 673914 581000 673920 581012
rect 673972 581000 673978 581052
rect 668578 580252 668584 580304
rect 668636 580292 668642 580304
rect 673914 580292 673920 580304
rect 668636 580264 673920 580292
rect 668636 580252 668642 580264
rect 673914 580252 673920 580264
rect 673972 580252 673978 580304
rect 669866 579844 669872 579896
rect 669924 579884 669930 579896
rect 673914 579884 673920 579896
rect 669924 579856 673920 579884
rect 669924 579844 669930 579856
rect 673914 579844 673920 579856
rect 673972 579844 673978 579896
rect 660298 579640 660304 579692
rect 660356 579680 660362 579692
rect 673546 579680 673552 579692
rect 660356 579652 673552 579680
rect 660356 579640 660362 579652
rect 673546 579640 673552 579652
rect 673604 579640 673610 579692
rect 669590 579368 669596 579420
rect 669648 579408 669654 579420
rect 673914 579408 673920 579420
rect 669648 579380 673920 579408
rect 669648 579368 669654 579380
rect 673914 579368 673920 579380
rect 673972 579368 673978 579420
rect 670234 579028 670240 579080
rect 670292 579068 670298 579080
rect 673914 579068 673920 579080
rect 670292 579040 673920 579068
rect 670292 579028 670298 579040
rect 673914 579028 673920 579040
rect 673972 579028 673978 579080
rect 670234 578552 670240 578604
rect 670292 578592 670298 578604
rect 673914 578592 673920 578604
rect 670292 578564 673920 578592
rect 670292 578552 670298 578564
rect 673914 578552 673920 578564
rect 673972 578552 673978 578604
rect 670050 578144 670056 578196
rect 670108 578184 670114 578196
rect 673914 578184 673920 578196
rect 670108 578156 673920 578184
rect 670108 578144 670114 578156
rect 673914 578144 673920 578156
rect 673972 578144 673978 578196
rect 669406 577736 669412 577788
rect 669464 577776 669470 577788
rect 673914 577776 673920 577788
rect 669464 577748 673920 577776
rect 669464 577736 669470 577748
rect 673914 577736 673920 577748
rect 673972 577736 673978 577788
rect 42426 577600 42432 577652
rect 42484 577600 42490 577652
rect 42444 577436 42472 577600
rect 42610 577532 42616 577584
rect 42668 577572 42674 577584
rect 42668 577544 42840 577572
rect 42668 577532 42674 577544
rect 42610 577436 42616 577448
rect 42444 577408 42616 577436
rect 42610 577396 42616 577408
rect 42668 577396 42674 577448
rect 42334 577260 42340 577312
rect 42392 577300 42398 577312
rect 42812 577300 42840 577544
rect 671430 577396 671436 577448
rect 671488 577436 671494 577448
rect 673914 577436 673920 577448
rect 671488 577408 673920 577436
rect 671488 577396 671494 577408
rect 673914 577396 673920 577408
rect 673972 577396 673978 577448
rect 42392 577272 42840 577300
rect 42392 577260 42398 577272
rect 671338 576920 671344 576972
rect 671396 576960 671402 576972
rect 673914 576960 673920 576972
rect 671396 576932 673920 576960
rect 671396 576920 671402 576932
rect 673914 576920 673920 576932
rect 673972 576920 673978 576972
rect 45094 575424 45100 575476
rect 45152 575464 45158 575476
rect 62390 575464 62396 575476
rect 45152 575436 62396 575464
rect 45152 575424 45158 575436
rect 62390 575424 62396 575436
rect 62448 575424 62454 575476
rect 671798 575356 671804 575408
rect 671856 575396 671862 575408
rect 673914 575396 673920 575408
rect 671856 575368 673920 575396
rect 671856 575356 671862 575368
rect 673914 575356 673920 575368
rect 673972 575356 673978 575408
rect 670418 574540 670424 574592
rect 670476 574580 670482 574592
rect 673546 574580 673552 574592
rect 670476 574552 673552 574580
rect 670476 574540 670482 574552
rect 673546 574540 673552 574552
rect 673604 574540 673610 574592
rect 671982 574268 671988 574320
rect 672040 574308 672046 574320
rect 673546 574308 673552 574320
rect 672040 574280 673552 574308
rect 672040 574268 672046 574280
rect 673546 574268 673552 574280
rect 673604 574268 673610 574320
rect 667014 574064 667020 574116
rect 667072 574104 667078 574116
rect 673914 574104 673920 574116
rect 667072 574076 673920 574104
rect 667072 574064 667078 574076
rect 673914 574064 673920 574076
rect 673972 574064 673978 574116
rect 45554 573996 45560 574048
rect 45612 574036 45618 574048
rect 62390 574036 62396 574048
rect 45612 574008 62396 574036
rect 45612 573996 45618 574008
rect 62390 573996 62396 574008
rect 62448 573996 62454 574048
rect 672534 573724 672540 573776
rect 672592 573764 672598 573776
rect 673914 573764 673920 573776
rect 672592 573736 673920 573764
rect 672592 573724 672598 573736
rect 673914 573724 673920 573736
rect 673972 573724 673978 573776
rect 671614 572092 671620 572144
rect 671672 572132 671678 572144
rect 673914 572132 673920 572144
rect 671672 572104 673920 572132
rect 671672 572092 671678 572104
rect 673914 572092 673920 572104
rect 673972 572092 673978 572144
rect 674650 571548 674656 571600
rect 674708 571588 674714 571600
rect 676214 571588 676220 571600
rect 674708 571560 676220 571588
rect 674708 571548 674714 571560
rect 676214 571548 676220 571560
rect 676272 571548 676278 571600
rect 671982 570800 671988 570852
rect 672040 570840 672046 570852
rect 673914 570840 673920 570852
rect 672040 570812 673920 570840
rect 672040 570800 672046 570812
rect 673914 570800 673920 570812
rect 673972 570800 673978 570852
rect 667198 570528 667204 570580
rect 667256 570568 667262 570580
rect 667658 570568 667664 570580
rect 667256 570540 667664 570568
rect 667256 570528 667262 570540
rect 667658 570528 667664 570540
rect 667716 570528 667722 570580
rect 667658 570188 667664 570240
rect 667716 570228 667722 570240
rect 673914 570228 673920 570240
rect 667716 570200 673920 570228
rect 667716 570188 667722 570200
rect 673914 570188 673920 570200
rect 673972 570188 673978 570240
rect 674650 569916 674656 569968
rect 674708 569956 674714 569968
rect 683114 569956 683120 569968
rect 674708 569928 683120 569956
rect 674708 569916 674714 569928
rect 683114 569916 683120 569928
rect 683172 569916 683178 569968
rect 669774 569576 669780 569628
rect 669832 569616 669838 569628
rect 673546 569616 673552 569628
rect 669832 569588 673552 569616
rect 669832 569576 669838 569588
rect 673546 569576 673552 569588
rect 673604 569576 673610 569628
rect 42426 569372 42432 569424
rect 42484 569372 42490 569424
rect 42444 569220 42472 569372
rect 42426 569168 42432 569220
rect 42484 569168 42490 569220
rect 653398 565836 653404 565888
rect 653456 565876 653462 565888
rect 673546 565876 673552 565888
rect 653456 565848 673552 565876
rect 653456 565836 653462 565848
rect 673546 565836 673552 565848
rect 673604 565836 673610 565888
rect 674650 558016 674656 558068
rect 674708 558056 674714 558068
rect 675294 558056 675300 558068
rect 674708 558028 675300 558056
rect 674708 558016 674714 558028
rect 675294 558016 675300 558028
rect 675352 558016 675358 558068
rect 657814 554752 657820 554804
rect 657872 554792 657878 554804
rect 674006 554792 674012 554804
rect 657872 554764 674012 554792
rect 657872 554752 657878 554764
rect 674006 554752 674012 554764
rect 674064 554752 674070 554804
rect 655146 553392 655152 553444
rect 655204 553432 655210 553444
rect 674006 553432 674012 553444
rect 655204 553404 674012 553432
rect 655204 553392 655210 553404
rect 674006 553392 674012 553404
rect 674064 553392 674070 553444
rect 40034 553324 40040 553376
rect 40092 553364 40098 553376
rect 41690 553364 41696 553376
rect 40092 553336 41696 553364
rect 40092 553324 40098 553336
rect 41690 553324 41696 553336
rect 41748 553324 41754 553376
rect 651466 552644 651472 552696
rect 651524 552684 651530 552696
rect 665818 552684 665824 552696
rect 651524 552656 665824 552684
rect 651524 552644 651530 552656
rect 665818 552644 665824 552656
rect 665876 552644 665882 552696
rect 41322 552100 41328 552152
rect 41380 552140 41386 552152
rect 41690 552140 41696 552152
rect 41380 552112 41696 552140
rect 41380 552100 41386 552112
rect 41690 552100 41696 552112
rect 41748 552100 41754 552152
rect 651466 550604 651472 550656
rect 651524 550644 651530 550656
rect 669958 550644 669964 550656
rect 651524 550616 669964 550644
rect 651524 550604 651530 550616
rect 669958 550604 669964 550616
rect 670016 550604 670022 550656
rect 41138 550536 41144 550588
rect 41196 550576 41202 550588
rect 41690 550576 41696 550588
rect 41196 550548 41696 550576
rect 41196 550536 41202 550548
rect 41690 550536 41696 550548
rect 41748 550536 41754 550588
rect 651374 550332 651380 550384
rect 651432 550372 651438 550384
rect 653398 550372 653404 550384
rect 651432 550344 653404 550372
rect 651432 550332 651438 550344
rect 653398 550332 653404 550344
rect 653456 550332 653462 550384
rect 675294 550060 675300 550112
rect 675352 550060 675358 550112
rect 674742 549964 674748 549976
rect 674576 549936 674748 549964
rect 674576 549284 674604 549936
rect 674742 549924 674748 549936
rect 674800 549924 674806 549976
rect 674834 549788 674840 549840
rect 674892 549828 674898 549840
rect 675312 549828 675340 550060
rect 674892 549800 675340 549828
rect 674892 549788 674898 549800
rect 674742 549284 674748 549296
rect 674576 549256 674748 549284
rect 674742 549244 674748 549256
rect 674800 549244 674806 549296
rect 651466 549176 651472 549228
rect 651524 549216 651530 549228
rect 657814 549216 657820 549228
rect 651524 549188 657820 549216
rect 651524 549176 651530 549188
rect 657814 549176 657820 549188
rect 657872 549176 657878 549228
rect 651466 548836 651472 548888
rect 651524 548876 651530 548888
rect 655146 548876 655152 548888
rect 651524 548848 655152 548876
rect 651524 548836 651530 548848
rect 655146 548836 655152 548848
rect 655204 548836 655210 548888
rect 674374 547272 674380 547324
rect 674432 547312 674438 547324
rect 683206 547312 683212 547324
rect 674432 547284 683212 547312
rect 674432 547272 674438 547284
rect 683206 547272 683212 547284
rect 683264 547272 683270 547324
rect 675294 546864 675300 546916
rect 675352 546904 675358 546916
rect 682378 546904 682384 546916
rect 675352 546876 682384 546904
rect 675352 546864 675358 546876
rect 682378 546864 682384 546876
rect 682436 546864 682442 546916
rect 672626 544552 672632 544604
rect 672684 544592 672690 544604
rect 672684 544564 672856 544592
rect 672684 544552 672690 544564
rect 672828 544400 672856 544564
rect 675018 544552 675024 544604
rect 675076 544592 675082 544604
rect 675386 544592 675392 544604
rect 675076 544564 675392 544592
rect 675076 544552 675082 544564
rect 675386 544552 675392 544564
rect 675444 544552 675450 544604
rect 29638 544348 29644 544400
rect 29696 544388 29702 544400
rect 41690 544388 41696 544400
rect 29696 544360 41696 544388
rect 29696 544348 29702 544360
rect 41690 544348 41696 544360
rect 41748 544348 41754 544400
rect 672810 544348 672816 544400
rect 672868 544348 672874 544400
rect 674282 537140 674288 537192
rect 674340 537180 674346 537192
rect 675478 537180 675484 537192
rect 674340 537152 675484 537180
rect 674340 537140 674346 537152
rect 675478 537140 675484 537152
rect 675536 537140 675542 537192
rect 673914 536392 673920 536444
rect 673972 536392 673978 536444
rect 673932 536172 673960 536392
rect 673914 536120 673920 536172
rect 673972 536120 673978 536172
rect 673730 535984 673736 536036
rect 673788 536024 673794 536036
rect 673788 535996 673960 536024
rect 673788 535984 673794 535996
rect 667382 535780 667388 535832
rect 667440 535820 667446 535832
rect 673730 535820 673736 535832
rect 667440 535792 673736 535820
rect 667440 535780 667446 535792
rect 673730 535780 673736 535792
rect 673788 535780 673794 535832
rect 661678 535440 661684 535492
rect 661736 535480 661742 535492
rect 673932 535480 673960 535996
rect 661736 535452 673960 535480
rect 661736 535440 661742 535452
rect 669590 534964 669596 535016
rect 669648 535004 669654 535016
rect 672626 535004 672632 535016
rect 669648 534976 672632 535004
rect 669648 534964 669654 534976
rect 672626 534964 672632 534976
rect 672684 534964 672690 535016
rect 670234 534284 670240 534336
rect 670292 534324 670298 534336
rect 672626 534324 672632 534336
rect 670292 534296 672632 534324
rect 670292 534284 670298 534296
rect 672626 534284 672632 534296
rect 672684 534284 672690 534336
rect 674282 534216 674288 534268
rect 674340 534256 674346 534268
rect 676214 534256 676220 534268
rect 674340 534228 676220 534256
rect 674340 534216 674346 534228
rect 676214 534216 676220 534228
rect 676272 534216 676278 534268
rect 658918 534080 658924 534132
rect 658976 534120 658982 534132
rect 673730 534120 673736 534132
rect 658976 534092 673736 534120
rect 658976 534080 658982 534092
rect 673730 534080 673736 534092
rect 673788 534080 673794 534132
rect 42242 533400 42248 533452
rect 42300 533440 42306 533452
rect 42978 533440 42984 533452
rect 42300 533412 42984 533440
rect 42300 533400 42306 533412
rect 42978 533400 42984 533412
rect 43036 533400 43042 533452
rect 669406 533332 669412 533384
rect 669464 533372 669470 533384
rect 672626 533372 672632 533384
rect 669464 533344 672632 533372
rect 669464 533332 669470 533344
rect 672626 533332 672632 533344
rect 672684 533332 672690 533384
rect 675478 533332 675484 533384
rect 675536 533372 675542 533384
rect 683574 533372 683580 533384
rect 675536 533344 683580 533372
rect 675536 533332 675542 533344
rect 683574 533332 683580 533344
rect 683632 533332 683638 533384
rect 674282 532788 674288 532840
rect 674340 532828 674346 532840
rect 676030 532828 676036 532840
rect 674340 532800 676036 532828
rect 674340 532788 674346 532800
rect 676030 532788 676036 532800
rect 676088 532788 676094 532840
rect 44726 531224 44732 531276
rect 44784 531264 44790 531276
rect 62298 531264 62304 531276
rect 44784 531236 62304 531264
rect 44784 531224 44790 531236
rect 62298 531224 62304 531236
rect 62356 531224 62362 531276
rect 53098 531088 53104 531140
rect 53156 531128 53162 531140
rect 62114 531128 62120 531140
rect 53156 531100 62120 531128
rect 53156 531088 53162 531100
rect 62114 531088 62120 531100
rect 62172 531088 62178 531140
rect 673178 530068 673184 530120
rect 673236 530108 673242 530120
rect 673730 530108 673736 530120
rect 673236 530080 673736 530108
rect 673236 530068 673242 530080
rect 673730 530068 673736 530080
rect 673788 530068 673794 530120
rect 668946 529932 668952 529984
rect 669004 529972 669010 529984
rect 673730 529972 673736 529984
rect 669004 529944 673736 529972
rect 669004 529932 669010 529944
rect 673730 529932 673736 529944
rect 673788 529932 673794 529984
rect 670970 529456 670976 529508
rect 671028 529496 671034 529508
rect 673730 529496 673736 529508
rect 671028 529468 673736 529496
rect 671028 529456 671034 529468
rect 673730 529456 673736 529468
rect 673788 529456 673794 529508
rect 671154 529184 671160 529236
rect 671212 529224 671218 529236
rect 673730 529224 673736 529236
rect 671212 529196 673736 529224
rect 671212 529184 671218 529196
rect 673730 529184 673736 529196
rect 673788 529184 673794 529236
rect 672994 528844 673000 528896
rect 673052 528884 673058 528896
rect 673052 528856 673454 528884
rect 673052 528844 673058 528856
rect 673426 528816 673454 528856
rect 673730 528816 673736 528828
rect 673426 528788 673736 528816
rect 673730 528776 673736 528788
rect 673788 528776 673794 528828
rect 45094 528572 45100 528624
rect 45152 528612 45158 528624
rect 62114 528612 62120 528624
rect 45152 528584 62120 528612
rect 45152 528572 45158 528584
rect 62114 528572 62120 528584
rect 62172 528572 62178 528624
rect 674374 527552 674380 527604
rect 674432 527592 674438 527604
rect 676214 527592 676220 527604
rect 674432 527564 676220 527592
rect 674432 527552 674438 527564
rect 676214 527552 676220 527564
rect 676272 527552 676278 527604
rect 54478 527076 54484 527128
rect 54536 527116 54542 527128
rect 62114 527116 62120 527128
rect 54536 527088 62120 527116
rect 54536 527076 54542 527088
rect 62114 527076 62120 527088
rect 62172 527076 62178 527128
rect 674282 526736 674288 526788
rect 674340 526776 674346 526788
rect 676030 526776 676036 526788
rect 674340 526748 676036 526776
rect 674340 526736 674346 526748
rect 676030 526736 676036 526748
rect 676088 526736 676094 526788
rect 674466 526328 674472 526380
rect 674524 526368 674530 526380
rect 676030 526368 676036 526380
rect 674524 526340 676036 526368
rect 674524 526328 674530 526340
rect 676030 526328 676036 526340
rect 676088 526328 676094 526380
rect 674282 524560 674288 524612
rect 674340 524600 674346 524612
rect 683114 524600 683120 524612
rect 674340 524572 683120 524600
rect 674340 524560 674346 524572
rect 683114 524560 683120 524572
rect 683172 524560 683178 524612
rect 670620 524504 673454 524532
rect 668762 524356 668768 524408
rect 668820 524396 668826 524408
rect 670620 524396 670648 524504
rect 673426 524464 673454 524504
rect 674006 524464 674012 524476
rect 673426 524436 674012 524464
rect 674006 524424 674012 524436
rect 674064 524424 674070 524476
rect 668820 524368 670648 524396
rect 668820 524356 668826 524368
rect 652202 520888 652208 520940
rect 652260 520928 652266 520940
rect 668762 520928 668768 520940
rect 652260 520900 668768 520928
rect 652260 520888 652266 520900
rect 668762 520888 668768 520900
rect 668820 520888 668826 520940
rect 675662 520208 675668 520260
rect 675720 520248 675726 520260
rect 680354 520248 680360 520260
rect 675720 520220 680360 520248
rect 675720 520208 675726 520220
rect 680354 520208 680360 520220
rect 680412 520208 680418 520260
rect 675478 520072 675484 520124
rect 675536 520112 675542 520124
rect 678974 520112 678980 520124
rect 675536 520084 678980 520112
rect 675536 520072 675542 520084
rect 678974 520072 678980 520084
rect 679032 520072 679038 520124
rect 674926 503820 674932 503872
rect 674984 503860 674990 503872
rect 678238 503860 678244 503872
rect 674984 503832 678244 503860
rect 674984 503820 674990 503832
rect 678238 503820 678244 503832
rect 678296 503820 678302 503872
rect 675110 503616 675116 503668
rect 675168 503656 675174 503668
rect 679618 503656 679624 503668
rect 675168 503628 679624 503656
rect 675168 503616 675174 503628
rect 679618 503616 679624 503628
rect 679676 503616 679682 503668
rect 675294 503480 675300 503532
rect 675352 503520 675358 503532
rect 680998 503520 681004 503532
rect 675352 503492 681004 503520
rect 675352 503480 675358 503492
rect 680998 503480 681004 503492
rect 681056 503480 681062 503532
rect 652018 493280 652024 493332
rect 652076 493320 652082 493332
rect 673178 493320 673184 493332
rect 652076 493292 673184 493320
rect 652076 493280 652082 493292
rect 673178 493280 673184 493292
rect 673236 493280 673242 493332
rect 669958 491444 669964 491496
rect 670016 491484 670022 491496
rect 673822 491484 673828 491496
rect 670016 491456 673828 491484
rect 670016 491444 670022 491456
rect 673822 491444 673828 491456
rect 673880 491444 673886 491496
rect 674282 491444 674288 491496
rect 674340 491484 674346 491496
rect 676030 491484 676036 491496
rect 674340 491456 676036 491484
rect 674340 491444 674346 491456
rect 676030 491444 676036 491456
rect 676088 491444 676094 491496
rect 665818 491308 665824 491360
rect 665876 491348 665882 491360
rect 674006 491348 674012 491360
rect 665876 491320 674012 491348
rect 665876 491308 665882 491320
rect 674006 491308 674012 491320
rect 674064 491308 674070 491360
rect 670786 490900 670792 490952
rect 670844 490940 670850 490952
rect 674006 490940 674012 490952
rect 670844 490912 674012 490940
rect 670844 490900 670850 490912
rect 674006 490900 674012 490912
rect 674064 490900 674070 490952
rect 672626 490084 672632 490136
rect 672684 490124 672690 490136
rect 674006 490124 674012 490136
rect 672684 490096 674012 490124
rect 672684 490084 672690 490096
rect 674006 490084 674012 490096
rect 674064 490084 674070 490136
rect 672626 489880 672632 489932
rect 672684 489920 672690 489932
rect 673178 489920 673184 489932
rect 672684 489892 673184 489920
rect 672684 489880 672690 489892
rect 673178 489880 673184 489892
rect 673236 489880 673242 489932
rect 672442 489608 672448 489660
rect 672500 489648 672506 489660
rect 674006 489648 674012 489660
rect 672500 489620 674012 489648
rect 672500 489608 672506 489620
rect 674006 489608 674012 489620
rect 674064 489608 674070 489660
rect 671522 489268 671528 489320
rect 671580 489308 671586 489320
rect 674006 489308 674012 489320
rect 671580 489280 674012 489308
rect 671580 489268 671586 489280
rect 674006 489268 674012 489280
rect 674064 489268 674070 489320
rect 671338 488452 671344 488504
rect 671396 488492 671402 488504
rect 674006 488492 674012 488504
rect 671396 488464 674012 488492
rect 671396 488452 671402 488464
rect 674006 488452 674012 488464
rect 674064 488452 674070 488504
rect 671798 486820 671804 486872
rect 671856 486860 671862 486872
rect 674006 486860 674012 486872
rect 671856 486832 674012 486860
rect 671856 486820 671862 486832
rect 674006 486820 674012 486832
rect 674064 486820 674070 486872
rect 672258 486004 672264 486056
rect 672316 486044 672322 486056
rect 674006 486044 674012 486056
rect 672316 486016 674012 486044
rect 672316 486004 672322 486016
rect 674006 486004 674012 486016
rect 674064 486004 674070 486056
rect 676030 485324 676036 485376
rect 676088 485364 676094 485376
rect 677134 485364 677140 485376
rect 676088 485336 677140 485364
rect 676088 485324 676094 485336
rect 677134 485324 677140 485336
rect 677192 485324 677198 485376
rect 674282 485120 674288 485172
rect 674340 485160 674346 485172
rect 676030 485160 676036 485172
rect 674340 485132 676036 485160
rect 674340 485120 674346 485132
rect 676030 485120 676036 485132
rect 676088 485120 676094 485172
rect 667014 484372 667020 484424
rect 667072 484412 667078 484424
rect 674006 484412 674012 484424
rect 667072 484384 674012 484412
rect 667072 484372 667078 484384
rect 674006 484372 674012 484384
rect 674064 484372 674070 484424
rect 674466 484372 674472 484424
rect 674524 484412 674530 484424
rect 675846 484412 675852 484424
rect 674524 484384 675852 484412
rect 674524 484372 674530 484384
rect 675846 484372 675852 484384
rect 675904 484372 675910 484424
rect 676214 484304 676220 484356
rect 676272 484344 676278 484356
rect 677410 484344 677416 484356
rect 676272 484316 677416 484344
rect 676272 484304 676278 484316
rect 677410 484304 677416 484316
rect 677468 484304 677474 484356
rect 674282 482468 674288 482520
rect 674340 482508 674346 482520
rect 676030 482508 676036 482520
rect 674340 482480 676036 482508
rect 674340 482468 674346 482480
rect 676030 482468 676036 482480
rect 676088 482468 676094 482520
rect 674006 482168 674012 482180
rect 669286 482140 674012 482168
rect 668394 481924 668400 481976
rect 668452 481964 668458 481976
rect 669286 481964 669314 482140
rect 674006 482128 674012 482140
rect 674064 482128 674070 482180
rect 674282 482060 674288 482112
rect 674340 482100 674346 482112
rect 676030 482100 676036 482112
rect 674340 482072 676036 482100
rect 674340 482060 674346 482072
rect 676030 482060 676036 482072
rect 676088 482060 676094 482112
rect 668452 481936 669314 481964
rect 668452 481924 668458 481936
rect 667566 481788 667572 481840
rect 667624 481828 667630 481840
rect 674006 481828 674012 481840
rect 667624 481800 674012 481828
rect 667624 481788 667630 481800
rect 674006 481788 674012 481800
rect 674064 481788 674070 481840
rect 658918 480904 658924 480956
rect 658976 480944 658982 480956
rect 670418 480944 670424 480956
rect 658976 480916 670424 480944
rect 658976 480904 658982 480916
rect 670418 480904 670424 480916
rect 670476 480944 670482 480956
rect 674006 480944 674012 480956
rect 670476 480916 674012 480944
rect 670476 480904 670482 480916
rect 674006 480904 674012 480916
rect 674064 480904 674070 480956
rect 674282 480360 674288 480412
rect 674340 480400 674346 480412
rect 683114 480400 683120 480412
rect 674340 480372 683120 480400
rect 674340 480360 674346 480372
rect 683114 480360 683120 480372
rect 683172 480360 683178 480412
rect 650638 476076 650644 476128
rect 650696 476116 650702 476128
rect 652202 476116 652208 476128
rect 650696 476088 652208 476116
rect 650696 476076 650702 476088
rect 652202 476076 652208 476088
rect 652260 476076 652266 476128
rect 673362 475464 673368 475516
rect 673420 475504 673426 475516
rect 674006 475504 674012 475516
rect 673420 475476 674012 475504
rect 673420 475464 673426 475476
rect 674006 475464 674012 475476
rect 674064 475464 674070 475516
rect 674282 475464 674288 475516
rect 674340 475504 674346 475516
rect 676214 475504 676220 475516
rect 674340 475476 676220 475504
rect 674340 475464 674346 475476
rect 676214 475464 676220 475476
rect 676272 475464 676278 475516
rect 676030 475124 676036 475176
rect 676088 475164 676094 475176
rect 680354 475164 680360 475176
rect 676088 475136 680360 475164
rect 676088 475124 676094 475136
rect 680354 475124 680360 475136
rect 680412 475124 680418 475176
rect 656158 466420 656164 466472
rect 656216 466460 656222 466472
rect 658918 466460 658924 466472
rect 656216 466432 658924 466460
rect 656216 466420 656222 466432
rect 658918 466420 658924 466432
rect 658976 466420 658982 466472
rect 651374 458396 651380 458448
rect 651432 458436 651438 458448
rect 656158 458436 656164 458448
rect 651432 458408 656164 458436
rect 651432 458396 651438 458408
rect 656158 458396 656164 458408
rect 656216 458396 656222 458448
rect 667842 456560 667848 456612
rect 667900 456600 667906 456612
rect 667900 456572 673988 456600
rect 667900 456560 667906 456572
rect 673960 456246 673988 456572
rect 674282 456084 674288 456136
rect 674340 456124 674346 456136
rect 676214 456124 676220 456136
rect 674340 456096 676220 456124
rect 674340 456084 674346 456096
rect 676214 456084 676220 456096
rect 676272 456084 676278 456136
rect 673828 456068 673880 456074
rect 673828 456010 673880 456016
rect 672810 455744 672816 455796
rect 672868 455784 672874 455796
rect 672868 455756 673762 455784
rect 672868 455744 672874 455756
rect 669222 455608 669228 455660
rect 669280 455648 669286 455660
rect 669280 455620 673624 455648
rect 669280 455608 669286 455620
rect 673270 455336 673276 455388
rect 673328 455336 673334 455388
rect 672074 455064 672080 455116
rect 672132 455104 672138 455116
rect 672132 455076 673204 455104
rect 672132 455064 672138 455076
rect 673176 454818 673204 455076
rect 673288 455022 673316 455336
rect 673388 455252 673440 455258
rect 673388 455194 673440 455200
rect 673506 455252 673558 455258
rect 673506 455194 673558 455200
rect 673040 454724 673046 454776
rect 673098 454724 673104 454776
rect 674282 454724 674288 454776
rect 674340 454764 674346 454776
rect 675662 454764 675668 454776
rect 674340 454736 675668 454764
rect 674340 454724 674346 454736
rect 675662 454724 675668 454736
rect 675720 454724 675726 454776
rect 673058 454614 673086 454724
rect 650822 454520 650828 454572
rect 650880 454560 650886 454572
rect 651374 454560 651380 454572
rect 650880 454532 651380 454560
rect 650880 454520 650886 454532
rect 651374 454520 651380 454532
rect 651432 454520 651438 454572
rect 674282 454452 674288 454504
rect 674340 454492 674346 454504
rect 675478 454492 675484 454504
rect 674340 454464 675484 454492
rect 674340 454452 674346 454464
rect 675478 454452 675484 454464
rect 675536 454452 675542 454504
rect 672954 454436 673006 454442
rect 672954 454378 673006 454384
rect 672816 454232 672868 454238
rect 674282 454180 674288 454232
rect 674340 454220 674346 454232
rect 675846 454220 675852 454232
rect 674340 454192 675852 454220
rect 674340 454180 674346 454192
rect 675846 454180 675852 454192
rect 675904 454180 675910 454232
rect 672816 454174 672868 454180
rect 672258 453908 672264 453960
rect 672316 453948 672322 453960
rect 672316 453920 672750 453948
rect 672316 453908 672322 453920
rect 674282 453908 674288 453960
rect 674340 453948 674346 453960
rect 676030 453948 676036 453960
rect 674340 453920 676036 453948
rect 674340 453908 674346 453920
rect 676030 453908 676036 453920
rect 676088 453908 676094 453960
rect 35802 429156 35808 429208
rect 35860 429196 35866 429208
rect 41322 429196 41328 429208
rect 35860 429168 41328 429196
rect 35860 429156 35866 429168
rect 41322 429156 41328 429168
rect 41380 429156 41386 429208
rect 41138 425348 41144 425400
rect 41196 425388 41202 425400
rect 41690 425388 41696 425400
rect 41196 425360 41696 425388
rect 41196 425348 41202 425360
rect 41690 425348 41696 425360
rect 41748 425348 41754 425400
rect 40954 420928 40960 420980
rect 41012 420968 41018 420980
rect 41690 420968 41696 420980
rect 41012 420940 41696 420968
rect 41012 420928 41018 420940
rect 41690 420928 41696 420940
rect 41748 420928 41754 420980
rect 33042 415896 33048 415948
rect 33100 415936 33106 415948
rect 40586 415936 40592 415948
rect 33100 415908 40592 415936
rect 33100 415896 33106 415908
rect 40586 415896 40592 415908
rect 40644 415896 40650 415948
rect 42242 406036 42248 406088
rect 42300 406036 42306 406088
rect 42260 405680 42288 406036
rect 42242 405628 42248 405680
rect 42300 405628 42306 405680
rect 45094 404268 45100 404320
rect 45152 404308 45158 404320
rect 62114 404308 62120 404320
rect 45152 404280 62120 404308
rect 45152 404268 45158 404280
rect 62114 404268 62120 404280
rect 62172 404268 62178 404320
rect 674558 403248 674564 403300
rect 674616 403288 674622 403300
rect 676214 403288 676220 403300
rect 674616 403260 676220 403288
rect 674616 403248 674622 403260
rect 676214 403248 676220 403260
rect 676272 403248 676278 403300
rect 46106 402908 46112 402960
rect 46164 402948 46170 402960
rect 62114 402948 62120 402960
rect 46164 402920 62120 402948
rect 46164 402908 46170 402920
rect 62114 402908 62120 402920
rect 62172 402908 62178 402960
rect 51074 400188 51080 400240
rect 51132 400228 51138 400240
rect 62114 400228 62120 400240
rect 51132 400200 62120 400228
rect 51132 400188 51138 400200
rect 62114 400188 62120 400200
rect 62172 400188 62178 400240
rect 47946 400052 47952 400104
rect 48004 400092 48010 400104
rect 62114 400092 62120 400104
rect 48004 400064 62120 400092
rect 48004 400052 48010 400064
rect 62114 400052 62120 400064
rect 62172 400052 62178 400104
rect 674926 398828 674932 398880
rect 674984 398868 674990 398880
rect 676030 398868 676036 398880
rect 674984 398840 676036 398868
rect 674984 398828 674990 398840
rect 676030 398828 676036 398840
rect 676088 398828 676094 398880
rect 54478 398760 54484 398812
rect 54536 398800 54542 398812
rect 62114 398800 62120 398812
rect 54536 398772 62120 398800
rect 54536 398760 54542 398772
rect 62114 398760 62120 398772
rect 62172 398760 62178 398812
rect 47578 397400 47584 397452
rect 47636 397440 47642 397452
rect 50706 397440 50712 397452
rect 47636 397412 50712 397440
rect 47636 397400 47642 397412
rect 50706 397400 50712 397412
rect 50764 397400 50770 397452
rect 674374 396040 674380 396092
rect 674432 396080 674438 396092
rect 676030 396080 676036 396092
rect 674432 396052 676036 396080
rect 674432 396040 674438 396052
rect 676030 396040 676036 396052
rect 676088 396040 676094 396092
rect 675018 395700 675024 395752
rect 675076 395740 675082 395752
rect 676214 395740 676220 395752
rect 675076 395712 676220 395740
rect 675076 395700 675082 395712
rect 676214 395700 676220 395712
rect 676272 395700 676278 395752
rect 674466 394272 674472 394324
rect 674524 394312 674530 394324
rect 676214 394312 676220 394324
rect 674524 394284 676220 394312
rect 674524 394272 674530 394284
rect 676214 394272 676220 394284
rect 676272 394272 676278 394324
rect 679618 386764 679624 386776
rect 675588 386736 679624 386764
rect 675588 386424 675616 386736
rect 679618 386724 679624 386736
rect 679676 386724 679682 386776
rect 675496 386396 675616 386424
rect 674834 386112 674840 386164
rect 674892 386152 674898 386164
rect 675294 386152 675300 386164
rect 674892 386124 675300 386152
rect 674892 386112 674898 386124
rect 675294 386112 675300 386124
rect 675352 386112 675358 386164
rect 675496 386028 675524 386396
rect 675478 385976 675484 386028
rect 675536 385976 675542 386028
rect 41322 382372 41328 382424
rect 41380 382412 41386 382424
rect 41690 382412 41696 382424
rect 41380 382384 41696 382412
rect 41380 382372 41386 382384
rect 41690 382372 41696 382384
rect 41748 382372 41754 382424
rect 674374 382168 674380 382220
rect 674432 382208 674438 382220
rect 675110 382208 675116 382220
rect 674432 382180 675116 382208
rect 674432 382168 674438 382180
rect 675110 382168 675116 382180
rect 675168 382168 675174 382220
rect 674558 378088 674564 378140
rect 674616 378128 674622 378140
rect 675110 378128 675116 378140
rect 674616 378100 675116 378128
rect 674616 378088 674622 378100
rect 675110 378088 675116 378100
rect 675168 378088 675174 378140
rect 674374 375300 674380 375352
rect 674432 375340 674438 375352
rect 675110 375340 675116 375352
rect 674432 375312 675116 375340
rect 674432 375300 674438 375312
rect 675110 375300 675116 375312
rect 675168 375300 675174 375352
rect 651466 373940 651472 373992
rect 651524 373980 651530 373992
rect 657538 373980 657544 373992
rect 651524 373952 657544 373980
rect 651524 373940 651530 373952
rect 657538 373940 657544 373952
rect 657596 373940 657602 373992
rect 32398 373260 32404 373312
rect 32456 373300 32462 373312
rect 41690 373300 41696 373312
rect 32456 373272 41696 373300
rect 32456 373260 32462 373272
rect 41690 373260 41696 373272
rect 41748 373260 41754 373312
rect 42058 373192 42064 373244
rect 42116 373232 42122 373244
rect 42610 373232 42616 373244
rect 42116 373204 42616 373232
rect 42116 373192 42122 373204
rect 42610 373192 42616 373204
rect 42668 373192 42674 373244
rect 674742 372512 674748 372564
rect 674800 372552 674806 372564
rect 675294 372552 675300 372564
rect 674800 372524 675300 372552
rect 674800 372512 674806 372524
rect 675294 372512 675300 372524
rect 675352 372512 675358 372564
rect 37918 372308 37924 372360
rect 37976 372348 37982 372360
rect 41690 372348 41696 372360
rect 37976 372320 41696 372348
rect 37976 372308 37982 372320
rect 41690 372308 41696 372320
rect 41748 372308 41754 372360
rect 651466 370948 651472 371000
rect 651524 370988 651530 371000
rect 654778 370988 654784 371000
rect 651524 370960 654784 370988
rect 651524 370948 651530 370960
rect 654778 370948 654784 370960
rect 654836 370948 654842 371000
rect 45370 361496 45376 361548
rect 45428 361536 45434 361548
rect 62114 361536 62120 361548
rect 45428 361508 62120 361536
rect 45428 361496 45434 361508
rect 62114 361496 62120 361508
rect 62172 361496 62178 361548
rect 46750 360136 46756 360188
rect 46808 360176 46814 360188
rect 62114 360176 62120 360188
rect 46808 360148 62120 360176
rect 46808 360136 46814 360148
rect 62114 360136 62120 360148
rect 62172 360136 62178 360188
rect 42150 359932 42156 359984
rect 42208 359972 42214 359984
rect 42794 359972 42800 359984
rect 42208 359944 42800 359972
rect 42208 359932 42214 359944
rect 42794 359932 42800 359944
rect 42852 359932 42858 359984
rect 44634 359048 44640 359100
rect 44692 359088 44698 359100
rect 45370 359088 45376 359100
rect 44692 359060 45376 359088
rect 44692 359048 44698 359060
rect 45370 359048 45376 359060
rect 45428 359048 45434 359100
rect 51718 357416 51724 357468
rect 51776 357456 51782 357468
rect 62114 357456 62120 357468
rect 51776 357428 62120 357456
rect 51776 357416 51782 357428
rect 62114 357416 62120 357428
rect 62172 357416 62178 357468
rect 47946 355988 47952 356040
rect 48004 356028 48010 356040
rect 62114 356028 62120 356040
rect 48004 356000 62120 356028
rect 48004 355988 48010 356000
rect 62114 355988 62120 356000
rect 62172 355988 62178 356040
rect 44634 354968 44640 355020
rect 44692 355008 44698 355020
rect 44692 354980 44895 355008
rect 44692 354968 44698 354980
rect 44640 354680 44692 354686
rect 44640 354622 44692 354628
rect 44732 354476 44784 354482
rect 44732 354418 44784 354424
rect 44867 354314 44895 354980
rect 45278 354396 45284 354408
rect 44974 354368 45284 354396
rect 44974 354110 45002 354368
rect 45278 354356 45284 354368
rect 45336 354356 45342 354408
rect 45278 353920 45284 353932
rect 45105 353892 45284 353920
rect 45278 353880 45284 353892
rect 45336 353880 45342 353932
rect 45297 353716 45303 353728
rect 45218 353688 45303 353716
rect 45297 353676 45303 353688
rect 45355 353676 45361 353728
rect 45830 353512 45836 353524
rect 45329 353484 45836 353512
rect 45830 353472 45836 353484
rect 45888 353472 45894 353524
rect 45422 353252 45474 353258
rect 45422 353194 45474 353200
rect 35802 344564 35808 344616
rect 35860 344604 35866 344616
rect 40034 344604 40040 344616
rect 35860 344576 40040 344604
rect 35860 344564 35866 344576
rect 40034 344564 40040 344576
rect 40092 344564 40098 344616
rect 35526 343748 35532 343800
rect 35584 343788 35590 343800
rect 39850 343788 39856 343800
rect 35584 343760 39856 343788
rect 35584 343748 35590 343760
rect 39850 343748 39856 343760
rect 39908 343748 39914 343800
rect 35802 342184 35808 342236
rect 35860 342224 35866 342236
rect 40218 342224 40224 342236
rect 35860 342196 40224 342224
rect 35860 342184 35866 342196
rect 40218 342184 40224 342196
rect 40276 342184 40282 342236
rect 45462 342184 45468 342236
rect 45520 342224 45526 342236
rect 62298 342224 62304 342236
rect 45520 342196 62304 342224
rect 45520 342184 45526 342196
rect 62298 342184 62304 342196
rect 62356 342184 62362 342236
rect 35802 341164 35808 341216
rect 35860 341204 35866 341216
rect 40218 341204 40224 341216
rect 35860 341176 40224 341204
rect 35860 341164 35866 341176
rect 40218 341164 40224 341176
rect 40276 341164 40282 341216
rect 35618 341028 35624 341080
rect 35676 341068 35682 341080
rect 39666 341068 39672 341080
rect 35676 341040 39672 341068
rect 35676 341028 35682 341040
rect 39666 341028 39672 341040
rect 39724 341028 39730 341080
rect 35526 339600 35532 339652
rect 35584 339640 35590 339652
rect 36538 339640 36544 339652
rect 35584 339612 36544 339640
rect 35584 339600 35590 339612
rect 36538 339600 36544 339612
rect 36596 339600 36602 339652
rect 35802 339464 35808 339516
rect 35860 339504 35866 339516
rect 38562 339504 38568 339516
rect 35860 339476 38568 339504
rect 35860 339464 35866 339476
rect 38562 339464 38568 339476
rect 38620 339464 38626 339516
rect 660298 338716 660304 338768
rect 660356 338756 660362 338768
rect 669314 338756 669320 338768
rect 660356 338728 669320 338756
rect 660356 338716 660362 338728
rect 669314 338716 669320 338728
rect 669372 338716 669378 338768
rect 674374 336676 674380 336728
rect 674432 336716 674438 336728
rect 675110 336716 675116 336728
rect 674432 336688 675116 336716
rect 674432 336676 674438 336688
rect 675110 336676 675116 336688
rect 675168 336676 675174 336728
rect 674374 336472 674380 336524
rect 674432 336512 674438 336524
rect 675294 336512 675300 336524
rect 674432 336484 675300 336512
rect 674432 336472 674438 336484
rect 675294 336472 675300 336484
rect 675352 336472 675358 336524
rect 35802 336200 35808 336252
rect 35860 336240 35866 336252
rect 40034 336240 40040 336252
rect 35860 336212 40040 336240
rect 35860 336200 35866 336212
rect 40034 336200 40040 336212
rect 40092 336200 40098 336252
rect 35526 335316 35532 335368
rect 35584 335356 35590 335368
rect 40218 335356 40224 335368
rect 35584 335328 40224 335356
rect 35584 335316 35590 335328
rect 40218 335316 40224 335328
rect 40276 335316 40282 335368
rect 35802 334092 35808 334144
rect 35860 334132 35866 334144
rect 39758 334132 39764 334144
rect 35860 334104 39764 334132
rect 35860 334092 35866 334104
rect 39758 334092 39764 334104
rect 39816 334092 39822 334144
rect 674466 331100 674472 331152
rect 674524 331140 674530 331152
rect 675294 331140 675300 331152
rect 674524 331112 675300 331140
rect 674524 331100 674530 331112
rect 675294 331100 675300 331112
rect 675352 331100 675358 331152
rect 651466 328380 651472 328432
rect 651524 328420 651530 328432
rect 667382 328420 667388 328432
rect 651524 328392 667388 328420
rect 651524 328380 651530 328392
rect 667382 328380 667388 328392
rect 667440 328380 667446 328432
rect 651374 325592 651380 325644
rect 651432 325632 651438 325644
rect 653398 325632 653404 325644
rect 651432 325604 653404 325632
rect 651432 325592 651438 325604
rect 653398 325592 653404 325604
rect 653456 325592 653462 325644
rect 42242 319880 42248 319932
rect 42300 319920 42306 319932
rect 43346 319920 43352 319932
rect 42300 319892 43352 319920
rect 42300 319880 42306 319892
rect 43346 319880 43352 319892
rect 43404 319880 43410 319932
rect 53834 317364 53840 317416
rect 53892 317404 53898 317416
rect 62114 317404 62120 317416
rect 53892 317376 62120 317404
rect 53892 317364 53898 317376
rect 62114 317364 62120 317376
rect 62172 317364 62178 317416
rect 53098 315936 53104 315988
rect 53156 315976 53162 315988
rect 62114 315976 62120 315988
rect 53156 315948 62120 315976
rect 53156 315936 53162 315948
rect 62114 315936 62120 315948
rect 62172 315936 62178 315988
rect 53834 314712 53840 314764
rect 53892 314752 53898 314764
rect 62114 314752 62120 314764
rect 53892 314724 62120 314752
rect 53892 314712 53898 314724
rect 62114 314712 62120 314724
rect 62172 314712 62178 314764
rect 652018 313896 652024 313948
rect 652076 313936 652082 313948
rect 660298 313936 660304 313948
rect 652076 313908 660304 313936
rect 652076 313896 652082 313908
rect 660298 313896 660304 313908
rect 660356 313896 660362 313948
rect 674558 311992 674564 312044
rect 674616 312032 674622 312044
rect 675478 312032 675484 312044
rect 674616 312004 675484 312032
rect 674616 311992 674622 312004
rect 675478 311992 675484 312004
rect 675536 311992 675542 312044
rect 674834 306348 674840 306400
rect 674892 306388 674898 306400
rect 675478 306388 675484 306400
rect 674892 306360 675484 306388
rect 674892 306348 674898 306360
rect 675478 306348 675484 306360
rect 675536 306348 675542 306400
rect 676214 306348 676220 306400
rect 676272 306388 676278 306400
rect 676858 306388 676864 306400
rect 676272 306360 676864 306388
rect 676272 306348 676278 306360
rect 676858 306348 676864 306360
rect 676916 306348 676922 306400
rect 675846 304852 675852 304904
rect 675904 304892 675910 304904
rect 676398 304892 676404 304904
rect 675904 304864 676404 304892
rect 675904 304852 675910 304864
rect 676398 304852 676404 304864
rect 676456 304852 676462 304904
rect 651466 302132 651472 302184
rect 651524 302172 651530 302184
rect 667382 302172 667388 302184
rect 651524 302144 667388 302172
rect 651524 302132 651530 302144
rect 667382 302132 667388 302144
rect 667440 302132 667446 302184
rect 47578 301724 47584 301776
rect 47636 301764 47642 301776
rect 51902 301764 51908 301776
rect 47636 301736 51908 301764
rect 47636 301724 47642 301736
rect 51902 301724 51908 301736
rect 51960 301724 51966 301776
rect 651466 300772 651472 300824
rect 651524 300812 651530 300824
rect 660298 300812 660304 300824
rect 651524 300784 660304 300812
rect 651524 300772 651530 300784
rect 660298 300772 660304 300784
rect 660356 300772 660362 300824
rect 35618 298732 35624 298784
rect 35676 298772 35682 298784
rect 41598 298772 41604 298784
rect 35676 298744 41604 298772
rect 35676 298732 35682 298744
rect 41598 298732 41604 298744
rect 41656 298732 41662 298784
rect 35802 298256 35808 298308
rect 35860 298296 35866 298308
rect 41598 298296 41604 298308
rect 35860 298268 41604 298296
rect 35860 298256 35866 298268
rect 41598 298256 41604 298268
rect 41656 298256 41662 298308
rect 676122 298052 676128 298104
rect 676180 298092 676186 298104
rect 678238 298092 678244 298104
rect 676180 298064 678244 298092
rect 676180 298052 676186 298064
rect 678238 298052 678244 298064
rect 678296 298052 678302 298104
rect 678974 298092 678980 298104
rect 678946 298052 678980 298092
rect 679032 298052 679038 298104
rect 675938 297916 675944 297968
rect 675996 297956 676002 297968
rect 678946 297956 678974 298052
rect 675996 297928 678974 297956
rect 675996 297916 676002 297928
rect 675018 297304 675024 297356
rect 675076 297304 675082 297356
rect 675036 297016 675064 297304
rect 675202 297100 675208 297152
rect 675260 297100 675266 297152
rect 675018 296964 675024 297016
rect 675076 296964 675082 297016
rect 674834 296828 674840 296880
rect 674892 296868 674898 296880
rect 675220 296868 675248 297100
rect 674892 296840 675248 296868
rect 674892 296828 674898 296840
rect 651742 296760 651748 296812
rect 651800 296800 651806 296812
rect 651800 296772 654134 296800
rect 651800 296760 651806 296772
rect 35802 296692 35808 296744
rect 35860 296732 35866 296744
rect 41598 296732 41604 296744
rect 35860 296704 41604 296732
rect 35860 296692 35866 296704
rect 41598 296692 41604 296704
rect 41656 296692 41662 296744
rect 654106 296732 654134 296772
rect 665818 296732 665824 296744
rect 654106 296704 665824 296732
rect 665818 296692 665824 296704
rect 665876 296692 665882 296744
rect 674466 295672 674472 295724
rect 674524 295712 674530 295724
rect 675478 295712 675484 295724
rect 674524 295684 675484 295712
rect 674524 295672 674530 295684
rect 675478 295672 675484 295684
rect 675536 295672 675542 295724
rect 35618 295468 35624 295520
rect 35676 295508 35682 295520
rect 39298 295508 39304 295520
rect 35676 295480 39304 295508
rect 35676 295468 35682 295480
rect 39298 295468 39304 295480
rect 39356 295468 39362 295520
rect 35802 295332 35808 295384
rect 35860 295372 35866 295384
rect 41322 295372 41328 295384
rect 35860 295344 41328 295372
rect 35860 295332 35866 295344
rect 41322 295332 41328 295344
rect 41380 295332 41386 295384
rect 51902 295060 51908 295112
rect 51960 295100 51966 295112
rect 56502 295100 56508 295112
rect 51960 295072 56508 295100
rect 51960 295060 51966 295072
rect 56502 295060 56508 295072
rect 56560 295060 56566 295112
rect 35434 294584 35440 294636
rect 35492 294624 35498 294636
rect 41690 294624 41696 294636
rect 35492 294596 41696 294624
rect 35492 294584 35498 294596
rect 41690 294584 41696 294596
rect 41748 294584 41754 294636
rect 35802 293972 35808 294024
rect 35860 294012 35866 294024
rect 40034 294012 40040 294024
rect 35860 293984 40040 294012
rect 35860 293972 35866 293984
rect 40034 293972 40040 293984
rect 40092 293972 40098 294024
rect 53098 293972 53104 294024
rect 53156 294012 53162 294024
rect 62206 294012 62212 294024
rect 53156 293984 62212 294012
rect 53156 293972 53162 293984
rect 62206 293972 62212 293984
rect 62264 293972 62270 294024
rect 651466 293972 651472 294024
rect 651524 294012 651530 294024
rect 664438 294012 664444 294024
rect 651524 293984 664444 294012
rect 651524 293972 651530 293984
rect 664438 293972 664444 293984
rect 664496 293972 664502 294024
rect 35802 292884 35808 292936
rect 35860 292924 35866 292936
rect 35860 292884 35894 292924
rect 35866 292856 35894 292884
rect 39850 292856 39856 292868
rect 35866 292828 39856 292856
rect 39850 292816 39856 292828
rect 39908 292816 39914 292868
rect 36004 292624 38654 292652
rect 35802 292544 35808 292596
rect 35860 292584 35866 292596
rect 36004 292584 36032 292624
rect 35860 292556 36032 292584
rect 35860 292544 35866 292556
rect 38626 292380 38654 292624
rect 54478 292544 54484 292596
rect 54536 292584 54542 292596
rect 62298 292584 62304 292596
rect 54536 292556 62304 292584
rect 54536 292544 54542 292556
rect 62298 292544 62304 292556
rect 62356 292544 62362 292596
rect 46198 292408 46204 292460
rect 46256 292448 46262 292460
rect 62114 292448 62120 292460
rect 46256 292420 62120 292448
rect 46256 292408 46262 292420
rect 62114 292408 62120 292420
rect 62172 292408 62178 292460
rect 41598 292380 41604 292392
rect 38626 292352 41604 292380
rect 41598 292340 41604 292352
rect 41656 292340 41662 292392
rect 40770 292068 40776 292120
rect 40828 292108 40834 292120
rect 41598 292108 41604 292120
rect 40828 292080 41604 292108
rect 40828 292068 40834 292080
rect 41598 292068 41604 292080
rect 41656 292068 41662 292120
rect 649258 291864 649264 291916
rect 649316 291904 649322 291916
rect 652018 291904 652024 291916
rect 649316 291876 652024 291904
rect 649316 291864 649322 291876
rect 652018 291864 652024 291876
rect 652076 291864 652082 291916
rect 40034 291320 40040 291372
rect 40092 291360 40098 291372
rect 41690 291360 41696 291372
rect 40092 291332 41696 291360
rect 40092 291320 40098 291332
rect 41690 291320 41696 291332
rect 41748 291320 41754 291372
rect 42150 291320 42156 291372
rect 42208 291360 42214 291372
rect 43346 291360 43352 291372
rect 42208 291332 43352 291360
rect 42208 291320 42214 291332
rect 43346 291320 43352 291332
rect 43404 291320 43410 291372
rect 42058 291184 42064 291236
rect 42116 291224 42122 291236
rect 42610 291224 42616 291236
rect 42116 291196 42616 291224
rect 42116 291184 42122 291196
rect 42610 291184 42616 291196
rect 42668 291184 42674 291236
rect 39850 291116 39856 291168
rect 39908 291156 39914 291168
rect 41598 291156 41604 291168
rect 39908 291128 41604 291156
rect 39908 291116 39914 291128
rect 41598 291116 41604 291128
rect 41656 291116 41662 291168
rect 59998 291116 60004 291168
rect 60056 291156 60062 291168
rect 62298 291156 62304 291168
rect 60056 291128 62304 291156
rect 60056 291116 60062 291128
rect 62298 291116 62304 291128
rect 62356 291116 62362 291168
rect 651466 289824 651472 289876
rect 651524 289864 651530 289876
rect 663058 289864 663064 289876
rect 651524 289836 663064 289864
rect 651524 289824 651530 289836
rect 663058 289824 663064 289836
rect 663116 289824 663122 289876
rect 56502 289756 56508 289808
rect 56560 289796 56566 289808
rect 58802 289796 58808 289808
rect 56560 289768 58808 289796
rect 56560 289756 56566 289768
rect 58802 289756 58808 289768
rect 58860 289756 58866 289808
rect 59998 288464 60004 288516
rect 60056 288504 60062 288516
rect 62114 288504 62120 288516
rect 60056 288476 62120 288504
rect 60056 288464 60062 288476
rect 62114 288464 62120 288476
rect 62172 288464 62178 288516
rect 651466 288396 651472 288448
rect 651524 288436 651530 288448
rect 672074 288436 672080 288448
rect 651524 288408 672080 288436
rect 651524 288396 651530 288408
rect 672074 288396 672080 288408
rect 672132 288396 672138 288448
rect 651650 287648 651656 287700
rect 651708 287688 651714 287700
rect 672442 287688 672448 287700
rect 651708 287660 672448 287688
rect 651708 287648 651714 287660
rect 672442 287648 672448 287660
rect 672500 287648 672506 287700
rect 31018 286288 31024 286340
rect 31076 286328 31082 286340
rect 41506 286328 41512 286340
rect 31076 286300 41512 286328
rect 31076 286288 31082 286300
rect 41506 286288 41512 286300
rect 41564 286288 41570 286340
rect 46198 285676 46204 285728
rect 46256 285716 46262 285728
rect 62114 285716 62120 285728
rect 46256 285688 62120 285716
rect 46256 285676 46262 285688
rect 62114 285676 62120 285688
rect 62172 285676 62178 285728
rect 651466 285676 651472 285728
rect 651524 285716 651530 285728
rect 672258 285716 672264 285728
rect 651524 285688 672264 285716
rect 651524 285676 651530 285688
rect 672258 285676 672264 285688
rect 672316 285676 672322 285728
rect 674650 285132 674656 285184
rect 674708 285132 674714 285184
rect 674668 284980 674696 285132
rect 35802 284928 35808 284980
rect 35860 284968 35866 284980
rect 41690 284968 41696 284980
rect 35860 284940 41696 284968
rect 35860 284928 35866 284940
rect 41690 284928 41696 284940
rect 41748 284928 41754 284980
rect 674650 284928 674656 284980
rect 674708 284928 674714 284980
rect 47578 284316 47584 284368
rect 47636 284356 47642 284368
rect 62942 284356 62948 284368
rect 47636 284328 62948 284356
rect 47636 284316 47642 284328
rect 62942 284316 62948 284328
rect 63000 284316 63006 284368
rect 651466 284316 651472 284368
rect 651524 284356 651530 284368
rect 672258 284356 672264 284368
rect 651524 284328 672264 284356
rect 651524 284316 651530 284328
rect 672258 284316 672264 284328
rect 672316 284316 672322 284368
rect 651466 282888 651472 282940
rect 651524 282928 651530 282940
rect 667382 282928 667388 282940
rect 651524 282900 667388 282928
rect 651524 282888 651530 282900
rect 667382 282888 667388 282900
rect 667440 282888 667446 282940
rect 651466 281528 651472 281580
rect 651524 281568 651530 281580
rect 667750 281568 667756 281580
rect 651524 281540 667756 281568
rect 651524 281528 651530 281540
rect 667750 281528 667756 281540
rect 667808 281528 667814 281580
rect 47946 280168 47952 280220
rect 48004 280208 48010 280220
rect 62114 280208 62120 280220
rect 48004 280180 62120 280208
rect 48004 280168 48010 280180
rect 62114 280168 62120 280180
rect 62172 280168 62178 280220
rect 651466 280168 651472 280220
rect 651524 280208 651530 280220
rect 667566 280208 667572 280220
rect 651524 280180 667572 280208
rect 651524 280168 651530 280180
rect 667566 280168 667572 280180
rect 667624 280168 667630 280220
rect 47762 278672 47768 278724
rect 47820 278712 47826 278724
rect 650822 278712 650828 278724
rect 47820 278684 650828 278712
rect 47820 278672 47826 278684
rect 650822 278672 650828 278684
rect 650880 278672 650886 278724
rect 62850 278536 62856 278588
rect 62908 278576 62914 278588
rect 672626 278576 672632 278588
rect 62908 278548 672632 278576
rect 62908 278536 62914 278548
rect 672626 278536 672632 278548
rect 672684 278536 672690 278588
rect 58802 278400 58808 278452
rect 58860 278440 58866 278452
rect 650638 278440 650644 278452
rect 58860 278412 650644 278440
rect 58860 278400 58866 278412
rect 650638 278400 650644 278412
rect 650696 278400 650702 278452
rect 50706 278264 50712 278316
rect 50764 278304 50770 278316
rect 649258 278304 649264 278316
rect 50764 278276 649264 278304
rect 50764 278264 50770 278276
rect 649258 278264 649264 278276
rect 649316 278264 649322 278316
rect 63218 278128 63224 278180
rect 63276 278168 63282 278180
rect 667198 278168 667204 278180
rect 63276 278140 667204 278168
rect 63276 278128 63282 278140
rect 667198 278128 667204 278140
rect 667256 278128 667262 278180
rect 503530 277380 503536 277432
rect 503588 277420 503594 277432
rect 587066 277420 587072 277432
rect 503588 277392 587072 277420
rect 503588 277380 503594 277392
rect 587066 277380 587072 277392
rect 587124 277380 587130 277432
rect 484026 277176 484032 277228
rect 484084 277216 484090 277228
rect 561122 277216 561128 277228
rect 484084 277188 561128 277216
rect 484084 277176 484090 277188
rect 561122 277176 561128 277188
rect 561180 277176 561186 277228
rect 485498 277040 485504 277092
rect 485556 277080 485562 277092
rect 562318 277080 562324 277092
rect 485556 277052 562324 277080
rect 485556 277040 485562 277052
rect 562318 277040 562324 277052
rect 562376 277040 562382 277092
rect 495066 276904 495072 276956
rect 495124 276944 495130 276956
rect 576486 276944 576492 276956
rect 495124 276916 576492 276944
rect 495124 276904 495130 276916
rect 576486 276904 576492 276916
rect 576544 276904 576550 276956
rect 514478 276768 514484 276820
rect 514536 276808 514542 276820
rect 603626 276808 603632 276820
rect 514536 276780 603632 276808
rect 514536 276768 514542 276780
rect 603626 276768 603632 276780
rect 603684 276768 603690 276820
rect 521102 276632 521108 276684
rect 521160 276672 521166 276684
rect 613102 276672 613108 276684
rect 521160 276644 613108 276672
rect 521160 276632 521166 276644
rect 613102 276632 613108 276644
rect 613160 276632 613166 276684
rect 479978 276496 479984 276548
rect 480036 276536 480042 276548
rect 554038 276536 554044 276548
rect 480036 276508 554044 276536
rect 480036 276496 480042 276508
rect 554038 276496 554044 276508
rect 554096 276496 554102 276548
rect 478506 276360 478512 276412
rect 478564 276400 478570 276412
rect 551646 276400 551652 276412
rect 478564 276372 551652 276400
rect 478564 276360 478570 276372
rect 551646 276360 551652 276372
rect 551704 276360 551710 276412
rect 470410 276224 470416 276276
rect 470468 276264 470474 276276
rect 539870 276264 539876 276276
rect 470468 276236 539876 276264
rect 470468 276224 470474 276236
rect 539870 276224 539876 276236
rect 539928 276224 539934 276276
rect 107194 275952 107200 276004
rect 107252 275992 107258 276004
rect 163498 275992 163504 276004
rect 107252 275964 163504 275992
rect 107252 275952 107258 275964
rect 163498 275952 163504 275964
rect 163556 275952 163562 276004
rect 167546 275952 167552 276004
rect 167604 275992 167610 276004
rect 178678 275992 178684 276004
rect 167604 275964 178684 275992
rect 167604 275952 167610 275964
rect 178678 275952 178684 275964
rect 178736 275952 178742 276004
rect 185210 275952 185216 276004
rect 185268 275992 185274 276004
rect 221274 275992 221280 276004
rect 185268 275964 221280 275992
rect 185268 275952 185274 275964
rect 221274 275952 221280 275964
rect 221332 275952 221338 276004
rect 410794 275952 410800 276004
rect 410852 275992 410858 276004
rect 455874 275992 455880 276004
rect 410852 275964 455880 275992
rect 410852 275952 410858 275964
rect 455874 275952 455880 275964
rect 455932 275952 455938 276004
rect 456426 275952 456432 276004
rect 456484 275992 456490 276004
rect 509050 275992 509056 276004
rect 456484 275964 509056 275992
rect 456484 275952 456490 275964
rect 509050 275952 509056 275964
rect 509108 275952 509114 276004
rect 513190 275952 513196 276004
rect 513248 275992 513254 276004
rect 601326 275992 601332 276004
rect 513248 275964 601332 275992
rect 513248 275952 513254 275964
rect 601326 275952 601332 275964
rect 601384 275952 601390 276004
rect 139118 275816 139124 275868
rect 139176 275856 139182 275868
rect 174262 275856 174268 275868
rect 139176 275828 174268 275856
rect 139176 275816 139182 275828
rect 174262 275816 174268 275828
rect 174320 275816 174326 275868
rect 178126 275816 178132 275868
rect 178184 275856 178190 275868
rect 216674 275856 216680 275868
rect 178184 275828 216680 275856
rect 178184 275816 178190 275828
rect 216674 275816 216680 275828
rect 216732 275816 216738 275868
rect 224218 275816 224224 275868
rect 224276 275856 224282 275868
rect 233050 275856 233056 275868
rect 224276 275828 233056 275856
rect 224276 275816 224282 275828
rect 233050 275816 233056 275828
rect 233108 275816 233114 275868
rect 236086 275816 236092 275868
rect 236144 275856 236150 275868
rect 250438 275856 250444 275868
rect 236144 275828 250444 275856
rect 236144 275816 236150 275828
rect 250438 275816 250444 275828
rect 250496 275816 250502 275868
rect 284570 275816 284576 275868
rect 284628 275856 284634 275868
rect 290090 275856 290096 275868
rect 284628 275828 290096 275856
rect 284628 275816 284634 275828
rect 290090 275816 290096 275828
rect 290148 275816 290154 275868
rect 430206 275816 430212 275868
rect 430264 275856 430270 275868
rect 484302 275856 484308 275868
rect 430264 275828 484308 275856
rect 430264 275816 430270 275828
rect 484302 275816 484308 275828
rect 484360 275816 484366 275868
rect 485038 275816 485044 275868
rect 485096 275856 485102 275868
rect 491386 275856 491392 275868
rect 485096 275828 491392 275856
rect 485096 275816 485102 275828
rect 491386 275816 491392 275828
rect 491444 275816 491450 275868
rect 522758 275816 522764 275868
rect 522816 275856 522822 275868
rect 615494 275856 615500 275868
rect 522816 275828 615500 275856
rect 522816 275816 522822 275828
rect 615494 275816 615500 275828
rect 615552 275816 615558 275868
rect 260926 275748 260932 275800
rect 260984 275788 260990 275800
rect 266354 275788 266360 275800
rect 260984 275760 266360 275788
rect 260984 275748 260990 275760
rect 266354 275748 266360 275760
rect 266412 275748 266418 275800
rect 93026 275680 93032 275732
rect 93084 275720 93090 275732
rect 152826 275720 152832 275732
rect 93084 275692 152832 275720
rect 93084 275680 93090 275692
rect 152826 275680 152832 275692
rect 152884 275680 152890 275732
rect 160462 275680 160468 275732
rect 160520 275720 160526 275732
rect 199378 275720 199384 275732
rect 160520 275692 199384 275720
rect 160520 275680 160526 275692
rect 199378 275680 199384 275692
rect 199436 275680 199442 275732
rect 217134 275680 217140 275732
rect 217192 275720 217198 275732
rect 224218 275720 224224 275732
rect 217192 275692 224224 275720
rect 217192 275680 217198 275692
rect 224218 275680 224224 275692
rect 224276 275680 224282 275732
rect 229002 275680 229008 275732
rect 229060 275720 229066 275732
rect 243722 275720 243728 275732
rect 229060 275692 243728 275720
rect 229060 275680 229066 275692
rect 243722 275680 243728 275692
rect 243780 275680 243786 275732
rect 250254 275680 250260 275732
rect 250312 275720 250318 275732
rect 259362 275720 259368 275732
rect 250312 275692 259368 275720
rect 250312 275680 250318 275692
rect 259362 275680 259368 275692
rect 259420 275680 259426 275732
rect 286870 275680 286876 275732
rect 286928 275720 286934 275732
rect 291838 275720 291844 275732
rect 286928 275692 291844 275720
rect 286928 275680 286934 275692
rect 291838 275680 291844 275692
rect 291896 275680 291902 275732
rect 416406 275680 416412 275732
rect 416464 275720 416470 275732
rect 462958 275720 462964 275732
rect 416464 275692 462964 275720
rect 416464 275680 416470 275692
rect 462958 275680 462964 275692
rect 463016 275680 463022 275732
rect 463142 275680 463148 275732
rect 463200 275720 463206 275732
rect 516226 275720 516232 275732
rect 463200 275692 516232 275720
rect 463200 275680 463206 275692
rect 516226 275680 516232 275692
rect 516284 275680 516290 275732
rect 528186 275680 528192 275732
rect 528244 275720 528250 275732
rect 622578 275720 622584 275732
rect 528244 275692 622584 275720
rect 528244 275680 528250 275692
rect 622578 275680 622584 275692
rect 622636 275680 622642 275732
rect 76466 275544 76472 275596
rect 76524 275584 76530 275596
rect 86218 275584 86224 275596
rect 76524 275556 86224 275584
rect 76524 275544 76530 275556
rect 86218 275544 86224 275556
rect 86276 275544 86282 275596
rect 90726 275544 90732 275596
rect 90784 275584 90790 275596
rect 154758 275584 154764 275596
rect 90784 275556 154764 275584
rect 90784 275544 90790 275556
rect 154758 275544 154764 275556
rect 154816 275544 154822 275596
rect 171042 275544 171048 275596
rect 171100 275584 171106 275596
rect 211430 275584 211436 275596
rect 171100 275556 211436 275584
rect 171100 275544 171106 275556
rect 211430 275544 211436 275556
rect 211488 275544 211494 275596
rect 218330 275544 218336 275596
rect 218388 275584 218394 275596
rect 233878 275584 233884 275596
rect 218388 275556 233884 275584
rect 218388 275544 218394 275556
rect 233878 275544 233884 275556
rect 233936 275544 233942 275596
rect 239582 275544 239588 275596
rect 239640 275584 239646 275596
rect 255958 275584 255964 275596
rect 239640 275556 255964 275584
rect 239640 275544 239646 275556
rect 255958 275544 255964 275556
rect 256016 275544 256022 275596
rect 257338 275544 257344 275596
rect 257396 275584 257402 275596
rect 262306 275584 262312 275596
rect 257396 275556 262312 275584
rect 257396 275544 257402 275556
rect 262306 275544 262312 275556
rect 262364 275544 262370 275596
rect 266814 275544 266820 275596
rect 266872 275584 266878 275596
rect 276474 275584 276480 275596
rect 266872 275556 276480 275584
rect 266872 275544 266878 275556
rect 276474 275544 276480 275556
rect 276532 275544 276538 275596
rect 363874 275544 363880 275596
rect 363932 275584 363938 275596
rect 388530 275584 388536 275596
rect 363932 275556 388536 275584
rect 363932 275544 363938 275556
rect 388530 275544 388536 275556
rect 388588 275544 388594 275596
rect 445018 275544 445024 275596
rect 445076 275584 445082 275596
rect 498470 275584 498476 275596
rect 445076 275556 498476 275584
rect 445076 275544 445082 275556
rect 498470 275544 498476 275556
rect 498528 275544 498534 275596
rect 498838 275544 498844 275596
rect 498896 275584 498902 275596
rect 505554 275584 505560 275596
rect 498896 275556 505560 275584
rect 498896 275544 498902 275556
rect 505554 275544 505560 275556
rect 505612 275544 505618 275596
rect 505738 275544 505744 275596
rect 505796 275584 505802 275596
rect 512638 275584 512644 275596
rect 505796 275556 512644 275584
rect 505796 275544 505802 275556
rect 512638 275544 512644 275556
rect 512696 275544 512702 275596
rect 516778 275544 516784 275596
rect 516836 275584 516842 275596
rect 526806 275584 526812 275596
rect 516836 275556 526812 275584
rect 516836 275544 516842 275556
rect 526806 275544 526812 275556
rect 526864 275544 526870 275596
rect 532326 275544 532332 275596
rect 532384 275584 532390 275596
rect 629662 275584 629668 275596
rect 532384 275556 629668 275584
rect 532384 275544 532390 275556
rect 629662 275544 629668 275556
rect 629720 275544 629726 275596
rect 277486 275476 277492 275528
rect 277544 275516 277550 275528
rect 285122 275516 285128 275528
rect 277544 275488 285128 275516
rect 277544 275476 277550 275488
rect 285122 275476 285128 275488
rect 285180 275476 285186 275528
rect 100110 275408 100116 275460
rect 100168 275448 100174 275460
rect 100168 275420 142154 275448
rect 100168 275408 100174 275420
rect 71774 275272 71780 275324
rect 71832 275312 71838 275324
rect 141050 275312 141056 275324
rect 71832 275284 141056 275312
rect 71832 275272 71838 275284
rect 141050 275272 141056 275284
rect 141108 275272 141114 275324
rect 142126 275312 142154 275420
rect 156874 275408 156880 275460
rect 156932 275448 156938 275460
rect 156932 275420 161474 275448
rect 156932 275408 156938 275420
rect 159450 275312 159456 275324
rect 142126 275284 159456 275312
rect 159450 275272 159456 275284
rect 159508 275272 159514 275324
rect 161446 275312 161474 275420
rect 163958 275408 163964 275460
rect 164016 275448 164022 275460
rect 206370 275448 206376 275460
rect 164016 275420 206376 275448
rect 164016 275408 164022 275420
rect 206370 275408 206376 275420
rect 206428 275408 206434 275460
rect 221918 275408 221924 275460
rect 221976 275448 221982 275460
rect 243538 275448 243544 275460
rect 221976 275420 243544 275448
rect 221976 275408 221982 275420
rect 243538 275408 243544 275420
rect 243596 275408 243602 275460
rect 256142 275408 256148 275460
rect 256200 275448 256206 275460
rect 269390 275448 269396 275460
rect 256200 275420 269396 275448
rect 256200 275408 256206 275420
rect 269390 275408 269396 275420
rect 269448 275408 269454 275460
rect 285674 275408 285680 275460
rect 285732 275448 285738 275460
rect 291194 275448 291200 275460
rect 285732 275420 291200 275448
rect 285732 275408 285738 275420
rect 291194 275408 291200 275420
rect 291252 275408 291258 275460
rect 358630 275408 358636 275460
rect 358688 275448 358694 275460
rect 381446 275448 381452 275460
rect 358688 275420 381452 275448
rect 358688 275408 358694 275420
rect 381446 275408 381452 275420
rect 381504 275408 381510 275460
rect 385954 275408 385960 275460
rect 386012 275448 386018 275460
rect 420454 275448 420460 275460
rect 386012 275420 420460 275448
rect 386012 275408 386018 275420
rect 420454 275408 420460 275420
rect 420512 275408 420518 275460
rect 435634 275408 435640 275460
rect 435692 275448 435698 275460
rect 485038 275448 485044 275460
rect 435692 275420 485044 275448
rect 435692 275408 435698 275420
rect 485038 275408 485044 275420
rect 485096 275408 485102 275460
rect 485774 275408 485780 275460
rect 485832 275448 485838 275460
rect 530394 275448 530400 275460
rect 485832 275420 530400 275448
rect 485832 275408 485838 275420
rect 530394 275408 530400 275420
rect 530452 275408 530458 275460
rect 537662 275408 537668 275460
rect 537720 275448 537726 275460
rect 636746 275448 636752 275460
rect 537720 275420 636752 275448
rect 537720 275408 537726 275420
rect 636746 275408 636752 275420
rect 636804 275408 636810 275460
rect 299934 275340 299940 275392
rect 299992 275380 299998 275392
rect 301130 275380 301136 275392
rect 299992 275352 301136 275380
rect 299992 275340 299998 275352
rect 301130 275340 301136 275352
rect 301188 275340 301194 275392
rect 200758 275312 200764 275324
rect 161446 275284 200764 275312
rect 200758 275272 200764 275284
rect 200816 275272 200822 275324
rect 214834 275272 214840 275324
rect 214892 275312 214898 275324
rect 239398 275312 239404 275324
rect 214892 275284 239404 275312
rect 214892 275272 214898 275284
rect 239398 275272 239404 275284
rect 239456 275272 239462 275324
rect 243170 275272 243176 275324
rect 243228 275312 243234 275324
rect 256694 275312 256700 275324
rect 243228 275284 256700 275312
rect 243228 275272 243234 275284
rect 256694 275272 256700 275284
rect 256752 275272 256758 275324
rect 263226 275272 263232 275324
rect 263284 275312 263290 275324
rect 273254 275312 273260 275324
rect 263284 275284 273260 275312
rect 263284 275272 263290 275284
rect 273254 275272 273260 275284
rect 273312 275272 273318 275324
rect 276290 275272 276296 275324
rect 276348 275312 276354 275324
rect 283098 275312 283104 275324
rect 276348 275284 283104 275312
rect 276348 275272 276354 275284
rect 283098 275272 283104 275284
rect 283156 275272 283162 275324
rect 291654 275272 291660 275324
rect 291712 275312 291718 275324
rect 295334 275312 295340 275324
rect 291712 275284 295340 275312
rect 291712 275272 291718 275284
rect 295334 275272 295340 275284
rect 295392 275272 295398 275324
rect 326430 275272 326436 275324
rect 326488 275312 326494 275324
rect 335354 275312 335360 275324
rect 326488 275284 335360 275312
rect 326488 275272 326494 275284
rect 335354 275272 335360 275284
rect 335412 275272 335418 275324
rect 371050 275272 371056 275324
rect 371108 275312 371114 275324
rect 399202 275312 399208 275324
rect 371108 275284 399208 275312
rect 371108 275272 371114 275284
rect 399202 275272 399208 275284
rect 399260 275272 399266 275324
rect 418798 275272 418804 275324
rect 418856 275312 418862 275324
rect 466546 275312 466552 275324
rect 418856 275284 466552 275312
rect 418856 275272 418862 275284
rect 466546 275272 466552 275284
rect 466604 275272 466610 275324
rect 467558 275272 467564 275324
rect 467616 275312 467622 275324
rect 537478 275312 537484 275324
rect 467616 275284 537484 275312
rect 467616 275272 467622 275284
rect 537478 275272 537484 275284
rect 537536 275272 537542 275324
rect 542078 275272 542084 275324
rect 542136 275312 542142 275324
rect 643830 275312 643836 275324
rect 542136 275284 643836 275312
rect 542136 275272 542142 275284
rect 643830 275272 643836 275284
rect 643888 275272 643894 275324
rect 298738 275204 298744 275256
rect 298796 275244 298802 275256
rect 300026 275244 300032 275256
rect 298796 275216 300032 275244
rect 298796 275204 298802 275216
rect 300026 275204 300032 275216
rect 300084 275204 300090 275256
rect 96614 275136 96620 275188
rect 96672 275176 96678 275188
rect 149974 275176 149980 275188
rect 96672 275148 149980 275176
rect 96672 275136 96678 275148
rect 149974 275136 149980 275148
rect 150032 275136 150038 275188
rect 153378 275136 153384 275188
rect 153436 275176 153442 275188
rect 169018 275176 169024 275188
rect 153436 275148 169024 275176
rect 153436 275136 153442 275148
rect 169018 275136 169024 275148
rect 169076 275136 169082 275188
rect 189994 275136 190000 275188
rect 190052 275176 190058 275188
rect 222930 275176 222936 275188
rect 190052 275148 222936 275176
rect 190052 275136 190058 275148
rect 222930 275136 222936 275148
rect 222988 275136 222994 275188
rect 232498 275136 232504 275188
rect 232556 275176 232562 275188
rect 240042 275176 240048 275188
rect 232556 275148 240048 275176
rect 232556 275136 232562 275148
rect 240042 275136 240048 275148
rect 240100 275136 240106 275188
rect 292850 275136 292856 275188
rect 292908 275176 292914 275188
rect 295794 275176 295800 275188
rect 292908 275148 295800 275176
rect 292908 275136 292914 275148
rect 295794 275136 295800 275148
rect 295852 275136 295858 275188
rect 427078 275136 427084 275188
rect 427136 275176 427142 275188
rect 477218 275176 477224 275188
rect 427136 275148 477224 275176
rect 427136 275136 427142 275148
rect 477218 275136 477224 275148
rect 477276 275136 477282 275188
rect 507486 275136 507492 275188
rect 507544 275176 507550 275188
rect 594242 275176 594248 275188
rect 507544 275148 594248 275176
rect 507544 275136 507550 275148
rect 594242 275136 594248 275148
rect 594300 275136 594306 275188
rect 269206 275068 269212 275120
rect 269264 275108 269270 275120
rect 274634 275108 274640 275120
rect 269264 275080 274640 275108
rect 269264 275068 269270 275080
rect 274634 275068 274640 275080
rect 274692 275068 274698 275120
rect 81250 275000 81256 275052
rect 81308 275040 81314 275052
rect 145282 275040 145288 275052
rect 81308 275012 145288 275040
rect 81308 275000 81314 275012
rect 145282 275000 145288 275012
rect 145340 275000 145346 275052
rect 149790 275000 149796 275052
rect 149848 275040 149854 275052
rect 189074 275040 189080 275052
rect 149848 275012 189080 275040
rect 149848 275000 149854 275012
rect 189074 275000 189080 275012
rect 189132 275000 189138 275052
rect 288066 275000 288072 275052
rect 288124 275040 288130 275052
rect 292850 275040 292856 275052
rect 288124 275012 292856 275040
rect 288124 275000 288130 275012
rect 292850 275000 292856 275012
rect 292908 275000 292914 275052
rect 420546 275000 420552 275052
rect 420604 275040 420610 275052
rect 470134 275040 470140 275052
rect 420604 275012 470140 275040
rect 420604 275000 420610 275012
rect 470134 275000 470140 275012
rect 470192 275000 470198 275052
rect 497918 275000 497924 275052
rect 497976 275040 497982 275052
rect 579982 275040 579988 275052
rect 497976 275012 579988 275040
rect 497976 275000 497982 275012
rect 579982 275000 579988 275012
rect 580040 275000 580046 275052
rect 293954 274932 293960 274984
rect 294012 274972 294018 274984
rect 297174 274972 297180 274984
rect 294012 274944 297180 274972
rect 294012 274932 294018 274944
rect 297174 274932 297180 274944
rect 297232 274932 297238 274984
rect 136818 274864 136824 274916
rect 136876 274904 136882 274916
rect 137646 274904 137652 274916
rect 136876 274876 137652 274904
rect 136876 274864 136882 274876
rect 137646 274864 137652 274876
rect 137704 274864 137710 274916
rect 146202 274864 146208 274916
rect 146260 274904 146266 274916
rect 185302 274904 185308 274916
rect 146260 274876 185308 274904
rect 146260 274864 146266 274876
rect 185302 274864 185308 274876
rect 185360 274864 185366 274916
rect 289262 274864 289268 274916
rect 289320 274904 289326 274916
rect 292666 274904 292672 274916
rect 289320 274876 292672 274904
rect 289320 274864 289326 274876
rect 292666 274864 292672 274876
rect 292724 274864 292730 274916
rect 473078 274864 473084 274916
rect 473136 274904 473142 274916
rect 544562 274904 544568 274916
rect 473136 274876 544568 274904
rect 473136 274864 473142 274876
rect 544562 274864 544568 274876
rect 544620 274864 544626 274916
rect 296346 274796 296352 274848
rect 296404 274836 296410 274848
rect 298370 274836 298376 274848
rect 296404 274808 298376 274836
rect 296404 274796 296410 274808
rect 298370 274796 298376 274808
rect 298428 274796 298434 274848
rect 128538 274728 128544 274780
rect 128596 274768 128602 274780
rect 166994 274768 167000 274780
rect 128596 274740 167000 274768
rect 128596 274728 128602 274740
rect 166994 274728 167000 274740
rect 167052 274728 167058 274780
rect 207750 274728 207756 274780
rect 207808 274768 207814 274780
rect 210694 274768 210700 274780
rect 207808 274740 210700 274768
rect 207808 274728 207814 274740
rect 210694 274728 210700 274740
rect 210752 274728 210758 274780
rect 476758 274728 476764 274780
rect 476816 274768 476822 274780
rect 523310 274768 523316 274780
rect 476816 274740 523316 274768
rect 476816 274728 476822 274740
rect 523310 274728 523316 274740
rect 523368 274728 523374 274780
rect 523678 274728 523684 274780
rect 523736 274768 523742 274780
rect 533890 274768 533896 274780
rect 523736 274740 533896 274768
rect 523736 274728 523742 274740
rect 533890 274728 533896 274740
rect 533948 274728 533954 274780
rect 534718 274728 534724 274780
rect 534776 274768 534782 274780
rect 540974 274768 540980 274780
rect 534776 274740 540980 274768
rect 534776 274728 534782 274740
rect 540974 274728 540980 274740
rect 541032 274728 541038 274780
rect 74166 274660 74172 274712
rect 74224 274700 74230 274712
rect 76834 274700 76840 274712
rect 74224 274672 76840 274700
rect 74224 274660 74230 274672
rect 76834 274660 76840 274672
rect 76892 274660 76898 274712
rect 85942 274660 85948 274712
rect 86000 274700 86006 274712
rect 90358 274700 90364 274712
rect 86000 274672 90364 274700
rect 86000 274660 86006 274672
rect 90358 274660 90364 274672
rect 90416 274660 90422 274712
rect 103698 274660 103704 274712
rect 103756 274700 103762 274712
rect 104802 274700 104808 274712
rect 103756 274672 104808 274700
rect 103756 274660 103762 274672
rect 104802 274660 104808 274672
rect 104860 274660 104866 274712
rect 110782 274660 110788 274712
rect 110840 274700 110846 274712
rect 111702 274700 111708 274712
rect 110840 274672 111708 274700
rect 110840 274660 110846 274672
rect 111702 274660 111708 274672
rect 111760 274660 111766 274712
rect 253842 274660 253848 274712
rect 253900 274700 253906 274712
rect 256878 274700 256884 274712
rect 253900 274672 256884 274700
rect 253900 274660 253906 274672
rect 256878 274660 256884 274672
rect 256936 274660 256942 274712
rect 275094 274660 275100 274712
rect 275152 274700 275158 274712
rect 278406 274700 278412 274712
rect 275152 274672 278412 274700
rect 275152 274660 275158 274672
rect 278406 274660 278412 274672
rect 278464 274660 278470 274712
rect 283374 274660 283380 274712
rect 283432 274700 283438 274712
rect 289170 274700 289176 274712
rect 283432 274672 289176 274700
rect 283432 274660 283438 274672
rect 289170 274660 289176 274672
rect 289228 274660 289234 274712
rect 290458 274660 290464 274712
rect 290516 274700 290522 274712
rect 294138 274700 294144 274712
rect 290516 274672 294144 274700
rect 290516 274660 290522 274672
rect 294138 274660 294144 274672
rect 294196 274660 294202 274712
rect 295150 274660 295156 274712
rect 295208 274700 295214 274712
rect 296806 274700 296812 274712
rect 295208 274672 296812 274700
rect 295208 274660 295214 274672
rect 296806 274660 296812 274672
rect 296864 274660 296870 274712
rect 297542 274660 297548 274712
rect 297600 274700 297606 274712
rect 299474 274700 299480 274712
rect 297600 274672 299480 274700
rect 297600 274660 297606 274672
rect 299474 274660 299480 274672
rect 299532 274660 299538 274712
rect 303430 274660 303436 274712
rect 303488 274700 303494 274712
rect 303982 274700 303988 274712
rect 303488 274672 303988 274700
rect 303488 274660 303494 274672
rect 303982 274660 303988 274672
rect 304040 274660 304046 274712
rect 321186 274660 321192 274712
rect 321244 274700 321250 274712
rect 328270 274700 328276 274712
rect 321244 274672 328276 274700
rect 321244 274660 321250 274672
rect 328270 274660 328276 274672
rect 328328 274660 328334 274712
rect 114370 274592 114376 274644
rect 114428 274632 114434 274644
rect 171594 274632 171600 274644
rect 114428 274604 171600 274632
rect 114428 274592 114434 274604
rect 171594 274592 171600 274604
rect 171652 274592 171658 274644
rect 179322 274592 179328 274644
rect 179380 274632 179386 274644
rect 214558 274632 214564 274644
rect 179380 274604 214564 274632
rect 179380 274592 179386 274604
rect 214558 274592 214564 274604
rect 214616 274592 214622 274644
rect 409782 274592 409788 274644
rect 409840 274632 409846 274644
rect 453574 274632 453580 274644
rect 409840 274604 453580 274632
rect 409840 274592 409846 274604
rect 453574 274592 453580 274604
rect 453632 274592 453638 274644
rect 460658 274632 460664 274644
rect 455892 274604 460664 274632
rect 101306 274456 101312 274508
rect 101364 274496 101370 274508
rect 160922 274496 160928 274508
rect 101364 274468 160928 274496
rect 101364 274456 101370 274468
rect 160922 274456 160928 274468
rect 160980 274456 160986 274508
rect 168742 274456 168748 274508
rect 168800 274496 168806 274508
rect 208394 274496 208400 274508
rect 168800 274468 208400 274496
rect 168800 274456 168806 274468
rect 208394 274456 208400 274468
rect 208452 274456 208458 274508
rect 381538 274456 381544 274508
rect 381596 274496 381602 274508
rect 392118 274496 392124 274508
rect 381596 274468 392124 274496
rect 381596 274456 381602 274468
rect 392118 274456 392124 274468
rect 392176 274456 392182 274508
rect 413830 274456 413836 274508
rect 413888 274496 413894 274508
rect 455892 274496 455920 274604
rect 460658 274592 460664 274604
rect 460716 274592 460722 274644
rect 464430 274592 464436 274644
rect 464488 274632 464494 274644
rect 480714 274632 480720 274644
rect 464488 274604 480720 274632
rect 464488 274592 464494 274604
rect 480714 274592 480720 274604
rect 480772 274592 480778 274644
rect 486786 274592 486792 274644
rect 486844 274632 486850 274644
rect 563422 274632 563428 274644
rect 486844 274604 563428 274632
rect 486844 274592 486850 274604
rect 563422 274592 563428 274604
rect 563480 274592 563486 274644
rect 413888 274468 455920 274496
rect 413888 274456 413894 274468
rect 456058 274456 456064 274508
rect 456116 274496 456122 274508
rect 465902 274496 465908 274508
rect 456116 274468 465908 274496
rect 456116 274456 456122 274468
rect 465902 274456 465908 274468
rect 465960 274456 465966 274508
rect 466086 274456 466092 274508
rect 466144 274496 466150 274508
rect 485774 274496 485780 274508
rect 466144 274468 485780 274496
rect 466144 274456 466150 274468
rect 485774 274456 485780 274468
rect 485832 274456 485838 274508
rect 488350 274456 488356 274508
rect 488408 274496 488414 274508
rect 567010 274496 567016 274508
rect 488408 274468 567016 274496
rect 488408 274456 488414 274468
rect 567010 274456 567016 274468
rect 567068 274456 567074 274508
rect 95418 274320 95424 274372
rect 95476 274360 95482 274372
rect 157610 274360 157616 274372
rect 95476 274332 157616 274360
rect 95476 274320 95482 274332
rect 157610 274320 157616 274332
rect 157668 274320 157674 274372
rect 159266 274320 159272 274372
rect 159324 274360 159330 274372
rect 202322 274360 202328 274372
rect 159324 274332 202328 274360
rect 159324 274320 159330 274332
rect 202322 274320 202328 274332
rect 202380 274320 202386 274372
rect 223114 274320 223120 274372
rect 223172 274360 223178 274372
rect 247218 274360 247224 274372
rect 223172 274332 247224 274360
rect 223172 274320 223178 274332
rect 247218 274320 247224 274332
rect 247276 274320 247282 274372
rect 368934 274320 368940 274372
rect 368992 274360 368998 274372
rect 387334 274360 387340 274372
rect 368992 274332 387340 274360
rect 368992 274320 368998 274332
rect 387334 274320 387340 274332
rect 387392 274320 387398 274372
rect 419074 274320 419080 274372
rect 419132 274360 419138 274372
rect 467742 274360 467748 274372
rect 419132 274332 467748 274360
rect 419132 274320 419138 274332
rect 467742 274320 467748 274332
rect 467800 274320 467806 274372
rect 474826 274360 474832 274372
rect 470566 274332 474832 274360
rect 331950 274252 331956 274304
rect 332008 274292 332014 274304
rect 337746 274292 337752 274304
rect 332008 274264 337752 274292
rect 332008 274252 332014 274264
rect 337746 274252 337752 274264
rect 337804 274252 337810 274304
rect 67082 274184 67088 274236
rect 67140 274224 67146 274236
rect 130378 274224 130384 274236
rect 67140 274196 130384 274224
rect 67140 274184 67146 274196
rect 130378 274184 130384 274196
rect 130436 274184 130442 274236
rect 130838 274184 130844 274236
rect 130896 274224 130902 274236
rect 182450 274224 182456 274236
rect 130896 274196 182456 274224
rect 130896 274184 130902 274196
rect 182450 274184 182456 274196
rect 182508 274184 182514 274236
rect 193490 274184 193496 274236
rect 193548 274224 193554 274236
rect 226426 274224 226432 274236
rect 193548 274196 226432 274224
rect 193548 274184 193554 274196
rect 226426 274184 226432 274196
rect 226484 274184 226490 274236
rect 240042 274184 240048 274236
rect 240100 274224 240106 274236
rect 253934 274224 253940 274236
rect 240100 274196 253940 274224
rect 240100 274184 240106 274196
rect 253934 274184 253940 274196
rect 253992 274184 253998 274236
rect 359458 274184 359464 274236
rect 359516 274224 359522 274236
rect 380250 274224 380256 274236
rect 359516 274196 380256 274224
rect 359516 274184 359522 274196
rect 380250 274184 380256 274196
rect 380308 274184 380314 274236
rect 388990 274184 388996 274236
rect 389048 274224 389054 274236
rect 425146 274224 425152 274236
rect 389048 274196 425152 274224
rect 389048 274184 389054 274196
rect 425146 274184 425152 274196
rect 425204 274184 425210 274236
rect 425698 274184 425704 274236
rect 425756 274224 425762 274236
rect 470566 274224 470594 274332
rect 474826 274320 474832 274332
rect 474884 274320 474890 274372
rect 506198 274320 506204 274372
rect 506256 274360 506262 274372
rect 591850 274360 591856 274372
rect 506256 274332 591856 274360
rect 506256 274320 506262 274332
rect 591850 274320 591856 274332
rect 591908 274320 591914 274372
rect 425756 274196 470594 274224
rect 425756 274184 425762 274196
rect 472250 274184 472256 274236
rect 472308 274224 472314 274236
rect 472308 274196 480254 274224
rect 472308 274184 472314 274196
rect 77662 274048 77668 274100
rect 77720 274088 77726 274100
rect 144914 274088 144920 274100
rect 77720 274060 144920 274088
rect 77720 274048 77726 274060
rect 144914 274048 144920 274060
rect 144972 274048 144978 274100
rect 154482 274048 154488 274100
rect 154540 274088 154546 274100
rect 198090 274088 198096 274100
rect 154540 274060 198096 274088
rect 154540 274048 154546 274060
rect 198090 274048 198096 274060
rect 198148 274048 198154 274100
rect 210050 274048 210056 274100
rect 210108 274088 210114 274100
rect 237834 274088 237840 274100
rect 210108 274060 237840 274088
rect 210108 274048 210114 274060
rect 237834 274048 237840 274060
rect 237892 274048 237898 274100
rect 249058 274048 249064 274100
rect 249116 274088 249122 274100
rect 265250 274088 265256 274100
rect 249116 274060 265256 274088
rect 249116 274048 249122 274060
rect 265250 274048 265256 274060
rect 265308 274048 265314 274100
rect 266354 274048 266360 274100
rect 266412 274088 266418 274100
rect 273530 274088 273536 274100
rect 266412 274060 273536 274088
rect 266412 274048 266418 274060
rect 273530 274048 273536 274060
rect 273588 274048 273594 274100
rect 278590 274048 278596 274100
rect 278648 274088 278654 274100
rect 285858 274088 285864 274100
rect 278648 274060 285864 274088
rect 278648 274048 278654 274060
rect 285858 274048 285864 274060
rect 285916 274048 285922 274100
rect 337746 274048 337752 274100
rect 337804 274088 337810 274100
rect 351914 274088 351920 274100
rect 337804 274060 351920 274088
rect 337804 274048 337810 274060
rect 351914 274048 351920 274060
rect 351972 274048 351978 274100
rect 353938 274048 353944 274100
rect 353996 274088 354002 274100
rect 369578 274088 369584 274100
rect 353996 274060 369584 274088
rect 353996 274048 354002 274060
rect 369578 274048 369584 274060
rect 369636 274048 369642 274100
rect 373258 274048 373264 274100
rect 373316 274088 373322 274100
rect 400306 274088 400312 274100
rect 373316 274060 400312 274088
rect 373316 274048 373322 274060
rect 400306 274048 400312 274060
rect 400364 274048 400370 274100
rect 401502 274048 401508 274100
rect 401560 274088 401566 274100
rect 442902 274088 442908 274100
rect 401560 274060 442908 274088
rect 401560 274048 401566 274060
rect 442902 274048 442908 274060
rect 442960 274048 442966 274100
rect 451182 274048 451188 274100
rect 451240 274088 451246 274100
rect 456058 274088 456064 274100
rect 451240 274060 456064 274088
rect 451240 274048 451246 274060
rect 456058 274048 456064 274060
rect 456116 274048 456122 274100
rect 456242 274048 456248 274100
rect 456300 274088 456306 274100
rect 480226 274088 480254 274196
rect 481358 274184 481364 274236
rect 481416 274224 481422 274236
rect 485314 274224 485320 274236
rect 481416 274196 485320 274224
rect 481416 274184 481422 274196
rect 485314 274184 485320 274196
rect 485372 274184 485378 274236
rect 511626 274184 511632 274236
rect 511684 274224 511690 274236
rect 598934 274224 598940 274236
rect 511684 274196 598940 274224
rect 511684 274184 511690 274196
rect 598934 274184 598940 274196
rect 598992 274184 598998 274236
rect 513834 274088 513840 274100
rect 456300 274060 474504 274088
rect 480226 274060 513840 274088
rect 456300 274048 456306 274060
rect 69382 273912 69388 273964
rect 69440 273952 69446 273964
rect 139394 273952 139400 273964
rect 69440 273924 139400 273952
rect 69440 273912 69446 273924
rect 139394 273912 139400 273924
rect 139452 273912 139458 273964
rect 148594 273912 148600 273964
rect 148652 273952 148658 273964
rect 194778 273952 194784 273964
rect 148652 273924 194784 273952
rect 148652 273912 148658 273924
rect 194778 273912 194784 273924
rect 194836 273912 194842 273964
rect 208854 273912 208860 273964
rect 208912 273952 208918 273964
rect 237374 273952 237380 273964
rect 208912 273924 237380 273952
rect 208912 273912 208918 273924
rect 237374 273912 237380 273924
rect 237432 273912 237438 273964
rect 238478 273912 238484 273964
rect 238536 273952 238542 273964
rect 238536 273924 238754 273952
rect 238536 273912 238542 273924
rect 88334 273776 88340 273828
rect 88392 273816 88398 273828
rect 119338 273816 119344 273828
rect 88392 273788 119344 273816
rect 88392 273776 88398 273788
rect 119338 273776 119344 273788
rect 119396 273776 119402 273828
rect 120258 273776 120264 273828
rect 120316 273816 120322 273828
rect 175274 273816 175280 273828
rect 120316 273788 175280 273816
rect 120316 273776 120322 273788
rect 175274 273776 175280 273788
rect 175332 273776 175338 273828
rect 192386 273776 192392 273828
rect 192444 273816 192450 273828
rect 224954 273816 224960 273828
rect 192444 273788 224960 273816
rect 192444 273776 192450 273788
rect 224954 273776 224960 273788
rect 225012 273776 225018 273828
rect 238726 273816 238754 273924
rect 271506 273912 271512 273964
rect 271564 273952 271570 273964
rect 280338 273952 280344 273964
rect 271564 273924 280344 273952
rect 271564 273912 271570 273924
rect 280338 273912 280344 273924
rect 280396 273912 280402 273964
rect 322750 273912 322756 273964
rect 322808 273952 322814 273964
rect 330570 273952 330576 273964
rect 322808 273924 330576 273952
rect 322808 273912 322814 273924
rect 330570 273912 330576 273924
rect 330628 273912 330634 273964
rect 335262 273912 335268 273964
rect 335320 273952 335326 273964
rect 348326 273952 348332 273964
rect 335320 273924 348332 273952
rect 335320 273912 335326 273924
rect 348326 273912 348332 273924
rect 348384 273912 348390 273964
rect 350350 273912 350356 273964
rect 350408 273952 350414 273964
rect 368474 273952 368480 273964
rect 350408 273924 368480 273952
rect 350408 273912 350414 273924
rect 368474 273912 368480 273924
rect 368532 273912 368538 273964
rect 377674 273912 377680 273964
rect 377732 273952 377738 273964
rect 408586 273952 408592 273964
rect 377732 273924 408592 273952
rect 377732 273912 377738 273924
rect 408586 273912 408592 273924
rect 408644 273912 408650 273964
rect 422110 273912 422116 273964
rect 422168 273952 422174 273964
rect 465718 273952 465724 273964
rect 422168 273924 465724 273952
rect 422168 273912 422174 273924
rect 465718 273912 465724 273924
rect 465776 273912 465782 273964
rect 465902 273912 465908 273964
rect 465960 273952 465966 273964
rect 472250 273952 472256 273964
rect 465960 273924 472256 273952
rect 465960 273912 465966 273924
rect 472250 273912 472256 273924
rect 472308 273912 472314 273964
rect 474476 273952 474504 274060
rect 513834 274048 513840 274060
rect 513892 274048 513898 274100
rect 536742 274048 536748 274100
rect 536800 274088 536806 274100
rect 634354 274088 634360 274100
rect 536800 274060 634360 274088
rect 536800 274048 536806 274060
rect 634354 274048 634360 274060
rect 634412 274048 634418 274100
rect 481910 273952 481916 273964
rect 474476 273924 481916 273952
rect 481910 273912 481916 273924
rect 481968 273912 481974 273964
rect 545758 273952 545764 273964
rect 485056 273924 545764 273952
rect 258074 273816 258080 273828
rect 238726 273788 258080 273816
rect 258074 273776 258080 273788
rect 258132 273776 258138 273828
rect 396994 273776 397000 273828
rect 397052 273816 397058 273828
rect 435818 273816 435824 273828
rect 397052 273788 435824 273816
rect 397052 273776 397058 273788
rect 435818 273776 435824 273788
rect 435876 273776 435882 273828
rect 438118 273776 438124 273828
rect 438176 273816 438182 273828
rect 473630 273816 473636 273828
rect 438176 273788 473636 273816
rect 438176 273776 438182 273788
rect 473630 273776 473636 273788
rect 473688 273776 473694 273828
rect 474642 273776 474648 273828
rect 474700 273816 474706 273828
rect 485056 273816 485084 273924
rect 545758 273912 545764 273924
rect 545816 273912 545822 273964
rect 545942 273912 545948 273964
rect 546000 273952 546006 273964
rect 639138 273952 639144 273964
rect 546000 273924 639144 273952
rect 546000 273912 546006 273924
rect 639138 273912 639144 273924
rect 639196 273912 639202 273964
rect 559926 273816 559932 273828
rect 474700 273788 485084 273816
rect 485148 273788 559932 273816
rect 474700 273776 474706 273788
rect 119062 273640 119068 273692
rect 119120 273680 119126 273692
rect 173250 273680 173256 273692
rect 119120 273652 173256 273680
rect 119120 273640 119126 273652
rect 173250 273640 173256 273652
rect 173308 273640 173314 273692
rect 440878 273640 440884 273692
rect 440936 273680 440942 273692
rect 440936 273652 464660 273680
rect 440936 273640 440942 273652
rect 132034 273504 132040 273556
rect 132092 273544 132098 273556
rect 153838 273544 153844 273556
rect 132092 273516 153844 273544
rect 132092 273504 132098 273516
rect 153838 273504 153844 273516
rect 153896 273504 153902 273556
rect 259362 273504 259368 273556
rect 259420 273544 259426 273556
rect 266354 273544 266360 273556
rect 259420 273516 266360 273544
rect 259420 273504 259426 273516
rect 266354 273504 266360 273516
rect 266412 273504 266418 273556
rect 447778 273504 447784 273556
rect 447836 273544 447842 273556
rect 456242 273544 456248 273556
rect 447836 273516 456248 273544
rect 447836 273504 447842 273516
rect 456242 273504 456248 273516
rect 456300 273504 456306 273556
rect 457438 273504 457444 273556
rect 457496 273544 457502 273556
rect 464430 273544 464436 273556
rect 457496 273516 464436 273544
rect 457496 273504 457502 273516
rect 464430 273504 464436 273516
rect 464488 273504 464494 273556
rect 464632 273544 464660 273652
rect 465718 273640 465724 273692
rect 465776 273680 465782 273692
rect 472434 273680 472440 273692
rect 465776 273652 472440 273680
rect 465776 273640 465782 273652
rect 472434 273640 472440 273652
rect 472492 273640 472498 273692
rect 484210 273640 484216 273692
rect 484268 273680 484274 273692
rect 485148 273680 485176 273788
rect 559926 273776 559932 273788
rect 559984 273776 559990 273828
rect 484268 273652 485176 273680
rect 484268 273640 484274 273652
rect 485314 273640 485320 273692
rect 485372 273680 485378 273692
rect 556338 273680 556344 273692
rect 485372 273652 556344 273680
rect 485372 273640 485378 273652
rect 556338 273640 556344 273652
rect 556396 273640 556402 273692
rect 556798 273640 556804 273692
rect 556856 273680 556862 273692
rect 590654 273680 590660 273692
rect 556856 273652 590660 273680
rect 556856 273640 556862 273652
rect 590654 273640 590660 273652
rect 590712 273640 590718 273692
rect 471238 273544 471244 273556
rect 464632 273516 471244 273544
rect 471238 273504 471244 273516
rect 471296 273504 471302 273556
rect 476022 273504 476028 273556
rect 476080 273544 476086 273556
rect 549254 273544 549260 273556
rect 476080 273516 549260 273544
rect 476080 273504 476086 273516
rect 549254 273504 549260 273516
rect 549312 273504 549318 273556
rect 551278 273504 551284 273556
rect 551336 273544 551342 273556
rect 583570 273544 583576 273556
rect 551336 273516 583576 273544
rect 551336 273504 551342 273516
rect 583570 273504 583576 273516
rect 583628 273504 583634 273556
rect 145282 273368 145288 273420
rect 145340 273408 145346 273420
rect 147858 273408 147864 273420
rect 145340 273380 147864 273408
rect 145340 273368 145346 273380
rect 147858 273368 147864 273380
rect 147916 273368 147922 273420
rect 463234 273368 463240 273420
rect 463292 273408 463298 273420
rect 466086 273408 466092 273420
rect 463292 273380 466092 273408
rect 463292 273368 463298 273380
rect 466086 273368 466092 273380
rect 466144 273368 466150 273420
rect 478690 273368 478696 273420
rect 478748 273408 478754 273420
rect 552842 273408 552848 273420
rect 478748 273380 552848 273408
rect 478748 273368 478754 273380
rect 552842 273368 552848 273380
rect 552900 273368 552906 273420
rect 327718 273232 327724 273284
rect 327776 273272 327782 273284
rect 329466 273272 329472 273284
rect 327776 273244 329472 273272
rect 327776 273232 327782 273244
rect 329466 273232 329472 273244
rect 329524 273232 329530 273284
rect 108390 273164 108396 273216
rect 108448 273204 108454 273216
rect 165890 273204 165896 273216
rect 108448 273176 165896 273204
rect 108448 273164 108454 273176
rect 165890 273164 165896 273176
rect 165948 273164 165954 273216
rect 186406 273164 186412 273216
rect 186464 273204 186470 273216
rect 218698 273204 218704 273216
rect 186464 273176 218704 273204
rect 186464 273164 186470 273176
rect 218698 273164 218704 273176
rect 218756 273164 218762 273216
rect 362770 273164 362776 273216
rect 362828 273204 362834 273216
rect 386138 273204 386144 273216
rect 362828 273176 386144 273204
rect 362828 273164 362834 273176
rect 386138 273164 386144 273176
rect 386196 273164 386202 273216
rect 400030 273164 400036 273216
rect 400088 273204 400094 273216
rect 439314 273204 439320 273216
rect 400088 273176 439320 273204
rect 400088 273164 400094 273176
rect 439314 273164 439320 273176
rect 439372 273164 439378 273216
rect 444006 273164 444012 273216
rect 444064 273204 444070 273216
rect 444064 273176 499712 273204
rect 444064 273164 444070 273176
rect 102502 273028 102508 273080
rect 102560 273068 102566 273080
rect 162854 273068 162860 273080
rect 102560 273040 162860 273068
rect 102560 273028 102566 273040
rect 162854 273028 162860 273040
rect 162912 273028 162918 273080
rect 172238 273028 172244 273080
rect 172296 273068 172302 273080
rect 209774 273068 209780 273080
rect 172296 273040 209780 273068
rect 172296 273028 172302 273040
rect 209774 273028 209780 273040
rect 209832 273028 209838 273080
rect 219526 273028 219532 273080
rect 219584 273068 219590 273080
rect 244550 273068 244556 273080
rect 219584 273040 244556 273068
rect 219584 273028 219590 273040
rect 244550 273028 244556 273040
rect 244608 273028 244614 273080
rect 280982 273028 280988 273080
rect 281040 273068 281046 273080
rect 286318 273068 286324 273080
rect 281040 273040 286324 273068
rect 281040 273028 281046 273040
rect 286318 273028 286324 273040
rect 286376 273028 286382 273080
rect 361206 273028 361212 273080
rect 361264 273068 361270 273080
rect 384942 273068 384948 273080
rect 361264 273040 384948 273068
rect 361264 273028 361270 273040
rect 384942 273028 384948 273040
rect 385000 273028 385006 273080
rect 385678 273028 385684 273080
rect 385736 273068 385742 273080
rect 395614 273068 395620 273080
rect 385736 273040 395620 273068
rect 385736 273028 385742 273040
rect 395614 273028 395620 273040
rect 395672 273028 395678 273080
rect 404170 273028 404176 273080
rect 404228 273068 404234 273080
rect 446490 273068 446496 273080
rect 404228 273040 446496 273068
rect 404228 273028 404234 273040
rect 446490 273028 446496 273040
rect 446548 273028 446554 273080
rect 446858 273028 446864 273080
rect 446916 273068 446922 273080
rect 499482 273068 499488 273080
rect 446916 273040 499488 273068
rect 446916 273028 446922 273040
rect 499482 273028 499488 273040
rect 499540 273028 499546 273080
rect 499684 273068 499712 273176
rect 499942 273164 499948 273216
rect 500000 273204 500006 273216
rect 511442 273204 511448 273216
rect 500000 273176 511448 273204
rect 500000 273164 500006 273176
rect 511442 273164 511448 273176
rect 511500 273164 511506 273216
rect 515214 273204 515220 273216
rect 511644 273176 515220 273204
rect 503162 273068 503168 273080
rect 499684 273040 503168 273068
rect 503162 273028 503168 273040
rect 503220 273028 503226 273080
rect 503346 273028 503352 273080
rect 503404 273068 503410 273080
rect 507946 273068 507952 273080
rect 503404 273040 507952 273068
rect 503404 273028 503410 273040
rect 507946 273028 507952 273040
rect 508004 273028 508010 273080
rect 509694 273028 509700 273080
rect 509752 273068 509758 273080
rect 511644 273068 511672 273176
rect 515214 273164 515220 273176
rect 515272 273164 515278 273216
rect 515398 273164 515404 273216
rect 515456 273204 515462 273216
rect 519722 273204 519728 273216
rect 515456 273176 519728 273204
rect 515456 273164 515462 273176
rect 519722 273164 519728 273176
rect 519780 273164 519786 273216
rect 521470 273164 521476 273216
rect 521528 273204 521534 273216
rect 614298 273204 614304 273216
rect 521528 273176 614304 273204
rect 521528 273164 521534 273176
rect 614298 273164 614304 273176
rect 614356 273164 614362 273216
rect 509752 273040 511672 273068
rect 509752 273028 509758 273040
rect 513558 273028 513564 273080
rect 513616 273068 513622 273080
rect 518526 273068 518532 273080
rect 513616 273040 518532 273068
rect 513616 273028 513622 273040
rect 518526 273028 518532 273040
rect 518584 273028 518590 273080
rect 562134 273068 562140 273080
rect 518866 273040 562140 273068
rect 94222 272892 94228 272944
rect 94280 272932 94286 272944
rect 155954 272932 155960 272944
rect 94280 272904 155960 272932
rect 94280 272892 94286 272904
rect 155954 272892 155960 272904
rect 156012 272892 156018 272944
rect 166350 272892 166356 272944
rect 166408 272932 166414 272944
rect 207290 272932 207296 272944
rect 166408 272904 207296 272932
rect 166408 272892 166414 272904
rect 207290 272892 207296 272904
rect 207348 272892 207354 272944
rect 211246 272892 211252 272944
rect 211304 272932 211310 272944
rect 220078 272932 220084 272944
rect 211304 272904 220084 272932
rect 211304 272892 211310 272904
rect 220078 272892 220084 272904
rect 220136 272892 220142 272944
rect 220722 272892 220728 272944
rect 220780 272932 220786 272944
rect 245746 272932 245752 272944
rect 220780 272904 245752 272932
rect 220780 272892 220786 272904
rect 245746 272892 245752 272904
rect 245804 272892 245810 272944
rect 247862 272892 247868 272944
rect 247920 272932 247926 272944
rect 264238 272932 264244 272944
rect 247920 272904 264244 272932
rect 247920 272892 247926 272904
rect 264238 272892 264244 272904
rect 264296 272892 264302 272944
rect 333790 272892 333796 272944
rect 333848 272932 333854 272944
rect 345934 272932 345940 272944
rect 333848 272904 345940 272932
rect 333848 272892 333854 272904
rect 345934 272892 345940 272904
rect 345992 272892 345998 272944
rect 348418 272892 348424 272944
rect 348476 272932 348482 272944
rect 362494 272932 362500 272944
rect 348476 272904 362500 272932
rect 348476 272892 348482 272904
rect 362494 272892 362500 272904
rect 362552 272892 362558 272944
rect 365438 272892 365444 272944
rect 365496 272932 365502 272944
rect 390922 272932 390928 272944
rect 365496 272904 390928 272932
rect 365496 272892 365502 272904
rect 390922 272892 390928 272904
rect 390980 272892 390986 272944
rect 405550 272892 405556 272944
rect 405608 272932 405614 272944
rect 448790 272932 448796 272944
rect 405608 272904 448796 272932
rect 405608 272892 405614 272904
rect 448790 272892 448796 272904
rect 448848 272892 448854 272944
rect 455322 272892 455328 272944
rect 455380 272932 455386 272944
rect 461394 272932 461400 272944
rect 455380 272904 461400 272932
rect 455380 272892 455386 272904
rect 461394 272892 461400 272904
rect 461452 272892 461458 272944
rect 515030 272932 515036 272944
rect 461596 272904 515036 272932
rect 82446 272756 82452 272808
rect 82504 272796 82510 272808
rect 148410 272796 148416 272808
rect 82504 272768 148416 272796
rect 82504 272756 82510 272768
rect 148410 272756 148416 272768
rect 148468 272756 148474 272808
rect 155678 272756 155684 272808
rect 155736 272796 155742 272808
rect 200114 272796 200120 272808
rect 155736 272768 200120 272796
rect 155736 272756 155742 272768
rect 200114 272756 200120 272768
rect 200172 272756 200178 272808
rect 205358 272756 205364 272808
rect 205416 272796 205422 272808
rect 234798 272796 234804 272808
rect 205416 272768 234804 272796
rect 205416 272756 205422 272768
rect 234798 272756 234804 272768
rect 234856 272756 234862 272808
rect 245378 272756 245384 272808
rect 245436 272796 245442 272808
rect 245436 272768 258074 272796
rect 245436 272756 245442 272768
rect 72970 272620 72976 272672
rect 73028 272660 73034 272672
rect 142154 272660 142160 272672
rect 73028 272632 142160 272660
rect 73028 272620 73034 272632
rect 142154 272620 142160 272632
rect 142212 272620 142218 272672
rect 142706 272620 142712 272672
rect 142764 272660 142770 272672
rect 145558 272660 145564 272672
rect 142764 272632 145564 272660
rect 142764 272620 142770 272632
rect 145558 272620 145564 272632
rect 145616 272620 145622 272672
rect 147398 272620 147404 272672
rect 147456 272660 147462 272672
rect 193214 272660 193220 272672
rect 147456 272632 193220 272660
rect 147456 272620 147462 272632
rect 193214 272620 193220 272632
rect 193272 272620 193278 272672
rect 195882 272620 195888 272672
rect 195940 272660 195946 272672
rect 227898 272660 227904 272672
rect 195940 272632 227904 272660
rect 195940 272620 195946 272632
rect 227898 272620 227904 272632
rect 227956 272620 227962 272672
rect 228082 272620 228088 272672
rect 228140 272660 228146 272672
rect 249058 272660 249064 272672
rect 228140 272632 249064 272660
rect 228140 272620 228146 272632
rect 249058 272620 249064 272632
rect 249116 272620 249122 272672
rect 258046 272660 258074 272768
rect 262306 272756 262312 272808
rect 262364 272796 262370 272808
rect 270954 272796 270960 272808
rect 262364 272768 270960 272796
rect 262364 272756 262370 272768
rect 270954 272756 270960 272768
rect 271012 272756 271018 272808
rect 273898 272756 273904 272808
rect 273956 272796 273962 272808
rect 282914 272796 282920 272808
rect 273956 272768 282920 272796
rect 273956 272756 273962 272768
rect 282914 272756 282920 272768
rect 282972 272756 282978 272808
rect 325326 272756 325332 272808
rect 325384 272796 325390 272808
rect 332962 272796 332968 272808
rect 325384 272768 332968 272796
rect 325384 272756 325390 272768
rect 332962 272756 332968 272768
rect 333020 272756 333026 272808
rect 344646 272756 344652 272808
rect 344704 272796 344710 272808
rect 361390 272796 361396 272808
rect 344704 272768 361396 272796
rect 344704 272756 344710 272768
rect 361390 272756 361396 272768
rect 361448 272756 361454 272808
rect 362218 272756 362224 272808
rect 362276 272796 362282 272808
rect 370774 272796 370780 272808
rect 362276 272768 370780 272796
rect 362276 272756 362282 272768
rect 370774 272756 370780 272768
rect 370832 272756 370838 272808
rect 396810 272796 396816 272808
rect 373966 272768 396816 272796
rect 262674 272660 262680 272672
rect 258046 272632 262680 272660
rect 262674 272620 262680 272632
rect 262732 272620 262738 272672
rect 264422 272620 264428 272672
rect 264480 272660 264486 272672
rect 269114 272660 269120 272672
rect 264480 272632 269120 272660
rect 264480 272620 264486 272632
rect 269114 272620 269120 272632
rect 269172 272620 269178 272672
rect 269390 272620 269396 272672
rect 269448 272660 269454 272672
rect 270586 272660 270592 272672
rect 269448 272632 270592 272660
rect 269448 272620 269454 272632
rect 270586 272620 270592 272632
rect 270644 272620 270650 272672
rect 324038 272620 324044 272672
rect 324096 272660 324102 272672
rect 331766 272660 331772 272672
rect 324096 272632 331772 272660
rect 324096 272620 324102 272632
rect 331766 272620 331772 272632
rect 331824 272620 331830 272672
rect 332318 272620 332324 272672
rect 332376 272660 332382 272672
rect 343634 272660 343640 272672
rect 332376 272632 343640 272660
rect 332376 272620 332382 272632
rect 343634 272620 343640 272632
rect 343692 272620 343698 272672
rect 346210 272620 346216 272672
rect 346268 272660 346274 272672
rect 363690 272660 363696 272672
rect 346268 272632 363696 272660
rect 346268 272620 346274 272632
rect 363690 272620 363696 272632
rect 363748 272620 363754 272672
rect 370498 272620 370504 272672
rect 370556 272660 370562 272672
rect 373966 272660 373994 272768
rect 396810 272756 396816 272768
rect 396868 272756 396874 272808
rect 406838 272756 406844 272808
rect 406896 272796 406902 272808
rect 449986 272796 449992 272808
rect 406896 272768 449992 272796
rect 406896 272756 406902 272768
rect 449986 272756 449992 272768
rect 450044 272756 450050 272808
rect 452286 272756 452292 272808
rect 452344 272796 452350 272808
rect 461596 272796 461624 272904
rect 515030 272892 515036 272904
rect 515088 272892 515094 272944
rect 515214 272892 515220 272944
rect 515272 272932 515278 272944
rect 518866 272932 518894 273040
rect 562134 273028 562140 273040
rect 562192 273028 562198 273080
rect 562318 273028 562324 273080
rect 562376 273068 562382 273080
rect 601142 273068 601148 273080
rect 562376 273040 601148 273068
rect 562376 273028 562382 273040
rect 601142 273028 601148 273040
rect 601200 273028 601206 273080
rect 624970 273068 624976 273080
rect 605806 273040 624976 273068
rect 515272 272904 518894 272932
rect 515272 272892 515278 272904
rect 532510 272892 532516 272944
rect 532568 272932 532574 272944
rect 532568 272904 538904 272932
rect 532568 272892 532574 272904
rect 513558 272796 513564 272808
rect 452344 272768 461624 272796
rect 461688 272768 513564 272796
rect 452344 272756 452350 272768
rect 370556 272632 373994 272660
rect 370556 272620 370562 272632
rect 376110 272620 376116 272672
rect 376168 272660 376174 272672
rect 406286 272660 406292 272672
rect 376168 272632 406292 272660
rect 376168 272620 376174 272632
rect 406286 272620 406292 272632
rect 406344 272620 406350 272672
rect 412266 272620 412272 272672
rect 412324 272660 412330 272672
rect 457070 272660 457076 272672
rect 412324 272632 457076 272660
rect 412324 272620 412330 272632
rect 457070 272620 457076 272632
rect 457128 272620 457134 272672
rect 457254 272620 457260 272672
rect 457312 272660 457318 272672
rect 461026 272660 461032 272672
rect 457312 272632 461032 272660
rect 457312 272620 457318 272632
rect 461026 272620 461032 272632
rect 461084 272620 461090 272672
rect 461394 272620 461400 272672
rect 461452 272660 461458 272672
rect 461688 272660 461716 272768
rect 513558 272756 513564 272768
rect 513616 272756 513622 272808
rect 513742 272756 513748 272808
rect 513800 272796 513806 272808
rect 525610 272796 525616 272808
rect 513800 272768 525616 272796
rect 513800 272756 513806 272768
rect 525610 272756 525616 272768
rect 525668 272756 525674 272808
rect 529842 272756 529848 272808
rect 529900 272796 529906 272808
rect 532878 272796 532884 272808
rect 529900 272768 532884 272796
rect 529900 272756 529906 272768
rect 532878 272756 532884 272768
rect 532936 272756 532942 272808
rect 533706 272756 533712 272808
rect 533764 272796 533770 272808
rect 538674 272796 538680 272808
rect 533764 272768 538680 272796
rect 533764 272756 533770 272768
rect 538674 272756 538680 272768
rect 538732 272756 538738 272808
rect 538876 272796 538904 272904
rect 539042 272892 539048 272944
rect 539100 272932 539106 272944
rect 605806 272932 605834 273040
rect 624970 273028 624976 273040
rect 625028 273028 625034 273080
rect 539100 272904 605834 272932
rect 539100 272892 539106 272904
rect 618438 272892 618444 272944
rect 618496 272932 618502 272944
rect 621382 272932 621388 272944
rect 618496 272904 621388 272932
rect 618496 272892 618502 272904
rect 621382 272892 621388 272904
rect 621440 272892 621446 272944
rect 628466 272796 628472 272808
rect 538876 272768 628472 272796
rect 628466 272756 628472 272768
rect 628524 272756 628530 272808
rect 461452 272632 461716 272660
rect 461452 272620 461458 272632
rect 461854 272620 461860 272672
rect 461912 272660 461918 272672
rect 461912 272632 463924 272660
rect 461912 272620 461918 272632
rect 319070 272552 319076 272604
rect 319128 272592 319134 272604
rect 319622 272592 319628 272604
rect 319128 272564 319628 272592
rect 319128 272552 319134 272564
rect 319622 272552 319628 272564
rect 319680 272552 319686 272604
rect 463896 272592 463924 272632
rect 466408 272620 466414 272672
rect 466466 272660 466472 272672
rect 522114 272660 522120 272672
rect 466466 272632 522120 272660
rect 466466 272620 466472 272632
rect 522114 272620 522120 272632
rect 522172 272620 522178 272672
rect 526806 272620 526812 272672
rect 526864 272660 526870 272672
rect 618438 272660 618444 272672
rect 526864 272632 618444 272660
rect 526864 272620 526870 272632
rect 618438 272620 618444 272632
rect 618496 272620 618502 272672
rect 620278 272620 620284 272672
rect 620336 272660 620342 272672
rect 635550 272660 635556 272672
rect 620336 272632 635556 272660
rect 620336 272620 620342 272632
rect 635550 272620 635556 272632
rect 635608 272620 635614 272672
rect 463896 272564 466316 272592
rect 65886 272484 65892 272536
rect 65944 272524 65950 272536
rect 136818 272524 136824 272536
rect 65944 272496 136824 272524
rect 65944 272484 65950 272496
rect 136818 272484 136824 272496
rect 136876 272484 136882 272536
rect 137922 272484 137928 272536
rect 137980 272524 137986 272536
rect 137980 272496 180794 272524
rect 137980 272484 137986 272496
rect 116670 272348 116676 272400
rect 116728 272388 116734 272400
rect 172514 272388 172520 272400
rect 116728 272360 172520 272388
rect 116728 272348 116734 272360
rect 172514 272348 172520 272360
rect 172572 272348 172578 272400
rect 180766 272388 180794 272496
rect 181714 272484 181720 272536
rect 181772 272524 181778 272536
rect 187142 272524 187148 272536
rect 181772 272496 187148 272524
rect 181772 272484 181778 272496
rect 187142 272484 187148 272496
rect 187200 272484 187206 272536
rect 189074 272484 189080 272536
rect 189132 272524 189138 272536
rect 196434 272524 196440 272536
rect 189132 272496 196440 272524
rect 189132 272484 189138 272496
rect 196434 272484 196440 272496
rect 196492 272484 196498 272536
rect 197078 272484 197084 272536
rect 197136 272524 197142 272536
rect 229094 272524 229100 272536
rect 197136 272496 229100 272524
rect 197136 272484 197142 272496
rect 229094 272484 229100 272496
rect 229152 272484 229158 272536
rect 233694 272484 233700 272536
rect 233752 272524 233758 272536
rect 254394 272524 254400 272536
rect 233752 272496 254400 272524
rect 233752 272484 233758 272496
rect 254394 272484 254400 272496
rect 254452 272484 254458 272536
rect 254946 272484 254952 272536
rect 255004 272524 255010 272536
rect 269298 272524 269304 272536
rect 255004 272496 269304 272524
rect 255004 272484 255010 272496
rect 269298 272484 269304 272496
rect 269356 272484 269362 272536
rect 270310 272484 270316 272536
rect 270368 272524 270374 272536
rect 280522 272524 280528 272536
rect 270368 272496 280528 272524
rect 270368 272484 270374 272496
rect 280522 272484 280528 272496
rect 280580 272484 280586 272536
rect 329742 272484 329748 272536
rect 329800 272524 329806 272536
rect 338850 272524 338856 272536
rect 329800 272496 338856 272524
rect 329800 272484 329806 272496
rect 338850 272484 338856 272496
rect 338908 272484 338914 272536
rect 339218 272484 339224 272536
rect 339276 272524 339282 272536
rect 354214 272524 354220 272536
rect 339276 272496 354220 272524
rect 339276 272484 339282 272496
rect 354214 272484 354220 272496
rect 354272 272484 354278 272536
rect 354490 272484 354496 272536
rect 354548 272524 354554 272536
rect 375558 272524 375564 272536
rect 354548 272496 375564 272524
rect 354548 272484 354554 272496
rect 375558 272484 375564 272496
rect 375616 272484 375622 272536
rect 379422 272484 379428 272536
rect 379480 272524 379486 272536
rect 410978 272524 410984 272536
rect 379480 272496 410984 272524
rect 379480 272484 379486 272496
rect 410978 272484 410984 272496
rect 411036 272484 411042 272536
rect 416590 272484 416596 272536
rect 416648 272524 416654 272536
rect 463694 272524 463700 272536
rect 416648 272496 463700 272524
rect 416648 272484 416654 272496
rect 463694 272484 463700 272496
rect 463752 272484 463758 272536
rect 466288 272524 466316 272564
rect 470548 272524 470554 272536
rect 466288 272496 470554 272524
rect 470548 272484 470554 272496
rect 470606 272484 470612 272536
rect 470686 272484 470692 272536
rect 470744 272524 470750 272536
rect 532694 272524 532700 272536
rect 470744 272496 532700 272524
rect 470744 272484 470750 272496
rect 532694 272484 532700 272496
rect 532752 272484 532758 272536
rect 532878 272484 532884 272536
rect 532936 272524 532942 272536
rect 538490 272524 538496 272536
rect 532936 272496 538496 272524
rect 532936 272484 532942 272496
rect 538490 272484 538496 272496
rect 538548 272484 538554 272536
rect 538674 272484 538680 272536
rect 538732 272524 538738 272536
rect 632054 272524 632060 272536
rect 538732 272496 632060 272524
rect 538732 272484 538738 272496
rect 632054 272484 632060 272496
rect 632112 272484 632118 272536
rect 634078 272484 634084 272536
rect 634136 272524 634142 272536
rect 640334 272524 640340 272536
rect 634136 272496 640340 272524
rect 634136 272484 634142 272496
rect 640334 272484 640340 272496
rect 640392 272484 640398 272536
rect 318702 272416 318708 272468
rect 318760 272456 318766 272468
rect 324682 272456 324688 272468
rect 318760 272428 324688 272456
rect 318760 272416 318766 272428
rect 324682 272416 324688 272428
rect 324740 272416 324746 272468
rect 187694 272388 187700 272400
rect 180766 272360 187700 272388
rect 187694 272348 187700 272360
rect 187752 272348 187758 272400
rect 194962 272348 194968 272400
rect 195020 272388 195026 272400
rect 227162 272388 227168 272400
rect 195020 272360 227168 272388
rect 195020 272348 195026 272360
rect 227162 272348 227168 272360
rect 227220 272348 227226 272400
rect 269114 272348 269120 272400
rect 269172 272388 269178 272400
rect 276014 272388 276020 272400
rect 269172 272360 276020 272388
rect 269172 272348 269178 272360
rect 276014 272348 276020 272360
rect 276072 272348 276078 272400
rect 395982 272348 395988 272400
rect 396040 272388 396046 272400
rect 434622 272388 434628 272400
rect 396040 272360 434628 272388
rect 396040 272348 396046 272360
rect 434622 272348 434628 272360
rect 434680 272348 434686 272400
rect 449710 272348 449716 272400
rect 449768 272388 449774 272400
rect 499482 272388 499488 272400
rect 449768 272360 499488 272388
rect 449768 272348 449774 272360
rect 499482 272348 499488 272360
rect 499540 272348 499546 272400
rect 499666 272348 499672 272400
rect 499724 272388 499730 272400
rect 513742 272388 513748 272400
rect 499724 272360 513748 272388
rect 499724 272348 499730 272360
rect 513742 272348 513748 272360
rect 513800 272348 513806 272400
rect 517422 272348 517428 272400
rect 517480 272388 517486 272400
rect 600958 272388 600964 272400
rect 517480 272360 600964 272388
rect 517480 272348 517486 272360
rect 600958 272348 600964 272360
rect 601016 272348 601022 272400
rect 601142 272348 601148 272400
rect 601200 272388 601206 272400
rect 620278 272388 620284 272400
rect 601200 272360 620284 272388
rect 601200 272348 601206 272360
rect 620278 272348 620284 272360
rect 620336 272348 620342 272400
rect 127342 272212 127348 272264
rect 127400 272252 127406 272264
rect 179874 272252 179880 272264
rect 127400 272224 179880 272252
rect 127400 272212 127406 272224
rect 179874 272212 179880 272224
rect 179932 272212 179938 272264
rect 391842 272212 391848 272264
rect 391900 272252 391906 272264
rect 428734 272252 428740 272264
rect 391900 272224 428740 272252
rect 391900 272212 391906 272224
rect 428734 272212 428740 272224
rect 428792 272212 428798 272264
rect 450538 272212 450544 272264
rect 450596 272252 450602 272264
rect 510246 272252 510252 272264
rect 450596 272224 510252 272252
rect 450596 272212 450602 272224
rect 510246 272212 510252 272224
rect 510304 272212 510310 272264
rect 520090 272212 520096 272264
rect 520148 272252 520154 272264
rect 610710 272252 610716 272264
rect 520148 272224 610716 272252
rect 520148 272212 520154 272224
rect 610710 272212 610716 272224
rect 610768 272212 610774 272264
rect 145098 272076 145104 272128
rect 145156 272116 145162 272128
rect 192386 272116 192392 272128
rect 145156 272088 192392 272116
rect 145156 272076 145162 272088
rect 192386 272076 192392 272088
rect 192444 272076 192450 272128
rect 384942 272076 384948 272128
rect 385000 272116 385006 272128
rect 418062 272116 418068 272128
rect 385000 272088 418068 272116
rect 385000 272076 385006 272088
rect 418062 272076 418068 272088
rect 418120 272076 418126 272128
rect 431678 272076 431684 272128
rect 431736 272116 431742 272128
rect 480162 272116 480168 272128
rect 431736 272088 480168 272116
rect 431736 272076 431742 272088
rect 480162 272076 480168 272088
rect 480220 272076 480226 272128
rect 489868 272116 489874 272128
rect 482756 272088 489874 272116
rect 124950 271940 124956 271992
rect 125008 271980 125014 271992
rect 151078 271980 151084 271992
rect 125008 271952 151084 271980
rect 125008 271940 125014 271952
rect 151078 271940 151084 271952
rect 151136 271940 151142 271992
rect 428458 271940 428464 271992
rect 428516 271980 428522 271992
rect 470548 271980 470554 271992
rect 428516 271952 470554 271980
rect 428516 271940 428522 271952
rect 470548 271940 470554 271952
rect 470606 271940 470612 271992
rect 470686 271940 470692 271992
rect 470744 271980 470750 271992
rect 482756 271980 482784 272088
rect 489868 272076 489874 272088
rect 489926 272076 489932 272128
rect 490006 272076 490012 272128
rect 490064 272116 490070 272128
rect 552290 272116 552296 272128
rect 490064 272088 552296 272116
rect 490064 272076 490070 272088
rect 552290 272076 552296 272088
rect 552348 272076 552354 272128
rect 562318 272116 562324 272128
rect 552676 272088 562324 272116
rect 552676 272048 552704 272088
rect 562318 272076 562324 272088
rect 562376 272076 562382 272128
rect 600958 272076 600964 272128
rect 601016 272116 601022 272128
rect 607214 272116 607220 272128
rect 601016 272088 607220 272116
rect 601016 272076 601022 272088
rect 607214 272076 607220 272088
rect 607272 272076 607278 272128
rect 552492 272020 552704 272048
rect 470744 271952 482784 271980
rect 470744 271940 470750 271952
rect 483198 271940 483204 271992
rect 483256 271980 483262 271992
rect 547506 271980 547512 271992
rect 483256 271952 547512 271980
rect 483256 271940 483262 271952
rect 547506 271940 547512 271952
rect 547564 271940 547570 271992
rect 547690 271940 547696 271992
rect 547748 271980 547754 271992
rect 552492 271980 552520 272020
rect 547748 271952 552520 271980
rect 547748 271940 547754 271952
rect 552842 271940 552848 271992
rect 552900 271980 552906 271992
rect 558730 271980 558736 271992
rect 552900 271952 558736 271980
rect 552900 271940 552906 271952
rect 558730 271940 558736 271952
rect 558788 271940 558794 271992
rect 562134 271940 562140 271992
rect 562192 271980 562198 271992
rect 569402 271980 569408 271992
rect 562192 271952 569408 271980
rect 562192 271940 562198 271952
rect 569402 271940 569408 271952
rect 569460 271940 569466 271992
rect 105998 271804 106004 271856
rect 106056 271844 106062 271856
rect 164970 271844 164976 271856
rect 106056 271816 164976 271844
rect 106056 271804 106062 271816
rect 164970 271804 164976 271816
rect 165028 271804 165034 271856
rect 174262 271804 174268 271856
rect 174320 271844 174326 271856
rect 189258 271844 189264 271856
rect 174320 271816 189264 271844
rect 174320 271804 174326 271816
rect 189258 271804 189264 271816
rect 189316 271804 189322 271856
rect 202966 271804 202972 271856
rect 203024 271844 203030 271856
rect 233234 271844 233240 271856
rect 203024 271816 233240 271844
rect 203024 271804 203030 271816
rect 233234 271804 233240 271816
rect 233292 271804 233298 271856
rect 274634 271804 274640 271856
rect 274692 271844 274698 271856
rect 279234 271844 279240 271856
rect 274692 271816 279240 271844
rect 274692 271804 274698 271816
rect 279234 271804 279240 271816
rect 279292 271804 279298 271856
rect 355318 271804 355324 271856
rect 355376 271844 355382 271856
rect 356606 271844 356612 271856
rect 355376 271816 356612 271844
rect 355376 271804 355382 271816
rect 356606 271804 356612 271816
rect 356664 271804 356670 271856
rect 375282 271804 375288 271856
rect 375340 271844 375346 271856
rect 403894 271844 403900 271856
rect 375340 271816 403900 271844
rect 375340 271804 375346 271816
rect 403894 271804 403900 271816
rect 403952 271804 403958 271856
rect 433150 271804 433156 271856
rect 433208 271844 433214 271856
rect 433208 271816 483428 271844
rect 433208 271804 433214 271816
rect 97810 271668 97816 271720
rect 97868 271708 97874 271720
rect 158806 271708 158812 271720
rect 97868 271680 158812 271708
rect 97868 271668 97874 271680
rect 158806 271668 158812 271680
rect 158864 271668 158870 271720
rect 169846 271668 169852 271720
rect 169904 271708 169910 271720
rect 209958 271708 209964 271720
rect 169904 271680 209964 271708
rect 169904 271668 169910 271680
rect 209958 271668 209964 271680
rect 210016 271668 210022 271720
rect 225414 271668 225420 271720
rect 225472 271708 225478 271720
rect 228358 271708 228364 271720
rect 225472 271680 228364 271708
rect 225472 271668 225478 271680
rect 228358 271668 228364 271680
rect 228416 271668 228422 271720
rect 351178 271668 351184 271720
rect 351236 271708 351242 271720
rect 366082 271708 366088 271720
rect 351236 271680 366088 271708
rect 351236 271668 351242 271680
rect 366082 271668 366088 271680
rect 366140 271668 366146 271720
rect 381998 271668 382004 271720
rect 382056 271708 382062 271720
rect 414566 271708 414572 271720
rect 382056 271680 414572 271708
rect 382056 271668 382062 271680
rect 414566 271668 414572 271680
rect 414624 271668 414630 271720
rect 421650 271708 421656 271720
rect 417160 271680 421656 271708
rect 87138 271532 87144 271584
rect 87196 271572 87202 271584
rect 151998 271572 152004 271584
rect 87196 271544 152004 271572
rect 87196 271532 87202 271544
rect 151998 271532 152004 271544
rect 152056 271532 152062 271584
rect 165154 271532 165160 271584
rect 165212 271572 165218 271584
rect 205634 271572 205640 271584
rect 165212 271544 205640 271572
rect 165212 271532 165218 271544
rect 205634 271532 205640 271544
rect 205692 271532 205698 271584
rect 215938 271532 215944 271584
rect 215996 271572 216002 271584
rect 242066 271572 242072 271584
rect 215996 271544 242072 271572
rect 215996 271532 216002 271544
rect 242066 271532 242072 271544
rect 242124 271532 242130 271584
rect 337930 271532 337936 271584
rect 337988 271572 337994 271584
rect 350718 271572 350724 271584
rect 337988 271544 350724 271572
rect 337988 271532 337994 271544
rect 350718 271532 350724 271544
rect 350776 271532 350782 271584
rect 360838 271532 360844 271584
rect 360896 271572 360902 271584
rect 377858 271572 377864 271584
rect 360896 271544 377864 271572
rect 360896 271532 360902 271544
rect 377858 271532 377864 271544
rect 377916 271532 377922 271584
rect 387702 271532 387708 271584
rect 387760 271572 387766 271584
rect 417160 271572 417188 271680
rect 421650 271668 421656 271680
rect 421708 271668 421714 271720
rect 430390 271668 430396 271720
rect 430448 271708 430454 271720
rect 483014 271708 483020 271720
rect 430448 271680 483020 271708
rect 430448 271668 430454 271680
rect 483014 271668 483020 271680
rect 483072 271668 483078 271720
rect 483400 271708 483428 271816
rect 485038 271804 485044 271856
rect 485096 271844 485102 271856
rect 490006 271844 490012 271856
rect 485096 271816 490012 271844
rect 485096 271804 485102 271816
rect 490006 271804 490012 271816
rect 490064 271804 490070 271856
rect 496538 271804 496544 271856
rect 496596 271844 496602 271856
rect 578878 271844 578884 271856
rect 496596 271816 578884 271844
rect 496596 271804 496602 271816
rect 578878 271804 578884 271816
rect 578936 271804 578942 271856
rect 486602 271708 486608 271720
rect 483400 271680 486608 271708
rect 486602 271668 486608 271680
rect 486660 271668 486666 271720
rect 494698 271668 494704 271720
rect 494756 271708 494762 271720
rect 501782 271708 501788 271720
rect 494756 271680 501788 271708
rect 494756 271668 494762 271680
rect 501782 271668 501788 271680
rect 501840 271668 501846 271720
rect 501966 271668 501972 271720
rect 502024 271708 502030 271720
rect 585962 271708 585968 271720
rect 502024 271680 585968 271708
rect 502024 271668 502030 271680
rect 585962 271668 585968 271680
rect 586020 271668 586026 271720
rect 387760 271544 417188 271572
rect 387760 271532 387766 271544
rect 420178 271532 420184 271584
rect 420236 271572 420242 271584
rect 431126 271572 431132 271584
rect 420236 271544 431132 271572
rect 420236 271532 420242 271544
rect 431126 271532 431132 271544
rect 431184 271532 431190 271584
rect 437198 271532 437204 271584
rect 437256 271572 437262 271584
rect 493686 271572 493692 271584
rect 437256 271544 493692 271572
rect 437256 271532 437262 271544
rect 493686 271532 493692 271544
rect 493744 271532 493750 271584
rect 499298 271532 499304 271584
rect 499356 271572 499362 271584
rect 582374 271572 582380 271584
rect 499356 271544 582380 271572
rect 499356 271532 499362 271544
rect 582374 271532 582380 271544
rect 582432 271532 582438 271584
rect 583018 271532 583024 271584
rect 583076 271572 583082 271584
rect 611630 271572 611636 271584
rect 583076 271544 611636 271572
rect 583076 271532 583082 271544
rect 611630 271532 611636 271544
rect 611688 271532 611694 271584
rect 611998 271532 612004 271584
rect 612056 271572 612062 271584
rect 618990 271572 618996 271584
rect 612056 271544 618996 271572
rect 612056 271532 612062 271544
rect 618990 271532 618996 271544
rect 619048 271532 619054 271584
rect 75362 271396 75368 271448
rect 75420 271436 75426 271448
rect 142706 271436 142712 271448
rect 75420 271408 142712 271436
rect 75420 271396 75426 271408
rect 142706 271396 142712 271408
rect 142764 271396 142770 271448
rect 162670 271396 162676 271448
rect 162728 271436 162734 271448
rect 204714 271436 204720 271448
rect 162728 271408 204720 271436
rect 162728 271396 162734 271408
rect 204714 271396 204720 271408
rect 204772 271396 204778 271448
rect 213638 271396 213644 271448
rect 213696 271436 213702 271448
rect 240410 271436 240416 271448
rect 213696 271408 240416 271436
rect 213696 271396 213702 271408
rect 240410 271396 240416 271408
rect 240468 271396 240474 271448
rect 240778 271396 240784 271448
rect 240836 271436 240842 271448
rect 259638 271436 259644 271448
rect 240836 271408 259644 271436
rect 240836 271396 240842 271408
rect 259638 271396 259644 271408
rect 259696 271396 259702 271448
rect 259822 271396 259828 271448
rect 259880 271436 259886 271448
rect 272610 271436 272616 271448
rect 259880 271408 272616 271436
rect 259880 271396 259886 271408
rect 272610 271396 272616 271408
rect 272668 271396 272674 271448
rect 325510 271396 325516 271448
rect 325568 271436 325574 271448
rect 334158 271436 334164 271448
rect 325568 271408 334164 271436
rect 325568 271396 325574 271408
rect 334158 271396 334164 271408
rect 334216 271396 334222 271448
rect 347682 271396 347688 271448
rect 347740 271436 347746 271448
rect 364886 271436 364892 271448
rect 347740 271408 364892 271436
rect 347740 271396 347746 271408
rect 364886 271396 364892 271408
rect 364944 271396 364950 271448
rect 366358 271396 366364 271448
rect 366416 271436 366422 271448
rect 383838 271436 383844 271448
rect 366416 271408 383844 271436
rect 366416 271396 366422 271408
rect 383838 271396 383844 271408
rect 383896 271396 383902 271448
rect 384758 271396 384764 271448
rect 384816 271436 384822 271448
rect 419258 271436 419264 271448
rect 384816 271408 419264 271436
rect 384816 271396 384822 271408
rect 419258 271396 419264 271408
rect 419316 271396 419322 271448
rect 426342 271436 426348 271448
rect 424336 271408 426348 271436
rect 76834 271260 76840 271312
rect 76892 271300 76898 271312
rect 143534 271300 143540 271312
rect 76892 271272 143540 271300
rect 76892 271260 76898 271272
rect 143534 271260 143540 271272
rect 143592 271260 143598 271312
rect 152182 271260 152188 271312
rect 152240 271300 152246 271312
rect 197354 271300 197360 271312
rect 152240 271272 197360 271300
rect 152240 271260 152246 271272
rect 197354 271260 197360 271272
rect 197412 271260 197418 271312
rect 198274 271260 198280 271312
rect 198332 271300 198338 271312
rect 229554 271300 229560 271312
rect 198332 271272 229560 271300
rect 198332 271260 198338 271272
rect 229554 271260 229560 271272
rect 229612 271260 229618 271312
rect 235258 271260 235264 271312
rect 235316 271300 235322 271312
rect 255314 271300 255320 271312
rect 235316 271272 255320 271300
rect 235316 271260 235322 271272
rect 255314 271260 255320 271272
rect 255372 271260 255378 271312
rect 256694 271260 256700 271312
rect 256752 271300 256758 271312
rect 261018 271300 261024 271312
rect 256752 271272 261024 271300
rect 256752 271260 256758 271272
rect 261018 271260 261024 271272
rect 261076 271260 261082 271312
rect 262030 271260 262036 271312
rect 262088 271300 262094 271312
rect 274634 271300 274640 271312
rect 262088 271272 274640 271300
rect 262088 271260 262094 271272
rect 274634 271260 274640 271272
rect 274692 271260 274698 271312
rect 329558 271260 329564 271312
rect 329616 271300 329622 271312
rect 340046 271300 340052 271312
rect 329616 271272 340052 271300
rect 329616 271260 329622 271272
rect 340046 271260 340052 271272
rect 340104 271260 340110 271312
rect 340598 271260 340604 271312
rect 340656 271300 340662 271312
rect 355134 271300 355140 271312
rect 340656 271272 355140 271300
rect 340656 271260 340662 271272
rect 355134 271260 355140 271272
rect 355192 271260 355198 271312
rect 357158 271260 357164 271312
rect 357216 271300 357222 271312
rect 379054 271300 379060 271312
rect 357216 271272 379060 271300
rect 357216 271260 357222 271272
rect 379054 271260 379060 271272
rect 379112 271260 379118 271312
rect 390278 271260 390284 271312
rect 390336 271300 390342 271312
rect 424336 271300 424364 271408
rect 426342 271396 426348 271408
rect 426400 271396 426406 271448
rect 439958 271396 439964 271448
rect 440016 271436 440022 271448
rect 497274 271436 497280 271448
rect 440016 271408 497280 271436
rect 440016 271396 440022 271408
rect 497274 271396 497280 271408
rect 497332 271396 497338 271448
rect 505002 271396 505008 271448
rect 505060 271436 505066 271448
rect 589458 271436 589464 271448
rect 505060 271408 589464 271436
rect 505060 271396 505066 271408
rect 589458 271396 589464 271408
rect 589516 271396 589522 271448
rect 589918 271396 589924 271448
rect 589976 271436 589982 271448
rect 633250 271436 633256 271448
rect 589976 271408 633256 271436
rect 589976 271396 589982 271408
rect 633250 271396 633256 271408
rect 633308 271396 633314 271448
rect 432230 271300 432236 271312
rect 390336 271272 424364 271300
rect 425992 271272 432236 271300
rect 390336 271260 390342 271272
rect 68186 271124 68192 271176
rect 68244 271164 68250 271176
rect 138474 271164 138480 271176
rect 68244 271136 138480 271164
rect 68244 271124 68250 271136
rect 138474 271124 138480 271136
rect 138532 271124 138538 271176
rect 141510 271124 141516 271176
rect 141568 271164 141574 271176
rect 189074 271164 189080 271176
rect 141568 271136 189080 271164
rect 141568 271124 141574 271136
rect 189074 271124 189080 271136
rect 189132 271124 189138 271176
rect 191190 271124 191196 271176
rect 191248 271164 191254 271176
rect 225138 271164 225144 271176
rect 191248 271136 225144 271164
rect 191248 271124 191254 271136
rect 225138 271124 225144 271136
rect 225196 271124 225202 271176
rect 230198 271124 230204 271176
rect 230256 271164 230262 271176
rect 252002 271164 252008 271176
rect 230256 271136 252008 271164
rect 230256 271124 230262 271136
rect 252002 271124 252008 271136
rect 252060 271124 252066 271176
rect 268010 271124 268016 271176
rect 268068 271164 268074 271176
rect 278866 271164 278872 271176
rect 268068 271136 278872 271164
rect 268068 271124 268074 271136
rect 278866 271124 278872 271136
rect 278924 271124 278930 271176
rect 279786 271124 279792 271176
rect 279844 271164 279850 271176
rect 287054 271164 287060 271176
rect 279844 271136 287060 271164
rect 279844 271124 279850 271136
rect 287054 271124 287060 271136
rect 287112 271124 287118 271176
rect 331122 271124 331128 271176
rect 331180 271164 331186 271176
rect 342438 271164 342444 271176
rect 331180 271136 342444 271164
rect 331180 271124 331186 271136
rect 342438 271124 342444 271136
rect 342496 271124 342502 271176
rect 343542 271124 343548 271176
rect 343600 271164 343606 271176
rect 360194 271164 360200 271176
rect 343600 271136 360200 271164
rect 343600 271124 343606 271136
rect 360194 271124 360200 271136
rect 360252 271124 360258 271176
rect 364150 271124 364156 271176
rect 364208 271164 364214 271176
rect 389726 271164 389732 271176
rect 364208 271136 389732 271164
rect 364208 271124 364214 271136
rect 389726 271124 389732 271136
rect 389784 271124 389790 271176
rect 394326 271124 394332 271176
rect 394384 271164 394390 271176
rect 425992 271164 426020 271272
rect 432230 271260 432236 271272
rect 432288 271260 432294 271312
rect 442902 271260 442908 271312
rect 442960 271300 442966 271312
rect 500862 271300 500868 271312
rect 442960 271272 500868 271300
rect 442960 271260 442966 271272
rect 500862 271260 500868 271272
rect 500920 271260 500926 271312
rect 507670 271260 507676 271312
rect 507728 271300 507734 271312
rect 593046 271300 593052 271312
rect 507728 271272 593052 271300
rect 507728 271260 507734 271272
rect 593046 271260 593052 271272
rect 593104 271260 593110 271312
rect 598198 271260 598204 271312
rect 598256 271300 598262 271312
rect 645026 271300 645032 271312
rect 598256 271272 645032 271300
rect 598256 271260 598262 271272
rect 645026 271260 645032 271272
rect 645084 271260 645090 271312
rect 437934 271164 437940 271176
rect 394384 271136 426020 271164
rect 427096 271136 437940 271164
rect 394384 271124 394390 271136
rect 113450 270988 113456 271040
rect 113508 271028 113514 271040
rect 169938 271028 169944 271040
rect 113508 271000 169944 271028
rect 113508 270988 113514 271000
rect 169938 270988 169944 271000
rect 169996 270988 170002 271040
rect 187418 270988 187424 271040
rect 187476 271028 187482 271040
rect 216122 271028 216128 271040
rect 187476 271000 216128 271028
rect 187476 270988 187482 271000
rect 216122 270988 216128 271000
rect 216180 270988 216186 271040
rect 251450 270988 251456 271040
rect 251508 271028 251514 271040
rect 266906 271028 266912 271040
rect 251508 271000 266912 271028
rect 251508 270988 251514 271000
rect 266906 270988 266912 271000
rect 266964 270988 266970 271040
rect 417418 270988 417424 271040
rect 417476 271028 417482 271040
rect 427096 271028 427124 271136
rect 437934 271124 437940 271136
rect 437992 271124 437998 271176
rect 441338 271124 441344 271176
rect 441396 271164 441402 271176
rect 445018 271164 445024 271176
rect 441396 271136 445024 271164
rect 441396 271124 441402 271136
rect 445018 271124 445024 271136
rect 445076 271124 445082 271176
rect 445662 271124 445668 271176
rect 445720 271164 445726 271176
rect 504358 271164 504364 271176
rect 445720 271136 504364 271164
rect 445720 271124 445726 271136
rect 504358 271124 504364 271136
rect 504416 271124 504422 271176
rect 524046 271124 524052 271176
rect 524104 271164 524110 271176
rect 617334 271164 617340 271176
rect 524104 271136 617340 271164
rect 524104 271124 524110 271136
rect 617334 271124 617340 271136
rect 617392 271124 617398 271176
rect 617518 271124 617524 271176
rect 617576 271164 617582 271176
rect 626074 271164 626080 271176
rect 617576 271136 626080 271164
rect 617576 271124 617582 271136
rect 626074 271124 626080 271136
rect 626132 271124 626138 271176
rect 417476 271000 427124 271028
rect 417476 270988 417482 271000
rect 427446 270988 427452 271040
rect 427504 271028 427510 271040
rect 479150 271028 479156 271040
rect 427504 271000 479156 271028
rect 427504 270988 427510 271000
rect 479150 270988 479156 271000
rect 479208 270988 479214 271040
rect 482278 270988 482284 271040
rect 482336 271028 482342 271040
rect 494698 271028 494704 271040
rect 482336 271000 494704 271028
rect 482336 270988 482342 271000
rect 494698 270988 494704 271000
rect 494756 270988 494762 271040
rect 495250 270988 495256 271040
rect 495308 271028 495314 271040
rect 575290 271028 575296 271040
rect 495308 271000 575296 271028
rect 495308 270988 495314 271000
rect 575290 270988 575296 271000
rect 575348 270988 575354 271040
rect 576118 270988 576124 271040
rect 576176 271028 576182 271040
rect 604822 271028 604828 271040
rect 576176 271000 604828 271028
rect 576176 270988 576182 271000
rect 604822 270988 604828 271000
rect 604880 270988 604886 271040
rect 123754 270852 123760 270904
rect 123812 270892 123818 270904
rect 177482 270892 177488 270904
rect 123812 270864 177488 270892
rect 123812 270852 123818 270864
rect 177482 270852 177488 270864
rect 177540 270852 177546 270904
rect 407758 270852 407764 270904
rect 407816 270892 407822 270904
rect 440510 270892 440516 270904
rect 407816 270864 440516 270892
rect 407816 270852 407822 270864
rect 440510 270852 440516 270864
rect 440568 270852 440574 270904
rect 449158 270852 449164 270904
rect 449216 270892 449222 270904
rect 490190 270892 490196 270904
rect 449216 270864 490196 270892
rect 449216 270852 449222 270864
rect 490190 270852 490196 270864
rect 490248 270852 490254 270904
rect 492490 270852 492496 270904
rect 492548 270892 492554 270904
rect 571702 270892 571708 270904
rect 492548 270864 571708 270892
rect 492548 270852 492554 270864
rect 571702 270852 571708 270864
rect 571760 270852 571766 270904
rect 134426 270716 134432 270768
rect 134484 270756 134490 270768
rect 185118 270756 185124 270768
rect 134484 270728 185124 270756
rect 134484 270716 134490 270728
rect 185118 270716 185124 270728
rect 185176 270716 185182 270768
rect 321370 270716 321376 270768
rect 321428 270756 321434 270768
rect 327074 270756 327080 270768
rect 321428 270728 327080 270756
rect 321428 270716 321434 270728
rect 327074 270716 327080 270728
rect 327132 270716 327138 270768
rect 414474 270716 414480 270768
rect 414532 270756 414538 270768
rect 450814 270756 450820 270768
rect 414532 270728 450820 270756
rect 414532 270716 414538 270728
rect 450814 270716 450820 270728
rect 450872 270716 450878 270768
rect 486970 270716 486976 270768
rect 487028 270756 487034 270768
rect 564618 270756 564624 270768
rect 487028 270728 564624 270756
rect 487028 270716 487034 270728
rect 564618 270716 564624 270728
rect 564676 270716 564682 270768
rect 567838 270716 567844 270768
rect 567896 270756 567902 270768
rect 597738 270756 597744 270768
rect 567896 270728 597744 270756
rect 567896 270716 567902 270728
rect 597738 270716 597744 270728
rect 597796 270716 597802 270768
rect 121454 270580 121460 270632
rect 121512 270620 121518 270632
rect 168098 270620 168104 270632
rect 121512 270592 168104 270620
rect 121512 270580 121518 270592
rect 168098 270580 168104 270592
rect 168156 270580 168162 270632
rect 403618 270580 403624 270632
rect 403676 270620 403682 270632
rect 433426 270620 433432 270632
rect 403676 270592 433432 270620
rect 403676 270580 403682 270592
rect 433426 270580 433432 270592
rect 433484 270580 433490 270632
rect 453298 270580 453304 270632
rect 453356 270620 453362 270632
rect 487798 270620 487804 270632
rect 453356 270592 487804 270620
rect 453356 270580 453362 270592
rect 487798 270580 487804 270592
rect 487856 270580 487862 270632
rect 489638 270580 489644 270632
rect 489696 270620 489702 270632
rect 568206 270620 568212 270632
rect 489696 270592 568212 270620
rect 489696 270580 489702 270592
rect 568206 270580 568212 270592
rect 568264 270580 568270 270632
rect 84102 270444 84108 270496
rect 84160 270484 84166 270496
rect 137462 270484 137468 270496
rect 84160 270456 137468 270484
rect 84160 270444 84166 270456
rect 137462 270444 137468 270456
rect 137520 270444 137526 270496
rect 137646 270444 137652 270496
rect 137704 270484 137710 270496
rect 186130 270484 186136 270496
rect 137704 270456 186136 270484
rect 137704 270444 137710 270456
rect 186130 270444 186136 270456
rect 186188 270444 186194 270496
rect 200758 270444 200764 270496
rect 200816 270484 200822 270496
rect 201862 270484 201868 270496
rect 200816 270456 201868 270484
rect 200816 270444 200822 270456
rect 201862 270444 201868 270456
rect 201920 270444 201926 270496
rect 206830 270444 206836 270496
rect 206888 270484 206894 270496
rect 235810 270484 235816 270496
rect 206888 270456 235816 270484
rect 206888 270444 206894 270456
rect 235810 270444 235816 270456
rect 235868 270444 235874 270496
rect 278406 270444 278412 270496
rect 278464 270484 278470 270496
rect 283834 270484 283840 270496
rect 278464 270456 283840 270484
rect 278464 270444 278470 270456
rect 283834 270444 283840 270456
rect 283892 270444 283898 270496
rect 400858 270444 400864 270496
rect 400916 270484 400922 270496
rect 441614 270484 441620 270496
rect 400916 270456 441620 270484
rect 400916 270444 400922 270456
rect 441614 270444 441620 270456
rect 441672 270444 441678 270496
rect 456426 270444 456432 270496
rect 456484 270484 456490 270496
rect 520274 270484 520280 270496
rect 456484 270456 520280 270484
rect 456484 270444 456490 270456
rect 520274 270444 520280 270456
rect 520332 270444 520338 270496
rect 523126 270444 523132 270496
rect 523184 270484 523190 270496
rect 532786 270484 532792 270496
rect 523184 270456 532792 270484
rect 523184 270444 523190 270456
rect 532786 270444 532792 270456
rect 532844 270444 532850 270496
rect 619634 270484 619640 270496
rect 533356 270456 619640 270484
rect 533356 270416 533384 270456
rect 619634 270444 619640 270456
rect 619692 270444 619698 270496
rect 533172 270388 533384 270416
rect 78858 270308 78864 270360
rect 78916 270348 78922 270360
rect 132494 270348 132500 270360
rect 78916 270320 132500 270348
rect 78916 270308 78922 270320
rect 132494 270308 132500 270320
rect 132552 270308 132558 270360
rect 133782 270308 133788 270360
rect 133840 270348 133846 270360
rect 183646 270348 183652 270360
rect 133840 270320 183652 270348
rect 133840 270308 133846 270320
rect 183646 270308 183652 270320
rect 183704 270308 183710 270360
rect 185302 270308 185308 270360
rect 185360 270348 185366 270360
rect 194410 270348 194416 270360
rect 185360 270320 194416 270348
rect 185360 270308 185366 270320
rect 194410 270308 194416 270320
rect 194468 270308 194474 270360
rect 199930 270308 199936 270360
rect 199988 270348 199994 270360
rect 230842 270348 230848 270360
rect 199988 270320 230848 270348
rect 199988 270308 199994 270320
rect 230842 270308 230848 270320
rect 230900 270308 230906 270360
rect 233050 270308 233056 270360
rect 233108 270348 233114 270360
rect 248230 270348 248236 270360
rect 233108 270320 248236 270348
rect 233108 270308 233114 270320
rect 248230 270308 248236 270320
rect 248288 270308 248294 270360
rect 283098 270308 283104 270360
rect 283156 270348 283162 270360
rect 284662 270348 284668 270360
rect 283156 270320 284668 270348
rect 283156 270308 283162 270320
rect 284662 270308 284668 270320
rect 284720 270308 284726 270360
rect 355042 270308 355048 270360
rect 355100 270348 355106 270360
rect 376938 270348 376944 270360
rect 355100 270320 376944 270348
rect 355100 270308 355106 270320
rect 376938 270308 376944 270320
rect 376996 270308 377002 270360
rect 380526 270308 380532 270360
rect 380584 270348 380590 270360
rect 404354 270348 404360 270360
rect 380584 270320 404360 270348
rect 380584 270308 380590 270320
rect 404354 270308 404360 270320
rect 404412 270308 404418 270360
rect 409598 270308 409604 270360
rect 409656 270348 409662 270360
rect 454034 270348 454040 270360
rect 409656 270320 454040 270348
rect 409656 270308 409662 270320
rect 454034 270308 454040 270320
rect 454092 270308 454098 270360
rect 458818 270308 458824 270360
rect 458876 270348 458882 270360
rect 524414 270348 524420 270360
rect 458876 270320 524420 270348
rect 458876 270308 458882 270320
rect 524414 270308 524420 270320
rect 524472 270308 524478 270360
rect 525610 270308 525616 270360
rect 525668 270348 525674 270360
rect 533172 270348 533200 270388
rect 525668 270320 533200 270348
rect 525668 270308 525674 270320
rect 533522 270308 533528 270360
rect 533580 270348 533586 270360
rect 626534 270348 626540 270360
rect 533580 270320 626540 270348
rect 533580 270308 533586 270320
rect 626534 270308 626540 270320
rect 626592 270308 626598 270360
rect 111978 270172 111984 270224
rect 112036 270212 112042 270224
rect 168742 270212 168748 270224
rect 112036 270184 168748 270212
rect 112036 270172 112042 270184
rect 168742 270172 168748 270184
rect 168800 270172 168806 270224
rect 184842 270172 184848 270224
rect 184900 270212 184906 270224
rect 219342 270212 219348 270224
rect 184900 270184 219348 270212
rect 184900 270172 184906 270184
rect 219342 270172 219348 270184
rect 219400 270172 219406 270224
rect 244366 270172 244372 270224
rect 244424 270212 244430 270224
rect 262306 270212 262312 270224
rect 244424 270184 262312 270212
rect 244424 270172 244430 270184
rect 262306 270172 262312 270184
rect 262364 270172 262370 270224
rect 334342 270172 334348 270224
rect 334400 270212 334406 270224
rect 346394 270212 346400 270224
rect 334400 270184 346400 270212
rect 334400 270172 334406 270184
rect 346394 270172 346400 270184
rect 346452 270172 346458 270224
rect 372246 270172 372252 270224
rect 372304 270212 372310 270224
rect 397454 270212 397460 270224
rect 372304 270184 397460 270212
rect 372304 270172 372310 270184
rect 397454 270172 397460 270184
rect 397512 270172 397518 270224
rect 397914 270172 397920 270224
rect 397972 270212 397978 270224
rect 412634 270212 412640 270224
rect 397972 270184 412640 270212
rect 397972 270172 397978 270184
rect 412634 270172 412640 270184
rect 412692 270172 412698 270224
rect 414658 270172 414664 270224
rect 414716 270212 414722 270224
rect 461210 270212 461216 270224
rect 414716 270184 461216 270212
rect 414716 270172 414722 270184
rect 461210 270172 461216 270184
rect 461268 270172 461274 270224
rect 461394 270172 461400 270224
rect 461452 270212 461458 270224
rect 527174 270212 527180 270224
rect 461452 270184 527180 270212
rect 461452 270172 461458 270184
rect 527174 270172 527180 270184
rect 527232 270172 527238 270224
rect 528370 270172 528376 270224
rect 528428 270212 528434 270224
rect 533246 270212 533252 270224
rect 528428 270184 533252 270212
rect 528428 270172 528434 270184
rect 533246 270172 533252 270184
rect 533304 270172 533310 270224
rect 533522 270172 533528 270224
rect 533580 270212 533586 270224
rect 623958 270212 623964 270224
rect 533580 270184 623964 270212
rect 533580 270172 533586 270184
rect 623958 270172 623964 270184
rect 624016 270172 624022 270224
rect 89622 270036 89628 270088
rect 89680 270076 89686 270088
rect 153010 270076 153016 270088
rect 89680 270048 153016 270076
rect 89680 270036 89686 270048
rect 153010 270036 153016 270048
rect 153068 270036 153074 270088
rect 176562 270036 176568 270088
rect 176620 270076 176626 270088
rect 211154 270076 211160 270088
rect 176620 270048 211160 270076
rect 176620 270036 176626 270048
rect 211154 270036 211160 270048
rect 211212 270036 211218 270088
rect 212442 270036 212448 270088
rect 212500 270076 212506 270088
rect 239950 270076 239956 270088
rect 212500 270048 239956 270076
rect 212500 270036 212506 270048
rect 239950 270036 239956 270048
rect 240008 270036 240014 270088
rect 241882 270036 241888 270088
rect 241940 270076 241946 270088
rect 260650 270076 260656 270088
rect 241940 270048 260656 270076
rect 241940 270036 241946 270048
rect 260650 270036 260656 270048
rect 260708 270036 260714 270088
rect 266170 270036 266176 270088
rect 266228 270076 266234 270088
rect 277210 270076 277216 270088
rect 266228 270048 277216 270076
rect 266228 270036 266234 270048
rect 277210 270036 277216 270048
rect 277268 270036 277274 270088
rect 345290 270036 345296 270088
rect 345348 270076 345354 270088
rect 358814 270076 358820 270088
rect 345348 270048 358820 270076
rect 345348 270036 345354 270048
rect 358814 270036 358820 270048
rect 358872 270036 358878 270088
rect 366634 270036 366640 270088
rect 366692 270076 366698 270088
rect 393314 270076 393320 270088
rect 366692 270048 393320 270076
rect 366692 270036 366698 270048
rect 393314 270036 393320 270048
rect 393372 270036 393378 270088
rect 394694 270036 394700 270088
rect 394752 270076 394758 270088
rect 408770 270076 408776 270088
rect 394752 270048 408776 270076
rect 394752 270036 394758 270048
rect 408770 270036 408776 270048
rect 408828 270036 408834 270088
rect 412450 270036 412456 270088
rect 412508 270076 412514 270088
rect 458174 270076 458180 270088
rect 412508 270048 458180 270076
rect 412508 270036 412514 270048
rect 458174 270036 458180 270048
rect 458232 270036 458238 270088
rect 463510 270036 463516 270088
rect 463568 270076 463574 270088
rect 530762 270076 530768 270088
rect 463568 270048 530768 270076
rect 463568 270036 463574 270048
rect 530762 270036 530768 270048
rect 530820 270036 530826 270088
rect 530946 270036 530952 270088
rect 531004 270076 531010 270088
rect 532970 270076 532976 270088
rect 531004 270048 532976 270076
rect 531004 270036 531010 270048
rect 532970 270036 532976 270048
rect 533028 270036 533034 270088
rect 538306 270076 538312 270088
rect 533356 270048 538312 270076
rect 85482 269900 85488 269952
rect 85540 269940 85546 269952
rect 149698 269940 149704 269952
rect 85540 269912 149704 269940
rect 85540 269900 85546 269912
rect 149698 269900 149704 269912
rect 149756 269900 149762 269952
rect 152826 269900 152832 269952
rect 152884 269940 152890 269952
rect 157150 269940 157156 269952
rect 152884 269912 157156 269940
rect 152884 269900 152890 269912
rect 157150 269900 157156 269912
rect 157208 269900 157214 269952
rect 173802 269900 173808 269952
rect 173860 269940 173866 269952
rect 212626 269940 212632 269952
rect 173860 269912 212632 269940
rect 173860 269900 173866 269912
rect 212626 269900 212632 269912
rect 212684 269900 212690 269952
rect 226610 269900 226616 269952
rect 226668 269940 226674 269952
rect 249886 269940 249892 269952
rect 226668 269912 249892 269940
rect 226668 269900 226674 269912
rect 249886 269900 249892 269912
rect 249944 269900 249950 269952
rect 256878 269900 256884 269952
rect 256936 269940 256942 269952
rect 268930 269940 268936 269952
rect 256936 269912 268936 269940
rect 256936 269900 256942 269912
rect 268930 269900 268936 269912
rect 268988 269900 268994 269952
rect 330202 269900 330208 269952
rect 330260 269940 330266 269952
rect 340874 269940 340880 269952
rect 330260 269912 340880 269940
rect 330260 269900 330266 269912
rect 340874 269900 340880 269912
rect 340932 269900 340938 269952
rect 341794 269900 341800 269952
rect 341852 269940 341858 269952
rect 357434 269940 357440 269952
rect 341852 269912 357440 269940
rect 341852 269900 341858 269912
rect 357434 269900 357440 269912
rect 357492 269900 357498 269952
rect 359182 269900 359188 269952
rect 359240 269940 359246 269952
rect 382274 269940 382280 269952
rect 359240 269912 382280 269940
rect 359240 269900 359246 269912
rect 382274 269900 382280 269912
rect 382332 269900 382338 269952
rect 383010 269900 383016 269952
rect 383068 269940 383074 269952
rect 411254 269940 411260 269952
rect 383068 269912 411260 269940
rect 383068 269900 383074 269912
rect 411254 269900 411260 269912
rect 411312 269900 411318 269952
rect 419626 269900 419632 269952
rect 419684 269940 419690 269952
rect 467926 269940 467932 269952
rect 419684 269912 467932 269940
rect 419684 269900 419690 269912
rect 467926 269900 467932 269912
rect 467984 269900 467990 269952
rect 468478 269900 468484 269952
rect 468536 269940 468542 269952
rect 533356 269940 533384 270048
rect 538306 270036 538312 270048
rect 538364 270036 538370 270088
rect 630674 270076 630680 270088
rect 538876 270048 630680 270076
rect 468536 269912 533384 269940
rect 468536 269900 468542 269912
rect 533982 269900 533988 269952
rect 534040 269940 534046 269952
rect 538876 269940 538904 270048
rect 630674 270036 630680 270048
rect 630732 270036 630738 270088
rect 534040 269912 538904 269940
rect 534040 269900 534046 269912
rect 540514 269900 540520 269952
rect 540572 269940 540578 269952
rect 640518 269940 640524 269952
rect 540572 269912 640524 269940
rect 540572 269900 540578 269912
rect 640518 269900 640524 269912
rect 640576 269900 640582 269952
rect 70578 269764 70584 269816
rect 70636 269804 70642 269816
rect 79318 269804 79324 269816
rect 70636 269776 79324 269804
rect 70636 269764 70642 269776
rect 79318 269764 79324 269776
rect 79376 269764 79382 269816
rect 80054 269764 80060 269816
rect 80112 269804 80118 269816
rect 146386 269804 146392 269816
rect 80112 269776 146392 269804
rect 80112 269764 80118 269776
rect 146386 269764 146392 269776
rect 146444 269764 146450 269816
rect 158622 269764 158628 269816
rect 158680 269804 158686 269816
rect 201034 269804 201040 269816
rect 158680 269776 201040 269804
rect 158680 269764 158686 269776
rect 201034 269764 201040 269776
rect 201092 269764 201098 269816
rect 201678 269764 201684 269816
rect 201736 269804 201742 269816
rect 232498 269804 232504 269816
rect 201736 269776 232504 269804
rect 201736 269764 201742 269776
rect 232498 269764 232504 269776
rect 232556 269764 232562 269816
rect 237190 269764 237196 269816
rect 237248 269804 237254 269816
rect 257338 269804 257344 269816
rect 237248 269776 257344 269804
rect 237248 269764 237254 269776
rect 257338 269764 257344 269776
rect 257396 269764 257402 269816
rect 258534 269764 258540 269816
rect 258592 269804 258598 269816
rect 272242 269804 272248 269816
rect 258592 269776 272248 269804
rect 258592 269764 258598 269776
rect 272242 269764 272248 269776
rect 272300 269764 272306 269816
rect 273070 269764 273076 269816
rect 273128 269804 273134 269816
rect 282178 269804 282184 269816
rect 273128 269776 282184 269804
rect 273128 269764 273134 269776
rect 282178 269764 282184 269776
rect 282236 269764 282242 269816
rect 326890 269764 326896 269816
rect 326948 269804 326954 269816
rect 335538 269804 335544 269816
rect 326948 269776 335544 269804
rect 326948 269764 326954 269776
rect 335538 269764 335544 269776
rect 335596 269764 335602 269816
rect 335998 269764 336004 269816
rect 336056 269804 336062 269816
rect 349154 269804 349160 269816
rect 336056 269776 349160 269804
rect 336056 269764 336062 269776
rect 349154 269764 349160 269776
rect 349212 269764 349218 269816
rect 351730 269764 351736 269816
rect 351788 269804 351794 269816
rect 371234 269804 371240 269816
rect 351788 269776 371240 269804
rect 351788 269764 351794 269776
rect 371234 269764 371240 269776
rect 371292 269764 371298 269816
rect 376570 269764 376576 269816
rect 376628 269804 376634 269816
rect 407114 269804 407120 269816
rect 376628 269776 407120 269804
rect 376628 269764 376634 269776
rect 407114 269764 407120 269776
rect 407172 269764 407178 269816
rect 417142 269764 417148 269816
rect 417200 269804 417206 269816
rect 465074 269804 465080 269816
rect 417200 269776 465080 269804
rect 417200 269764 417206 269776
rect 465074 269764 465080 269776
rect 465132 269764 465138 269816
rect 465994 269764 466000 269816
rect 466052 269804 466058 269816
rect 532234 269804 532240 269816
rect 466052 269776 532240 269804
rect 466052 269764 466058 269776
rect 532234 269764 532240 269776
rect 532292 269764 532298 269816
rect 538858 269804 538864 269816
rect 532436 269776 538864 269804
rect 122742 269628 122748 269680
rect 122800 269668 122806 269680
rect 176194 269668 176200 269680
rect 122800 269640 176200 269668
rect 122800 269628 122806 269640
rect 176194 269628 176200 269640
rect 176252 269628 176258 269680
rect 183462 269628 183468 269680
rect 183520 269668 183526 269680
rect 205450 269668 205456 269680
rect 183520 269640 205456 269668
rect 183520 269628 183526 269640
rect 205450 269628 205456 269640
rect 205508 269628 205514 269680
rect 392026 269628 392032 269680
rect 392084 269668 392090 269680
rect 401686 269668 401692 269680
rect 392084 269640 401692 269668
rect 392084 269628 392090 269640
rect 401686 269628 401692 269640
rect 401744 269628 401750 269680
rect 404354 269628 404360 269680
rect 404412 269668 404418 269680
rect 423674 269668 423680 269680
rect 404412 269640 423680 269668
rect 404412 269628 404418 269640
rect 423674 269628 423680 269640
rect 423732 269628 423738 269680
rect 423858 269628 423864 269680
rect 423916 269668 423922 269680
rect 451366 269668 451372 269680
rect 423916 269640 451372 269668
rect 423916 269628 423922 269640
rect 451366 269628 451372 269640
rect 451424 269628 451430 269680
rect 453574 269628 453580 269680
rect 453632 269668 453638 269680
rect 509234 269668 509240 269680
rect 453632 269640 509240 269668
rect 453632 269628 453638 269640
rect 509234 269628 509240 269640
rect 509292 269628 509298 269680
rect 532436 269668 532464 269776
rect 538858 269764 538864 269776
rect 538916 269764 538922 269816
rect 539042 269764 539048 269816
rect 539100 269804 539106 269816
rect 541618 269804 541624 269816
rect 539100 269776 541624 269804
rect 539100 269764 539106 269776
rect 541618 269764 541624 269776
rect 541676 269764 541682 269816
rect 541802 269764 541808 269816
rect 541860 269804 541866 269816
rect 637574 269804 637580 269816
rect 541860 269776 637580 269804
rect 541860 269764 541866 269776
rect 637574 269764 637580 269776
rect 637632 269764 637638 269816
rect 509712 269640 532464 269668
rect 129642 269492 129648 269544
rect 129700 269532 129706 269544
rect 181162 269532 181168 269544
rect 129700 269504 181168 269532
rect 129700 269492 129706 269504
rect 181162 269492 181168 269504
rect 181220 269492 181226 269544
rect 204162 269492 204168 269544
rect 204220 269532 204226 269544
rect 223482 269532 223488 269544
rect 204220 269504 223488 269532
rect 204220 269492 204226 269504
rect 223482 269492 223488 269504
rect 223540 269492 223546 269544
rect 401686 269492 401692 269544
rect 401744 269532 401750 269544
rect 416774 269532 416780 269544
rect 401744 269504 416780 269532
rect 401744 269492 401750 269504
rect 416774 269492 416780 269504
rect 416832 269492 416838 269544
rect 424594 269492 424600 269544
rect 424652 269532 424658 269544
rect 475010 269532 475016 269544
rect 424652 269504 475016 269532
rect 424652 269492 424658 269504
rect 475010 269492 475016 269504
rect 475068 269492 475074 269544
rect 492766 269492 492772 269544
rect 492824 269532 492830 269544
rect 509712 269532 509740 269640
rect 532786 269628 532792 269680
rect 532844 269668 532850 269680
rect 615678 269668 615684 269680
rect 532844 269640 615684 269668
rect 532844 269628 532850 269640
rect 615678 269628 615684 269640
rect 615736 269628 615742 269680
rect 492824 269504 509740 269532
rect 492824 269492 492830 269504
rect 509878 269492 509884 269544
rect 509936 269532 509942 269544
rect 596174 269532 596180 269544
rect 509936 269504 596180 269532
rect 509936 269492 509942 269504
rect 596174 269492 596180 269504
rect 596232 269492 596238 269544
rect 126882 269356 126888 269408
rect 126940 269396 126946 269408
rect 178310 269396 178316 269408
rect 126940 269368 178316 269396
rect 126940 269356 126946 269368
rect 178310 269356 178316 269368
rect 178368 269356 178374 269408
rect 408310 269356 408316 269408
rect 408368 269396 408374 269408
rect 426526 269396 426532 269408
rect 408368 269368 426532 269396
rect 408368 269356 408374 269368
rect 426526 269356 426532 269368
rect 426584 269356 426590 269408
rect 441614 269356 441620 269408
rect 441672 269396 441678 269408
rect 458450 269396 458456 269408
rect 441672 269368 458456 269396
rect 441672 269356 441678 269368
rect 458450 269356 458456 269368
rect 458508 269356 458514 269408
rect 470962 269356 470968 269408
rect 471020 269396 471026 269408
rect 538674 269396 538680 269408
rect 471020 269368 538680 269396
rect 471020 269356 471026 269368
rect 538674 269356 538680 269368
rect 538732 269356 538738 269408
rect 538858 269356 538864 269408
rect 538916 269396 538922 269408
rect 572714 269396 572720 269408
rect 538916 269368 572720 269396
rect 538916 269356 538922 269368
rect 572714 269356 572720 269368
rect 572772 269356 572778 269408
rect 143902 269220 143908 269272
rect 143960 269260 143966 269272
rect 191098 269260 191104 269272
rect 143960 269232 191104 269260
rect 143960 269220 143966 269232
rect 191098 269220 191104 269232
rect 191156 269220 191162 269272
rect 282730 269220 282736 269272
rect 282788 269260 282794 269272
rect 288802 269260 288808 269272
rect 282788 269232 288808 269260
rect 282788 269220 282794 269232
rect 288802 269220 288808 269232
rect 288860 269220 288866 269272
rect 474274 269220 474280 269272
rect 474332 269260 474338 269272
rect 546494 269260 546500 269272
rect 474332 269232 546500 269260
rect 474332 269220 474338 269232
rect 546494 269220 546500 269232
rect 546552 269220 546558 269272
rect 319438 269084 319444 269136
rect 319496 269124 319502 269136
rect 325694 269124 325700 269136
rect 319496 269096 325700 269124
rect 319496 269084 319502 269096
rect 325694 269084 325700 269096
rect 325752 269084 325758 269136
rect 118602 269016 118608 269068
rect 118660 269056 118666 269068
rect 174538 269056 174544 269068
rect 118660 269028 174544 269056
rect 118660 269016 118666 269028
rect 174538 269016 174544 269028
rect 174596 269016 174602 269068
rect 175090 269016 175096 269068
rect 175148 269056 175154 269068
rect 177666 269056 177672 269068
rect 175148 269028 177672 269056
rect 175148 269016 175154 269028
rect 177666 269016 177672 269028
rect 177724 269016 177730 269068
rect 273254 269016 273260 269068
rect 273312 269056 273318 269068
rect 275554 269056 275560 269068
rect 273312 269028 275560 269056
rect 273312 269016 273318 269028
rect 275554 269016 275560 269028
rect 275612 269016 275618 269068
rect 436554 269016 436560 269068
rect 436612 269056 436618 269068
rect 491662 269056 491668 269068
rect 436612 269028 491668 269056
rect 436612 269016 436618 269028
rect 491662 269016 491668 269028
rect 491720 269016 491726 269068
rect 493318 269016 493324 269068
rect 493376 269056 493382 269068
rect 574094 269056 574100 269068
rect 493376 269028 574100 269056
rect 493376 269016 493382 269028
rect 574094 269016 574100 269028
rect 574152 269016 574158 269068
rect 115842 268880 115848 268932
rect 115900 268920 115906 268932
rect 115900 268892 166304 268920
rect 115900 268880 115906 268892
rect 110322 268744 110328 268796
rect 110380 268784 110386 268796
rect 110380 268756 164740 268784
rect 110380 268744 110386 268756
rect 104986 268608 104992 268660
rect 105044 268648 105050 268660
rect 163774 268648 163780 268660
rect 105044 268620 163780 268648
rect 105044 268608 105050 268620
rect 163774 268608 163780 268620
rect 163832 268608 163838 268660
rect 99282 268472 99288 268524
rect 99340 268512 99346 268524
rect 160462 268512 160468 268524
rect 99340 268484 160468 268512
rect 99340 268472 99346 268484
rect 160462 268472 160468 268484
rect 160520 268472 160526 268524
rect 164712 268512 164740 268756
rect 166276 268648 166304 268892
rect 188890 268880 188896 268932
rect 188948 268920 188954 268932
rect 190546 268920 190552 268932
rect 188948 268892 190552 268920
rect 188948 268880 188954 268892
rect 190546 268880 190552 268892
rect 190604 268880 190610 268932
rect 382366 268880 382372 268932
rect 382424 268920 382430 268932
rect 415394 268920 415400 268932
rect 382424 268892 415400 268920
rect 382424 268880 382430 268892
rect 415394 268880 415400 268892
rect 415452 268880 415458 268932
rect 433702 268880 433708 268932
rect 433760 268920 433766 268932
rect 488534 268920 488540 268932
rect 433760 268892 488540 268920
rect 433760 268880 433766 268892
rect 488534 268880 488540 268892
rect 488592 268880 488598 268932
rect 498286 268880 498292 268932
rect 498344 268920 498350 268932
rect 580994 268920 581000 268932
rect 498344 268892 581000 268920
rect 498344 268880 498350 268892
rect 580994 268880 581000 268892
rect 581052 268880 581058 268932
rect 166994 268744 167000 268796
rect 167052 268784 167058 268796
rect 181990 268784 181996 268796
rect 167052 268756 181996 268784
rect 167052 268744 167058 268756
rect 181990 268744 181996 268756
rect 182048 268744 182054 268796
rect 200574 268744 200580 268796
rect 200632 268784 200638 268796
rect 231302 268784 231308 268796
rect 200632 268756 231308 268784
rect 200632 268744 200638 268756
rect 231302 268744 231308 268756
rect 231360 268744 231366 268796
rect 387334 268744 387340 268796
rect 387392 268784 387398 268796
rect 422294 268784 422300 268796
rect 387392 268756 422300 268784
rect 387392 268744 387398 268756
rect 422294 268744 422300 268756
rect 422352 268744 422358 268796
rect 438670 268744 438676 268796
rect 438728 268784 438734 268796
rect 495434 268784 495440 268796
rect 438728 268756 495440 268784
rect 438728 268744 438734 268756
rect 495434 268744 495440 268756
rect 495492 268744 495498 268796
rect 500770 268744 500776 268796
rect 500828 268784 500834 268796
rect 583754 268784 583760 268796
rect 500828 268756 583760 268784
rect 500828 268744 500834 268756
rect 583754 268744 583760 268756
rect 583812 268744 583818 268796
rect 171226 268648 171232 268660
rect 166276 268620 171232 268648
rect 171226 268608 171232 268620
rect 171284 268608 171290 268660
rect 176930 268608 176936 268660
rect 176988 268648 176994 268660
rect 215110 268648 215116 268660
rect 176988 268620 215116 268648
rect 176988 268608 176994 268620
rect 215110 268608 215116 268620
rect 215168 268608 215174 268660
rect 224218 268608 224224 268660
rect 224276 268648 224282 268660
rect 243262 268648 243268 268660
rect 224276 268620 243268 268648
rect 224276 268608 224282 268620
rect 243262 268608 243268 268620
rect 243320 268608 243326 268660
rect 352558 268608 352564 268660
rect 352616 268648 352622 268660
rect 372614 268648 372620 268660
rect 352616 268620 372620 268648
rect 352616 268608 352622 268620
rect 372614 268608 372620 268620
rect 372672 268608 372678 268660
rect 393314 268608 393320 268660
rect 393372 268648 393378 268660
rect 429194 268648 429200 268660
rect 393372 268620 429200 268648
rect 393372 268608 393378 268620
rect 429194 268608 429200 268620
rect 429252 268608 429258 268660
rect 441154 268608 441160 268660
rect 441212 268648 441218 268660
rect 500126 268648 500132 268660
rect 441212 268620 500132 268648
rect 441212 268608 441218 268620
rect 500126 268608 500132 268620
rect 500184 268608 500190 268660
rect 503254 268608 503260 268660
rect 503312 268648 503318 268660
rect 587894 268648 587900 268660
rect 503312 268620 587900 268648
rect 503312 268608 503318 268620
rect 587894 268608 587900 268620
rect 587952 268608 587958 268660
rect 167914 268512 167920 268524
rect 164712 268484 167920 268512
rect 167914 268472 167920 268484
rect 167972 268472 167978 268524
rect 180610 268472 180616 268524
rect 180668 268512 180674 268524
rect 217594 268512 217600 268524
rect 180668 268484 217600 268512
rect 180668 268472 180674 268484
rect 217594 268472 217600 268484
rect 217652 268472 217658 268524
rect 231670 268472 231676 268524
rect 231728 268512 231734 268524
rect 253198 268512 253204 268524
rect 231728 268484 253204 268512
rect 231728 268472 231734 268484
rect 253198 268472 253204 268484
rect 253256 268472 253262 268524
rect 338482 268472 338488 268524
rect 338540 268512 338546 268524
rect 352098 268512 352104 268524
rect 338540 268484 352104 268512
rect 338540 268472 338546 268484
rect 352098 268472 352104 268484
rect 352156 268472 352162 268524
rect 367462 268472 367468 268524
rect 367520 268512 367526 268524
rect 393498 268512 393504 268524
rect 367520 268484 393504 268512
rect 367520 268472 367526 268484
rect 393498 268472 393504 268484
rect 393556 268472 393562 268524
rect 397270 268472 397276 268524
rect 397328 268512 397334 268524
rect 436094 268512 436100 268524
rect 397328 268484 436100 268512
rect 397328 268472 397334 268484
rect 436094 268472 436100 268484
rect 436152 268472 436158 268524
rect 446122 268472 446128 268524
rect 446180 268512 446186 268524
rect 506474 268512 506480 268524
rect 446180 268484 506480 268512
rect 446180 268472 446186 268484
rect 506474 268472 506480 268484
rect 506532 268472 506538 268524
rect 508222 268472 508228 268524
rect 508280 268512 508286 268524
rect 594794 268512 594800 268524
rect 508280 268484 594800 268512
rect 508280 268472 508286 268484
rect 594794 268472 594800 268484
rect 594852 268472 594858 268524
rect 92382 268336 92388 268388
rect 92440 268376 92446 268388
rect 155494 268376 155500 268388
rect 92440 268348 155500 268376
rect 92440 268336 92446 268348
rect 155494 268336 155500 268348
rect 155552 268336 155558 268388
rect 161566 268336 161572 268388
rect 161624 268376 161630 268388
rect 203518 268376 203524 268388
rect 161624 268348 203524 268376
rect 161624 268336 161630 268348
rect 203518 268336 203524 268348
rect 203576 268336 203582 268388
rect 210694 268336 210700 268388
rect 210752 268376 210758 268388
rect 236638 268376 236644 268388
rect 210752 268348 236644 268376
rect 210752 268336 210758 268348
rect 236638 268336 236644 268348
rect 236696 268336 236702 268388
rect 252646 268336 252652 268388
rect 252704 268376 252710 268388
rect 268102 268376 268108 268388
rect 252704 268348 268108 268376
rect 252704 268336 252710 268348
rect 268102 268336 268108 268348
rect 268160 268336 268166 268388
rect 348786 268336 348792 268388
rect 348844 268376 348850 268388
rect 367094 268376 367100 268388
rect 348844 268348 367100 268376
rect 348844 268336 348850 268348
rect 367094 268336 367100 268348
rect 367152 268336 367158 268388
rect 372430 268336 372436 268388
rect 372488 268376 372494 268388
rect 400490 268376 400496 268388
rect 372488 268348 400496 268376
rect 372488 268336 372494 268348
rect 400490 268336 400496 268348
rect 400548 268336 400554 268388
rect 402238 268336 402244 268388
rect 402296 268376 402302 268388
rect 443086 268376 443092 268388
rect 402296 268348 443092 268376
rect 402296 268336 402302 268348
rect 443086 268336 443092 268348
rect 443144 268336 443150 268388
rect 461854 268336 461860 268388
rect 461912 268376 461918 268388
rect 528554 268376 528560 268388
rect 461912 268348 528560 268376
rect 461912 268336 461918 268348
rect 528554 268336 528560 268348
rect 528612 268336 528618 268388
rect 541342 268336 541348 268388
rect 541400 268376 541406 268388
rect 641714 268376 641720 268388
rect 541400 268348 641720 268376
rect 541400 268336 541406 268348
rect 641714 268336 641720 268348
rect 641772 268336 641778 268388
rect 140682 268200 140688 268252
rect 140740 268240 140746 268252
rect 188614 268240 188620 268252
rect 140740 268212 188620 268240
rect 140740 268200 140746 268212
rect 188614 268200 188620 268212
rect 188672 268200 188678 268252
rect 416222 268200 416228 268252
rect 416280 268240 416286 268252
rect 447134 268240 447140 268252
rect 416280 268212 447140 268240
rect 416280 268200 416286 268212
rect 447134 268200 447140 268212
rect 447192 268200 447198 268252
rect 448422 268200 448428 268252
rect 448480 268240 448486 268252
rect 494054 268240 494060 268252
rect 448480 268212 494060 268240
rect 448480 268200 448486 268212
rect 494054 268200 494060 268212
rect 494112 268200 494118 268252
rect 495802 268200 495808 268252
rect 495860 268240 495866 268252
rect 576854 268240 576860 268252
rect 495860 268212 576860 268240
rect 495860 268200 495866 268212
rect 576854 268200 576860 268212
rect 576912 268200 576918 268252
rect 151722 268064 151728 268116
rect 151780 268104 151786 268116
rect 196066 268104 196072 268116
rect 151780 268076 196072 268104
rect 151780 268064 151786 268076
rect 196066 268064 196072 268076
rect 196124 268064 196130 268116
rect 422294 268064 422300 268116
rect 422352 268104 422358 268116
rect 444374 268104 444380 268116
rect 422352 268076 444380 268104
rect 422352 268064 422358 268076
rect 444374 268064 444380 268076
rect 444432 268064 444438 268116
rect 527174 268064 527180 268116
rect 527232 268104 527238 268116
rect 607398 268104 607404 268116
rect 527232 268076 607404 268104
rect 527232 268064 527238 268076
rect 607398 268064 607404 268076
rect 607456 268064 607462 268116
rect 490834 267928 490840 267980
rect 490892 267968 490898 267980
rect 569954 267968 569960 267980
rect 490892 267940 569960 267968
rect 490892 267928 490898 267940
rect 569954 267928 569960 267940
rect 570012 267928 570018 267980
rect 135622 267792 135628 267844
rect 135680 267832 135686 267844
rect 135680 267804 139440 267832
rect 135680 267792 135686 267804
rect 130378 267656 130384 267708
rect 130436 267696 130442 267708
rect 138106 267696 138112 267708
rect 130436 267668 138112 267696
rect 130436 267656 130442 267668
rect 138106 267656 138112 267668
rect 138164 267656 138170 267708
rect 139412 267696 139440 267804
rect 276474 267724 276480 267776
rect 276532 267764 276538 267776
rect 278038 267764 278044 267776
rect 276532 267736 278044 267764
rect 276532 267724 276538 267736
rect 278038 267724 278044 267736
rect 278096 267724 278102 267776
rect 186958 267696 186964 267708
rect 139412 267668 186964 267696
rect 186958 267656 186964 267668
rect 187016 267656 187022 267708
rect 187142 267656 187148 267708
rect 187200 267696 187206 267708
rect 195238 267696 195244 267708
rect 187200 267668 195244 267696
rect 187200 267656 187206 267668
rect 195238 267656 195244 267668
rect 195296 267656 195302 267708
rect 353386 267656 353392 267708
rect 353444 267696 353450 267708
rect 374454 267696 374460 267708
rect 353444 267668 374460 267696
rect 353444 267656 353450 267668
rect 374454 267656 374460 267668
rect 374512 267656 374518 267708
rect 378226 267656 378232 267708
rect 378284 267696 378290 267708
rect 394694 267696 394700 267708
rect 378284 267668 394700 267696
rect 378284 267656 378290 267668
rect 394694 267656 394700 267668
rect 394752 267656 394758 267708
rect 408034 267656 408040 267708
rect 408092 267696 408098 267708
rect 423858 267696 423864 267708
rect 408092 267668 423864 267696
rect 408092 267656 408098 267668
rect 423858 267656 423864 267668
rect 423916 267656 423922 267708
rect 445294 267656 445300 267708
rect 445352 267696 445358 267708
rect 498838 267696 498844 267708
rect 445352 267668 498844 267696
rect 445352 267656 445358 267668
rect 498838 267656 498844 267668
rect 498896 267656 498902 267708
rect 509878 267656 509884 267708
rect 509936 267696 509942 267708
rect 567838 267696 567844 267708
rect 509936 267668 567844 267696
rect 509936 267656 509942 267668
rect 567838 267656 567844 267668
rect 567896 267656 567902 267708
rect 111702 267520 111708 267572
rect 111760 267560 111766 267572
rect 169570 267560 169576 267572
rect 111760 267532 169576 267560
rect 111760 267520 111766 267532
rect 169570 267520 169576 267532
rect 169628 267520 169634 267572
rect 178678 267520 178684 267572
rect 178736 267560 178742 267572
rect 209314 267560 209320 267572
rect 178736 267532 209320 267560
rect 178736 267520 178742 267532
rect 209314 267520 209320 267532
rect 209372 267520 209378 267572
rect 368290 267520 368296 267572
rect 368348 267560 368354 267572
rect 385678 267560 385684 267572
rect 368348 267532 385684 267560
rect 368348 267520 368354 267532
rect 385678 267520 385684 267532
rect 385736 267520 385742 267572
rect 403066 267520 403072 267572
rect 403124 267560 403130 267572
rect 422294 267560 422300 267572
rect 403124 267532 422300 267560
rect 403124 267520 403130 267532
rect 422294 267520 422300 267532
rect 422352 267520 422358 267572
rect 428734 267520 428740 267572
rect 428792 267560 428798 267572
rect 447778 267560 447784 267572
rect 428792 267532 447784 267560
rect 428792 267520 428798 267532
rect 447778 267520 447784 267532
rect 447836 267520 447842 267572
rect 450262 267520 450268 267572
rect 450320 267560 450326 267572
rect 505738 267560 505744 267572
rect 450320 267532 505744 267560
rect 450320 267520 450326 267532
rect 505738 267520 505744 267532
rect 505796 267520 505802 267572
rect 514846 267520 514852 267572
rect 514904 267560 514910 267572
rect 576118 267560 576124 267572
rect 514904 267532 576124 267560
rect 514904 267520 514910 267532
rect 576118 267520 576124 267532
rect 576176 267520 576182 267572
rect 86218 267384 86224 267436
rect 86276 267424 86282 267436
rect 144730 267424 144736 267436
rect 86276 267396 144736 267424
rect 86276 267384 86282 267396
rect 144730 267384 144736 267396
rect 144788 267384 144794 267436
rect 153838 267384 153844 267436
rect 153896 267424 153902 267436
rect 184474 267424 184480 267436
rect 153896 267396 184480 267424
rect 153896 267384 153902 267396
rect 184474 267384 184480 267396
rect 184532 267384 184538 267436
rect 190546 267384 190552 267436
rect 190604 267424 190610 267436
rect 190604 267396 192156 267424
rect 190604 267384 190610 267396
rect 104802 267248 104808 267300
rect 104860 267288 104866 267300
rect 164602 267288 164608 267300
rect 104860 267260 164608 267288
rect 104860 267248 104866 267260
rect 164602 267248 164608 267260
rect 164660 267248 164666 267300
rect 191926 267288 191932 267300
rect 180766 267260 191932 267288
rect 79318 267112 79324 267164
rect 79376 267152 79382 267164
rect 140590 267152 140596 267164
rect 79376 267124 140596 267152
rect 79376 267112 79382 267124
rect 140590 267112 140596 267124
rect 140648 267112 140654 267164
rect 145558 267112 145564 267164
rect 145616 267152 145622 267164
rect 180766 267152 180794 267260
rect 191926 267248 191932 267260
rect 191984 267248 191990 267300
rect 192128 267288 192156 267396
rect 195238 267384 195244 267436
rect 195296 267424 195302 267436
rect 219250 267424 219256 267436
rect 195296 267396 219256 267424
rect 195296 267384 195302 267396
rect 219250 267384 219256 267396
rect 219308 267384 219314 267436
rect 223482 267384 223488 267436
rect 223540 267424 223546 267436
rect 234154 267424 234160 267436
rect 223540 267396 234160 267424
rect 223540 267384 223546 267396
rect 234154 267384 234160 267396
rect 234212 267384 234218 267436
rect 243722 267384 243728 267436
rect 243780 267424 243786 267436
rect 251542 267424 251548 267436
rect 243780 267396 251548 267424
rect 243780 267384 243786 267396
rect 251542 267384 251548 267396
rect 251600 267384 251606 267436
rect 315298 267384 315304 267436
rect 315356 267424 315362 267436
rect 319070 267424 319076 267436
rect 315356 267396 319076 267424
rect 315356 267384 315362 267396
rect 319070 267384 319076 267396
rect 319128 267384 319134 267436
rect 340966 267384 340972 267436
rect 341024 267424 341030 267436
rect 355318 267424 355324 267436
rect 341024 267396 355324 267424
rect 341024 267384 341030 267396
rect 355318 267384 355324 267396
rect 355376 267384 355382 267436
rect 371602 267384 371608 267436
rect 371660 267424 371666 267436
rect 373258 267424 373264 267436
rect 371660 267396 373264 267424
rect 371660 267384 371666 267396
rect 373258 267384 373264 267396
rect 373316 267384 373322 267436
rect 380710 267384 380716 267436
rect 380768 267424 380774 267436
rect 397914 267424 397920 267436
rect 380768 267396 397920 267424
rect 380768 267384 380774 267396
rect 397914 267384 397920 267396
rect 397972 267384 397978 267436
rect 404722 267384 404728 267436
rect 404780 267424 404786 267436
rect 416222 267424 416228 267436
rect 404780 267396 416228 267424
rect 404780 267384 404786 267396
rect 416222 267384 416228 267396
rect 416280 267384 416286 267436
rect 421282 267384 421288 267436
rect 421340 267424 421346 267436
rect 440878 267424 440884 267436
rect 421340 267396 440884 267424
rect 421340 267384 421346 267396
rect 440878 267384 440884 267396
rect 440936 267384 440942 267436
rect 447778 267384 447784 267436
rect 447836 267424 447842 267436
rect 456058 267424 456064 267436
rect 447836 267396 456064 267424
rect 447836 267384 447842 267396
rect 456058 267384 456064 267396
rect 456116 267384 456122 267436
rect 460198 267384 460204 267436
rect 460256 267424 460262 267436
rect 516778 267424 516784 267436
rect 460256 267396 516784 267424
rect 460256 267384 460262 267396
rect 516778 267384 516784 267396
rect 516836 267384 516842 267436
rect 519814 267384 519820 267436
rect 519872 267424 519878 267436
rect 583018 267424 583024 267436
rect 519872 267396 583024 267424
rect 519872 267384 519878 267396
rect 583018 267384 583024 267396
rect 583076 267384 583082 267436
rect 224218 267288 224224 267300
rect 192128 267260 224224 267288
rect 224218 267248 224224 267260
rect 224276 267248 224282 267300
rect 233878 267248 233884 267300
rect 233936 267288 233942 267300
rect 244090 267288 244096 267300
rect 233936 267260 244096 267288
rect 233936 267248 233942 267260
rect 244090 267248 244096 267260
rect 244148 267248 244154 267300
rect 249058 267248 249064 267300
rect 249116 267288 249122 267300
rect 250714 267288 250720 267300
rect 249116 267260 250720 267288
rect 249116 267248 249122 267260
rect 250714 267248 250720 267260
rect 250772 267248 250778 267300
rect 321922 267248 321928 267300
rect 321980 267288 321986 267300
rect 327718 267288 327724 267300
rect 321980 267260 327724 267288
rect 321980 267248 321986 267260
rect 327718 267248 327724 267260
rect 327776 267248 327782 267300
rect 350902 267248 350908 267300
rect 350960 267288 350966 267300
rect 362218 267288 362224 267300
rect 350960 267260 362224 267288
rect 350960 267248 350966 267260
rect 362218 267248 362224 267260
rect 362276 267248 362282 267300
rect 373258 267248 373264 267300
rect 373316 267288 373322 267300
rect 392026 267288 392032 267300
rect 373316 267260 392032 267288
rect 373316 267248 373322 267260
rect 392026 267248 392032 267260
rect 392084 267248 392090 267300
rect 398098 267248 398104 267300
rect 398156 267288 398162 267300
rect 417418 267288 417424 267300
rect 398156 267260 417424 267288
rect 398156 267248 398162 267260
rect 417418 267248 417424 267260
rect 417476 267248 417482 267300
rect 432874 267248 432880 267300
rect 432932 267288 432938 267300
rect 453298 267288 453304 267300
rect 432932 267260 453304 267288
rect 432932 267248 432938 267260
rect 453298 267248 453304 267260
rect 453356 267248 453362 267300
rect 459370 267248 459376 267300
rect 459428 267288 459434 267300
rect 460842 267288 460848 267300
rect 459428 267260 460848 267288
rect 459428 267248 459434 267260
rect 460842 267248 460848 267260
rect 460900 267248 460906 267300
rect 465166 267248 465172 267300
rect 465224 267288 465230 267300
rect 523678 267288 523684 267300
rect 465224 267260 523684 267288
rect 465224 267248 465230 267260
rect 523678 267248 523684 267260
rect 523736 267248 523742 267300
rect 524782 267248 524788 267300
rect 524840 267288 524846 267300
rect 611998 267288 612004 267300
rect 524840 267260 612004 267288
rect 524840 267248 524846 267260
rect 611998 267248 612004 267260
rect 612056 267248 612062 267300
rect 145616 267124 180794 267152
rect 145616 267112 145622 267124
rect 199378 267112 199384 267164
rect 199436 267152 199442 267164
rect 204346 267152 204352 267164
rect 199436 267124 204352 267152
rect 199436 267112 199442 267124
rect 204346 267112 204352 267124
rect 204404 267112 204410 267164
rect 205450 267112 205456 267164
rect 205508 267152 205514 267164
rect 218422 267152 218428 267164
rect 205508 267124 218428 267152
rect 205508 267112 205514 267124
rect 218422 267112 218428 267124
rect 218480 267112 218486 267164
rect 220078 267112 220084 267164
rect 220136 267152 220142 267164
rect 239122 267152 239128 267164
rect 220136 267124 239128 267152
rect 220136 267112 220142 267124
rect 239122 267112 239128 267124
rect 239180 267112 239186 267164
rect 246942 267112 246948 267164
rect 247000 267152 247006 267164
rect 263962 267152 263968 267164
rect 247000 267124 263968 267152
rect 247000 267112 247006 267124
rect 263962 267112 263968 267124
rect 264020 267112 264026 267164
rect 313642 267112 313648 267164
rect 313700 267152 313706 267164
rect 317414 267152 317420 267164
rect 313700 267124 317420 267152
rect 313700 267112 313706 267124
rect 317414 267112 317420 267124
rect 317472 267112 317478 267164
rect 365806 267112 365812 267164
rect 365864 267152 365870 267164
rect 381538 267152 381544 267164
rect 365864 267124 381544 267152
rect 365864 267112 365870 267124
rect 381538 267112 381544 267124
rect 381596 267112 381602 267164
rect 383194 267112 383200 267164
rect 383252 267152 383258 267164
rect 401686 267152 401692 267164
rect 383252 267124 401692 267152
rect 383252 267112 383258 267124
rect 401686 267112 401692 267124
rect 401744 267112 401750 267164
rect 413002 267112 413008 267164
rect 413060 267152 413066 267164
rect 441614 267152 441620 267164
rect 413060 267124 441620 267152
rect 413060 267112 413066 267124
rect 441614 267112 441620 267124
rect 441672 267112 441678 267164
rect 455138 267112 455144 267164
rect 455196 267152 455202 267164
rect 515398 267152 515404 267164
rect 455196 267124 515404 267152
rect 455196 267112 455202 267124
rect 515398 267112 515404 267124
rect 515456 267112 515462 267164
rect 517238 267112 517244 267164
rect 517296 267152 517302 267164
rect 527174 267152 527180 267164
rect 517296 267124 527180 267152
rect 517296 267112 517302 267124
rect 527174 267112 527180 267124
rect 527232 267112 527238 267164
rect 529658 267112 529664 267164
rect 529716 267152 529722 267164
rect 617518 267152 617524 267164
rect 529716 267124 617524 267152
rect 529716 267112 529722 267124
rect 617518 267112 617524 267124
rect 617576 267112 617582 267164
rect 90358 266976 90364 267028
rect 90416 267016 90422 267028
rect 151354 267016 151360 267028
rect 90416 266988 151360 267016
rect 90416 266976 90422 266988
rect 151354 266976 151360 266988
rect 151412 266976 151418 267028
rect 159450 266976 159456 267028
rect 159508 267016 159514 267028
rect 162118 267016 162124 267028
rect 159508 266988 162124 267016
rect 159508 266976 159514 266988
rect 162118 266976 162124 266988
rect 162176 266976 162182 267028
rect 168098 266976 168104 267028
rect 168156 267016 168162 267028
rect 177022 267016 177028 267028
rect 168156 266988 177028 267016
rect 168156 266976 168162 266988
rect 177022 266976 177028 266988
rect 177080 266976 177086 267028
rect 177666 266976 177672 267028
rect 177724 267016 177730 267028
rect 214282 267016 214288 267028
rect 177724 266988 214288 267016
rect 177724 266976 177730 266988
rect 214282 266976 214288 266988
rect 214340 266976 214346 267028
rect 218698 266976 218704 267028
rect 218756 267016 218762 267028
rect 220906 267016 220912 267028
rect 218756 266988 220912 267016
rect 218756 266976 218762 266988
rect 220906 266976 220912 266988
rect 220964 266976 220970 267028
rect 228358 266976 228364 267028
rect 228416 267016 228422 267028
rect 249058 267016 249064 267028
rect 228416 266988 249064 267016
rect 228416 266976 228422 266988
rect 249058 266976 249064 266988
rect 249116 266976 249122 267028
rect 255958 266976 255964 267028
rect 256016 267016 256022 267028
rect 258994 267016 259000 267028
rect 256016 266988 259000 267016
rect 256016 266976 256022 266988
rect 258994 266976 259000 266988
rect 259052 266976 259058 267028
rect 286318 266976 286324 267028
rect 286376 267016 286382 267028
rect 287974 267016 287980 267028
rect 286376 266988 287980 267016
rect 286376 266976 286382 266988
rect 287974 266976 287980 266988
rect 288032 266976 288038 267028
rect 312814 266976 312820 267028
rect 312872 267016 312878 267028
rect 316034 267016 316040 267028
rect 312872 266988 316040 267016
rect 312872 266976 312878 266988
rect 316034 266976 316040 266988
rect 316092 266976 316098 267028
rect 317782 266976 317788 267028
rect 317840 267016 317846 267028
rect 322934 267016 322940 267028
rect 317840 266988 322940 267016
rect 317840 266976 317846 266988
rect 322934 266976 322940 266988
rect 322992 266976 322998 267028
rect 393130 266976 393136 267028
rect 393188 267016 393194 267028
rect 420178 267016 420184 267028
rect 393188 266988 420184 267016
rect 393188 266976 393194 266988
rect 420178 266976 420184 266988
rect 420236 266976 420242 267028
rect 434346 266976 434352 267028
rect 434404 267016 434410 267028
rect 457438 267016 457444 267028
rect 434404 266988 457444 267016
rect 434404 266976 434410 266988
rect 457438 266976 457444 266988
rect 457496 266976 457502 267028
rect 469306 266976 469312 267028
rect 469364 267016 469370 267028
rect 470410 267016 470416 267028
rect 469364 266988 470416 267016
rect 469364 266976 469370 266988
rect 470410 266976 470416 266988
rect 470468 266976 470474 267028
rect 470594 266976 470600 267028
rect 470652 267016 470658 267028
rect 534718 267016 534724 267028
rect 470652 266988 534724 267016
rect 470652 266976 470658 266988
rect 534718 266976 534724 266988
rect 534776 266976 534782 267028
rect 535546 266976 535552 267028
rect 535604 267016 535610 267028
rect 536742 267016 536748 267028
rect 535604 266988 536748 267016
rect 535604 266976 535610 266988
rect 536742 266976 536748 266988
rect 536800 266976 536806 267028
rect 539686 266976 539692 267028
rect 539744 267016 539750 267028
rect 634078 267016 634084 267028
rect 539744 266988 634084 267016
rect 539744 266976 539750 266988
rect 634078 266976 634084 266988
rect 634136 266976 634142 267028
rect 119338 266840 119344 266892
rect 119396 266880 119402 266892
rect 153838 266880 153844 266892
rect 119396 266852 153844 266880
rect 119396 266840 119402 266852
rect 153838 266840 153844 266852
rect 153896 266840 153902 266892
rect 169018 266840 169024 266892
rect 169076 266880 169082 266892
rect 199378 266880 199384 266892
rect 169076 266852 199384 266880
rect 169076 266840 169082 266852
rect 199378 266840 199384 266852
rect 199436 266840 199442 266892
rect 216122 266840 216128 266892
rect 216180 266880 216186 266892
rect 222562 266880 222568 266892
rect 216180 266852 222568 266880
rect 216180 266840 216186 266852
rect 222562 266840 222568 266852
rect 222620 266840 222626 266892
rect 314470 266840 314476 266892
rect 314528 266880 314534 266892
rect 319254 266880 319260 266892
rect 314528 266852 319260 266880
rect 314528 266840 314534 266852
rect 319254 266840 319260 266852
rect 319312 266840 319318 266892
rect 332686 266840 332692 266892
rect 332744 266880 332750 266892
rect 343818 266880 343824 266892
rect 332744 266852 343824 266880
rect 332744 266840 332750 266852
rect 343818 266840 343824 266852
rect 343876 266840 343882 266892
rect 362494 266840 362500 266892
rect 362552 266880 362558 266892
rect 368934 266880 368940 266892
rect 362552 266852 368940 266880
rect 362552 266840 362558 266852
rect 368934 266840 368940 266852
rect 368992 266840 368998 266892
rect 390646 266840 390652 266892
rect 390704 266880 390710 266892
rect 408310 266880 408316 266892
rect 390704 266852 408316 266880
rect 390704 266840 390710 266852
rect 408310 266840 408316 266852
rect 408368 266840 408374 266892
rect 422938 266840 422944 266892
rect 422996 266880 423002 266892
rect 438118 266880 438124 266892
rect 422996 266852 438124 266880
rect 422996 266840 423002 266852
rect 438118 266840 438124 266852
rect 438176 266840 438182 266892
rect 442718 266840 442724 266892
rect 442776 266880 442782 266892
rect 442776 266852 480254 266880
rect 442776 266840 442782 266852
rect 137462 266704 137468 266756
rect 137520 266744 137526 266756
rect 150526 266744 150532 266756
rect 137520 266716 150532 266744
rect 137520 266704 137526 266716
rect 150526 266704 150532 266716
rect 150584 266704 150590 266756
rect 151078 266704 151084 266756
rect 151136 266744 151142 266756
rect 179506 266744 179512 266756
rect 151136 266716 179512 266744
rect 151136 266704 151142 266716
rect 179506 266704 179512 266716
rect 179564 266704 179570 266756
rect 347498 266704 347504 266756
rect 347556 266744 347562 266756
rect 351178 266744 351184 266756
rect 347556 266716 351184 266744
rect 347556 266704 347562 266716
rect 351178 266704 351184 266716
rect 351236 266704 351242 266756
rect 360010 266704 360016 266756
rect 360068 266744 360074 266756
rect 366358 266744 366364 266756
rect 360068 266716 366364 266744
rect 360068 266704 360074 266716
rect 366358 266704 366364 266716
rect 366416 266704 366422 266756
rect 388162 266704 388168 266756
rect 388220 266744 388226 266756
rect 404354 266744 404360 266756
rect 388220 266716 404360 266744
rect 388220 266704 388226 266716
rect 404354 266704 404360 266716
rect 404412 266704 404418 266756
rect 407206 266704 407212 266756
rect 407264 266744 407270 266756
rect 414474 266744 414480 266756
rect 407264 266716 414480 266744
rect 407264 266704 407270 266716
rect 414474 266704 414480 266716
rect 414532 266704 414538 266756
rect 434530 266704 434536 266756
rect 434588 266744 434594 266756
rect 449158 266744 449164 266756
rect 434588 266716 449164 266744
rect 434588 266704 434594 266716
rect 449158 266704 449164 266716
rect 449216 266704 449222 266756
rect 457714 266704 457720 266756
rect 457772 266744 457778 266756
rect 476758 266744 476764 266756
rect 457772 266716 476764 266744
rect 457772 266704 457778 266716
rect 476758 266704 476764 266716
rect 476816 266704 476822 266756
rect 308674 266636 308680 266688
rect 308732 266676 308738 266688
rect 310606 266676 310612 266688
rect 308732 266648 310612 266676
rect 308732 266636 308738 266648
rect 310606 266636 310612 266648
rect 310664 266636 310670 266688
rect 316954 266636 316960 266688
rect 317012 266676 317018 266688
rect 321554 266676 321560 266688
rect 317012 266648 321560 266676
rect 317012 266636 317018 266648
rect 321554 266636 321560 266648
rect 321612 266636 321618 266688
rect 427906 266636 427912 266688
rect 427964 266676 427970 266688
rect 434346 266676 434352 266688
rect 427964 266648 434352 266676
rect 427964 266636 427970 266648
rect 434346 266636 434352 266648
rect 434404 266636 434410 266688
rect 132494 266568 132500 266620
rect 132552 266608 132558 266620
rect 147214 266608 147220 266620
rect 132552 266580 147220 266608
rect 132552 266568 132558 266580
rect 147214 266568 147220 266580
rect 147272 266568 147278 266620
rect 149974 266568 149980 266620
rect 150032 266608 150038 266620
rect 159634 266608 159640 266620
rect 150032 266580 159640 266608
rect 150032 266568 150038 266580
rect 159634 266568 159640 266580
rect 159692 266568 159698 266620
rect 345106 266568 345112 266620
rect 345164 266608 345170 266620
rect 348418 266608 348424 266620
rect 345164 266580 348424 266608
rect 345164 266568 345170 266580
rect 348418 266568 348424 266580
rect 348476 266568 348482 266620
rect 399754 266568 399760 266620
rect 399812 266608 399818 266620
rect 407758 266608 407764 266620
rect 399812 266580 407764 266608
rect 399812 266568 399818 266580
rect 407758 266568 407764 266580
rect 407816 266568 407822 266620
rect 437842 266568 437848 266620
rect 437900 266608 437906 266620
rect 448422 266608 448428 266620
rect 437900 266580 448428 266608
rect 437900 266568 437906 266580
rect 448422 266568 448428 266580
rect 448480 266568 448486 266620
rect 480226 266608 480254 266852
rect 499942 266840 499948 266892
rect 500000 266880 500006 266892
rect 507854 266880 507860 266892
rect 500000 266852 507860 266880
rect 500000 266840 500006 266852
rect 507854 266840 507860 266852
rect 507912 266840 507918 266892
rect 534718 266840 534724 266892
rect 534776 266880 534782 266892
rect 589918 266880 589924 266892
rect 534776 266852 589924 266880
rect 534776 266840 534782 266852
rect 589918 266840 589924 266852
rect 589976 266840 589982 266892
rect 490006 266704 490012 266756
rect 490064 266744 490070 266756
rect 509694 266744 509700 266756
rect 490064 266716 509700 266744
rect 490064 266704 490070 266716
rect 509694 266704 509700 266716
rect 509752 266704 509758 266756
rect 510706 266704 510712 266756
rect 510764 266744 510770 266756
rect 511626 266744 511632 266756
rect 510764 266716 511632 266744
rect 510764 266704 510770 266716
rect 511626 266704 511632 266716
rect 511684 266704 511690 266756
rect 512362 266704 512368 266756
rect 512420 266744 512426 266756
rect 513190 266744 513196 266756
rect 512420 266716 513196 266744
rect 512420 266704 512426 266716
rect 513190 266704 513196 266716
rect 513248 266704 513254 266756
rect 516502 266704 516508 266756
rect 516560 266744 516566 266756
rect 517422 266744 517428 266756
rect 516560 266716 517428 266744
rect 516560 266704 516566 266716
rect 517422 266704 517428 266716
rect 517480 266704 517486 266756
rect 518986 266704 518992 266756
rect 519044 266744 519050 266756
rect 520090 266744 520096 266756
rect 519044 266716 520096 266744
rect 519044 266704 519050 266716
rect 520090 266704 520096 266716
rect 520148 266704 520154 266756
rect 527266 266704 527272 266756
rect 527324 266744 527330 266756
rect 528186 266744 528192 266756
rect 527324 266716 528192 266744
rect 527324 266704 527330 266716
rect 528186 266704 528192 266716
rect 528244 266704 528250 266756
rect 528922 266704 528928 266756
rect 528980 266744 528986 266756
rect 529842 266744 529848 266756
rect 528980 266716 529848 266744
rect 528980 266704 528986 266716
rect 529842 266704 529848 266716
rect 529900 266704 529906 266756
rect 531406 266704 531412 266756
rect 531464 266744 531470 266756
rect 532602 266744 532608 266756
rect 531464 266716 532608 266744
rect 531464 266704 531470 266716
rect 532602 266704 532608 266716
rect 532660 266704 532666 266756
rect 533062 266704 533068 266756
rect 533120 266744 533126 266756
rect 533982 266744 533988 266756
rect 533120 266716 533988 266744
rect 533120 266704 533126 266716
rect 533982 266704 533988 266716
rect 534040 266704 534046 266756
rect 542998 266704 543004 266756
rect 543056 266744 543062 266756
rect 598198 266744 598204 266756
rect 543056 266716 598204 266744
rect 543056 266704 543062 266716
rect 598198 266704 598204 266716
rect 598256 266704 598262 266756
rect 482278 266608 482284 266620
rect 480226 266580 482284 266608
rect 482278 266568 482284 266580
rect 482336 266568 482342 266620
rect 482554 266568 482560 266620
rect 482612 266608 482618 266620
rect 485038 266608 485044 266620
rect 482612 266580 485044 266608
rect 482612 266568 482618 266580
rect 485038 266568 485044 266580
rect 485096 266568 485102 266620
rect 504818 266568 504824 266620
rect 504876 266608 504882 266620
rect 556798 266608 556804 266620
rect 504876 266580 556804 266608
rect 504876 266568 504882 266580
rect 556798 266568 556804 266580
rect 556856 266568 556862 266620
rect 310330 266500 310336 266552
rect 310388 266540 310394 266552
rect 311894 266540 311900 266552
rect 310388 266512 311900 266540
rect 310388 266500 310394 266512
rect 311894 266500 311900 266512
rect 311952 266500 311958 266552
rect 312354 266500 312360 266552
rect 312412 266540 312418 266552
rect 314654 266540 314660 266552
rect 312412 266512 314660 266540
rect 312412 266500 312418 266512
rect 314654 266500 314660 266512
rect 314712 266500 314718 266552
rect 316126 266500 316132 266552
rect 316184 266540 316190 266552
rect 320174 266540 320180 266552
rect 316184 266512 320180 266540
rect 316184 266500 316190 266512
rect 320174 266500 320180 266512
rect 320232 266500 320238 266552
rect 327718 266500 327724 266552
rect 327776 266540 327782 266552
rect 331950 266540 331956 266552
rect 327776 266512 331956 266540
rect 327776 266500 327782 266512
rect 331950 266500 331956 266512
rect 332008 266500 332014 266552
rect 350074 266500 350080 266552
rect 350132 266540 350138 266552
rect 353938 266540 353944 266552
rect 350132 266512 353944 266540
rect 350132 266500 350138 266512
rect 353938 266500 353944 266512
rect 353996 266500 354002 266552
rect 355870 266500 355876 266552
rect 355928 266540 355934 266552
rect 360838 266540 360844 266552
rect 355928 266512 360844 266540
rect 355928 266500 355934 266512
rect 360838 266500 360844 266512
rect 360896 266500 360902 266552
rect 369946 266500 369952 266552
rect 370004 266540 370010 266552
rect 372246 266540 372252 266552
rect 370004 266512 372252 266540
rect 370004 266500 370010 266512
rect 372246 266500 372252 266512
rect 372304 266500 372310 266552
rect 374914 266500 374920 266552
rect 374972 266540 374978 266552
rect 380526 266540 380532 266552
rect 374972 266512 380532 266540
rect 374972 266500 374978 266512
rect 380526 266500 380532 266512
rect 380584 266500 380590 266552
rect 423766 266500 423772 266552
rect 423824 266540 423830 266552
rect 425698 266540 425704 266552
rect 423824 266512 425704 266540
rect 423824 266500 423830 266512
rect 425698 266500 425704 266512
rect 425756 266500 425762 266552
rect 426250 266500 426256 266552
rect 426308 266540 426314 266552
rect 428458 266540 428464 266552
rect 426308 266512 428464 266540
rect 426308 266500 426314 266512
rect 428458 266500 428464 266512
rect 428516 266500 428522 266552
rect 452746 266500 452752 266552
rect 452804 266540 452810 266552
rect 462958 266540 462964 266552
rect 452804 266512 462964 266540
rect 452804 266500 452810 266512
rect 462958 266500 462964 266512
rect 463016 266500 463022 266552
rect 475102 266500 475108 266552
rect 475160 266540 475166 266552
rect 479518 266540 479524 266552
rect 475160 266512 479524 266540
rect 475160 266500 475166 266512
rect 479518 266500 479524 266512
rect 479576 266500 479582 266552
rect 342622 266432 342628 266484
rect 342680 266472 342686 266484
rect 345290 266472 345296 266484
rect 342680 266444 345296 266472
rect 342680 266432 342686 266444
rect 345290 266432 345296 266444
rect 345348 266432 345354 266484
rect 403618 266472 403624 266484
rect 400232 266444 403624 266472
rect 163498 266364 163504 266416
rect 163556 266404 163562 266416
rect 167086 266404 167092 266416
rect 163556 266376 167092 266404
rect 163556 266364 163562 266376
rect 167086 266364 167092 266376
rect 167144 266364 167150 266416
rect 211154 266364 211160 266416
rect 211212 266404 211218 266416
rect 213454 266404 213460 266416
rect 211212 266376 213460 266404
rect 211212 266364 211218 266376
rect 213454 266364 213460 266376
rect 213512 266364 213518 266416
rect 214558 266364 214564 266416
rect 214616 266404 214622 266416
rect 215938 266404 215944 266416
rect 214616 266376 215944 266404
rect 214616 266364 214622 266376
rect 215938 266364 215944 266376
rect 215996 266364 216002 266416
rect 239398 266364 239404 266416
rect 239456 266404 239462 266416
rect 241606 266404 241612 266416
rect 239456 266376 241612 266404
rect 239456 266364 239462 266376
rect 241606 266364 241612 266376
rect 241664 266364 241670 266416
rect 243538 266364 243544 266416
rect 243596 266404 243602 266416
rect 246574 266404 246580 266416
rect 243596 266376 246580 266404
rect 243596 266364 243602 266376
rect 246574 266364 246580 266376
rect 246632 266364 246638 266416
rect 250438 266364 250444 266416
rect 250496 266404 250502 266416
rect 256510 266404 256516 266416
rect 250496 266376 256516 266404
rect 250496 266364 250502 266376
rect 256510 266364 256516 266376
rect 256568 266364 256574 266416
rect 300946 266364 300952 266416
rect 301004 266404 301010 266416
rect 302050 266404 302056 266416
rect 301004 266376 302056 266404
rect 301004 266364 301010 266376
rect 302050 266364 302056 266376
rect 302108 266364 302114 266416
rect 303706 266364 303712 266416
rect 303764 266404 303770 266416
rect 304534 266404 304540 266416
rect 303764 266376 304540 266404
rect 303764 266364 303770 266376
rect 304534 266364 304540 266376
rect 304592 266364 304598 266416
rect 307846 266364 307852 266416
rect 307904 266404 307910 266416
rect 309134 266404 309140 266416
rect 307904 266376 309140 266404
rect 307904 266364 307910 266376
rect 309134 266364 309140 266376
rect 309192 266364 309198 266416
rect 309502 266364 309508 266416
rect 309560 266404 309566 266416
rect 310974 266404 310980 266416
rect 309560 266376 310980 266404
rect 309560 266364 309566 266376
rect 310974 266364 310980 266376
rect 311032 266364 311038 266416
rect 311158 266364 311164 266416
rect 311216 266404 311222 266416
rect 313274 266404 313280 266416
rect 311216 266376 313280 266404
rect 311216 266364 311222 266376
rect 313274 266364 313280 266376
rect 313332 266364 313338 266416
rect 320266 266364 320272 266416
rect 320324 266404 320330 266416
rect 321370 266404 321376 266416
rect 320324 266376 321376 266404
rect 320324 266364 320330 266376
rect 321370 266364 321376 266376
rect 321428 266364 321434 266416
rect 324406 266364 324412 266416
rect 324464 266404 324470 266416
rect 325326 266404 325332 266416
rect 324464 266376 325332 266404
rect 324464 266364 324470 266376
rect 325326 266364 325332 266376
rect 325384 266364 325390 266416
rect 328546 266364 328552 266416
rect 328604 266404 328610 266416
rect 329742 266404 329748 266416
rect 328604 266376 329748 266404
rect 328604 266364 328610 266376
rect 329742 266364 329748 266376
rect 329800 266364 329806 266416
rect 336826 266364 336832 266416
rect 336884 266404 336890 266416
rect 337930 266404 337936 266416
rect 336884 266376 337936 266404
rect 336884 266364 336890 266376
rect 337930 266364 337936 266376
rect 337988 266364 337994 266416
rect 346762 266364 346768 266416
rect 346820 266404 346826 266416
rect 347682 266404 347688 266416
rect 346820 266376 347688 266404
rect 346820 266364 346826 266376
rect 347682 266364 347688 266376
rect 347740 266364 347746 266416
rect 349246 266364 349252 266416
rect 349304 266404 349310 266416
rect 350350 266404 350356 266416
rect 349304 266376 350356 266404
rect 349304 266364 349310 266376
rect 350350 266364 350356 266376
rect 350408 266364 350414 266416
rect 357526 266364 357532 266416
rect 357584 266404 357590 266416
rect 359458 266404 359464 266416
rect 357584 266376 359464 266404
rect 357584 266364 357590 266376
rect 359458 266364 359464 266376
rect 359516 266364 359522 266416
rect 361666 266364 361672 266416
rect 361724 266404 361730 266416
rect 362770 266404 362776 266416
rect 361724 266376 362776 266404
rect 361724 266364 361730 266376
rect 362770 266364 362776 266376
rect 362828 266364 362834 266416
rect 369118 266364 369124 266416
rect 369176 266404 369182 266416
rect 370498 266404 370504 266416
rect 369176 266376 370504 266404
rect 369176 266364 369182 266376
rect 370498 266364 370504 266376
rect 370556 266364 370562 266416
rect 374086 266364 374092 266416
rect 374144 266404 374150 266416
rect 375282 266404 375288 266416
rect 374144 266376 375288 266404
rect 374144 266364 374150 266376
rect 375282 266364 375288 266376
rect 375340 266364 375346 266416
rect 379882 266364 379888 266416
rect 379940 266404 379946 266416
rect 383010 266404 383016 266416
rect 379940 266376 383016 266404
rect 379940 266364 379946 266376
rect 383010 266364 383016 266376
rect 383068 266364 383074 266416
rect 384022 266364 384028 266416
rect 384080 266404 384086 266416
rect 384942 266404 384948 266416
rect 384080 266376 384948 266404
rect 384080 266364 384086 266376
rect 384942 266364 384948 266376
rect 385000 266364 385006 266416
rect 386506 266364 386512 266416
rect 386564 266404 386570 266416
rect 387702 266404 387708 266416
rect 386564 266376 387708 266404
rect 386564 266364 386570 266376
rect 387702 266364 387708 266376
rect 387760 266364 387766 266416
rect 392302 266364 392308 266416
rect 392360 266404 392366 266416
rect 393314 266404 393320 266416
rect 392360 266376 393320 266404
rect 392360 266364 392366 266376
rect 393314 266364 393320 266376
rect 393372 266364 393378 266416
rect 394786 266364 394792 266416
rect 394844 266404 394850 266416
rect 394844 266376 398788 266404
rect 394844 266364 394850 266376
rect 398760 266268 398788 266376
rect 398926 266364 398932 266416
rect 398984 266404 398990 266416
rect 400030 266404 400036 266416
rect 398984 266376 400036 266404
rect 398984 266364 398990 266376
rect 400030 266364 400036 266376
rect 400088 266364 400094 266416
rect 400232 266268 400260 266444
rect 403618 266432 403624 266444
rect 403676 266432 403682 266484
rect 483382 266432 483388 266484
rect 483440 266472 483446 266484
rect 484210 266472 484216 266484
rect 483440 266444 484216 266472
rect 483440 266432 483446 266444
rect 484210 266432 484216 266444
rect 484268 266432 484274 266484
rect 485866 266432 485872 266484
rect 485924 266472 485930 266484
rect 486786 266472 486792 266484
rect 485924 266444 486792 266472
rect 485924 266432 485930 266444
rect 486786 266432 486792 266444
rect 486844 266432 486850 266484
rect 491662 266432 491668 266484
rect 491720 266472 491726 266484
rect 492398 266472 492404 266484
rect 491720 266444 492404 266472
rect 491720 266432 491726 266444
rect 492398 266432 492404 266444
rect 492456 266432 492462 266484
rect 494146 266432 494152 266484
rect 494204 266472 494210 266484
rect 495250 266472 495256 266484
rect 494204 266444 495256 266472
rect 494204 266432 494210 266444
rect 495250 266432 495256 266444
rect 495308 266432 495314 266484
rect 502426 266432 502432 266484
rect 502484 266472 502490 266484
rect 503530 266472 503536 266484
rect 502484 266444 503536 266472
rect 502484 266432 502490 266444
rect 503530 266432 503536 266444
rect 503588 266432 503594 266484
rect 504082 266432 504088 266484
rect 504140 266472 504146 266484
rect 505002 266472 505008 266484
rect 504140 266444 505008 266472
rect 504140 266432 504146 266444
rect 505002 266432 505008 266444
rect 505060 266432 505066 266484
rect 506566 266432 506572 266484
rect 506624 266472 506630 266484
rect 507670 266472 507676 266484
rect 506624 266444 507676 266472
rect 506624 266432 506630 266444
rect 507670 266432 507676 266444
rect 507728 266432 507734 266484
rect 507854 266432 507860 266484
rect 507912 266472 507918 266484
rect 551278 266472 551284 266484
rect 507912 266444 551284 266472
rect 507912 266432 507918 266444
rect 551278 266432 551284 266444
rect 551336 266432 551342 266484
rect 408862 266364 408868 266416
rect 408920 266404 408926 266416
rect 409782 266404 409788 266416
rect 408920 266376 409788 266404
rect 408920 266364 408926 266376
rect 409782 266364 409788 266376
rect 409840 266364 409846 266416
rect 411346 266364 411352 266416
rect 411404 266404 411410 266416
rect 412266 266404 412272 266416
rect 411404 266376 412272 266404
rect 411404 266364 411410 266376
rect 412266 266364 412272 266376
rect 412324 266364 412330 266416
rect 415486 266364 415492 266416
rect 415544 266404 415550 266416
rect 416406 266404 416412 266416
rect 415544 266376 416412 266404
rect 415544 266364 415550 266376
rect 416406 266364 416412 266376
rect 416464 266364 416470 266416
rect 417970 266364 417976 266416
rect 418028 266404 418034 266416
rect 418798 266404 418804 266416
rect 418028 266376 418804 266404
rect 418028 266364 418034 266376
rect 418798 266364 418804 266376
rect 418856 266364 418862 266416
rect 425422 266364 425428 266416
rect 425480 266404 425486 266416
rect 427078 266404 427084 266416
rect 425480 266376 427084 266404
rect 425480 266364 425486 266376
rect 427078 266364 427084 266376
rect 427136 266364 427142 266416
rect 429562 266364 429568 266416
rect 429620 266404 429626 266416
rect 430390 266404 430396 266416
rect 429620 266376 430396 266404
rect 429620 266364 429626 266376
rect 430390 266364 430396 266376
rect 430448 266364 430454 266416
rect 432046 266364 432052 266416
rect 432104 266404 432110 266416
rect 433150 266404 433156 266416
rect 432104 266376 433156 266404
rect 432104 266364 432110 266376
rect 433150 266364 433156 266376
rect 433208 266364 433214 266416
rect 440326 266364 440332 266416
rect 440384 266404 440390 266416
rect 441338 266404 441344 266416
rect 440384 266376 441344 266404
rect 440384 266364 440390 266376
rect 441338 266364 441344 266376
rect 441396 266364 441402 266416
rect 441982 266364 441988 266416
rect 442040 266404 442046 266416
rect 442902 266404 442908 266416
rect 442040 266376 442908 266404
rect 442040 266364 442046 266376
rect 442902 266364 442908 266376
rect 442960 266364 442966 266416
rect 444466 266364 444472 266416
rect 444524 266404 444530 266416
rect 445662 266404 445668 266416
rect 444524 266376 445668 266404
rect 444524 266364 444530 266376
rect 445662 266364 445668 266376
rect 445720 266364 445726 266416
rect 448606 266364 448612 266416
rect 448664 266404 448670 266416
rect 450538 266404 450544 266416
rect 448664 266376 450544 266404
rect 448664 266364 448670 266376
rect 450538 266364 450544 266376
rect 450596 266364 450602 266416
rect 454402 266364 454408 266416
rect 454460 266404 454466 266416
rect 455322 266404 455328 266416
rect 454460 266376 455328 266404
rect 454460 266364 454466 266376
rect 455322 266364 455328 266376
rect 455380 266364 455386 266416
rect 473446 266364 473452 266416
rect 473504 266404 473510 266416
rect 474642 266404 474648 266416
rect 473504 266376 474648 266404
rect 473504 266364 473510 266376
rect 474642 266364 474648 266376
rect 474700 266364 474706 266416
rect 477586 266364 477592 266416
rect 477644 266404 477650 266416
rect 478506 266404 478512 266416
rect 477644 266376 478512 266404
rect 477644 266364 477650 266376
rect 478506 266364 478512 266376
rect 478564 266364 478570 266416
rect 480070 266296 480076 266348
rect 480128 266336 480134 266348
rect 554774 266336 554780 266348
rect 480128 266308 554780 266336
rect 480128 266296 480134 266308
rect 554774 266296 554780 266308
rect 554832 266296 554838 266348
rect 398760 266240 400260 266268
rect 487522 266160 487528 266212
rect 487580 266200 487586 266212
rect 565814 266200 565820 266212
rect 487580 266172 565820 266200
rect 487580 266160 487586 266172
rect 565814 266160 565820 266172
rect 565872 266160 565878 266212
rect 511534 266024 511540 266076
rect 511592 266064 511598 266076
rect 599118 266064 599124 266076
rect 511592 266036 599124 266064
rect 511592 266024 511598 266036
rect 599118 266024 599124 266036
rect 599176 266024 599182 266076
rect 513190 265888 513196 265940
rect 513248 265928 513254 265940
rect 601694 265928 601700 265940
rect 513248 265900 601700 265928
rect 513248 265888 513254 265900
rect 601694 265888 601700 265900
rect 601752 265888 601758 265940
rect 515674 265752 515680 265804
rect 515732 265792 515738 265804
rect 605834 265792 605840 265804
rect 515732 265764 605840 265792
rect 515732 265752 515738 265764
rect 605834 265752 605840 265764
rect 605892 265752 605898 265804
rect 189074 265616 189080 265668
rect 189132 265656 189138 265668
rect 189902 265656 189908 265668
rect 189132 265628 189908 265656
rect 189132 265616 189138 265628
rect 189902 265616 189908 265628
rect 189960 265616 189966 265668
rect 209774 265616 209780 265668
rect 209832 265656 209838 265668
rect 210694 265656 210700 265668
rect 209832 265628 210700 265656
rect 209832 265616 209838 265628
rect 210694 265616 210700 265628
rect 210752 265616 210758 265668
rect 224954 265616 224960 265668
rect 225012 265656 225018 265668
rect 225598 265656 225604 265668
rect 225012 265628 225604 265656
rect 225012 265616 225018 265628
rect 225598 265616 225604 265628
rect 225656 265616 225662 265668
rect 280338 265616 280344 265668
rect 280396 265656 280402 265668
rect 280982 265656 280988 265668
rect 280396 265628 280988 265656
rect 280396 265616 280402 265628
rect 280982 265616 280988 265628
rect 281040 265616 281046 265668
rect 292666 265616 292672 265668
rect 292724 265656 292730 265668
rect 293494 265656 293500 265668
rect 292724 265628 293500 265656
rect 292724 265616 292730 265628
rect 293494 265616 293500 265628
rect 293552 265616 293558 265668
rect 296806 265616 296812 265668
rect 296864 265656 296870 265668
rect 297542 265656 297548 265668
rect 296864 265628 297548 265656
rect 296864 265616 296870 265628
rect 297542 265616 297548 265628
rect 297600 265616 297606 265668
rect 518158 265616 518164 265668
rect 518216 265656 518222 265668
rect 608594 265656 608600 265668
rect 518216 265628 608600 265656
rect 518216 265616 518222 265628
rect 608594 265616 608600 265628
rect 608652 265616 608658 265668
rect 481726 265480 481732 265532
rect 481784 265520 481790 265532
rect 557534 265520 557540 265532
rect 481784 265492 557540 265520
rect 481784 265480 481790 265492
rect 557534 265480 557540 265492
rect 557592 265480 557598 265532
rect 476758 265344 476764 265396
rect 476816 265384 476822 265396
rect 549438 265384 549444 265396
rect 476816 265356 549444 265384
rect 476816 265344 476822 265356
rect 549438 265344 549444 265356
rect 549496 265344 549502 265396
rect 471790 265208 471796 265260
rect 471848 265248 471854 265260
rect 542354 265248 542360 265260
rect 471848 265220 542360 265248
rect 471848 265208 471854 265220
rect 542354 265208 542360 265220
rect 542412 265208 542418 265260
rect 466822 265072 466828 265124
rect 466880 265112 466886 265124
rect 535730 265112 535736 265124
rect 466880 265084 535736 265112
rect 466880 265072 466886 265084
rect 535730 265072 535736 265084
rect 535788 265072 535794 265124
rect 570598 261468 570604 261520
rect 570656 261508 570662 261520
rect 645854 261508 645860 261520
rect 570656 261480 645860 261508
rect 570656 261468 570662 261480
rect 645854 261468 645860 261480
rect 645912 261468 645918 261520
rect 554406 260856 554412 260908
rect 554464 260896 554470 260908
rect 568574 260896 568580 260908
rect 554464 260868 568580 260896
rect 554464 260856 554470 260868
rect 568574 260856 568580 260868
rect 568632 260856 568638 260908
rect 554314 259428 554320 259480
rect 554372 259468 554378 259480
rect 560938 259468 560944 259480
rect 554372 259440 560944 259468
rect 554372 259428 554378 259440
rect 560938 259428 560944 259440
rect 560996 259428 561002 259480
rect 675846 259428 675852 259480
rect 675904 259468 675910 259480
rect 676398 259468 676404 259480
rect 675904 259440 676404 259468
rect 675904 259428 675910 259440
rect 676398 259428 676404 259440
rect 676456 259428 676462 259480
rect 35802 256708 35808 256760
rect 35860 256748 35866 256760
rect 40678 256748 40684 256760
rect 35860 256720 40684 256748
rect 35860 256708 35866 256720
rect 40678 256708 40684 256720
rect 40736 256708 40742 256760
rect 553946 256708 553952 256760
rect 554004 256748 554010 256760
rect 563698 256748 563704 256760
rect 554004 256720 563704 256748
rect 554004 256708 554010 256720
rect 563698 256708 563704 256720
rect 563756 256708 563762 256760
rect 553486 255552 553492 255604
rect 553544 255592 553550 255604
rect 555418 255592 555424 255604
rect 553544 255564 555424 255592
rect 553544 255552 553550 255564
rect 555418 255552 555424 255564
rect 555476 255552 555482 255604
rect 35802 255416 35808 255468
rect 35860 255456 35866 255468
rect 39390 255456 39396 255468
rect 35860 255428 39396 255456
rect 35860 255416 35866 255428
rect 39390 255416 39396 255428
rect 39448 255416 39454 255468
rect 35802 254192 35808 254244
rect 35860 254232 35866 254244
rect 39390 254232 39396 254244
rect 35860 254204 39396 254232
rect 35860 254192 35866 254204
rect 39390 254192 39396 254204
rect 39448 254192 39454 254244
rect 42058 253988 42064 254040
rect 42116 254028 42122 254040
rect 43162 254028 43168 254040
rect 42116 254000 43168 254028
rect 42116 253988 42122 254000
rect 43162 253988 43168 254000
rect 43220 253988 43226 254040
rect 35526 253920 35532 253972
rect 35584 253960 35590 253972
rect 41690 253960 41696 253972
rect 35584 253932 41696 253960
rect 35584 253920 35590 253932
rect 41690 253920 41696 253932
rect 41748 253920 41754 253972
rect 35802 252764 35808 252816
rect 35860 252804 35866 252816
rect 35860 252764 35894 252804
rect 35866 252736 35894 252764
rect 41690 252736 41696 252748
rect 35866 252708 41696 252736
rect 41690 252696 41696 252708
rect 41748 252696 41754 252748
rect 42058 252696 42064 252748
rect 42116 252736 42122 252748
rect 42702 252736 42708 252748
rect 42116 252708 42708 252736
rect 42116 252696 42122 252708
rect 42702 252696 42708 252708
rect 42760 252696 42766 252748
rect 35802 252560 35808 252612
rect 35860 252600 35866 252612
rect 41690 252600 41696 252612
rect 35860 252572 41696 252600
rect 35860 252560 35866 252572
rect 41690 252560 41696 252572
rect 41748 252560 41754 252612
rect 554406 252560 554412 252612
rect 554464 252600 554470 252612
rect 562318 252600 562324 252612
rect 554464 252572 562324 252600
rect 554464 252560 554470 252572
rect 562318 252560 562324 252572
rect 562376 252560 562382 252612
rect 675846 252492 675852 252544
rect 675904 252532 675910 252544
rect 679618 252532 679624 252544
rect 675904 252504 679624 252532
rect 675904 252492 675910 252504
rect 679618 252492 679624 252504
rect 679676 252492 679682 252544
rect 675478 251336 675484 251388
rect 675536 251336 675542 251388
rect 554130 251200 554136 251252
rect 554188 251240 554194 251252
rect 556798 251240 556804 251252
rect 554188 251212 556804 251240
rect 554188 251200 554194 251212
rect 556798 251200 556804 251212
rect 556856 251200 556862 251252
rect 675496 250776 675524 251336
rect 675478 250724 675484 250776
rect 675536 250724 675542 250776
rect 674834 250588 674840 250640
rect 674892 250628 674898 250640
rect 675294 250628 675300 250640
rect 674892 250600 675300 250628
rect 674892 250588 674898 250600
rect 675294 250588 675300 250600
rect 675352 250588 675358 250640
rect 35802 249908 35808 249960
rect 35860 249948 35866 249960
rect 39574 249948 39580 249960
rect 35860 249920 39580 249948
rect 35860 249908 35866 249920
rect 39574 249908 39580 249920
rect 39632 249908 39638 249960
rect 35802 248480 35808 248532
rect 35860 248520 35866 248532
rect 40310 248520 40316 248532
rect 35860 248492 40316 248520
rect 35860 248480 35866 248492
rect 40310 248480 40316 248492
rect 40368 248480 40374 248532
rect 35802 247188 35808 247240
rect 35860 247228 35866 247240
rect 40954 247228 40960 247240
rect 35860 247200 40960 247228
rect 35860 247188 35866 247200
rect 40954 247188 40960 247200
rect 41012 247188 41018 247240
rect 35802 247052 35808 247104
rect 35860 247092 35866 247104
rect 39390 247092 39396 247104
rect 35860 247064 39396 247092
rect 35860 247052 35866 247064
rect 39390 247052 39396 247064
rect 39448 247052 39454 247104
rect 558178 246304 558184 246356
rect 558236 246344 558242 246356
rect 647234 246344 647240 246356
rect 558236 246316 647240 246344
rect 558236 246304 558242 246316
rect 647234 246304 647240 246316
rect 647292 246304 647298 246356
rect 553854 245624 553860 245676
rect 553912 245664 553918 245676
rect 596818 245664 596824 245676
rect 553912 245636 596824 245664
rect 553912 245624 553918 245636
rect 596818 245624 596824 245636
rect 596876 245624 596882 245676
rect 554498 244264 554504 244316
rect 554556 244304 554562 244316
rect 573358 244304 573364 244316
rect 554556 244276 573364 244304
rect 554556 244264 554562 244276
rect 573358 244264 573364 244276
rect 573416 244264 573422 244316
rect 674466 243652 674472 243704
rect 674524 243692 674530 243704
rect 675202 243692 675208 243704
rect 674524 243664 675208 243692
rect 674524 243652 674530 243664
rect 675202 243652 675208 243664
rect 675260 243652 675266 243704
rect 674374 242836 674380 242888
rect 674432 242876 674438 242888
rect 675202 242876 675208 242888
rect 674432 242848 675208 242876
rect 674432 242836 674438 242848
rect 675202 242836 675208 242848
rect 675260 242836 675266 242888
rect 576118 242156 576124 242208
rect 576176 242196 576182 242208
rect 648614 242196 648620 242208
rect 576176 242168 648620 242196
rect 576176 242156 576182 242168
rect 648614 242156 648620 242168
rect 648672 242156 648678 242208
rect 553670 241476 553676 241528
rect 553728 241516 553734 241528
rect 629938 241516 629944 241528
rect 553728 241488 629944 241516
rect 553728 241476 553734 241488
rect 629938 241476 629944 241488
rect 629996 241476 630002 241528
rect 554498 240116 554504 240168
rect 554556 240156 554562 240168
rect 577498 240156 577504 240168
rect 554556 240128 577504 240156
rect 554556 240116 554562 240128
rect 577498 240116 577504 240128
rect 577556 240116 577562 240168
rect 554314 238688 554320 238740
rect 554372 238728 554378 238740
rect 576118 238728 576124 238740
rect 554372 238700 576124 238728
rect 554372 238688 554378 238700
rect 576118 238688 576124 238700
rect 576176 238688 576182 238740
rect 672074 236988 672080 237040
rect 672132 237028 672138 237040
rect 672756 237028 672784 237082
rect 672132 237000 672784 237028
rect 672132 236988 672138 237000
rect 671890 236852 671896 236904
rect 671948 236892 671954 236904
rect 671948 236864 672888 236892
rect 671948 236852 671954 236864
rect 672954 236768 673006 236774
rect 672954 236710 673006 236716
rect 672966 236524 673118 236552
rect 672966 236212 672994 236524
rect 673184 236496 673236 236502
rect 673184 236438 673236 236444
rect 673086 236212 673092 236224
rect 672966 236184 673092 236212
rect 673086 236172 673092 236184
rect 673144 236172 673150 236224
rect 554498 236036 554504 236088
rect 554556 236076 554562 236088
rect 558178 236076 558184 236088
rect 554556 236048 558184 236076
rect 554556 236036 554562 236048
rect 558178 236036 558184 236048
rect 558236 236036 558242 236088
rect 672276 236048 673330 236076
rect 671062 235900 671068 235952
rect 671120 235940 671126 235952
rect 672276 235940 672304 236048
rect 671120 235912 672304 235940
rect 672368 235912 673440 235940
rect 671120 235900 671126 235912
rect 671246 235764 671252 235816
rect 671304 235804 671310 235816
rect 672368 235804 672396 235912
rect 671304 235776 672396 235804
rect 671304 235764 671310 235776
rect 673426 235708 673554 235736
rect 669314 235560 669320 235612
rect 669372 235600 669378 235612
rect 673426 235600 673454 235708
rect 669372 235572 673454 235600
rect 669372 235560 669378 235572
rect 673540 235504 673670 235532
rect 670878 235424 670884 235476
rect 670936 235464 670942 235476
rect 673540 235464 673568 235504
rect 670936 235436 673568 235464
rect 670936 235424 670942 235436
rect 669774 235084 669780 235136
rect 669832 235124 669838 235136
rect 669832 235096 673454 235124
rect 669832 235084 669838 235096
rect 673426 235056 673454 235096
rect 673764 235056 673792 235314
rect 673426 235028 673792 235056
rect 672074 234812 672080 234864
rect 672132 234852 672138 234864
rect 673886 234852 673914 235110
rect 672132 234824 673914 234852
rect 672132 234812 672138 234824
rect 554406 234540 554412 234592
rect 554464 234580 554470 234592
rect 570598 234580 570604 234592
rect 554464 234552 570604 234580
rect 554464 234540 554470 234552
rect 570598 234540 570604 234552
rect 570656 234540 570662 234592
rect 668210 234540 668216 234592
rect 668268 234580 668274 234592
rect 673978 234580 674006 234906
rect 668268 234552 674006 234580
rect 668268 234540 668274 234552
rect 668026 234404 668032 234456
rect 668084 234444 668090 234456
rect 674100 234444 674128 234702
rect 668084 234416 674128 234444
rect 668084 234404 668090 234416
rect 670326 234132 670332 234184
rect 670384 234172 670390 234184
rect 674208 234172 674236 234498
rect 670384 234144 674236 234172
rect 670384 234132 670390 234144
rect 683298 234036 683304 234048
rect 678946 234008 683304 234036
rect 42242 233928 42248 233980
rect 42300 233968 42306 233980
rect 43254 233968 43260 233980
rect 42300 233940 43260 233968
rect 42300 233928 42306 233940
rect 43254 233928 43260 233940
rect 43312 233928 43318 233980
rect 675846 233928 675852 233980
rect 675904 233968 675910 233980
rect 678946 233968 678974 234008
rect 683298 233996 683304 234008
rect 683356 233996 683362 234048
rect 675904 233940 678974 233968
rect 675904 233928 675910 233940
rect 652386 233860 652392 233912
rect 652444 233900 652450 233912
rect 675478 233900 675484 233912
rect 652444 233872 675484 233900
rect 652444 233860 652450 233872
rect 675478 233860 675484 233872
rect 675536 233860 675542 233912
rect 675846 233724 675852 233776
rect 675904 233764 675910 233776
rect 678238 233764 678244 233776
rect 675904 233736 678244 233764
rect 675904 233724 675910 233736
rect 678238 233724 678244 233736
rect 678296 233724 678302 233776
rect 669590 233180 669596 233232
rect 669648 233220 669654 233232
rect 672074 233220 672080 233232
rect 669648 233192 672080 233220
rect 669648 233180 669654 233192
rect 672074 233180 672080 233192
rect 672132 233180 672138 233232
rect 675478 232744 675484 232756
rect 663766 232716 675484 232744
rect 663058 232636 663064 232688
rect 663116 232676 663122 232688
rect 663766 232676 663794 232716
rect 675478 232704 675484 232716
rect 675536 232704 675542 232756
rect 663116 232648 663794 232676
rect 663116 232636 663122 232648
rect 675846 232636 675852 232688
rect 675904 232676 675910 232688
rect 683666 232676 683672 232688
rect 675904 232648 683672 232676
rect 675904 232636 675910 232648
rect 683666 232636 683672 232648
rect 683724 232636 683730 232688
rect 652202 232500 652208 232552
rect 652260 232540 652266 232552
rect 652260 232512 663794 232540
rect 652260 232500 652266 232512
rect 663766 232404 663794 232512
rect 675478 232404 675484 232416
rect 663766 232376 675484 232404
rect 675478 232364 675484 232376
rect 675536 232364 675542 232416
rect 675846 232364 675852 232416
rect 675904 232404 675910 232416
rect 679250 232404 679256 232416
rect 675904 232376 679256 232404
rect 675904 232364 675910 232376
rect 679250 232364 679256 232376
rect 679308 232364 679314 232416
rect 137922 231752 137928 231804
rect 137980 231792 137986 231804
rect 152366 231792 152372 231804
rect 137980 231764 152372 231792
rect 137980 231752 137986 231764
rect 152366 231752 152372 231764
rect 152424 231752 152430 231804
rect 91738 231616 91744 231668
rect 91796 231656 91802 231668
rect 168558 231656 168564 231668
rect 91796 231628 168564 231656
rect 91796 231616 91802 231628
rect 168558 231616 168564 231628
rect 168616 231616 168622 231668
rect 662322 231616 662328 231668
rect 662380 231656 662386 231668
rect 668394 231656 668400 231668
rect 662380 231628 668400 231656
rect 662380 231616 662386 231628
rect 668394 231616 668400 231628
rect 668452 231616 668458 231668
rect 669130 231616 669136 231668
rect 669188 231656 669194 231668
rect 675386 231656 675392 231668
rect 669188 231628 675392 231656
rect 669188 231616 669194 231628
rect 675386 231616 675392 231628
rect 675444 231616 675450 231668
rect 128262 231480 128268 231532
rect 128320 231520 128326 231532
rect 195882 231520 195888 231532
rect 128320 231492 195888 231520
rect 128320 231480 128326 231492
rect 195882 231480 195888 231492
rect 195940 231480 195946 231532
rect 596818 231480 596824 231532
rect 596876 231520 596882 231532
rect 633618 231520 633624 231532
rect 596876 231492 633624 231520
rect 596876 231480 596882 231492
rect 633618 231480 633624 231492
rect 633676 231480 633682 231532
rect 664990 231480 664996 231532
rect 665048 231520 665054 231532
rect 665048 231492 675340 231520
rect 665048 231480 665054 231492
rect 57238 231344 57244 231396
rect 57296 231384 57302 231396
rect 669130 231384 669136 231396
rect 57296 231356 669136 231384
rect 57296 231344 57302 231356
rect 669130 231344 669136 231356
rect 669188 231344 669194 231396
rect 675312 231384 675340 231492
rect 675220 231356 675340 231384
rect 64138 231208 64144 231260
rect 64196 231248 64202 231260
rect 667198 231248 667204 231260
rect 64196 231220 667204 231248
rect 64196 231208 64202 231220
rect 667198 231208 667204 231220
rect 667256 231208 667262 231260
rect 675220 231180 675248 231356
rect 675220 231152 675326 231180
rect 58618 231072 58624 231124
rect 58676 231112 58682 231124
rect 674926 231112 674932 231124
rect 58676 231084 674932 231112
rect 58676 231072 58682 231084
rect 674926 231072 674932 231084
rect 674984 231072 674990 231124
rect 668394 230936 668400 230988
rect 668452 230976 668458 230988
rect 668452 230948 675142 230976
rect 668452 230936 668458 230948
rect 97902 230868 97908 230920
rect 97960 230908 97966 230920
rect 173986 230908 173992 230920
rect 97960 230880 173992 230908
rect 97960 230868 97966 230880
rect 173986 230868 173992 230880
rect 174044 230868 174050 230920
rect 668394 230800 668400 230852
rect 668452 230840 668458 230852
rect 668946 230840 668952 230852
rect 668452 230812 668952 230840
rect 668452 230800 668458 230812
rect 668946 230800 668952 230812
rect 669004 230800 669010 230852
rect 672074 230800 672080 230852
rect 672132 230840 672138 230852
rect 672132 230812 674982 230840
rect 672132 230800 672138 230812
rect 110322 230732 110328 230784
rect 110380 230772 110386 230784
rect 184290 230772 184296 230784
rect 110380 230744 184296 230772
rect 110380 230732 110386 230744
rect 184290 230732 184296 230744
rect 184348 230732 184354 230784
rect 118602 230596 118608 230648
rect 118660 230636 118666 230648
rect 188154 230636 188160 230648
rect 118660 230608 188160 230636
rect 118660 230596 118666 230608
rect 188154 230596 188160 230608
rect 188212 230596 188218 230648
rect 195054 230596 195060 230648
rect 195112 230636 195118 230648
rect 196894 230636 196900 230648
rect 195112 230608 196900 230636
rect 195112 230596 195118 230608
rect 196894 230596 196900 230608
rect 196952 230596 196958 230648
rect 665818 230596 665824 230648
rect 665876 230636 665882 230648
rect 665876 230608 674820 230636
rect 665876 230596 665882 230608
rect 439314 230528 439320 230580
rect 439372 230568 439378 230580
rect 439372 230540 439544 230568
rect 439372 230528 439378 230540
rect 152366 230460 152372 230512
rect 152424 230500 152430 230512
rect 203610 230500 203616 230512
rect 152424 230472 203616 230500
rect 152424 230460 152430 230472
rect 203610 230460 203616 230472
rect 203668 230460 203674 230512
rect 130378 230392 130384 230444
rect 130436 230432 130442 230444
rect 142614 230432 142620 230444
rect 130436 230404 142620 230432
rect 130436 230392 130442 230404
rect 142614 230392 142620 230404
rect 142672 230392 142678 230444
rect 142798 230392 142804 230444
rect 142856 230432 142862 230444
rect 150802 230432 150808 230444
rect 142856 230404 150808 230432
rect 142856 230392 142862 230404
rect 150802 230392 150808 230404
rect 150860 230392 150866 230444
rect 206278 230392 206284 230444
rect 206336 230432 206342 230444
rect 256418 230432 256424 230444
rect 206336 230404 256424 230432
rect 206336 230392 206342 230404
rect 256418 230392 256424 230404
rect 256476 230392 256482 230444
rect 276290 230392 276296 230444
rect 276348 230432 276354 230444
rect 292482 230432 292488 230444
rect 276348 230404 292488 230432
rect 276348 230392 276354 230404
rect 292482 230392 292488 230404
rect 292540 230392 292546 230444
rect 308398 230392 308404 230444
rect 308456 230432 308462 230444
rect 334986 230432 334992 230444
rect 308456 230404 334992 230432
rect 308456 230392 308462 230404
rect 334986 230392 334992 230404
rect 335044 230392 335050 230444
rect 439516 230432 439544 230540
rect 440694 230432 440700 230444
rect 439516 230404 440700 230432
rect 440694 230392 440700 230404
rect 440752 230392 440758 230444
rect 441890 230392 441896 230444
rect 441948 230432 441954 230444
rect 443454 230432 443460 230444
rect 441948 230404 443460 230432
rect 441948 230392 441954 230404
rect 443454 230392 443460 230404
rect 443512 230392 443518 230444
rect 526898 230392 526904 230444
rect 526956 230432 526962 230444
rect 536098 230432 536104 230444
rect 526956 230404 536104 230432
rect 526956 230392 526962 230404
rect 536098 230392 536104 230404
rect 536156 230392 536162 230444
rect 673454 230392 673460 230444
rect 673512 230432 673518 230444
rect 673512 230404 674702 230432
rect 673512 230392 673518 230404
rect 42150 230324 42156 230376
rect 42208 230364 42214 230376
rect 43070 230364 43076 230376
rect 42208 230336 43076 230364
rect 42208 230324 42214 230336
rect 43070 230324 43076 230336
rect 43128 230324 43134 230376
rect 387426 230324 387432 230376
rect 387484 230364 387490 230376
rect 388438 230364 388444 230376
rect 387484 230336 388444 230364
rect 387484 230324 387490 230336
rect 388438 230324 388444 230336
rect 388496 230324 388502 230376
rect 398098 230324 398104 230376
rect 398156 230364 398162 230376
rect 399386 230364 399392 230376
rect 398156 230336 399392 230364
rect 398156 230324 398162 230336
rect 399386 230324 399392 230336
rect 399444 230324 399450 230376
rect 438670 230324 438676 230376
rect 438728 230364 438734 230376
rect 439314 230364 439320 230376
rect 438728 230336 439320 230364
rect 438728 230324 438734 230336
rect 439314 230324 439320 230336
rect 439372 230324 439378 230376
rect 443822 230324 443828 230376
rect 443880 230364 443886 230376
rect 444834 230364 444840 230376
rect 443880 230336 444840 230364
rect 443880 230324 443886 230336
rect 444834 230324 444840 230336
rect 444892 230324 444898 230376
rect 449618 230324 449624 230376
rect 449676 230364 449682 230376
rect 450538 230364 450544 230376
rect 449676 230336 450544 230364
rect 449676 230324 449682 230336
rect 450538 230324 450544 230336
rect 450596 230324 450602 230376
rect 452838 230324 452844 230376
rect 452896 230364 452902 230376
rect 454310 230364 454316 230376
rect 452896 230336 454316 230364
rect 452896 230324 452902 230336
rect 454310 230324 454316 230336
rect 454368 230324 454374 230376
rect 455414 230324 455420 230376
rect 455472 230364 455478 230376
rect 457162 230364 457168 230376
rect 455472 230336 457168 230364
rect 455472 230324 455478 230336
rect 457162 230324 457168 230336
rect 457220 230324 457226 230376
rect 463786 230324 463792 230376
rect 463844 230364 463850 230376
rect 465718 230364 465724 230376
rect 463844 230336 465724 230364
rect 463844 230324 463850 230336
rect 465718 230324 465724 230336
rect 465776 230324 465782 230376
rect 470870 230324 470876 230376
rect 470928 230364 470934 230376
rect 471882 230364 471888 230376
rect 470928 230336 471888 230364
rect 470928 230324 470934 230336
rect 471882 230324 471888 230336
rect 471940 230324 471946 230376
rect 472158 230324 472164 230376
rect 472216 230364 472222 230376
rect 473170 230364 473176 230376
rect 472216 230336 473176 230364
rect 472216 230324 472222 230336
rect 473170 230324 473176 230336
rect 473228 230324 473234 230376
rect 487614 230324 487620 230376
rect 487672 230364 487678 230376
rect 488442 230364 488448 230376
rect 487672 230336 488448 230364
rect 487672 230324 487678 230336
rect 488442 230324 488448 230336
rect 488500 230324 488506 230376
rect 493410 230324 493416 230376
rect 493468 230364 493474 230376
rect 496354 230364 496360 230376
rect 493468 230336 496360 230364
rect 493468 230324 493474 230336
rect 496354 230324 496360 230336
rect 496412 230324 496418 230376
rect 497274 230324 497280 230376
rect 497332 230364 497338 230376
rect 498102 230364 498108 230376
rect 497332 230336 498108 230364
rect 497332 230324 497338 230336
rect 498102 230324 498108 230336
rect 498160 230324 498166 230376
rect 510798 230324 510804 230376
rect 510856 230364 510862 230376
rect 511902 230364 511908 230376
rect 510856 230336 511908 230364
rect 510856 230324 510862 230336
rect 511902 230324 511908 230336
rect 511960 230324 511966 230376
rect 133782 230256 133788 230308
rect 133840 230296 133846 230308
rect 202322 230296 202328 230308
rect 133840 230268 202328 230296
rect 133840 230256 133846 230268
rect 202322 230256 202328 230268
rect 202380 230256 202386 230308
rect 210418 230256 210424 230308
rect 210476 230296 210482 230308
rect 261570 230296 261576 230308
rect 210476 230268 261576 230296
rect 210476 230256 210482 230268
rect 261570 230256 261576 230268
rect 261628 230256 261634 230308
rect 275646 230256 275652 230308
rect 275704 230296 275710 230308
rect 313090 230296 313096 230308
rect 275704 230268 313096 230296
rect 275704 230256 275710 230268
rect 313090 230256 313096 230268
rect 313148 230256 313154 230308
rect 436094 230256 436100 230308
rect 436152 230296 436158 230308
rect 436830 230296 436836 230308
rect 436152 230268 436836 230296
rect 436152 230256 436158 230268
rect 436830 230256 436836 230268
rect 436888 230256 436894 230308
rect 528830 230256 528836 230308
rect 528888 230296 528894 230308
rect 539594 230296 539600 230308
rect 528888 230268 539600 230296
rect 528888 230256 528894 230268
rect 539594 230256 539600 230268
rect 539652 230256 539658 230308
rect 388438 230188 388444 230240
rect 388496 230228 388502 230240
rect 391658 230228 391664 230240
rect 388496 230200 391664 230228
rect 388496 230188 388502 230200
rect 391658 230188 391664 230200
rect 391716 230188 391722 230240
rect 444466 230188 444472 230240
rect 444524 230228 444530 230240
rect 447594 230228 447600 230240
rect 444524 230200 447600 230228
rect 444524 230188 444530 230200
rect 447594 230188 447600 230200
rect 447652 230188 447658 230240
rect 451550 230188 451556 230240
rect 451608 230228 451614 230240
rect 453298 230228 453304 230240
rect 451608 230200 453304 230228
rect 451608 230188 451614 230200
rect 453298 230188 453304 230200
rect 453356 230188 453362 230240
rect 453482 230188 453488 230240
rect 453540 230228 453546 230240
rect 455782 230228 455788 230240
rect 453540 230200 455788 230228
rect 453540 230188 453546 230200
rect 455782 230188 455788 230200
rect 455840 230188 455846 230240
rect 468294 230188 468300 230240
rect 468352 230228 468358 230240
rect 469122 230228 469128 230240
rect 468352 230200 469128 230228
rect 468352 230188 468358 230200
rect 469122 230188 469128 230200
rect 469180 230188 469186 230240
rect 490190 230188 490196 230240
rect 490248 230228 490254 230240
rect 493778 230228 493784 230240
rect 490248 230200 493784 230228
rect 490248 230188 490254 230200
rect 493778 230188 493784 230200
rect 493836 230188 493842 230240
rect 511442 230188 511448 230240
rect 511500 230228 511506 230240
rect 517514 230228 517520 230240
rect 511500 230200 517520 230228
rect 511500 230188 511506 230200
rect 517514 230188 517520 230200
rect 517572 230188 517578 230240
rect 674282 230188 674288 230240
rect 674340 230228 674346 230240
rect 674340 230200 674590 230228
rect 674340 230188 674346 230200
rect 95234 230120 95240 230172
rect 95292 230160 95298 230172
rect 157288 230160 157294 230172
rect 95292 230132 157294 230160
rect 95292 230120 95298 230132
rect 157288 230120 157294 230132
rect 157346 230120 157352 230172
rect 157426 230120 157432 230172
rect 157484 230160 157490 230172
rect 161106 230160 161112 230172
rect 157484 230132 161112 230160
rect 157484 230120 157490 230132
rect 161106 230120 161112 230132
rect 161164 230120 161170 230172
rect 176746 230120 176752 230172
rect 176804 230160 176810 230172
rect 235810 230160 235816 230172
rect 176804 230132 235816 230160
rect 176804 230120 176810 230132
rect 235810 230120 235816 230132
rect 235868 230120 235874 230172
rect 264238 230120 264244 230172
rect 264296 230160 264302 230172
rect 302786 230160 302792 230172
rect 264296 230132 302792 230160
rect 264296 230120 264302 230132
rect 302786 230120 302792 230132
rect 302844 230120 302850 230172
rect 302970 230120 302976 230172
rect 303028 230160 303034 230172
rect 329834 230160 329840 230172
rect 303028 230132 329840 230160
rect 303028 230120 303034 230132
rect 329834 230120 329840 230132
rect 329892 230120 329898 230172
rect 334250 230120 334256 230172
rect 334308 230160 334314 230172
rect 355594 230160 355600 230172
rect 334308 230132 355600 230160
rect 334308 230120 334314 230132
rect 355594 230120 355600 230132
rect 355652 230120 355658 230172
rect 521102 230120 521108 230172
rect 521160 230160 521166 230172
rect 529198 230160 529204 230172
rect 521160 230132 529204 230160
rect 521160 230120 521166 230132
rect 529198 230120 529204 230132
rect 529256 230120 529262 230172
rect 532694 230120 532700 230172
rect 532752 230160 532758 230172
rect 547138 230160 547144 230172
rect 532752 230132 547144 230160
rect 532752 230120 532758 230132
rect 547138 230120 547144 230132
rect 547196 230120 547202 230172
rect 454126 230052 454132 230104
rect 454184 230092 454190 230104
rect 455322 230092 455328 230104
rect 454184 230064 455328 230092
rect 454184 230052 454190 230064
rect 455322 230052 455328 230064
rect 455380 230052 455386 230104
rect 491478 230052 491484 230104
rect 491536 230092 491542 230104
rect 492490 230092 492496 230104
rect 491536 230064 492496 230092
rect 491536 230052 491542 230064
rect 492490 230052 492496 230064
rect 492548 230052 492554 230104
rect 126882 229984 126888 230036
rect 126940 230024 126946 230036
rect 195054 230024 195060 230036
rect 126940 229996 195060 230024
rect 126940 229984 126946 229996
rect 195054 229984 195060 229996
rect 195112 229984 195118 230036
rect 195422 229984 195428 230036
rect 195480 230024 195486 230036
rect 214742 230024 214748 230036
rect 195480 229996 214748 230024
rect 195480 229984 195486 229996
rect 214742 229984 214748 229996
rect 214800 229984 214806 230036
rect 219986 229984 219992 230036
rect 220044 230024 220050 230036
rect 230658 230024 230664 230036
rect 220044 229996 230664 230024
rect 220044 229984 220050 229996
rect 230658 229984 230664 229996
rect 230716 229984 230722 230036
rect 242526 229984 242532 230036
rect 242584 230024 242590 230036
rect 287330 230024 287336 230036
rect 242584 229996 287336 230024
rect 242584 229984 242590 229996
rect 287330 229984 287336 229996
rect 287388 229984 287394 230036
rect 287514 229984 287520 230036
rect 287572 230024 287578 230036
rect 307938 230024 307944 230036
rect 287572 229996 307944 230024
rect 287572 229984 287578 229996
rect 307938 229984 307944 229996
rect 307996 229984 308002 230036
rect 312630 229984 312636 230036
rect 312688 230024 312694 230036
rect 340138 230024 340144 230036
rect 312688 229996 340144 230024
rect 312688 229984 312694 229996
rect 340138 229984 340144 229996
rect 340196 229984 340202 230036
rect 354950 229984 354956 230036
rect 355008 230024 355014 230036
rect 371050 230024 371056 230036
rect 355008 229996 371056 230024
rect 355008 229984 355014 229996
rect 371050 229984 371056 229996
rect 371108 229984 371114 230036
rect 457346 229984 457352 230036
rect 457404 230024 457410 230036
rect 463878 230024 463884 230036
rect 457404 229996 463884 230024
rect 457404 229984 457410 229996
rect 463878 229984 463884 229996
rect 463936 229984 463942 230036
rect 515306 229984 515312 230036
rect 515364 230024 515370 230036
rect 524598 230024 524604 230036
rect 515364 229996 524604 230024
rect 515364 229984 515370 229996
rect 524598 229984 524604 229996
rect 524656 229984 524662 230036
rect 534626 229984 534632 230036
rect 534684 230024 534690 230036
rect 549254 230024 549260 230036
rect 534684 229996 549260 230024
rect 534684 229984 534690 229996
rect 549254 229984 549260 229996
rect 549312 229984 549318 230036
rect 674098 229984 674104 230036
rect 674156 229984 674162 230036
rect 86218 229848 86224 229900
rect 86276 229888 86282 229900
rect 156690 229888 156696 229900
rect 86276 229860 156696 229888
rect 86276 229848 86282 229860
rect 156690 229848 156696 229860
rect 156748 229848 156754 229900
rect 158530 229888 158536 229900
rect 157168 229860 158536 229888
rect 68278 229712 68284 229764
rect 68336 229752 68342 229764
rect 142798 229752 142804 229764
rect 68336 229724 142804 229752
rect 68336 229712 68342 229724
rect 142798 229712 142804 229724
rect 142856 229712 142862 229764
rect 142982 229712 142988 229764
rect 143040 229752 143046 229764
rect 145650 229752 145656 229764
rect 143040 229724 145656 229752
rect 143040 229712 143046 229724
rect 145650 229712 145656 229724
rect 145708 229712 145714 229764
rect 145834 229712 145840 229764
rect 145892 229752 145898 229764
rect 157168 229752 157196 229860
rect 158530 229848 158536 229860
rect 158588 229848 158594 229900
rect 158714 229848 158720 229900
rect 158772 229888 158778 229900
rect 163682 229888 163688 229900
rect 158772 229860 163688 229888
rect 158772 229848 158778 229860
rect 163682 229848 163688 229860
rect 163740 229848 163746 229900
rect 163958 229848 163964 229900
rect 164016 229888 164022 229900
rect 225506 229888 225512 229900
rect 164016 229860 225512 229888
rect 164016 229848 164022 229860
rect 225506 229848 225512 229860
rect 225564 229848 225570 229900
rect 230474 229848 230480 229900
rect 230532 229888 230538 229900
rect 277026 229888 277032 229900
rect 230532 229860 277032 229888
rect 230532 229848 230538 229860
rect 277026 229848 277032 229860
rect 277084 229848 277090 229900
rect 282546 229848 282552 229900
rect 282604 229888 282610 229900
rect 318242 229888 318248 229900
rect 282604 229860 318248 229888
rect 282604 229848 282610 229860
rect 318242 229848 318248 229860
rect 318300 229848 318306 229900
rect 324222 229848 324228 229900
rect 324280 229888 324286 229900
rect 350442 229888 350448 229900
rect 324280 229860 350448 229888
rect 324280 229848 324286 229860
rect 350442 229848 350448 229860
rect 350500 229848 350506 229900
rect 366726 229848 366732 229900
rect 366784 229888 366790 229900
rect 383930 229888 383936 229900
rect 366784 229860 383936 229888
rect 366784 229848 366790 229860
rect 383930 229848 383936 229860
rect 383988 229848 383994 229900
rect 467006 229848 467012 229900
rect 467064 229888 467070 229900
rect 473998 229888 474004 229900
rect 467064 229860 474004 229888
rect 467064 229848 467070 229860
rect 473998 229848 474004 229860
rect 474056 229848 474062 229900
rect 476666 229848 476672 229900
rect 476724 229888 476730 229900
rect 481634 229888 481640 229900
rect 476724 229860 481640 229888
rect 476724 229848 476730 229860
rect 481634 229848 481640 229860
rect 481692 229848 481698 229900
rect 481818 229848 481824 229900
rect 481876 229888 481882 229900
rect 489914 229888 489920 229900
rect 481876 229860 489920 229888
rect 481876 229848 481882 229860
rect 489914 229848 489920 229860
rect 489972 229848 489978 229900
rect 495986 229848 495992 229900
rect 496044 229888 496050 229900
rect 507118 229888 507124 229900
rect 496044 229860 507124 229888
rect 496044 229848 496050 229860
rect 507118 229848 507124 229860
rect 507176 229848 507182 229900
rect 509510 229848 509516 229900
rect 509568 229888 509574 229900
rect 515398 229888 515404 229900
rect 509568 229860 515404 229888
rect 509568 229848 509574 229860
rect 515398 229848 515404 229860
rect 515456 229848 515462 229900
rect 517238 229848 517244 229900
rect 517296 229888 517302 229900
rect 526438 229888 526444 229900
rect 517296 229860 526444 229888
rect 517296 229848 517302 229860
rect 526438 229848 526444 229860
rect 526496 229848 526502 229900
rect 536558 229848 536564 229900
rect 536616 229888 536622 229900
rect 559558 229888 559564 229900
rect 536616 229860 559564 229888
rect 536616 229848 536622 229860
rect 559558 229848 559564 229860
rect 559616 229848 559622 229900
rect 433518 229780 433524 229832
rect 433576 229820 433582 229832
rect 434162 229820 434168 229832
rect 433576 229792 434168 229820
rect 433576 229780 433582 229792
rect 434162 229780 434168 229792
rect 434220 229780 434226 229832
rect 145892 229724 157196 229752
rect 145892 229712 145898 229724
rect 157288 229712 157294 229764
rect 157346 229752 157352 229764
rect 166258 229752 166264 229764
rect 157346 229724 166264 229752
rect 157346 229712 157352 229724
rect 166258 229712 166264 229724
rect 166316 229712 166322 229764
rect 171042 229712 171048 229764
rect 171100 229752 171106 229764
rect 219986 229752 219992 229764
rect 171100 229724 219992 229752
rect 171100 229712 171106 229724
rect 219986 229712 219992 229724
rect 220044 229712 220050 229764
rect 246114 229752 246120 229764
rect 224926 229724 246120 229752
rect 82078 229576 82084 229628
rect 82136 229616 82142 229628
rect 82136 229588 147904 229616
rect 82136 229576 82142 229588
rect 102134 229440 102140 229492
rect 102192 229480 102198 229492
rect 139854 229480 139860 229492
rect 102192 229452 139860 229480
rect 102192 229440 102198 229452
rect 139854 229440 139860 229452
rect 139912 229440 139918 229492
rect 147876 229480 147904 229588
rect 149054 229576 149060 229628
rect 149112 229616 149118 229628
rect 153378 229616 153384 229628
rect 149112 229588 153384 229616
rect 149112 229576 149118 229588
rect 153378 229576 153384 229588
rect 153436 229576 153442 229628
rect 153838 229576 153844 229628
rect 153896 229616 153902 229628
rect 157702 229616 157708 229628
rect 153896 229588 157708 229616
rect 153896 229576 153902 229588
rect 157702 229576 157708 229588
rect 157760 229576 157766 229628
rect 157978 229576 157984 229628
rect 158036 229616 158042 229628
rect 158036 229588 214604 229616
rect 158036 229576 158042 229588
rect 149606 229480 149612 229492
rect 140148 229452 147168 229480
rect 147876 229452 149612 229480
rect 140148 229412 140176 229452
rect 140056 229384 140176 229412
rect 111058 229304 111064 229356
rect 111116 229344 111122 229356
rect 140056 229344 140084 229384
rect 111116 229316 140084 229344
rect 111116 229304 111122 229316
rect 140314 229304 140320 229356
rect 140372 229344 140378 229356
rect 142982 229344 142988 229356
rect 140372 229316 142988 229344
rect 140372 229304 140378 229316
rect 142982 229304 142988 229316
rect 143040 229304 143046 229356
rect 144178 229304 144184 229356
rect 144236 229344 144242 229356
rect 146938 229344 146944 229356
rect 144236 229316 146944 229344
rect 144236 229304 144242 229316
rect 146938 229304 146944 229316
rect 146996 229304 147002 229356
rect 147140 229344 147168 229452
rect 149606 229440 149612 229452
rect 149664 229440 149670 229492
rect 149974 229440 149980 229492
rect 150032 229480 150038 229492
rect 210050 229480 210056 229492
rect 150032 229452 210056 229480
rect 150032 229440 150038 229452
rect 210050 229440 210056 229452
rect 210108 229440 210114 229492
rect 214576 229480 214604 229588
rect 214742 229576 214748 229628
rect 214800 229616 214806 229628
rect 224926 229616 224954 229724
rect 246114 229712 246120 229724
rect 246172 229712 246178 229764
rect 256510 229712 256516 229764
rect 256568 229752 256574 229764
rect 297634 229752 297640 229764
rect 256568 229724 297640 229752
rect 256568 229712 256574 229724
rect 297634 229712 297640 229724
rect 297692 229712 297698 229764
rect 318058 229712 318064 229764
rect 318116 229752 318122 229764
rect 318116 229724 335354 229752
rect 318116 229712 318122 229724
rect 266722 229616 266728 229628
rect 214800 229588 224954 229616
rect 229066 229588 266728 229616
rect 214800 229576 214806 229588
rect 220354 229480 220360 229492
rect 214576 229452 220360 229480
rect 220354 229440 220360 229452
rect 220412 229440 220418 229492
rect 220722 229440 220728 229492
rect 220780 229480 220786 229492
rect 229066 229480 229094 229588
rect 266722 229576 266728 229588
rect 266780 229576 266786 229628
rect 296990 229576 296996 229628
rect 297048 229616 297054 229628
rect 323394 229616 323400 229628
rect 297048 229588 323400 229616
rect 297048 229576 297054 229588
rect 323394 229576 323400 229588
rect 323452 229576 323458 229628
rect 335326 229616 335354 229724
rect 345014 229712 345020 229764
rect 345072 229752 345078 229764
rect 360746 229752 360752 229764
rect 345072 229724 360752 229752
rect 345072 229712 345078 229724
rect 360746 229712 360752 229724
rect 360804 229712 360810 229764
rect 361206 229712 361212 229764
rect 361264 229752 361270 229764
rect 378778 229752 378784 229764
rect 361264 229724 378784 229752
rect 361264 229712 361270 229724
rect 378778 229712 378784 229724
rect 378836 229712 378842 229764
rect 391198 229712 391204 229764
rect 391256 229752 391262 229764
rect 398742 229752 398748 229764
rect 391256 229724 398748 229752
rect 391256 229712 391262 229724
rect 398742 229712 398748 229724
rect 398800 229712 398806 229764
rect 399846 229712 399852 229764
rect 399904 229752 399910 229764
rect 409690 229752 409696 229764
rect 399904 229724 409696 229752
rect 399904 229712 399910 229724
rect 409690 229712 409696 229724
rect 409748 229712 409754 229764
rect 410886 229712 410892 229764
rect 410944 229752 410950 229764
rect 417418 229752 417424 229764
rect 410944 229724 417424 229752
rect 410944 229712 410950 229724
rect 417418 229712 417424 229724
rect 417476 229712 417482 229764
rect 465442 229712 465448 229764
rect 465500 229752 465506 229764
rect 467466 229752 467472 229764
rect 465500 229724 467472 229752
rect 465500 229712 465506 229724
rect 467466 229712 467472 229724
rect 467524 229712 467530 229764
rect 469582 229712 469588 229764
rect 469640 229752 469646 229764
rect 476758 229752 476764 229764
rect 469640 229724 476764 229752
rect 469640 229712 469646 229724
rect 476758 229712 476764 229724
rect 476816 229712 476822 229764
rect 479242 229712 479248 229764
rect 479300 229752 479306 229764
rect 488074 229752 488080 229764
rect 479300 229724 488080 229752
rect 479300 229712 479306 229724
rect 488074 229712 488080 229724
rect 488132 229712 488138 229764
rect 492122 229712 492128 229764
rect 492180 229752 492186 229764
rect 505094 229752 505100 229764
rect 492180 229724 505100 229752
rect 492180 229712 492186 229724
rect 505094 229712 505100 229724
rect 505152 229712 505158 229764
rect 507578 229712 507584 229764
rect 507636 229752 507642 229764
rect 516778 229752 516784 229764
rect 507636 229724 516784 229752
rect 507636 229712 507642 229724
rect 516778 229712 516784 229724
rect 516836 229712 516842 229764
rect 523034 229712 523040 229764
rect 523092 229752 523098 229764
rect 534810 229752 534816 229764
rect 523092 229724 534816 229752
rect 523092 229712 523098 229724
rect 534810 229712 534816 229724
rect 534868 229712 534874 229764
rect 538490 229712 538496 229764
rect 538548 229752 538554 229764
rect 566458 229752 566464 229764
rect 538548 229724 566464 229752
rect 538548 229712 538554 229724
rect 566458 229712 566464 229724
rect 566516 229712 566522 229764
rect 660942 229712 660948 229764
rect 661000 229752 661006 229764
rect 672074 229752 672080 229764
rect 661000 229724 672080 229752
rect 661000 229712 661006 229724
rect 672074 229712 672080 229724
rect 672132 229712 672138 229764
rect 674116 229752 674144 229984
rect 674452 229968 674504 229974
rect 674452 229910 674504 229916
rect 674334 229832 674386 229838
rect 674334 229774 674386 229780
rect 673978 229724 674144 229752
rect 345290 229616 345296 229628
rect 335326 229588 345296 229616
rect 345290 229576 345296 229588
rect 345348 229576 345354 229628
rect 530118 229576 530124 229628
rect 530176 229616 530182 229628
rect 531130 229616 531136 229628
rect 530176 229588 531136 229616
rect 530176 229576 530182 229588
rect 531130 229576 531136 229588
rect 531188 229576 531194 229628
rect 538306 229616 538312 229628
rect 538186 229588 538312 229616
rect 384298 229508 384304 229560
rect 384356 229548 384362 229560
rect 389082 229548 389088 229560
rect 384356 229520 389088 229548
rect 384356 229508 384362 229520
rect 389082 229508 389088 229520
rect 389140 229508 389146 229560
rect 448974 229508 448980 229560
rect 449032 229548 449038 229560
rect 451918 229548 451924 229560
rect 449032 229520 451924 229548
rect 449032 229508 449038 229520
rect 451918 229508 451924 229520
rect 451976 229508 451982 229560
rect 220780 229452 229094 229480
rect 220780 229440 220786 229452
rect 231118 229440 231124 229492
rect 231176 229480 231182 229492
rect 271874 229480 271880 229492
rect 231176 229452 271880 229480
rect 231176 229440 231182 229452
rect 271874 229440 271880 229452
rect 271932 229440 271938 229492
rect 476022 229440 476028 229492
rect 476080 229480 476086 229492
rect 478598 229480 478604 229492
rect 476080 229452 478604 229480
rect 476080 229440 476086 229452
rect 478598 229440 478604 229452
rect 478656 229440 478662 229492
rect 530762 229440 530768 229492
rect 530820 229480 530826 229492
rect 538186 229480 538214 229588
rect 538306 229576 538312 229588
rect 538364 229576 538370 229628
rect 530820 229452 538214 229480
rect 530820 229440 530826 229452
rect 446398 229372 446404 229424
rect 446456 229412 446462 229424
rect 448790 229412 448796 229424
rect 446456 229384 448796 229412
rect 446456 229372 446462 229384
rect 448790 229372 448796 229384
rect 448848 229372 448854 229424
rect 450906 229372 450912 229424
rect 450964 229412 450970 229424
rect 453022 229412 453028 229424
rect 450964 229384 453028 229412
rect 450964 229372 450970 229384
rect 453022 229372 453028 229384
rect 453080 229372 453086 229424
rect 505646 229372 505652 229424
rect 505704 229412 505710 229424
rect 510982 229412 510988 229424
rect 505704 229384 510988 229412
rect 505704 229372 505710 229384
rect 510982 229372 510988 229384
rect 511040 229372 511046 229424
rect 673978 229412 674006 229724
rect 674242 229560 674294 229566
rect 674242 229502 674294 229508
rect 673978 229384 674130 229412
rect 147858 229344 147864 229356
rect 147140 229316 147864 229344
rect 147858 229304 147864 229316
rect 147916 229304 147922 229356
rect 151170 229304 151176 229356
rect 151228 229344 151234 229356
rect 151228 229316 156184 229344
rect 151228 229304 151234 229316
rect 123478 229168 123484 229220
rect 123536 229208 123542 229220
rect 149054 229208 149060 229220
rect 123536 229180 149060 229208
rect 123536 229168 123542 229180
rect 149054 229168 149060 229180
rect 149112 229168 149118 229220
rect 149606 229168 149612 229220
rect 149664 229208 149670 229220
rect 155954 229208 155960 229220
rect 149664 229180 155960 229208
rect 149664 229168 149670 229180
rect 155954 229168 155960 229180
rect 156012 229168 156018 229220
rect 156156 229208 156184 229316
rect 156322 229304 156328 229356
rect 156380 229344 156386 229356
rect 215202 229344 215208 229356
rect 156380 229316 215208 229344
rect 156380 229304 156386 229316
rect 215202 229304 215208 229316
rect 215260 229304 215266 229356
rect 246482 229304 246488 229356
rect 246540 229344 246546 229356
rect 282178 229344 282184 229356
rect 246540 229316 282184 229344
rect 246540 229304 246546 229316
rect 282178 229304 282184 229316
rect 282236 229304 282242 229356
rect 413830 229304 413836 229356
rect 413888 229344 413894 229356
rect 419994 229344 420000 229356
rect 413888 229316 420000 229344
rect 413888 229304 413894 229316
rect 419994 229304 420000 229316
rect 420052 229304 420058 229356
rect 450262 229236 450268 229288
rect 450320 229276 450326 229288
rect 451734 229276 451740 229288
rect 450320 229248 451740 229276
rect 450320 229236 450326 229248
rect 451734 229236 451740 229248
rect 451792 229236 451798 229288
rect 488258 229236 488264 229288
rect 488316 229276 488322 229288
rect 490374 229276 490380 229288
rect 488316 229248 490380 229276
rect 488316 229236 488322 229248
rect 490374 229236 490380 229248
rect 490432 229236 490438 229288
rect 495342 229236 495348 229288
rect 495400 229276 495406 229288
rect 500218 229276 500224 229288
rect 495400 229248 500224 229276
rect 495400 229236 495406 229248
rect 500218 229236 500224 229248
rect 500276 229236 500282 229288
rect 513374 229236 513380 229288
rect 513432 229276 513438 229288
rect 519354 229276 519360 229288
rect 513432 229248 519360 229276
rect 513432 229236 513438 229248
rect 519354 229236 519360 229248
rect 519412 229236 519418 229288
rect 161750 229208 161756 229220
rect 156156 229180 161756 229208
rect 161750 229168 161756 229180
rect 161808 229168 161814 229220
rect 164602 229168 164608 229220
rect 164660 229208 164666 229220
rect 174262 229208 174268 229220
rect 164660 229180 174268 229208
rect 164660 229168 164666 229180
rect 174262 229168 174268 229180
rect 174320 229168 174326 229220
rect 184658 229168 184664 229220
rect 184716 229208 184722 229220
rect 240962 229208 240968 229220
rect 184716 229180 240968 229208
rect 184716 229168 184722 229180
rect 240962 229168 240968 229180
rect 241020 229168 241026 229220
rect 423490 229100 423496 229152
rect 423548 229140 423554 229152
rect 427722 229140 427728 229152
rect 423548 229112 427728 229140
rect 423548 229100 423554 229112
rect 427722 229100 427728 229112
rect 427780 229100 427786 229152
rect 441246 229100 441252 229152
rect 441304 229140 441310 229152
rect 442074 229140 442080 229152
rect 441304 229112 442080 229140
rect 441304 229100 441310 229112
rect 442074 229100 442080 229112
rect 442132 229100 442138 229152
rect 503714 229100 503720 229152
rect 503772 229140 503778 229152
rect 509878 229140 509884 229152
rect 503772 229112 509884 229140
rect 503772 229100 503778 229112
rect 509878 229100 509884 229112
rect 509936 229100 509942 229152
rect 519170 229100 519176 229152
rect 519228 229140 519234 229152
rect 519228 229112 521654 229140
rect 519228 229100 519234 229112
rect 100662 229032 100668 229084
rect 100720 229072 100726 229084
rect 100720 229044 103514 229072
rect 100720 229032 100726 229044
rect 103486 228936 103514 229044
rect 106182 229032 106188 229084
rect 106240 229072 106246 229084
rect 142982 229072 142988 229084
rect 106240 229044 142988 229072
rect 106240 229032 106246 229044
rect 142982 229032 142988 229044
rect 143040 229032 143046 229084
rect 143442 229032 143448 229084
rect 143500 229072 143506 229084
rect 147122 229072 147128 229084
rect 143500 229044 147128 229072
rect 143500 229032 143506 229044
rect 147122 229032 147128 229044
rect 147180 229032 147186 229084
rect 147306 229032 147312 229084
rect 147364 229072 147370 229084
rect 202874 229072 202880 229084
rect 147364 229044 166948 229072
rect 147364 229032 147370 229044
rect 166920 229004 166948 229044
rect 167104 229044 202880 229072
rect 167104 229004 167132 229044
rect 202874 229032 202880 229044
rect 202932 229032 202938 229084
rect 204714 229032 204720 229084
rect 204772 229072 204778 229084
rect 212350 229072 212356 229084
rect 204772 229044 212356 229072
rect 204772 229032 204778 229044
rect 212350 229032 212356 229044
rect 212408 229032 212414 229084
rect 214374 229032 214380 229084
rect 214432 229072 214438 229084
rect 257062 229072 257068 229084
rect 214432 229044 257068 229072
rect 214432 229032 214438 229044
rect 257062 229032 257068 229044
rect 257120 229032 257126 229084
rect 257522 229032 257528 229084
rect 257580 229072 257586 229084
rect 296346 229072 296352 229084
rect 257580 229044 296352 229072
rect 257580 229032 257586 229044
rect 296346 229032 296352 229044
rect 296404 229032 296410 229084
rect 302142 229032 302148 229084
rect 302200 229072 302206 229084
rect 331122 229072 331128 229084
rect 302200 229044 331128 229072
rect 302200 229032 302206 229044
rect 331122 229032 331128 229044
rect 331180 229032 331186 229084
rect 166920 228976 167132 229004
rect 521626 229004 521654 229112
rect 524966 229100 524972 229152
rect 525024 229140 525030 229152
rect 529934 229140 529940 229152
rect 525024 229112 529940 229140
rect 525024 229100 525030 229112
rect 529934 229100 529940 229112
rect 529992 229100 529998 229152
rect 673730 229100 673736 229152
rect 673788 229140 673794 229152
rect 673788 229112 674038 229140
rect 673788 229100 673794 229112
rect 521626 228976 528554 229004
rect 164602 228936 164608 228948
rect 103486 228908 164608 228936
rect 164602 228896 164608 228908
rect 164660 228896 164666 228948
rect 167362 228896 167368 228948
rect 167420 228936 167426 228948
rect 169478 228936 169484 228948
rect 167420 228908 169484 228936
rect 167420 228896 167426 228908
rect 169478 228896 169484 228908
rect 169536 228896 169542 228948
rect 179782 228936 179788 228948
rect 171980 228908 179788 228936
rect 171980 228868 172008 228908
rect 179782 228896 179788 228908
rect 179840 228896 179846 228948
rect 180150 228896 180156 228948
rect 180208 228936 180214 228948
rect 180208 228908 220124 228936
rect 180208 228896 180214 228908
rect 171888 228840 172008 228868
rect 93762 228760 93768 228812
rect 93820 228800 93826 228812
rect 166810 228800 166816 228812
rect 93820 228772 166816 228800
rect 93820 228760 93826 228772
rect 166810 228760 166816 228772
rect 166868 228760 166874 228812
rect 166948 228760 166954 228812
rect 167006 228800 167012 228812
rect 171888 228800 171916 228840
rect 167006 228772 171916 228800
rect 167006 228760 167012 228772
rect 174814 228760 174820 228812
rect 174872 228800 174878 228812
rect 219802 228800 219808 228812
rect 174872 228772 219808 228800
rect 174872 228760 174878 228772
rect 219802 228760 219808 228772
rect 219860 228760 219866 228812
rect 220096 228800 220124 228908
rect 220354 228896 220360 228948
rect 220412 228936 220418 228948
rect 246758 228936 246764 228948
rect 220412 228908 246764 228936
rect 220412 228896 220418 228908
rect 246758 228896 246764 228908
rect 246816 228896 246822 228948
rect 257706 228896 257712 228948
rect 257764 228936 257770 228948
rect 299566 228936 299572 228948
rect 257764 228908 299572 228936
rect 257764 228896 257770 228908
rect 299566 228896 299572 228908
rect 299624 228896 299630 228948
rect 300670 228896 300676 228948
rect 300728 228936 300734 228948
rect 330478 228936 330484 228948
rect 300728 228908 330484 228936
rect 300728 228896 300734 228908
rect 330478 228896 330484 228908
rect 330536 228896 330542 228948
rect 517698 228936 517704 228948
rect 509206 228908 517704 228936
rect 226150 228800 226156 228812
rect 220096 228772 226156 228800
rect 226150 228760 226156 228772
rect 226208 228760 226214 228812
rect 238570 228760 238576 228812
rect 238628 228800 238634 228812
rect 282822 228800 282828 228812
rect 238628 228772 282828 228800
rect 238628 228760 238634 228772
rect 282822 228760 282828 228772
rect 282880 228760 282886 228812
rect 296622 228760 296628 228812
rect 296680 228800 296686 228812
rect 329190 228800 329196 228812
rect 296680 228772 329196 228800
rect 296680 228760 296686 228772
rect 329190 228760 329196 228772
rect 329248 228760 329254 228812
rect 336458 228760 336464 228812
rect 336516 228800 336522 228812
rect 358814 228800 358820 228812
rect 336516 228772 358820 228800
rect 336516 228760 336522 228772
rect 358814 228760 358820 228772
rect 358872 228760 358878 228812
rect 359918 228760 359924 228812
rect 359976 228800 359982 228812
rect 376846 228800 376852 228812
rect 359976 228772 376852 228800
rect 359976 228760 359982 228772
rect 376846 228760 376852 228772
rect 376904 228760 376910 228812
rect 478874 228760 478880 228812
rect 478932 228800 478938 228812
rect 490190 228800 490196 228812
rect 478932 228772 490196 228800
rect 478932 228760 478938 228772
rect 490190 228760 490196 228772
rect 490248 228760 490254 228812
rect 499850 228760 499856 228812
rect 499908 228800 499914 228812
rect 509206 228800 509234 228908
rect 517698 228896 517704 228908
rect 517756 228896 517762 228948
rect 528526 228936 528554 228976
rect 543182 228936 543188 228948
rect 528526 228908 543188 228936
rect 543182 228896 543188 228908
rect 543240 228896 543246 228948
rect 515766 228800 515772 228812
rect 499908 228772 509234 228800
rect 511920 228772 515772 228800
rect 499908 228760 499914 228772
rect 67542 228624 67548 228676
rect 67600 228664 67606 228676
rect 67600 228636 142844 228664
rect 67600 228624 67606 228636
rect 61654 228488 61660 228540
rect 61712 228528 61718 228540
rect 142430 228528 142436 228540
rect 61712 228500 142436 228528
rect 61712 228488 61718 228500
rect 142430 228488 142436 228500
rect 142488 228488 142494 228540
rect 57238 228352 57244 228404
rect 57296 228392 57302 228404
rect 141142 228392 141148 228404
rect 57296 228364 141148 228392
rect 57296 228352 57302 228364
rect 141142 228352 141148 228364
rect 141200 228352 141206 228404
rect 142816 228392 142844 228636
rect 142982 228624 142988 228676
rect 143040 228664 143046 228676
rect 152458 228664 152464 228676
rect 143040 228636 152464 228664
rect 143040 228624 143046 228636
rect 152458 228624 152464 228636
rect 152516 228624 152522 228676
rect 153102 228624 153108 228676
rect 153160 228664 153166 228676
rect 153160 228636 212212 228664
rect 153160 228624 153166 228636
rect 146110 228488 146116 228540
rect 146168 228528 146174 228540
rect 210694 228528 210700 228540
rect 146168 228500 210700 228528
rect 146168 228488 146174 228500
rect 210694 228488 210700 228500
rect 210752 228488 210758 228540
rect 212184 228528 212212 228636
rect 212350 228624 212356 228676
rect 212408 228664 212414 228676
rect 220354 228664 220360 228676
rect 212408 228636 220360 228664
rect 212408 228624 212414 228636
rect 220354 228624 220360 228636
rect 220412 228624 220418 228676
rect 220538 228624 220544 228676
rect 220596 228664 220602 228676
rect 264790 228664 264796 228676
rect 220596 228636 264796 228664
rect 220596 228624 220602 228636
rect 264790 228624 264796 228636
rect 264848 228624 264854 228676
rect 285490 228624 285496 228676
rect 285548 228664 285554 228676
rect 318886 228664 318892 228676
rect 285548 228636 318892 228664
rect 285548 228624 285554 228636
rect 318886 228624 318892 228636
rect 318944 228624 318950 228676
rect 325510 228624 325516 228676
rect 325568 228664 325574 228676
rect 349154 228664 349160 228676
rect 325568 228636 349160 228664
rect 325568 228624 325574 228636
rect 349154 228624 349160 228636
rect 349212 228624 349218 228676
rect 350166 228624 350172 228676
rect 350224 228664 350230 228676
rect 369118 228664 369124 228676
rect 350224 228636 369124 228664
rect 350224 228624 350230 228636
rect 369118 228624 369124 228636
rect 369176 228624 369182 228676
rect 377766 228624 377772 228676
rect 377824 228664 377830 228676
rect 390370 228664 390376 228676
rect 377824 228636 390376 228664
rect 377824 228624 377830 228636
rect 390370 228624 390376 228636
rect 390428 228624 390434 228676
rect 498562 228624 498568 228676
rect 498620 228664 498626 228676
rect 511920 228664 511948 228772
rect 515766 228760 515772 228772
rect 515824 228760 515830 228812
rect 518526 228760 518532 228812
rect 518584 228800 518590 228812
rect 541618 228800 541624 228812
rect 518584 228772 541624 228800
rect 518584 228760 518590 228772
rect 541618 228760 541624 228772
rect 541676 228760 541682 228812
rect 498620 228636 511948 228664
rect 498620 228624 498626 228636
rect 512086 228624 512092 228676
rect 512144 228664 512150 228676
rect 512144 228636 514156 228664
rect 512144 228624 512150 228636
rect 215846 228528 215852 228540
rect 212184 228500 215852 228528
rect 215846 228488 215852 228500
rect 215904 228488 215910 228540
rect 216214 228488 216220 228540
rect 216272 228528 216278 228540
rect 219618 228528 219624 228540
rect 216272 228500 219624 228528
rect 216272 228488 216278 228500
rect 219618 228488 219624 228500
rect 219676 228488 219682 228540
rect 219986 228488 219992 228540
rect 220044 228528 220050 228540
rect 260282 228528 260288 228540
rect 220044 228500 260288 228528
rect 220044 228488 220050 228500
rect 260282 228488 260288 228500
rect 260340 228488 260346 228540
rect 268930 228488 268936 228540
rect 268988 228528 268994 228540
rect 306006 228528 306012 228540
rect 268988 228500 306012 228528
rect 268988 228488 268994 228500
rect 306006 228488 306012 228500
rect 306064 228488 306070 228540
rect 313918 228488 313924 228540
rect 313976 228528 313982 228540
rect 320818 228528 320824 228540
rect 313976 228500 320824 228528
rect 313976 228488 313982 228500
rect 320818 228488 320824 228500
rect 320876 228488 320882 228540
rect 326890 228488 326896 228540
rect 326948 228528 326954 228540
rect 351086 228528 351092 228540
rect 326948 228500 351092 228528
rect 326948 228488 326954 228500
rect 351086 228488 351092 228500
rect 351144 228488 351150 228540
rect 354582 228488 354588 228540
rect 354640 228528 354646 228540
rect 372338 228528 372344 228540
rect 354640 228500 372344 228528
rect 354640 228488 354646 228500
rect 372338 228488 372344 228500
rect 372396 228488 372402 228540
rect 373442 228488 373448 228540
rect 373500 228528 373506 228540
rect 387150 228528 387156 228540
rect 373500 228500 387156 228528
rect 373500 228488 373506 228500
rect 387150 228488 387156 228500
rect 387208 228488 387214 228540
rect 390462 228488 390468 228540
rect 390520 228528 390526 228540
rect 400030 228528 400036 228540
rect 390520 228500 400036 228528
rect 390520 228488 390526 228500
rect 400030 228488 400036 228500
rect 400088 228488 400094 228540
rect 407758 228528 407764 228540
rect 400232 228500 407764 228528
rect 148870 228392 148876 228404
rect 142816 228364 148876 228392
rect 148870 228352 148876 228364
rect 148928 228352 148934 228404
rect 152458 228352 152464 228404
rect 152516 228392 152522 228404
rect 166810 228392 166816 228404
rect 152516 228364 166816 228392
rect 152516 228352 152522 228364
rect 166810 228352 166816 228364
rect 166868 228352 166874 228404
rect 166948 228352 166954 228404
rect 167006 228392 167012 228404
rect 214558 228392 214564 228404
rect 167006 228364 214564 228392
rect 167006 228352 167012 228364
rect 214558 228352 214564 228364
rect 214616 228352 214622 228404
rect 217502 228352 217508 228404
rect 217560 228392 217566 228404
rect 221458 228392 221464 228404
rect 217560 228364 221464 228392
rect 217560 228352 217566 228364
rect 221458 228352 221464 228364
rect 221516 228352 221522 228404
rect 224586 228352 224592 228404
rect 224644 228392 224650 228404
rect 273806 228392 273812 228404
rect 224644 228364 273812 228392
rect 224644 228352 224650 228364
rect 273806 228352 273812 228364
rect 273864 228352 273870 228404
rect 274266 228352 274272 228404
rect 274324 228392 274330 228404
rect 312446 228392 312452 228404
rect 274324 228364 312452 228392
rect 274324 228352 274330 228364
rect 312446 228352 312452 228364
rect 312504 228352 312510 228404
rect 320082 228352 320088 228404
rect 320140 228392 320146 228404
rect 346854 228392 346860 228404
rect 320140 228364 346860 228392
rect 320140 228352 320146 228364
rect 346854 228352 346860 228364
rect 346912 228352 346918 228404
rect 347038 228352 347044 228404
rect 347096 228392 347102 228404
rect 365898 228392 365904 228404
rect 347096 228364 365904 228392
rect 347096 228352 347102 228364
rect 365898 228352 365904 228364
rect 365956 228352 365962 228404
rect 371142 228352 371148 228404
rect 371200 228392 371206 228404
rect 385218 228392 385224 228404
rect 371200 228364 385224 228392
rect 371200 228352 371206 228364
rect 385218 228352 385224 228364
rect 385276 228352 385282 228404
rect 386230 228352 386236 228404
rect 386288 228392 386294 228404
rect 397454 228392 397460 228404
rect 386288 228364 397460 228392
rect 386288 228352 386294 228364
rect 397454 228352 397460 228364
rect 397512 228352 397518 228404
rect 112806 228216 112812 228268
rect 112864 228256 112870 228268
rect 184934 228256 184940 228268
rect 112864 228228 184940 228256
rect 112864 228216 112870 228228
rect 184934 228216 184940 228228
rect 184992 228216 184998 228268
rect 189718 228216 189724 228268
rect 189776 228256 189782 228268
rect 239030 228256 239036 228268
rect 189776 228228 239036 228256
rect 189776 228216 189782 228228
rect 239030 228216 239036 228228
rect 239088 228216 239094 228268
rect 254946 228216 254952 228268
rect 255004 228256 255010 228268
rect 295702 228256 295708 228268
rect 255004 228228 295708 228256
rect 255004 228216 255010 228228
rect 295702 228216 295708 228228
rect 295760 228216 295766 228268
rect 400232 228256 400260 228500
rect 407758 228488 407764 228500
rect 407816 228488 407822 228540
rect 409782 228488 409788 228540
rect 409840 228528 409846 228540
rect 415486 228528 415492 228540
rect 409840 228500 415492 228528
rect 409840 228488 409846 228500
rect 415486 228488 415492 228500
rect 415544 228488 415550 228540
rect 485682 228488 485688 228540
rect 485740 228528 485746 228540
rect 498286 228528 498292 228540
rect 485740 228500 498292 228528
rect 485740 228488 485746 228500
rect 498286 228488 498292 228500
rect 498344 228488 498350 228540
rect 502426 228488 502432 228540
rect 502484 228528 502490 228540
rect 502484 228500 514064 228528
rect 502484 228488 502490 228500
rect 402790 228352 402796 228404
rect 402848 228392 402854 228404
rect 411622 228392 411628 228404
rect 402848 228364 411628 228392
rect 402848 228352 402854 228364
rect 411622 228352 411628 228364
rect 411680 228352 411686 228404
rect 474458 228352 474464 228404
rect 474516 228392 474522 228404
rect 484578 228392 484584 228404
rect 474516 228364 484584 228392
rect 474516 228352 474522 228364
rect 484578 228352 484584 228364
rect 484636 228352 484642 228404
rect 485038 228352 485044 228404
rect 485096 228392 485102 228404
rect 498562 228392 498568 228404
rect 485096 228364 498568 228392
rect 485096 228352 485102 228364
rect 498562 228352 498568 228364
rect 498620 228352 498626 228404
rect 507118 228352 507124 228404
rect 507176 228392 507182 228404
rect 512730 228392 512736 228404
rect 507176 228364 512736 228392
rect 507176 228352 507182 228364
rect 512730 228352 512736 228364
rect 512788 228352 512794 228404
rect 400140 228228 400260 228256
rect 514036 228256 514064 228500
rect 514128 228392 514156 228636
rect 517882 228624 517888 228676
rect 517940 228664 517946 228676
rect 539410 228664 539416 228676
rect 517940 228636 539416 228664
rect 517940 228624 517946 228636
rect 539410 228624 539416 228636
rect 539468 228624 539474 228676
rect 539594 228624 539600 228676
rect 539652 228664 539658 228676
rect 555970 228664 555976 228676
rect 539652 228636 555976 228664
rect 539652 228624 539658 228636
rect 555970 228624 555976 228636
rect 556028 228624 556034 228676
rect 527542 228488 527548 228540
rect 527600 228528 527606 228540
rect 553302 228528 553308 228540
rect 527600 228500 553308 228528
rect 527600 228488 527606 228500
rect 553302 228488 553308 228500
rect 553360 228488 553366 228540
rect 555418 228488 555424 228540
rect 555476 228528 555482 228540
rect 571334 228528 571340 228540
rect 555476 228500 571340 228528
rect 555476 228488 555482 228500
rect 571334 228488 571340 228500
rect 571392 228488 571398 228540
rect 533338 228392 533344 228404
rect 514128 228364 533344 228392
rect 533338 228352 533344 228364
rect 533396 228352 533402 228404
rect 537202 228352 537208 228404
rect 537260 228392 537266 228404
rect 565630 228392 565636 228404
rect 537260 228364 565636 228392
rect 537260 228352 537266 228364
rect 565630 228352 565636 228364
rect 565688 228352 565694 228404
rect 520918 228256 520924 228268
rect 514036 228228 520924 228256
rect 400140 228132 400168 228228
rect 520918 228216 520924 228228
rect 520976 228216 520982 228268
rect 539410 228216 539416 228268
rect 539468 228256 539474 228268
rect 540790 228256 540796 228268
rect 539468 228228 540796 228256
rect 539468 228216 539474 228228
rect 540790 228216 540796 228228
rect 540848 228216 540854 228268
rect 119982 228080 119988 228132
rect 120040 228120 120046 228132
rect 190086 228120 190092 228132
rect 120040 228092 190092 228120
rect 120040 228080 120046 228092
rect 190086 228080 190092 228092
rect 190144 228080 190150 228132
rect 193030 228080 193036 228132
rect 193088 228120 193094 228132
rect 204714 228120 204720 228132
rect 193088 228092 204720 228120
rect 193088 228080 193094 228092
rect 204714 228080 204720 228092
rect 204772 228080 204778 228132
rect 214558 228080 214564 228132
rect 214616 228120 214622 228132
rect 214616 228092 215294 228120
rect 214616 228080 214622 228092
rect 126698 227944 126704 227996
rect 126756 227984 126762 227996
rect 195238 227984 195244 227996
rect 126756 227956 195244 227984
rect 126756 227944 126762 227956
rect 195238 227944 195244 227956
rect 195296 227944 195302 227996
rect 205450 227944 205456 227996
rect 205508 227984 205514 227996
rect 214374 227984 214380 227996
rect 205508 227956 214380 227984
rect 205508 227944 205514 227956
rect 214374 227944 214380 227956
rect 214432 227944 214438 227996
rect 215266 227984 215294 228092
rect 219802 228080 219808 228132
rect 219860 228120 219866 228132
rect 231302 228120 231308 228132
rect 219860 228092 231308 228120
rect 219860 228080 219866 228092
rect 231302 228080 231308 228092
rect 231360 228080 231366 228132
rect 233878 228080 233884 228132
rect 233936 228120 233942 228132
rect 272518 228120 272524 228132
rect 233936 228092 272524 228120
rect 233936 228080 233942 228092
rect 272518 228080 272524 228092
rect 272576 228080 272582 228132
rect 400122 228080 400128 228132
rect 400180 228080 400186 228132
rect 415026 228012 415032 228064
rect 415084 228052 415090 228064
rect 421926 228052 421932 228064
rect 415084 228024 421932 228052
rect 415084 228012 415090 228024
rect 421926 228012 421932 228024
rect 421984 228012 421990 228064
rect 220998 227984 221004 227996
rect 215266 227956 221004 227984
rect 220998 227944 221004 227956
rect 221056 227944 221062 227996
rect 221458 227944 221464 227996
rect 221516 227984 221522 227996
rect 251266 227984 251272 227996
rect 221516 227956 251272 227984
rect 221516 227944 221522 227956
rect 251266 227944 251272 227956
rect 251324 227944 251330 227996
rect 416682 227876 416688 227928
rect 416740 227916 416746 227928
rect 420638 227916 420644 227928
rect 416740 227888 420644 227916
rect 416740 227876 416746 227888
rect 420638 227876 420644 227888
rect 420696 227876 420702 227928
rect 447042 227876 447048 227928
rect 447100 227916 447106 227928
rect 450538 227916 450544 227928
rect 447100 227888 450544 227916
rect 447100 227876 447106 227888
rect 450538 227876 450544 227888
rect 450596 227876 450602 227928
rect 88242 227808 88248 227860
rect 88300 227848 88306 227860
rect 95234 227848 95240 227860
rect 88300 227820 95240 227848
rect 88300 227808 88306 227820
rect 95234 227808 95240 227820
rect 95292 227808 95298 227860
rect 133506 227808 133512 227860
rect 133564 227848 133570 227860
rect 200390 227848 200396 227860
rect 133564 227820 200396 227848
rect 133564 227808 133570 227820
rect 200390 227808 200396 227820
rect 200448 227808 200454 227860
rect 203518 227808 203524 227860
rect 203576 227848 203582 227860
rect 203576 227820 205128 227848
rect 203576 227808 203582 227820
rect 64782 227672 64788 227724
rect 64840 227712 64846 227724
rect 111058 227712 111064 227724
rect 64840 227684 111064 227712
rect 64840 227672 64846 227684
rect 111058 227672 111064 227684
rect 111116 227672 111122 227724
rect 117222 227672 117228 227724
rect 117280 227712 117286 227724
rect 117280 227684 184152 227712
rect 117280 227672 117286 227684
rect 110138 227536 110144 227588
rect 110196 227576 110202 227588
rect 182358 227576 182364 227588
rect 110196 227548 182364 227576
rect 110196 227536 110202 227548
rect 182358 227536 182364 227548
rect 182416 227536 182422 227588
rect 184124 227576 184152 227684
rect 185394 227672 185400 227724
rect 185452 227712 185458 227724
rect 192662 227712 192668 227724
rect 185452 227684 192668 227712
rect 185452 227672 185458 227684
rect 192662 227672 192668 227684
rect 192720 227672 192726 227724
rect 200022 227672 200028 227724
rect 200080 227712 200086 227724
rect 204898 227712 204904 227724
rect 200080 227684 204904 227712
rect 200080 227672 200086 227684
rect 204898 227672 204904 227684
rect 204956 227672 204962 227724
rect 205100 227712 205128 227820
rect 210970 227808 210976 227860
rect 211028 227848 211034 227860
rect 219986 227848 219992 227860
rect 211028 227820 219992 227848
rect 211028 227808 211034 227820
rect 219986 227808 219992 227820
rect 220044 227808 220050 227860
rect 226150 227808 226156 227860
rect 226208 227848 226214 227860
rect 233878 227848 233884 227860
rect 226208 227820 233884 227848
rect 226208 227808 226214 227820
rect 233878 227808 233884 227820
rect 233936 227808 233942 227860
rect 239306 227808 239312 227860
rect 239364 227848 239370 227860
rect 243538 227848 243544 227860
rect 239364 227820 243544 227848
rect 239364 227808 239370 227820
rect 243538 227808 243544 227820
rect 243596 227808 243602 227860
rect 246298 227808 246304 227860
rect 246356 227848 246362 227860
rect 248690 227848 248696 227860
rect 246356 227820 248696 227848
rect 246356 227808 246362 227820
rect 248690 227808 248696 227820
rect 248748 227808 248754 227860
rect 249058 227808 249064 227860
rect 249116 227848 249122 227860
rect 253842 227848 253848 227860
rect 249116 227820 253848 227848
rect 249116 227808 249122 227820
rect 253842 227808 253848 227820
rect 253900 227808 253906 227860
rect 331030 227740 331036 227792
rect 331088 227780 331094 227792
rect 334250 227780 334256 227792
rect 331088 227752 334256 227780
rect 331088 227740 331094 227752
rect 334250 227740 334256 227752
rect 334308 227740 334314 227792
rect 351086 227740 351092 227792
rect 351144 227780 351150 227792
rect 353018 227780 353024 227792
rect 351144 227752 353024 227780
rect 351144 227740 351150 227752
rect 353018 227740 353024 227752
rect 353076 227740 353082 227792
rect 371786 227740 371792 227792
rect 371844 227780 371850 227792
rect 373626 227780 373632 227792
rect 371844 227752 373632 227780
rect 371844 227740 371850 227752
rect 373626 227740 373632 227752
rect 373684 227740 373690 227792
rect 409046 227740 409052 227792
rect 409104 227780 409110 227792
rect 410334 227780 410340 227792
rect 409104 227752 410340 227780
rect 409104 227740 409110 227752
rect 410334 227740 410340 227752
rect 410392 227740 410398 227792
rect 411898 227740 411904 227792
rect 411956 227780 411962 227792
rect 413554 227780 413560 227792
rect 411956 227752 413560 227780
rect 411956 227740 411962 227752
rect 413554 227740 413560 227752
rect 413612 227740 413618 227792
rect 420638 227740 420644 227792
rect 420696 227780 420702 227792
rect 423858 227780 423864 227792
rect 420696 227752 423864 227780
rect 420696 227740 420702 227752
rect 423858 227740 423864 227752
rect 423916 227740 423922 227792
rect 471514 227740 471520 227792
rect 471572 227780 471578 227792
rect 479518 227780 479524 227792
rect 471572 227752 479524 227780
rect 471572 227740 471578 227752
rect 479518 227740 479524 227752
rect 479576 227740 479582 227792
rect 489914 227740 489920 227792
rect 489972 227780 489978 227792
rect 494698 227780 494704 227792
rect 489972 227752 494704 227780
rect 489972 227740 489978 227752
rect 494698 227740 494704 227752
rect 494756 227740 494762 227792
rect 664898 227740 664904 227792
rect 664956 227780 664962 227792
rect 665266 227780 665272 227792
rect 664956 227752 665272 227780
rect 664956 227740 664962 227752
rect 665266 227740 665272 227752
rect 665324 227740 665330 227792
rect 669130 227740 669136 227792
rect 669188 227780 669194 227792
rect 673638 227780 673644 227792
rect 669188 227752 673644 227780
rect 669188 227740 669194 227752
rect 673638 227740 673644 227752
rect 673696 227740 673702 227792
rect 217778 227712 217784 227724
rect 205100 227684 217784 227712
rect 217778 227672 217784 227684
rect 217836 227672 217842 227724
rect 219802 227672 219808 227724
rect 219860 227712 219866 227724
rect 228726 227712 228732 227724
rect 219860 227684 228732 227712
rect 219860 227672 219866 227684
rect 228726 227672 228732 227684
rect 228784 227672 228790 227724
rect 228910 227672 228916 227724
rect 228968 227712 228974 227724
rect 268010 227712 268016 227724
rect 228968 227684 268016 227712
rect 228968 227672 228974 227684
rect 268010 227672 268016 227684
rect 268068 227672 268074 227724
rect 293770 227672 293776 227724
rect 293828 227712 293834 227724
rect 325326 227712 325332 227724
rect 293828 227684 325332 227712
rect 293828 227672 293834 227684
rect 325326 227672 325332 227684
rect 325384 227672 325390 227724
rect 465902 227604 465908 227656
rect 465960 227644 465966 227656
rect 469858 227644 469864 227656
rect 465960 227616 469864 227644
rect 465960 227604 465966 227616
rect 469858 227604 469864 227616
rect 469916 227604 469922 227656
rect 187510 227576 187516 227588
rect 184124 227548 187516 227576
rect 187510 227536 187516 227548
rect 187568 227536 187574 227588
rect 214742 227576 214748 227588
rect 188356 227548 214748 227576
rect 60642 227400 60648 227452
rect 60700 227440 60706 227452
rect 102134 227440 102140 227452
rect 60700 227412 102140 227440
rect 60700 227400 60706 227412
rect 102134 227400 102140 227412
rect 102192 227400 102198 227452
rect 103422 227400 103428 227452
rect 103480 227440 103486 227452
rect 171226 227440 171232 227452
rect 103480 227412 171232 227440
rect 103480 227400 103486 227412
rect 171226 227400 171232 227412
rect 171284 227400 171290 227452
rect 172146 227400 172152 227452
rect 172204 227440 172210 227452
rect 177206 227440 177212 227452
rect 172204 227412 177212 227440
rect 172204 227400 172210 227412
rect 177206 227400 177212 227412
rect 177264 227400 177270 227452
rect 181346 227400 181352 227452
rect 181404 227440 181410 227452
rect 181404 227412 185900 227440
rect 181404 227400 181410 227412
rect 96430 227264 96436 227316
rect 96488 227304 96494 227316
rect 169478 227304 169484 227316
rect 96488 227276 157196 227304
rect 96488 227264 96494 227276
rect 157168 227236 157196 227276
rect 157444 227276 169484 227304
rect 157168 227208 157288 227236
rect 89622 227128 89628 227180
rect 89680 227168 89686 227180
rect 156690 227168 156696 227180
rect 89680 227140 156696 227168
rect 89680 227128 89686 227140
rect 156690 227128 156696 227140
rect 156748 227128 156754 227180
rect 157260 227168 157288 227208
rect 157444 227168 157472 227276
rect 169478 227264 169484 227276
rect 169536 227264 169542 227316
rect 185578 227304 185584 227316
rect 171336 227276 185584 227304
rect 157260 227140 157472 227168
rect 160186 227128 160192 227180
rect 160244 227168 160250 227180
rect 171336 227168 171364 227276
rect 185578 227264 185584 227276
rect 185636 227264 185642 227316
rect 185872 227304 185900 227412
rect 186130 227400 186136 227452
rect 186188 227440 186194 227452
rect 188356 227440 188384 227548
rect 214742 227536 214748 227548
rect 214800 227536 214806 227588
rect 214926 227536 214932 227588
rect 214984 227576 214990 227588
rect 262214 227576 262220 227588
rect 214984 227548 262220 227576
rect 214984 227536 214990 227548
rect 262214 227536 262220 227548
rect 262272 227536 262278 227588
rect 281350 227536 281356 227588
rect 281408 227576 281414 227588
rect 317598 227576 317604 227588
rect 281408 227548 317604 227576
rect 281408 227536 281414 227548
rect 317598 227536 317604 227548
rect 317656 227536 317662 227588
rect 337746 227536 337752 227588
rect 337804 227576 337810 227588
rect 345014 227576 345020 227588
rect 337804 227548 345020 227576
rect 337804 227536 337810 227548
rect 345014 227536 345020 227548
rect 345072 227536 345078 227588
rect 524598 227536 524604 227588
rect 524656 227576 524662 227588
rect 537478 227576 537484 227588
rect 524656 227548 537484 227576
rect 524656 227536 524662 227548
rect 537478 227536 537484 227548
rect 537536 227536 537542 227588
rect 186188 227412 188384 227440
rect 186188 227400 186194 227412
rect 189902 227400 189908 227452
rect 189960 227440 189966 227452
rect 204714 227440 204720 227452
rect 189960 227412 204720 227440
rect 189960 227400 189966 227412
rect 204714 227400 204720 227412
rect 204772 227400 204778 227452
rect 204898 227400 204904 227452
rect 204956 227440 204962 227452
rect 251910 227440 251916 227452
rect 204956 227412 251916 227440
rect 204956 227400 204962 227412
rect 251910 227400 251916 227412
rect 251968 227400 251974 227452
rect 264790 227400 264796 227452
rect 264848 227440 264854 227452
rect 304718 227440 304724 227452
rect 264848 227412 304724 227440
rect 264848 227400 264854 227412
rect 304718 227400 304724 227412
rect 304776 227400 304782 227452
rect 315482 227400 315488 227452
rect 315540 227440 315546 227452
rect 341426 227440 341432 227452
rect 315540 227412 341432 227440
rect 315540 227400 315546 227412
rect 341426 227400 341432 227412
rect 341484 227400 341490 227452
rect 352558 227400 352564 227452
rect 352616 227440 352622 227452
rect 363322 227440 363328 227452
rect 352616 227412 363328 227440
rect 352616 227400 352622 227412
rect 363322 227400 363328 227412
rect 363380 227400 363386 227452
rect 495066 227400 495072 227452
rect 495124 227440 495130 227452
rect 511166 227440 511172 227452
rect 495124 227412 511172 227440
rect 495124 227400 495130 227412
rect 511166 227400 511172 227412
rect 511224 227400 511230 227452
rect 514018 227400 514024 227452
rect 514076 227440 514082 227452
rect 535730 227440 535736 227452
rect 514076 227412 535736 227440
rect 514076 227400 514082 227412
rect 535730 227400 535736 227412
rect 535788 227400 535794 227452
rect 536098 227400 536104 227452
rect 536156 227440 536162 227452
rect 552474 227440 552480 227452
rect 536156 227412 552480 227440
rect 536156 227400 536162 227412
rect 552474 227400 552480 227412
rect 552532 227400 552538 227452
rect 219526 227304 219532 227316
rect 185872 227276 219532 227304
rect 219526 227264 219532 227276
rect 219584 227264 219590 227316
rect 219986 227264 219992 227316
rect 220044 227304 220050 227316
rect 241606 227304 241612 227316
rect 220044 227276 241612 227304
rect 220044 227264 220050 227276
rect 241606 227264 241612 227276
rect 241664 227264 241670 227316
rect 249426 227264 249432 227316
rect 249484 227304 249490 227316
rect 290550 227304 290556 227316
rect 249484 227276 290556 227304
rect 249484 227264 249490 227276
rect 290550 227264 290556 227276
rect 290608 227264 290614 227316
rect 291010 227264 291016 227316
rect 291068 227304 291074 227316
rect 322106 227304 322112 227316
rect 291068 227276 322112 227304
rect 291068 227264 291074 227276
rect 322106 227264 322112 227276
rect 322164 227264 322170 227316
rect 322290 227264 322296 227316
rect 322348 227304 322354 227316
rect 332410 227304 332416 227316
rect 322348 227276 332416 227304
rect 322348 227264 322354 227276
rect 332410 227264 332416 227276
rect 332468 227264 332474 227316
rect 333882 227264 333888 227316
rect 333940 227304 333946 227316
rect 356238 227304 356244 227316
rect 333940 227276 356244 227304
rect 333940 227264 333946 227276
rect 356238 227264 356244 227276
rect 356296 227264 356302 227316
rect 357250 227264 357256 227316
rect 357308 227304 357314 227316
rect 374270 227304 374276 227316
rect 357308 227276 374276 227304
rect 357308 227264 357314 227276
rect 374270 227264 374276 227276
rect 374328 227264 374334 227316
rect 382090 227264 382096 227316
rect 382148 227304 382154 227316
rect 392946 227304 392952 227316
rect 382148 227276 392952 227304
rect 382148 227264 382154 227276
rect 392946 227264 392952 227276
rect 393004 227264 393010 227316
rect 402606 227304 402612 227316
rect 393286 227276 402612 227304
rect 160244 227140 171364 227168
rect 160244 227128 160250 227140
rect 171594 227128 171600 227180
rect 171652 227168 171658 227180
rect 219802 227168 219808 227180
rect 171652 227140 219808 227168
rect 171652 227128 171658 227140
rect 219802 227128 219808 227140
rect 219860 227128 219866 227180
rect 233694 227168 233700 227180
rect 220096 227140 233700 227168
rect 56502 226992 56508 227044
rect 56560 227032 56566 227044
rect 142154 227032 142160 227044
rect 56560 227004 142160 227032
rect 56560 226992 56566 227004
rect 142154 226992 142160 227004
rect 142212 226992 142218 227044
rect 143258 226992 143264 227044
rect 143316 227032 143322 227044
rect 204070 227032 204076 227044
rect 143316 227004 204076 227032
rect 143316 226992 143322 227004
rect 204070 226992 204076 227004
rect 204128 226992 204134 227044
rect 214098 227032 214104 227044
rect 204916 227004 214104 227032
rect 122742 226856 122748 226908
rect 122800 226896 122806 226908
rect 185394 226896 185400 226908
rect 122800 226868 185400 226896
rect 122800 226856 122806 226868
rect 185394 226856 185400 226868
rect 185452 226856 185458 226908
rect 185578 226856 185584 226908
rect 185636 226896 185642 226908
rect 204916 226896 204944 227004
rect 214098 226992 214104 227004
rect 214156 226992 214162 227044
rect 220096 227032 220124 227140
rect 233694 227128 233700 227140
rect 233752 227128 233758 227180
rect 241146 227128 241152 227180
rect 241204 227168 241210 227180
rect 286686 227168 286692 227180
rect 241204 227140 286692 227168
rect 241204 227128 241210 227140
rect 286686 227128 286692 227140
rect 286744 227128 286750 227180
rect 306190 227128 306196 227180
rect 306248 227168 306254 227180
rect 336918 227168 336924 227180
rect 306248 227140 336924 227168
rect 306248 227128 306254 227140
rect 336918 227128 336924 227140
rect 336976 227128 336982 227180
rect 340690 227128 340696 227180
rect 340748 227168 340754 227180
rect 361390 227168 361396 227180
rect 340748 227140 361396 227168
rect 340748 227128 340754 227140
rect 361390 227128 361396 227140
rect 361448 227128 361454 227180
rect 363506 227128 363512 227180
rect 363564 227168 363570 227180
rect 368474 227168 368480 227180
rect 363564 227140 368480 227168
rect 363564 227128 363570 227140
rect 368474 227128 368480 227140
rect 368532 227128 368538 227180
rect 376662 227128 376668 227180
rect 376720 227168 376726 227180
rect 389726 227168 389732 227180
rect 376720 227140 389732 227168
rect 376720 227128 376726 227140
rect 389726 227128 389732 227140
rect 389784 227128 389790 227180
rect 393130 227128 393136 227180
rect 393188 227168 393194 227180
rect 393286 227168 393314 227276
rect 402606 227264 402612 227276
rect 402664 227264 402670 227316
rect 510982 227264 510988 227316
rect 511040 227304 511046 227316
rect 524414 227304 524420 227316
rect 511040 227276 524420 227304
rect 511040 227264 511046 227276
rect 524414 227264 524420 227276
rect 524472 227264 524478 227316
rect 526254 227264 526260 227316
rect 526312 227304 526318 227316
rect 551554 227304 551560 227316
rect 526312 227276 551560 227304
rect 526312 227264 526318 227276
rect 551554 227264 551560 227276
rect 551612 227264 551618 227316
rect 393188 227140 393314 227168
rect 393188 227128 393194 227140
rect 402238 227128 402244 227180
rect 402296 227168 402302 227180
rect 408402 227168 408408 227180
rect 402296 227140 408408 227168
rect 402296 227128 402302 227140
rect 408402 227128 408408 227140
rect 408460 227128 408466 227180
rect 478598 227128 478604 227180
rect 478656 227168 478662 227180
rect 486786 227168 486792 227180
rect 478656 227140 486792 227168
rect 478656 227128 478662 227140
rect 486786 227128 486792 227140
rect 486844 227128 486850 227180
rect 490374 227128 490380 227180
rect 490432 227168 490438 227180
rect 503162 227168 503168 227180
rect 490432 227140 503168 227168
rect 490432 227128 490438 227140
rect 503162 227128 503168 227140
rect 503220 227128 503226 227180
rect 504910 227128 504916 227180
rect 504968 227168 504974 227180
rect 523034 227168 523040 227180
rect 504968 227140 523040 227168
rect 504968 227128 504974 227140
rect 523034 227128 523040 227140
rect 523092 227128 523098 227180
rect 523678 227128 523684 227180
rect 523736 227168 523742 227180
rect 548518 227168 548524 227180
rect 523736 227140 548524 227168
rect 523736 227128 523742 227140
rect 548518 227128 548524 227140
rect 548576 227128 548582 227180
rect 556798 227128 556804 227180
rect 556856 227168 556862 227180
rect 570598 227168 570604 227180
rect 556856 227140 570604 227168
rect 556856 227128 556862 227140
rect 570598 227128 570604 227140
rect 570656 227128 570662 227180
rect 214576 227004 220124 227032
rect 214576 226896 214604 227004
rect 221826 226992 221832 227044
rect 221884 227032 221890 227044
rect 271230 227032 271236 227044
rect 221884 227004 271236 227032
rect 221884 226992 221890 227004
rect 271230 226992 271236 227004
rect 271288 226992 271294 227044
rect 271782 226992 271788 227044
rect 271840 227032 271846 227044
rect 308582 227032 308588 227044
rect 271840 227004 308588 227032
rect 271840 226992 271846 227004
rect 308582 226992 308588 227004
rect 308640 226992 308646 227044
rect 310330 226992 310336 227044
rect 310388 227032 310394 227044
rect 338206 227032 338212 227044
rect 310388 227004 338212 227032
rect 310388 226992 310394 227004
rect 338206 226992 338212 227004
rect 338264 226992 338270 227044
rect 338666 226992 338672 227044
rect 338724 227032 338730 227044
rect 360102 227032 360108 227044
rect 338724 227004 360108 227032
rect 338724 226992 338730 227004
rect 360102 226992 360108 227004
rect 360160 226992 360166 227044
rect 362770 226992 362776 227044
rect 362828 227032 362834 227044
rect 379054 227032 379060 227044
rect 362828 227004 379060 227032
rect 362828 226992 362834 227004
rect 379054 226992 379060 227004
rect 379112 226992 379118 227044
rect 391750 226992 391756 227044
rect 391808 227032 391814 227044
rect 403526 227032 403532 227044
rect 391808 227004 403532 227032
rect 391808 226992 391814 227004
rect 403526 226992 403532 227004
rect 403584 226992 403590 227044
rect 412542 226992 412548 227044
rect 412600 227032 412606 227044
rect 419350 227032 419356 227044
rect 412600 227004 419356 227032
rect 412600 226992 412606 227004
rect 419350 226992 419356 227004
rect 419408 226992 419414 227044
rect 486970 226992 486976 227044
rect 487028 227032 487034 227044
rect 500954 227032 500960 227044
rect 487028 227004 500960 227032
rect 487028 226992 487034 227004
rect 500954 226992 500960 227004
rect 501012 226992 501018 227044
rect 506290 226992 506296 227044
rect 506348 227032 506354 227044
rect 526622 227032 526628 227044
rect 506348 227004 526628 227032
rect 506348 226992 506354 227004
rect 526622 226992 526628 227004
rect 526680 226992 526686 227044
rect 533706 226992 533712 227044
rect 533764 227032 533770 227044
rect 560754 227032 560760 227044
rect 533764 227004 560760 227032
rect 533764 226992 533770 227004
rect 560754 226992 560760 227004
rect 560812 226992 560818 227044
rect 652018 226992 652024 227044
rect 652076 227032 652082 227044
rect 652076 227004 663794 227032
rect 652076 226992 652082 227004
rect 185636 226868 204944 226896
rect 209746 226868 214604 226896
rect 185636 226856 185642 226868
rect 129550 226720 129556 226772
rect 129608 226760 129614 226772
rect 197446 226760 197452 226772
rect 129608 226732 197452 226760
rect 129608 226720 129614 226732
rect 197446 226720 197452 226732
rect 197504 226720 197510 226772
rect 204714 226720 204720 226772
rect 204772 226760 204778 226772
rect 209746 226760 209774 226868
rect 214742 226856 214748 226908
rect 214800 226896 214806 226908
rect 219986 226896 219992 226908
rect 214800 226868 219992 226896
rect 214800 226856 214806 226868
rect 219986 226856 219992 226868
rect 220044 226856 220050 226908
rect 267366 226896 267372 226908
rect 229066 226868 267372 226896
rect 204772 226732 209774 226760
rect 204772 226720 204778 226732
rect 214098 226720 214104 226772
rect 214156 226760 214162 226772
rect 218422 226760 218428 226772
rect 214156 226732 218428 226760
rect 214156 226720 214162 226732
rect 218422 226720 218428 226732
rect 218480 226720 218486 226772
rect 219342 226720 219348 226772
rect 219400 226760 219406 226772
rect 229066 226760 229094 226868
rect 267366 226856 267372 226868
rect 267424 226856 267430 226908
rect 378778 226788 378784 226840
rect 378836 226828 378842 226840
rect 385862 226828 385868 226840
rect 378836 226800 385868 226828
rect 378836 226788 378842 226800
rect 385862 226788 385868 226800
rect 385920 226788 385926 226840
rect 663766 226828 663794 227004
rect 668946 226992 668952 227044
rect 669004 227032 669010 227044
rect 673454 227032 673460 227044
rect 669004 227004 673460 227032
rect 669004 226992 669010 227004
rect 673454 226992 673460 227004
rect 673512 226992 673518 227044
rect 673546 226828 673552 226840
rect 663766 226800 673552 226828
rect 673546 226788 673552 226800
rect 673604 226788 673610 226840
rect 676030 226788 676036 226840
rect 676088 226828 676094 226840
rect 678238 226828 678244 226840
rect 676088 226800 678244 226828
rect 676088 226788 676094 226800
rect 678238 226788 678244 226800
rect 678296 226788 678302 226840
rect 219400 226732 229094 226760
rect 219400 226720 219406 226732
rect 235810 226720 235816 226772
rect 235868 226760 235874 226772
rect 280246 226760 280252 226772
rect 235868 226732 280252 226760
rect 235868 226720 235874 226732
rect 280246 226720 280252 226732
rect 280304 226720 280310 226772
rect 136542 226584 136548 226636
rect 136600 226624 136606 226636
rect 203150 226624 203156 226636
rect 136600 226596 203156 226624
rect 136600 226584 136606 226596
rect 203150 226584 203156 226596
rect 203208 226584 203214 226636
rect 204070 226584 204076 226636
rect 204128 226624 204134 226636
rect 208118 226624 208124 226636
rect 204128 226596 208124 226624
rect 204128 226584 204134 226596
rect 208118 226584 208124 226596
rect 208176 226584 208182 226636
rect 212166 226584 212172 226636
rect 212224 226624 212230 226636
rect 214926 226624 214932 226636
rect 212224 226596 214932 226624
rect 212224 226584 212230 226596
rect 214926 226584 214932 226596
rect 214984 226584 214990 226636
rect 219526 226584 219532 226636
rect 219584 226624 219590 226636
rect 223574 226624 223580 226636
rect 219584 226596 223580 226624
rect 219584 226584 219590 226596
rect 223574 226584 223580 226596
rect 223632 226584 223638 226636
rect 225598 226584 225604 226636
rect 225656 226624 225662 226636
rect 238386 226624 238392 226636
rect 225656 226596 238392 226624
rect 225656 226584 225662 226596
rect 238386 226584 238392 226596
rect 238444 226584 238450 226636
rect 259362 226584 259368 226636
rect 259420 226624 259426 226636
rect 298278 226624 298284 226636
rect 259420 226596 298284 226624
rect 259420 226584 259426 226596
rect 298278 226584 298284 226596
rect 298336 226584 298342 226636
rect 673730 226556 673736 226568
rect 672842 226528 673736 226556
rect 673730 226516 673736 226528
rect 673788 226516 673794 226568
rect 106918 226448 106924 226500
rect 106976 226488 106982 226500
rect 146294 226488 146300 226500
rect 106976 226460 146300 226488
rect 106976 226448 106982 226460
rect 146294 226448 146300 226460
rect 146352 226448 146358 226500
rect 150066 226448 150072 226500
rect 150124 226488 150130 226500
rect 213270 226488 213276 226500
rect 150124 226460 213276 226488
rect 150124 226448 150130 226460
rect 213270 226448 213276 226460
rect 213328 226448 213334 226500
rect 216398 226448 216404 226500
rect 216456 226488 216462 226500
rect 220538 226488 220544 226500
rect 216456 226460 220544 226488
rect 216456 226448 216462 226460
rect 220538 226448 220544 226460
rect 220596 226448 220602 226500
rect 220722 226448 220728 226500
rect 220780 226488 220786 226500
rect 228910 226488 228916 226500
rect 220780 226460 228916 226488
rect 220780 226448 220786 226460
rect 228910 226448 228916 226460
rect 228968 226448 228974 226500
rect 369118 226448 369124 226500
rect 369176 226488 369182 226500
rect 376202 226488 376208 226500
rect 369176 226460 376208 226488
rect 369176 226448 369182 226460
rect 376202 226448 376208 226460
rect 376260 226448 376266 226500
rect 403986 226448 403992 226500
rect 404044 226488 404050 226500
rect 412266 226488 412272 226500
rect 404044 226460 412272 226488
rect 404044 226448 404050 226460
rect 412266 226448 412272 226460
rect 412324 226448 412330 226500
rect 474734 226448 474740 226500
rect 474792 226488 474798 226500
rect 482738 226488 482744 226500
rect 474792 226460 482744 226488
rect 474792 226448 474798 226460
rect 482738 226448 482744 226460
rect 482796 226448 482802 226500
rect 672724 226432 672776 226438
rect 386046 226380 386052 226432
rect 386104 226420 386110 226432
rect 391198 226420 391204 226432
rect 386104 226392 391204 226420
rect 386104 226380 386110 226392
rect 391198 226380 391204 226392
rect 391256 226380 391262 226432
rect 672724 226374 672776 226380
rect 407758 226312 407764 226364
rect 407816 226352 407822 226364
rect 408678 226352 408684 226364
rect 407816 226324 408684 226352
rect 407816 226312 407822 226324
rect 408678 226312 408684 226324
rect 408736 226312 408742 226364
rect 481634 226312 481640 226364
rect 481692 226352 481698 226364
rect 487798 226352 487804 226364
rect 481692 226324 487804 226352
rect 481692 226312 481698 226324
rect 487798 226312 487804 226324
rect 487856 226312 487862 226364
rect 488074 226312 488080 226364
rect 488132 226352 488138 226364
rect 490006 226352 490012 226364
rect 488132 226324 490012 226352
rect 488132 226312 488138 226324
rect 490006 226312 490012 226324
rect 490064 226312 490070 226364
rect 122558 226244 122564 226296
rect 122616 226284 122622 226296
rect 193950 226284 193956 226296
rect 122616 226256 193956 226284
rect 122616 226244 122622 226256
rect 193950 226244 193956 226256
rect 194008 226244 194014 226296
rect 195238 226244 195244 226296
rect 195296 226284 195302 226296
rect 201678 226284 201684 226296
rect 195296 226256 201684 226284
rect 195296 226244 195302 226256
rect 201678 226244 201684 226256
rect 201736 226244 201742 226296
rect 203150 226244 203156 226296
rect 203208 226284 203214 226296
rect 209406 226284 209412 226296
rect 203208 226256 209412 226284
rect 203208 226244 203214 226256
rect 209406 226244 209412 226256
rect 209464 226244 209470 226296
rect 209590 226244 209596 226296
rect 209648 226284 209654 226296
rect 255130 226284 255136 226296
rect 209648 226256 255136 226284
rect 209648 226244 209654 226256
rect 255130 226244 255136 226256
rect 255188 226244 255194 226296
rect 260650 226244 260656 226296
rect 260708 226284 260714 226296
rect 298922 226284 298928 226296
rect 260708 226256 298928 226284
rect 260708 226244 260714 226256
rect 298922 226244 298928 226256
rect 298980 226244 298986 226296
rect 308858 226244 308864 226296
rect 308916 226284 308922 226296
rect 336274 226284 336280 226296
rect 308916 226256 336280 226284
rect 308916 226244 308922 226256
rect 336274 226244 336280 226256
rect 336332 226244 336338 226296
rect 388622 226244 388628 226296
rect 388680 226284 388686 226296
rect 394234 226284 394240 226296
rect 388680 226256 394240 226284
rect 388680 226244 388686 226256
rect 394234 226244 394240 226256
rect 394292 226244 394298 226296
rect 458634 226244 458640 226296
rect 458692 226284 458698 226296
rect 462958 226284 462964 226296
rect 458692 226256 462964 226284
rect 458692 226244 458698 226256
rect 462958 226244 462964 226256
rect 463016 226244 463022 226296
rect 539962 226284 539968 226296
rect 528526 226256 539968 226284
rect 72418 226108 72424 226160
rect 72476 226148 72482 226160
rect 141142 226148 141148 226160
rect 72476 226120 141148 226148
rect 72476 226108 72482 226120
rect 141142 226108 141148 226120
rect 141200 226108 141206 226160
rect 141510 226108 141516 226160
rect 141568 226148 141574 226160
rect 145006 226148 145012 226160
rect 141568 226120 145012 226148
rect 141568 226108 141574 226120
rect 145006 226108 145012 226120
rect 145064 226108 145070 226160
rect 145190 226108 145196 226160
rect 145248 226148 145254 226160
rect 147490 226148 147496 226160
rect 145248 226120 147496 226148
rect 145248 226108 145254 226120
rect 147490 226108 147496 226120
rect 147548 226108 147554 226160
rect 148962 226108 148968 226160
rect 149020 226148 149026 226160
rect 214558 226148 214564 226160
rect 149020 226120 214564 226148
rect 149020 226108 149026 226120
rect 214558 226108 214564 226120
rect 214616 226108 214622 226160
rect 222010 226108 222016 226160
rect 222068 226148 222074 226160
rect 269942 226148 269948 226160
rect 222068 226120 269948 226148
rect 222068 226108 222074 226120
rect 269942 226108 269948 226120
rect 270000 226108 270006 226160
rect 270218 226108 270224 226160
rect 270276 226148 270282 226160
rect 287514 226148 287520 226160
rect 270276 226120 287520 226148
rect 270276 226108 270282 226120
rect 287514 226108 287520 226120
rect 287572 226108 287578 226160
rect 288066 226108 288072 226160
rect 288124 226148 288130 226160
rect 322750 226148 322756 226160
rect 288124 226120 322756 226148
rect 288124 226108 288130 226120
rect 322750 226108 322756 226120
rect 322808 226108 322814 226160
rect 526438 226108 526444 226160
rect 526496 226148 526502 226160
rect 528526 226148 528554 226256
rect 539962 226244 539968 226256
rect 540020 226244 540026 226296
rect 563698 226244 563704 226296
rect 563756 226284 563762 226296
rect 568114 226284 568120 226296
rect 563756 226256 568120 226284
rect 563756 226244 563762 226256
rect 568114 226244 568120 226256
rect 568172 226244 568178 226296
rect 672604 226160 672656 226166
rect 538490 226148 538496 226160
rect 526496 226120 528554 226148
rect 538186 226120 538496 226148
rect 526496 226108 526502 226120
rect 83458 225972 83464 226024
rect 83516 226012 83522 226024
rect 163038 226012 163044 226024
rect 83516 225984 163044 226012
rect 83516 225972 83522 225984
rect 163038 225972 163044 225984
rect 163096 225972 163102 226024
rect 193766 225972 193772 226024
rect 193824 226012 193830 226024
rect 199286 226012 199292 226024
rect 193824 225984 199292 226012
rect 193824 225972 193830 225984
rect 199286 225972 199292 225984
rect 199344 225972 199350 226024
rect 199470 225972 199476 226024
rect 199528 226012 199534 226024
rect 236454 226012 236460 226024
rect 199528 225984 236460 226012
rect 199528 225972 199534 225984
rect 236454 225972 236460 225984
rect 236512 225972 236518 226024
rect 252462 225972 252468 226024
rect 252520 226012 252526 226024
rect 293126 226012 293132 226024
rect 252520 225984 293132 226012
rect 252520 225972 252526 225984
rect 293126 225972 293132 225984
rect 293184 225972 293190 226024
rect 299382 225972 299388 226024
rect 299440 226012 299446 226024
rect 328546 226012 328552 226024
rect 299440 225984 328552 226012
rect 299440 225972 299446 225984
rect 328546 225972 328552 225984
rect 328604 225972 328610 226024
rect 335170 225972 335176 226024
rect 335228 226012 335234 226024
rect 356882 226012 356888 226024
rect 335228 225984 356888 226012
rect 335228 225972 335234 225984
rect 356882 225972 356888 225984
rect 356940 225972 356946 226024
rect 361206 225972 361212 226024
rect 361264 226012 361270 226024
rect 377490 226012 377496 226024
rect 361264 225984 377496 226012
rect 361264 225972 361270 225984
rect 377490 225972 377496 225984
rect 377548 225972 377554 226024
rect 498102 225972 498108 226024
rect 498160 226012 498166 226024
rect 514294 226012 514300 226024
rect 498160 225984 514300 226012
rect 498160 225972 498166 225984
rect 514294 225972 514300 225984
rect 514352 225972 514358 226024
rect 516594 225972 516600 226024
rect 516652 226012 516658 226024
rect 538186 226012 538214 226120
rect 538490 226108 538496 226120
rect 538548 226108 538554 226160
rect 672604 226102 672656 226108
rect 671246 226040 671252 226092
rect 671304 226080 671310 226092
rect 671304 226052 672520 226080
rect 671304 226040 671310 226052
rect 516652 225984 538214 226012
rect 516652 225972 516658 225984
rect 538306 225972 538312 226024
rect 538364 226012 538370 226024
rect 556154 226012 556160 226024
rect 538364 225984 556160 226012
rect 538364 225972 538370 225984
rect 556154 225972 556160 225984
rect 556212 226012 556218 226024
rect 557442 226012 557448 226024
rect 556212 225984 557448 226012
rect 556212 225972 556218 225984
rect 557442 225972 557448 225984
rect 557500 225972 557506 226024
rect 76558 225836 76564 225888
rect 76616 225876 76622 225888
rect 158254 225876 158260 225888
rect 76616 225848 158260 225876
rect 76616 225836 76622 225848
rect 158254 225836 158260 225848
rect 158312 225836 158318 225888
rect 169662 225836 169668 225888
rect 169720 225876 169726 225888
rect 171594 225876 171600 225888
rect 169720 225848 171600 225876
rect 169720 225836 169726 225848
rect 171594 225836 171600 225848
rect 171652 225836 171658 225888
rect 171778 225836 171784 225888
rect 171836 225876 171842 225888
rect 204530 225876 204536 225888
rect 171836 225848 204536 225876
rect 171836 225836 171842 225848
rect 204530 225836 204536 225848
rect 204588 225836 204594 225888
rect 204714 225836 204720 225888
rect 204772 225876 204778 225888
rect 249242 225876 249248 225888
rect 204772 225848 249248 225876
rect 204772 225836 204778 225848
rect 249242 225836 249248 225848
rect 249300 225836 249306 225888
rect 261846 225836 261852 225888
rect 261904 225876 261910 225888
rect 300854 225876 300860 225888
rect 261904 225848 300860 225876
rect 261904 225836 261910 225848
rect 300854 225836 300860 225848
rect 300912 225836 300918 225888
rect 312906 225836 312912 225888
rect 312964 225876 312970 225888
rect 341702 225876 341708 225888
rect 312964 225848 341708 225876
rect 312964 225836 312970 225848
rect 341702 225836 341708 225848
rect 341760 225836 341766 225888
rect 341978 225836 341984 225888
rect 342036 225876 342042 225888
rect 365254 225876 365260 225888
rect 342036 225848 365260 225876
rect 342036 225836 342042 225848
rect 365254 225836 365260 225848
rect 365312 225836 365318 225888
rect 375006 225836 375012 225888
rect 375064 225876 375070 225888
rect 387794 225876 387800 225888
rect 375064 225848 387800 225876
rect 375064 225836 375070 225848
rect 387794 225836 387800 225848
rect 387852 225836 387858 225888
rect 394326 225836 394332 225888
rect 394384 225876 394390 225888
rect 403250 225876 403256 225888
rect 394384 225848 403256 225876
rect 394384 225836 394390 225848
rect 403250 225836 403256 225848
rect 403308 225836 403314 225888
rect 501138 225836 501144 225888
rect 501196 225876 501202 225888
rect 519170 225876 519176 225888
rect 501196 225848 519176 225876
rect 501196 225836 501202 225848
rect 519170 225836 519176 225848
rect 519228 225836 519234 225888
rect 521746 225836 521752 225888
rect 521804 225876 521810 225888
rect 545758 225876 545764 225888
rect 521804 225848 545764 225876
rect 521804 225836 521810 225848
rect 545758 225836 545764 225848
rect 545816 225836 545822 225888
rect 672258 225836 672264 225888
rect 672316 225876 672322 225888
rect 672316 225848 672406 225876
rect 672316 225836 672322 225848
rect 66162 225700 66168 225752
rect 66220 225740 66226 225752
rect 149790 225740 149796 225752
rect 66220 225712 149796 225740
rect 66220 225700 66226 225712
rect 149790 225700 149796 225712
rect 149848 225700 149854 225752
rect 151262 225700 151268 225752
rect 151320 225740 151326 225752
rect 151320 225712 203380 225740
rect 151320 225700 151326 225712
rect 58986 225564 58992 225616
rect 59044 225604 59050 225616
rect 141510 225604 141516 225616
rect 59044 225576 141516 225604
rect 59044 225564 59050 225576
rect 141510 225564 141516 225576
rect 141568 225564 141574 225616
rect 141786 225564 141792 225616
rect 141844 225604 141850 225616
rect 203150 225604 203156 225616
rect 141844 225576 203156 225604
rect 141844 225564 141850 225576
rect 203150 225564 203156 225576
rect 203208 225564 203214 225616
rect 203352 225604 203380 225712
rect 204898 225700 204904 225752
rect 204956 225740 204962 225752
rect 244182 225740 244188 225752
rect 204956 225712 244188 225740
rect 204956 225700 204962 225712
rect 244182 225700 244188 225712
rect 244240 225700 244246 225752
rect 251082 225700 251088 225752
rect 251140 225740 251146 225752
rect 294414 225740 294420 225752
rect 251140 225712 294420 225740
rect 251140 225700 251146 225712
rect 294414 225700 294420 225712
rect 294472 225700 294478 225752
rect 296438 225700 296444 225752
rect 296496 225740 296502 225752
rect 327902 225740 327908 225752
rect 296496 225712 327908 225740
rect 296496 225700 296502 225712
rect 327902 225700 327908 225712
rect 327960 225700 327966 225752
rect 329742 225700 329748 225752
rect 329800 225740 329806 225752
rect 353662 225740 353668 225752
rect 329800 225712 353668 225740
rect 329800 225700 329806 225712
rect 353662 225700 353668 225712
rect 353720 225700 353726 225752
rect 365346 225700 365352 225752
rect 365404 225740 365410 225752
rect 383286 225740 383292 225752
rect 365404 225712 383292 225740
rect 365404 225700 365410 225712
rect 383286 225700 383292 225712
rect 383344 225700 383350 225752
rect 387702 225700 387708 225752
rect 387760 225740 387766 225752
rect 397822 225740 397828 225752
rect 387760 225712 397828 225740
rect 387760 225700 387766 225712
rect 397822 225700 397828 225712
rect 397880 225700 397886 225752
rect 481174 225700 481180 225752
rect 481232 225740 481238 225752
rect 492674 225740 492680 225752
rect 481232 225712 492680 225740
rect 481232 225700 481238 225712
rect 492674 225700 492680 225712
rect 492732 225700 492738 225752
rect 493778 225700 493784 225752
rect 493836 225740 493842 225752
rect 505278 225740 505284 225752
rect 493836 225712 505284 225740
rect 493836 225700 493842 225712
rect 505278 225700 505284 225712
rect 505336 225700 505342 225752
rect 508866 225700 508872 225752
rect 508924 225740 508930 225752
rect 529198 225740 529204 225752
rect 508924 225712 529204 225740
rect 508924 225700 508930 225712
rect 529198 225700 529204 225712
rect 529256 225700 529262 225752
rect 535914 225700 535920 225752
rect 535972 225740 535978 225752
rect 563054 225740 563060 225752
rect 535972 225712 563060 225740
rect 535972 225700 535978 225712
rect 563054 225700 563060 225712
rect 563112 225700 563118 225752
rect 217134 225604 217140 225616
rect 203352 225576 217140 225604
rect 217134 225564 217140 225576
rect 217192 225564 217198 225616
rect 219986 225564 219992 225616
rect 220044 225604 220050 225616
rect 266078 225604 266084 225616
rect 220044 225576 266084 225604
rect 220044 225564 220050 225576
rect 266078 225564 266084 225576
rect 266136 225564 266142 225616
rect 266998 225564 267004 225616
rect 267056 225604 267062 225616
rect 274450 225604 274456 225616
rect 267056 225576 274456 225604
rect 267056 225564 267062 225576
rect 274450 225564 274456 225576
rect 274508 225564 274514 225616
rect 278406 225564 278412 225616
rect 278464 225604 278470 225616
rect 313274 225604 313280 225616
rect 278464 225576 313280 225604
rect 278464 225564 278470 225576
rect 313274 225564 313280 225576
rect 313332 225564 313338 225616
rect 327718 225564 327724 225616
rect 327776 225604 327782 225616
rect 352374 225604 352380 225616
rect 327776 225576 352380 225604
rect 327776 225564 327782 225576
rect 352374 225564 352380 225576
rect 352432 225564 352438 225616
rect 352926 225564 352932 225616
rect 352984 225604 352990 225616
rect 371602 225604 371608 225616
rect 352984 225576 371608 225604
rect 352984 225564 352990 225576
rect 371602 225564 371608 225576
rect 371660 225564 371666 225616
rect 382918 225564 382924 225616
rect 382976 225604 382982 225616
rect 396166 225604 396172 225616
rect 382976 225576 396172 225604
rect 382976 225564 382982 225576
rect 396166 225564 396172 225576
rect 396224 225564 396230 225616
rect 410978 225564 410984 225616
rect 411036 225604 411042 225616
rect 416130 225604 416136 225616
rect 411036 225576 416136 225604
rect 411036 225564 411042 225576
rect 416130 225564 416136 225576
rect 416188 225564 416194 225616
rect 467650 225564 467656 225616
rect 467708 225604 467714 225616
rect 476574 225604 476580 225616
rect 467708 225576 476580 225604
rect 467708 225564 467714 225576
rect 476574 225564 476580 225576
rect 476632 225564 476638 225616
rect 477310 225564 477316 225616
rect 477368 225604 477374 225616
rect 488718 225604 488724 225616
rect 477368 225576 488724 225604
rect 477368 225564 477374 225576
rect 488718 225564 488724 225576
rect 488776 225564 488782 225616
rect 489362 225564 489368 225616
rect 489420 225604 489426 225616
rect 502978 225604 502984 225616
rect 489420 225576 502984 225604
rect 489420 225564 489426 225576
rect 502978 225564 502984 225576
rect 503036 225564 503042 225616
rect 510154 225564 510160 225616
rect 510212 225604 510218 225616
rect 530946 225604 530952 225616
rect 510212 225576 530952 225604
rect 510212 225564 510218 225576
rect 530946 225564 530952 225576
rect 531004 225564 531010 225616
rect 531406 225564 531412 225616
rect 531464 225604 531470 225616
rect 558178 225604 558184 225616
rect 531464 225576 558184 225604
rect 531464 225564 531470 225576
rect 558178 225564 558184 225576
rect 558236 225564 558242 225616
rect 672264 225548 672316 225554
rect 672264 225490 672316 225496
rect 125226 225428 125232 225480
rect 125284 225468 125290 225480
rect 196158 225468 196164 225480
rect 125284 225440 196164 225468
rect 125284 225428 125290 225440
rect 196158 225428 196164 225440
rect 196216 225428 196222 225480
rect 197998 225428 198004 225480
rect 198056 225468 198062 225480
rect 204714 225468 204720 225480
rect 198056 225440 204720 225468
rect 198056 225428 198062 225440
rect 204714 225428 204720 225440
rect 204772 225428 204778 225480
rect 205082 225428 205088 225480
rect 205140 225468 205146 225480
rect 209314 225468 209320 225480
rect 205140 225440 209320 225468
rect 205140 225428 205146 225440
rect 209314 225428 209320 225440
rect 209372 225428 209378 225480
rect 209498 225428 209504 225480
rect 209556 225468 209562 225480
rect 259638 225468 259644 225480
rect 209556 225440 259644 225468
rect 209556 225428 209562 225440
rect 259638 225428 259644 225440
rect 259696 225428 259702 225480
rect 297358 225428 297364 225480
rect 297416 225468 297422 225480
rect 310514 225468 310520 225480
rect 297416 225440 310520 225468
rect 297416 225428 297422 225440
rect 310514 225428 310520 225440
rect 310572 225428 310578 225480
rect 463142 225360 463148 225412
rect 463200 225400 463206 225412
rect 467282 225400 467288 225412
rect 463200 225372 467288 225400
rect 463200 225360 463206 225372
rect 467282 225360 467288 225372
rect 467340 225360 467346 225412
rect 672156 225344 672208 225350
rect 129366 225292 129372 225344
rect 129424 225332 129430 225344
rect 199102 225332 199108 225344
rect 129424 225304 199108 225332
rect 129424 225292 129430 225304
rect 199102 225292 199108 225304
rect 199160 225292 199166 225344
rect 199286 225292 199292 225344
rect 199344 225332 199350 225344
rect 204898 225332 204904 225344
rect 199344 225304 204904 225332
rect 199344 225292 199350 225304
rect 204898 225292 204904 225304
rect 204956 225292 204962 225344
rect 222930 225332 222936 225344
rect 205100 225304 222936 225332
rect 62022 225156 62028 225208
rect 62080 225196 62086 225208
rect 130378 225196 130384 225208
rect 62080 225168 130384 225196
rect 62080 225156 62086 225168
rect 130378 225156 130384 225168
rect 130436 225156 130442 225208
rect 132402 225156 132408 225208
rect 132460 225196 132466 225208
rect 195238 225196 195244 225208
rect 132460 225168 195244 225196
rect 132460 225156 132466 225168
rect 195238 225156 195244 225168
rect 195296 225156 195302 225208
rect 196618 225156 196624 225208
rect 196676 225196 196682 225208
rect 199470 225196 199476 225208
rect 196676 225168 199476 225196
rect 196676 225156 196682 225168
rect 199470 225156 199476 225168
rect 199528 225156 199534 225208
rect 202782 225156 202788 225208
rect 202840 225196 202846 225208
rect 202840 225168 204484 225196
rect 202840 225156 202846 225168
rect 135162 225020 135168 225072
rect 135220 225060 135226 225072
rect 204254 225060 204260 225072
rect 135220 225032 204260 225060
rect 135220 225020 135226 225032
rect 204254 225020 204260 225032
rect 204312 225020 204318 225072
rect 204456 225060 204484 225168
rect 204622 225156 204628 225208
rect 204680 225196 204686 225208
rect 205100 225196 205128 225304
rect 222930 225292 222936 225304
rect 222988 225292 222994 225344
rect 242894 225292 242900 225344
rect 242952 225332 242958 225344
rect 285030 225332 285036 225344
rect 242952 225304 285036 225332
rect 242952 225292 242958 225304
rect 285030 225292 285036 225304
rect 285088 225292 285094 225344
rect 672156 225286 672208 225292
rect 672034 225276 672086 225282
rect 672034 225218 672086 225224
rect 254486 225196 254492 225208
rect 204680 225168 205128 225196
rect 209746 225168 254492 225196
rect 204680 225156 204686 225168
rect 209746 225060 209774 225168
rect 254486 225156 254492 225168
rect 254544 225156 254550 225208
rect 204456 225032 209774 225060
rect 215202 225020 215208 225072
rect 215260 225060 215266 225072
rect 219986 225060 219992 225072
rect 215260 225032 219992 225060
rect 215260 225020 215266 225032
rect 219986 225020 219992 225032
rect 220044 225020 220050 225072
rect 666462 225020 666468 225072
rect 666520 225060 666526 225072
rect 666520 225032 671968 225060
rect 666520 225020 666526 225032
rect 355226 224952 355232 225004
rect 355284 224992 355290 225004
rect 358170 224992 358176 225004
rect 355284 224964 358176 224992
rect 355284 224952 355290 224964
rect 358170 224952 358176 224964
rect 358228 224952 358234 225004
rect 404170 224952 404176 225004
rect 404228 224992 404234 225004
rect 410610 224992 410616 225004
rect 404228 224964 410616 224992
rect 404228 224952 404234 224964
rect 410610 224952 410616 224964
rect 410668 224952 410674 225004
rect 416498 224952 416504 225004
rect 416556 224992 416562 225004
rect 422202 224992 422208 225004
rect 416556 224964 422208 224992
rect 416556 224952 416562 224964
rect 422202 224952 422208 224964
rect 422260 224952 422266 225004
rect 96246 224884 96252 224936
rect 96304 224924 96310 224936
rect 172974 224924 172980 224936
rect 96304 224896 172980 224924
rect 96304 224884 96310 224896
rect 172974 224884 172980 224896
rect 173032 224884 173038 224936
rect 176838 224884 176844 224936
rect 176896 224924 176902 224936
rect 176896 224896 178724 224924
rect 176896 224884 176902 224896
rect 89438 224748 89444 224800
rect 89496 224788 89502 224800
rect 168190 224788 168196 224800
rect 89496 224760 168196 224788
rect 89496 224748 89502 224760
rect 168190 224748 168196 224760
rect 168248 224748 168254 224800
rect 170858 224748 170864 224800
rect 170916 224788 170922 224800
rect 178494 224788 178500 224800
rect 170916 224760 178500 224788
rect 170916 224748 170922 224760
rect 178494 224748 178500 224760
rect 178552 224748 178558 224800
rect 178696 224788 178724 224896
rect 179322 224884 179328 224936
rect 179380 224924 179386 224936
rect 185578 224924 185584 224936
rect 179380 224896 185584 224924
rect 179380 224884 179386 224896
rect 185578 224884 185584 224896
rect 185636 224884 185642 224936
rect 185762 224884 185768 224936
rect 185820 224924 185826 224936
rect 199746 224924 199752 224936
rect 185820 224896 199752 224924
rect 185820 224884 185826 224896
rect 199746 224884 199752 224896
rect 199804 224884 199810 224936
rect 199930 224884 199936 224936
rect 199988 224924 199994 224936
rect 248046 224924 248052 224936
rect 199988 224896 248052 224924
rect 199988 224884 199994 224896
rect 248046 224884 248052 224896
rect 248104 224884 248110 224936
rect 272518 224884 272524 224936
rect 272576 224924 272582 224936
rect 309870 224924 309876 224936
rect 272576 224896 309876 224924
rect 272576 224884 272582 224896
rect 309870 224884 309876 224896
rect 309928 224884 309934 224936
rect 319806 224884 319812 224936
rect 319864 224924 319870 224936
rect 345934 224924 345940 224936
rect 319864 224896 345940 224924
rect 319864 224884 319870 224896
rect 345934 224884 345940 224896
rect 345992 224884 345998 224936
rect 460566 224884 460572 224936
rect 460624 224924 460630 224936
rect 463142 224924 463148 224936
rect 460624 224896 463148 224924
rect 460624 224884 460630 224896
rect 463142 224884 463148 224896
rect 463200 224884 463206 224936
rect 519354 224884 519360 224936
rect 519412 224924 519418 224936
rect 534994 224924 535000 224936
rect 519412 224896 535000 224924
rect 519412 224884 519418 224896
rect 534994 224884 535000 224896
rect 535052 224924 535058 224936
rect 621014 224924 621020 224936
rect 535052 224896 621020 224924
rect 535052 224884 535058 224896
rect 621014 224884 621020 224896
rect 621072 224884 621078 224936
rect 350350 224816 350356 224868
rect 350408 224856 350414 224868
rect 354950 224856 354956 224868
rect 350408 224828 354956 224856
rect 350408 224816 350414 224828
rect 354950 224816 354956 224828
rect 355008 224816 355014 224868
rect 670694 224816 670700 224868
rect 670752 224856 670758 224868
rect 670752 224828 671846 224856
rect 670752 224816 670758 224828
rect 232590 224788 232596 224800
rect 178696 224760 232596 224788
rect 232590 224748 232596 224760
rect 232648 224748 232654 224800
rect 245470 224748 245476 224800
rect 245528 224788 245534 224800
rect 287698 224788 287704 224800
rect 245528 224760 287704 224788
rect 245528 224748 245534 224760
rect 287698 224748 287704 224760
rect 287756 224748 287762 224800
rect 311526 224748 311532 224800
rect 311584 224788 311590 224800
rect 338850 224788 338856 224800
rect 311584 224760 338856 224788
rect 311584 224748 311590 224760
rect 338850 224748 338856 224760
rect 338908 224748 338914 224800
rect 462498 224748 462504 224800
rect 462556 224788 462562 224800
rect 469306 224788 469312 224800
rect 462556 224760 469312 224788
rect 462556 224748 462562 224760
rect 469306 224748 469312 224760
rect 469364 224748 469370 224800
rect 506934 224748 506940 224800
rect 506992 224788 506998 224800
rect 526346 224788 526352 224800
rect 506992 224760 526352 224788
rect 506992 224748 506998 224760
rect 526346 224748 526352 224760
rect 526404 224748 526410 224800
rect 529934 224748 529940 224800
rect 529992 224788 529998 224800
rect 542998 224788 543004 224800
rect 529992 224760 543004 224788
rect 529992 224748 529998 224760
rect 542998 224748 543004 224760
rect 543056 224748 543062 224800
rect 543182 224748 543188 224800
rect 543240 224788 543246 224800
rect 548610 224788 548616 224800
rect 543240 224760 548616 224788
rect 543240 224748 543246 224760
rect 548610 224748 548616 224760
rect 548668 224748 548674 224800
rect 548978 224748 548984 224800
rect 549036 224788 549042 224800
rect 549990 224788 549996 224800
rect 549036 224760 549996 224788
rect 549036 224748 549042 224760
rect 549990 224748 549996 224760
rect 550048 224788 550054 224800
rect 550048 224760 553394 224788
rect 550048 224748 550054 224760
rect 85482 224612 85488 224664
rect 85540 224652 85546 224664
rect 165614 224652 165620 224664
rect 85540 224624 165620 224652
rect 85540 224612 85546 224624
rect 165614 224612 165620 224624
rect 165672 224612 165678 224664
rect 171778 224652 171784 224664
rect 165908 224624 171784 224652
rect 79962 224476 79968 224528
rect 80020 224516 80026 224528
rect 160462 224516 160468 224528
rect 80020 224488 160468 224516
rect 80020 224476 80026 224488
rect 160462 224476 160468 224488
rect 160520 224476 160526 224528
rect 165522 224476 165528 224528
rect 165580 224516 165586 224528
rect 165908 224516 165936 224624
rect 171778 224612 171784 224624
rect 171836 224612 171842 224664
rect 171962 224612 171968 224664
rect 172020 224652 172026 224664
rect 185394 224652 185400 224664
rect 172020 224624 185400 224652
rect 172020 224612 172026 224624
rect 185394 224612 185400 224624
rect 185452 224612 185458 224664
rect 185578 224612 185584 224664
rect 185636 224652 185642 224664
rect 237742 224652 237748 224664
rect 185636 224624 237748 224652
rect 185636 224612 185642 224624
rect 237742 224612 237748 224624
rect 237800 224612 237806 224664
rect 248322 224612 248328 224664
rect 248380 224652 248386 224664
rect 291838 224652 291844 224664
rect 248380 224624 291844 224652
rect 248380 224612 248386 224624
rect 291838 224612 291844 224624
rect 291896 224612 291902 224664
rect 294874 224612 294880 224664
rect 294932 224652 294938 224664
rect 325970 224652 325976 224664
rect 294932 224624 325976 224652
rect 294932 224612 294938 224624
rect 325970 224612 325976 224624
rect 326028 224612 326034 224664
rect 346302 224612 346308 224664
rect 346360 224652 346366 224664
rect 366542 224652 366548 224664
rect 346360 224624 366548 224652
rect 346360 224612 346366 224624
rect 366542 224612 366548 224624
rect 366600 224612 366606 224664
rect 494054 224612 494060 224664
rect 494112 224652 494118 224664
rect 510154 224652 510160 224664
rect 494112 224624 510160 224652
rect 494112 224612 494118 224624
rect 510154 224612 510160 224624
rect 510212 224612 510218 224664
rect 520458 224612 520464 224664
rect 520516 224652 520522 224664
rect 544562 224652 544568 224664
rect 520516 224624 544568 224652
rect 520516 224612 520522 224624
rect 544562 224612 544568 224624
rect 544620 224612 544626 224664
rect 548058 224612 548064 224664
rect 548116 224652 548122 224664
rect 550634 224652 550640 224664
rect 548116 224624 550640 224652
rect 548116 224612 548122 224624
rect 550634 224612 550640 224624
rect 550692 224612 550698 224664
rect 553366 224652 553394 224760
rect 554958 224748 554964 224800
rect 555016 224788 555022 224800
rect 555970 224788 555976 224800
rect 555016 224760 555976 224788
rect 555016 224748 555022 224760
rect 555970 224748 555976 224760
rect 556028 224788 556034 224800
rect 557258 224788 557264 224800
rect 556028 224760 557264 224788
rect 556028 224748 556034 224760
rect 557258 224748 557264 224760
rect 557316 224748 557322 224800
rect 557442 224748 557448 224800
rect 557500 224788 557506 224800
rect 557500 224760 558316 224788
rect 557500 224748 557506 224760
rect 558288 224652 558316 224760
rect 558546 224748 558552 224800
rect 558604 224788 558610 224800
rect 561398 224788 561404 224800
rect 558604 224760 561404 224788
rect 558604 224748 558610 224760
rect 561398 224748 561404 224760
rect 561456 224748 561462 224800
rect 562686 224748 562692 224800
rect 562744 224788 562750 224800
rect 571702 224788 571708 224800
rect 562744 224760 571708 224788
rect 562744 224748 562750 224760
rect 571702 224748 571708 224760
rect 571760 224748 571766 224800
rect 670896 224692 671384 224720
rect 626534 224652 626540 224664
rect 553366 224624 558224 224652
rect 558288 224624 626540 224652
rect 224862 224516 224868 224528
rect 165580 224488 165936 224516
rect 166000 224488 224868 224516
rect 165580 224476 165586 224488
rect 73706 224340 73712 224392
rect 73764 224380 73770 224392
rect 155310 224380 155316 224392
rect 73764 224352 155316 224380
rect 73764 224340 73770 224352
rect 155310 224340 155316 224352
rect 155368 224340 155374 224392
rect 157242 224340 157248 224392
rect 157300 224380 157306 224392
rect 157978 224380 157984 224392
rect 157300 224352 157984 224380
rect 157300 224340 157306 224352
rect 157978 224340 157984 224352
rect 158036 224340 158042 224392
rect 162762 224340 162768 224392
rect 162820 224380 162826 224392
rect 166000 224380 166028 224488
rect 224862 224476 224868 224488
rect 224920 224476 224926 224528
rect 228726 224476 228732 224528
rect 228784 224516 228790 224528
rect 274910 224516 274916 224528
rect 228784 224488 274916 224516
rect 228784 224476 228790 224488
rect 274910 224476 274916 224488
rect 274968 224476 274974 224528
rect 275094 224476 275100 224528
rect 275152 224516 275158 224528
rect 311158 224516 311164 224528
rect 275152 224488 311164 224516
rect 275152 224476 275158 224488
rect 311158 224476 311164 224488
rect 311216 224476 311222 224528
rect 322842 224476 322848 224528
rect 322900 224516 322906 224528
rect 349798 224516 349804 224528
rect 322900 224488 349804 224516
rect 322900 224476 322906 224488
rect 349798 224476 349804 224488
rect 349856 224476 349862 224528
rect 359458 224476 359464 224528
rect 359516 224516 359522 224528
rect 378134 224516 378140 224528
rect 359516 224488 378140 224516
rect 359516 224476 359522 224488
rect 378134 224476 378140 224488
rect 378192 224476 378198 224528
rect 379238 224476 379244 224528
rect 379296 224516 379302 224528
rect 393590 224516 393596 224528
rect 379296 224488 393596 224516
rect 379296 224476 379302 224488
rect 393590 224476 393596 224488
rect 393648 224476 393654 224528
rect 456058 224476 456064 224528
rect 456116 224516 456122 224528
rect 459738 224516 459744 224528
rect 456116 224488 459744 224516
rect 456116 224476 456122 224488
rect 459738 224476 459744 224488
rect 459796 224476 459802 224528
rect 491294 224476 491300 224528
rect 491352 224516 491358 224528
rect 506014 224516 506020 224528
rect 491352 224488 506020 224516
rect 491352 224476 491358 224488
rect 506014 224476 506020 224488
rect 506072 224476 506078 224528
rect 515950 224476 515956 224528
rect 516008 224516 516014 224528
rect 539502 224516 539508 224528
rect 516008 224488 539508 224516
rect 516008 224476 516014 224488
rect 539502 224476 539508 224488
rect 539560 224476 539566 224528
rect 542998 224476 543004 224528
rect 543056 224516 543062 224528
rect 548978 224516 548984 224528
rect 543056 224488 548984 224516
rect 543056 224476 543062 224488
rect 548978 224476 548984 224488
rect 549036 224476 549042 224528
rect 549254 224476 549260 224528
rect 549312 224516 549318 224528
rect 555786 224516 555792 224528
rect 549312 224488 555792 224516
rect 549312 224476 549318 224488
rect 555786 224476 555792 224488
rect 555844 224476 555850 224528
rect 558196 224516 558224 224624
rect 626534 224612 626540 224624
rect 626592 224612 626598 224664
rect 562594 224516 562600 224528
rect 555988 224488 557580 224516
rect 558196 224488 562600 224516
rect 162820 224352 166028 224380
rect 162820 224340 162826 224352
rect 166166 224340 166172 224392
rect 166224 224380 166230 224392
rect 166224 224352 166994 224380
rect 166224 224340 166230 224352
rect 68922 224204 68928 224256
rect 68980 224244 68986 224256
rect 152734 224244 152740 224256
rect 68980 224216 152740 224244
rect 68980 224204 68986 224216
rect 152734 224204 152740 224216
rect 152792 224204 152798 224256
rect 155862 224204 155868 224256
rect 155920 224244 155926 224256
rect 160186 224244 160192 224256
rect 155920 224216 160192 224244
rect 155920 224204 155926 224216
rect 160186 224204 160192 224216
rect 160244 224204 160250 224256
rect 166966 224244 166994 224352
rect 168006 224340 168012 224392
rect 168064 224380 168070 224392
rect 171548 224380 171554 224392
rect 168064 224352 171554 224380
rect 168064 224340 168070 224352
rect 171548 224340 171554 224352
rect 171606 224340 171612 224392
rect 172146 224340 172152 224392
rect 172204 224380 172210 224392
rect 227438 224380 227444 224392
rect 172204 224352 227444 224380
rect 172204 224340 172210 224352
rect 227438 224340 227444 224352
rect 227496 224340 227502 224392
rect 233142 224340 233148 224392
rect 233200 224380 233206 224392
rect 277670 224380 277676 224392
rect 233200 224352 277676 224380
rect 233200 224340 233206 224352
rect 277670 224340 277676 224352
rect 277728 224340 277734 224392
rect 286318 224340 286324 224392
rect 286376 224380 286382 224392
rect 289906 224380 289912 224392
rect 286376 224352 289912 224380
rect 286376 224340 286382 224352
rect 289906 224340 289912 224352
rect 289964 224340 289970 224392
rect 290826 224340 290832 224392
rect 290884 224380 290890 224392
rect 324038 224380 324044 224392
rect 290884 224352 324044 224380
rect 290884 224340 290890 224352
rect 324038 224340 324044 224352
rect 324096 224340 324102 224392
rect 342162 224340 342168 224392
rect 342220 224380 342226 224392
rect 362034 224380 362040 224392
rect 342220 224352 362040 224380
rect 342220 224340 342226 224352
rect 362034 224340 362040 224352
rect 362092 224340 362098 224392
rect 366726 224340 366732 224392
rect 366784 224380 366790 224392
rect 381630 224380 381636 224392
rect 366784 224352 381636 224380
rect 366784 224340 366790 224352
rect 381630 224340 381636 224352
rect 381688 224340 381694 224392
rect 394510 224340 394516 224392
rect 394568 224380 394574 224392
rect 404538 224380 404544 224392
rect 394568 224352 404544 224380
rect 394568 224340 394574 224352
rect 404538 224340 404544 224352
rect 404596 224340 404602 224392
rect 480530 224340 480536 224392
rect 480588 224380 480594 224392
rect 492858 224380 492864 224392
rect 480588 224352 492864 224380
rect 480588 224340 480594 224352
rect 492858 224340 492864 224352
rect 492916 224340 492922 224392
rect 499206 224340 499212 224392
rect 499264 224380 499270 224392
rect 516594 224380 516600 224392
rect 499264 224352 516600 224380
rect 499264 224340 499270 224352
rect 516594 224340 516600 224352
rect 516652 224340 516658 224392
rect 525610 224340 525616 224392
rect 525668 224380 525674 224392
rect 548058 224380 548064 224392
rect 525668 224352 548064 224380
rect 525668 224340 525674 224352
rect 548058 224340 548064 224352
rect 548116 224340 548122 224392
rect 548610 224340 548616 224392
rect 548668 224380 548674 224392
rect 555988 224380 556016 224488
rect 548668 224352 556016 224380
rect 548668 224340 548674 224352
rect 556154 224340 556160 224392
rect 556212 224380 556218 224392
rect 557350 224380 557356 224392
rect 556212 224352 557356 224380
rect 556212 224340 556218 224352
rect 557350 224340 557356 224352
rect 557408 224340 557414 224392
rect 557552 224380 557580 224488
rect 562594 224476 562600 224488
rect 562652 224476 562658 224528
rect 563146 224476 563152 224528
rect 563204 224516 563210 224528
rect 625246 224516 625252 224528
rect 563204 224488 625252 224516
rect 563204 224476 563210 224488
rect 625246 224476 625252 224488
rect 625304 224476 625310 224528
rect 562778 224380 562784 224392
rect 557552 224352 562784 224380
rect 562778 224340 562784 224352
rect 562836 224340 562842 224392
rect 625982 224380 625988 224392
rect 572686 224352 625988 224380
rect 565170 224272 565176 224324
rect 565228 224312 565234 224324
rect 572686 224312 572714 224352
rect 625982 224340 625988 224352
rect 626040 224340 626046 224392
rect 667014 224340 667020 224392
rect 667072 224380 667078 224392
rect 670896 224380 670924 224692
rect 671356 224584 671384 224692
rect 671476 224612 671482 224664
rect 671534 224652 671540 224664
rect 671534 224624 671738 224652
rect 671534 224612 671540 224624
rect 671356 224556 671412 224584
rect 671384 224516 671412 224556
rect 671384 224488 671476 224516
rect 671448 224448 671476 224488
rect 671448 224420 671622 224448
rect 667072 224352 670924 224380
rect 667072 224340 667078 224352
rect 565228 224284 572714 224312
rect 565228 224272 565234 224284
rect 171962 224244 171968 224256
rect 166966 224216 171968 224244
rect 171962 224204 171968 224216
rect 172020 224204 172026 224256
rect 172146 224204 172152 224256
rect 172204 224244 172210 224256
rect 176286 224244 176292 224256
rect 172204 224216 176292 224244
rect 172204 224204 172210 224216
rect 176286 224204 176292 224216
rect 176344 224204 176350 224256
rect 230014 224244 230020 224256
rect 176626 224216 230020 224244
rect 102042 224068 102048 224120
rect 102100 224108 102106 224120
rect 170858 224108 170864 224120
rect 102100 224080 170864 224108
rect 102100 224068 102106 224080
rect 170858 224068 170864 224080
rect 170916 224068 170922 224120
rect 171778 224068 171784 224120
rect 171836 224108 171842 224120
rect 176626 224108 176654 224216
rect 230014 224204 230020 224216
rect 230072 224204 230078 224256
rect 231670 224204 231676 224256
rect 231728 224244 231734 224256
rect 278958 224244 278964 224256
rect 231728 224216 278964 224244
rect 231728 224204 231734 224216
rect 278958 224204 278964 224216
rect 279016 224204 279022 224256
rect 289630 224204 289636 224256
rect 289688 224244 289694 224256
rect 296990 224244 296996 224256
rect 289688 224216 296996 224244
rect 289688 224204 289694 224216
rect 296990 224204 296996 224216
rect 297048 224204 297054 224256
rect 299106 224204 299112 224256
rect 299164 224244 299170 224256
rect 331766 224244 331772 224256
rect 299164 224216 331772 224244
rect 299164 224204 299170 224216
rect 331766 224204 331772 224216
rect 331824 224204 331830 224256
rect 339402 224204 339408 224256
rect 339460 224244 339466 224256
rect 362310 224244 362316 224256
rect 339460 224216 362316 224244
rect 339460 224204 339466 224216
rect 362310 224204 362316 224216
rect 362368 224204 362374 224256
rect 372522 224204 372528 224256
rect 372580 224244 372586 224256
rect 387426 224244 387432 224256
rect 372580 224216 387432 224244
rect 372580 224204 372586 224216
rect 387426 224204 387432 224216
rect 387484 224204 387490 224256
rect 390186 224204 390192 224256
rect 390244 224244 390250 224256
rect 401962 224244 401968 224256
rect 390244 224216 401968 224244
rect 390244 224204 390250 224216
rect 401962 224204 401968 224216
rect 402020 224204 402026 224256
rect 405550 224204 405556 224256
rect 405608 224244 405614 224256
rect 414198 224244 414204 224256
rect 405608 224216 414204 224244
rect 405608 224204 405614 224216
rect 414198 224204 414204 224216
rect 414256 224204 414262 224256
rect 470226 224204 470232 224256
rect 470284 224244 470290 224256
rect 480346 224244 480352 224256
rect 470284 224216 480352 224244
rect 470284 224204 470290 224216
rect 480346 224204 480352 224216
rect 480404 224204 480410 224256
rect 483750 224204 483756 224256
rect 483808 224244 483814 224256
rect 496906 224244 496912 224256
rect 483808 224216 496912 224244
rect 483808 224204 483814 224216
rect 496906 224204 496912 224216
rect 496964 224204 496970 224256
rect 523494 224244 523500 224256
rect 505066 224216 523500 224244
rect 171836 224080 176654 224108
rect 171836 224068 171842 224080
rect 177482 224068 177488 224120
rect 177540 224108 177546 224120
rect 177540 224080 185256 224108
rect 177540 224068 177546 224080
rect 105998 223932 106004 223984
rect 106056 223972 106062 223984
rect 181070 223972 181076 223984
rect 106056 223944 181076 223972
rect 106056 223932 106062 223944
rect 181070 223932 181076 223944
rect 181128 223932 181134 223984
rect 185228 223972 185256 224080
rect 185394 224068 185400 224120
rect 185452 224108 185458 224120
rect 194594 224108 194600 224120
rect 185452 224080 194600 224108
rect 185452 224068 185458 224080
rect 194594 224068 194600 224080
rect 194652 224068 194658 224120
rect 195882 224068 195888 224120
rect 195940 224108 195946 224120
rect 250622 224108 250628 224120
rect 195940 224080 250628 224108
rect 195940 224068 195946 224080
rect 250622 224068 250628 224080
rect 250680 224068 250686 224120
rect 266262 224068 266268 224120
rect 266320 224108 266326 224120
rect 303430 224108 303436 224120
rect 266320 224080 303436 224108
rect 266320 224068 266326 224080
rect 303430 224068 303436 224080
rect 303488 224068 303494 224120
rect 304258 224068 304264 224120
rect 304316 224108 304322 224120
rect 315298 224108 315304 224120
rect 304316 224080 315304 224108
rect 304316 224068 304322 224080
rect 315298 224068 315304 224080
rect 315356 224068 315362 224120
rect 504358 224068 504364 224120
rect 504416 224108 504422 224120
rect 505066 224108 505094 224216
rect 523494 224204 523500 224216
rect 523552 224204 523558 224256
rect 535270 224204 535276 224256
rect 535328 224244 535334 224256
rect 562686 224244 562692 224256
rect 535328 224216 562692 224244
rect 535328 224204 535334 224216
rect 562686 224204 562692 224216
rect 562744 224204 562750 224256
rect 671172 224216 671508 224244
rect 562870 224136 562876 224188
rect 562928 224176 562934 224188
rect 610434 224176 610440 224188
rect 562928 224148 610440 224176
rect 562928 224136 562934 224148
rect 610434 224136 610440 224148
rect 610492 224136 610498 224188
rect 610618 224136 610624 224188
rect 610676 224176 610682 224188
rect 617058 224176 617064 224188
rect 610676 224148 617064 224176
rect 610676 224136 610682 224148
rect 617058 224136 617064 224148
rect 617116 224136 617122 224188
rect 670786 224136 670792 224188
rect 670844 224176 670850 224188
rect 671172 224176 671200 224216
rect 670844 224148 671200 224176
rect 670844 224136 670850 224148
rect 504416 224080 505094 224108
rect 504416 224068 504422 224080
rect 524414 224000 524420 224052
rect 524472 224040 524478 224052
rect 525058 224040 525064 224052
rect 524472 224012 525064 224040
rect 524472 224000 524478 224012
rect 525058 224000 525064 224012
rect 525116 224040 525122 224052
rect 619634 224040 619640 224052
rect 525116 224012 619640 224040
rect 525116 224000 525122 224012
rect 619634 224000 619640 224012
rect 619692 224000 619698 224052
rect 666830 224000 666836 224052
rect 666888 224040 666894 224052
rect 666888 224012 671398 224040
rect 666888 224000 666894 224012
rect 185762 223972 185768 223984
rect 185228 223944 185768 223972
rect 185762 223932 185768 223944
rect 185820 223932 185826 223984
rect 191558 223932 191564 223984
rect 191616 223972 191622 223984
rect 199838 223972 199844 223984
rect 191616 223944 199844 223972
rect 191616 223932 191622 223944
rect 199838 223932 199844 223944
rect 199896 223932 199902 223984
rect 201402 223932 201408 223984
rect 201460 223972 201466 223984
rect 255774 223972 255780 223984
rect 201460 223944 255780 223972
rect 201460 223932 201466 223944
rect 255774 223932 255780 223944
rect 255832 223932 255838 223984
rect 331858 223932 331864 223984
rect 331916 223972 331922 223984
rect 337562 223972 337568 223984
rect 331916 223944 337568 223972
rect 331916 223932 331922 223944
rect 337562 223932 337568 223944
rect 337620 223932 337626 223984
rect 279418 223864 279424 223916
rect 279476 223904 279482 223916
rect 284754 223904 284760 223916
rect 279476 223876 284760 223904
rect 279476 223864 279482 223876
rect 284754 223864 284760 223876
rect 284812 223864 284818 223916
rect 517698 223864 517704 223916
rect 517756 223904 517762 223916
rect 610618 223904 610624 223916
rect 517756 223876 610624 223904
rect 517756 223864 517762 223876
rect 610618 223864 610624 223876
rect 610676 223864 610682 223916
rect 610802 223864 610808 223916
rect 610860 223904 610866 223916
rect 622486 223904 622492 223916
rect 610860 223876 622492 223904
rect 610860 223864 610866 223876
rect 622486 223864 622492 223876
rect 622544 223864 622550 223916
rect 108666 223796 108672 223848
rect 108724 223836 108730 223848
rect 183830 223836 183836 223848
rect 108724 223808 183836 223836
rect 108724 223796 108730 223808
rect 183830 223796 183836 223808
rect 183888 223796 183894 223848
rect 184382 223796 184388 223848
rect 184440 223836 184446 223848
rect 207474 223836 207480 223848
rect 184440 223808 207480 223836
rect 184440 223796 184446 223808
rect 207474 223796 207480 223808
rect 207532 223796 207538 223848
rect 227530 223796 227536 223848
rect 227588 223836 227594 223848
rect 273162 223836 273168 223848
rect 227588 223808 273168 223836
rect 227588 223796 227594 223808
rect 273162 223796 273168 223808
rect 273220 223796 273226 223848
rect 670712 223808 671278 223836
rect 505094 223728 505100 223780
rect 505152 223768 505158 223780
rect 507670 223768 507676 223780
rect 505152 223740 507676 223768
rect 505152 223728 505158 223740
rect 507670 223728 507676 223740
rect 507728 223728 507734 223780
rect 539962 223728 539968 223780
rect 540020 223768 540026 223780
rect 622670 223768 622676 223780
rect 540020 223740 622676 223768
rect 540020 223728 540026 223740
rect 622670 223728 622676 223740
rect 622728 223728 622734 223780
rect 667014 223728 667020 223780
rect 667072 223768 667078 223780
rect 670712 223768 670740 223808
rect 667072 223740 670740 223768
rect 667072 223728 667078 223740
rect 115290 223660 115296 223712
rect 115348 223700 115354 223712
rect 188798 223700 188804 223712
rect 115348 223672 188804 223700
rect 115348 223660 115354 223672
rect 188798 223660 188804 223672
rect 188856 223660 188862 223712
rect 207658 223660 207664 223712
rect 207716 223700 207722 223712
rect 228082 223700 228088 223712
rect 207716 223672 228088 223700
rect 207716 223660 207722 223672
rect 228082 223660 228088 223672
rect 228140 223660 228146 223712
rect 505278 223592 505284 223644
rect 505336 223632 505342 223644
rect 614942 223632 614948 223644
rect 505336 223604 614948 223632
rect 505336 223592 505342 223604
rect 614942 223592 614948 223604
rect 615000 223592 615006 223644
rect 670786 223592 670792 223644
rect 670844 223632 670850 223644
rect 670844 223604 671186 223632
rect 670844 223592 670850 223604
rect 87966 223524 87972 223576
rect 88024 223564 88030 223576
rect 164970 223564 164976 223576
rect 88024 223536 164976 223564
rect 88024 223524 88030 223536
rect 164970 223524 164976 223536
rect 165028 223524 165034 223576
rect 171778 223524 171784 223576
rect 171836 223564 171842 223576
rect 181714 223564 181720 223576
rect 171836 223536 181720 223564
rect 171836 223524 171842 223536
rect 181714 223524 181720 223536
rect 181772 223524 181778 223576
rect 183186 223524 183192 223576
rect 183244 223564 183250 223576
rect 184658 223564 184664 223576
rect 183244 223536 184664 223564
rect 183244 223524 183250 223536
rect 184658 223524 184664 223536
rect 184716 223524 184722 223576
rect 184842 223524 184848 223576
rect 184900 223564 184906 223576
rect 239674 223564 239680 223576
rect 184900 223536 239680 223564
rect 184900 223524 184906 223536
rect 239674 223524 239680 223536
rect 239732 223524 239738 223576
rect 249426 223524 249432 223576
rect 249484 223564 249490 223576
rect 276290 223564 276296 223576
rect 249484 223536 276296 223564
rect 249484 223524 249490 223536
rect 276290 223524 276296 223536
rect 276348 223524 276354 223576
rect 278590 223524 278596 223576
rect 278648 223564 278654 223576
rect 315022 223564 315028 223576
rect 278648 223536 315028 223564
rect 278648 223524 278654 223536
rect 315022 223524 315028 223536
rect 315080 223524 315086 223576
rect 406746 223524 406752 223576
rect 406804 223564 406810 223576
rect 414842 223564 414848 223576
rect 406804 223536 414848 223564
rect 406804 223524 406810 223536
rect 414842 223524 414848 223536
rect 414900 223524 414906 223576
rect 454862 223524 454868 223576
rect 454920 223564 454926 223576
rect 460474 223564 460480 223576
rect 454920 223536 460480 223564
rect 454920 223524 454926 223536
rect 460474 223524 460480 223536
rect 460532 223524 460538 223576
rect 473446 223524 473452 223576
rect 473504 223564 473510 223576
rect 475562 223564 475568 223576
rect 473504 223536 475568 223564
rect 473504 223524 473510 223536
rect 475562 223524 475568 223536
rect 475620 223524 475626 223576
rect 670804 223468 671048 223496
rect 99282 223388 99288 223440
rect 99340 223428 99346 223440
rect 176010 223428 176016 223440
rect 99340 223400 176016 223428
rect 99340 223388 99346 223400
rect 176010 223388 176016 223400
rect 176068 223388 176074 223440
rect 187326 223388 187332 223440
rect 187384 223428 187390 223440
rect 242250 223428 242256 223440
rect 187384 223400 242256 223428
rect 187384 223388 187390 223400
rect 242250 223388 242256 223400
rect 242308 223388 242314 223440
rect 244090 223388 244096 223440
rect 244148 223428 244154 223440
rect 286042 223428 286048 223440
rect 244148 223400 286048 223428
rect 244148 223388 244154 223400
rect 286042 223388 286048 223400
rect 286100 223388 286106 223440
rect 291194 223428 291200 223440
rect 287026 223400 291200 223428
rect 81342 223252 81348 223304
rect 81400 223292 81406 223304
rect 151906 223292 151912 223304
rect 81400 223264 151912 223292
rect 81400 223252 81406 223264
rect 151906 223252 151912 223264
rect 151964 223252 151970 223304
rect 156414 223292 156420 223304
rect 152108 223264 156420 223292
rect 68738 223116 68744 223168
rect 68796 223156 68802 223168
rect 146478 223156 146484 223168
rect 68796 223128 146484 223156
rect 68796 223116 68802 223128
rect 146478 223116 146484 223128
rect 146536 223116 146542 223168
rect 146662 223116 146668 223168
rect 146720 223156 146726 223168
rect 152108 223156 152136 223264
rect 156414 223252 156420 223264
rect 156472 223252 156478 223304
rect 156598 223252 156604 223304
rect 156656 223292 156662 223304
rect 161934 223292 161940 223304
rect 156656 223264 161940 223292
rect 156656 223252 156662 223264
rect 161934 223252 161940 223264
rect 161992 223252 161998 223304
rect 162118 223252 162124 223304
rect 162176 223292 162182 223304
rect 186866 223292 186872 223304
rect 162176 223264 186872 223292
rect 162176 223252 162182 223264
rect 186866 223252 186872 223264
rect 186924 223252 186930 223304
rect 188890 223252 188896 223304
rect 188948 223292 188954 223304
rect 245102 223292 245108 223304
rect 188948 223264 245108 223292
rect 188948 223252 188954 223264
rect 245102 223252 245108 223264
rect 245160 223252 245166 223304
rect 250898 223252 250904 223304
rect 250956 223292 250962 223304
rect 287026 223292 287054 223400
rect 291194 223388 291200 223400
rect 291252 223388 291258 223440
rect 316678 223388 316684 223440
rect 316736 223428 316742 223440
rect 327258 223428 327264 223440
rect 316736 223400 327264 223428
rect 316736 223388 316742 223400
rect 327258 223388 327264 223400
rect 327316 223388 327322 223440
rect 517514 223388 517520 223440
rect 517572 223428 517578 223440
rect 532510 223428 532516 223440
rect 517572 223400 532516 223428
rect 517572 223388 517578 223400
rect 532510 223388 532516 223400
rect 532568 223388 532574 223440
rect 534810 223388 534816 223440
rect 534868 223428 534874 223440
rect 547414 223428 547420 223440
rect 534868 223400 547420 223428
rect 534868 223388 534874 223400
rect 547414 223388 547420 223400
rect 547472 223388 547478 223440
rect 297542 223320 297548 223372
rect 297600 223360 297606 223372
rect 305362 223360 305368 223372
rect 297600 223332 305368 223360
rect 297600 223320 297606 223332
rect 305362 223320 305368 223332
rect 305420 223320 305426 223372
rect 670804 223360 670832 223468
rect 670620 223332 670832 223360
rect 250956 223264 287054 223292
rect 250956 223252 250962 223264
rect 288986 223252 288992 223304
rect 289044 223292 289050 223304
rect 295058 223292 295064 223304
rect 289044 223264 295064 223292
rect 289044 223252 289050 223264
rect 295058 223252 295064 223264
rect 295116 223252 295122 223304
rect 307662 223252 307668 223304
rect 307720 223292 307726 223304
rect 335630 223292 335636 223304
rect 307720 223264 335636 223292
rect 307720 223252 307726 223264
rect 335630 223252 335636 223264
rect 335688 223252 335694 223304
rect 337930 223252 337936 223304
rect 337988 223292 337994 223304
rect 359182 223292 359188 223304
rect 337988 223264 359188 223292
rect 337988 223252 337994 223264
rect 359182 223252 359188 223264
rect 359240 223252 359246 223304
rect 493042 223252 493048 223304
rect 493100 223292 493106 223304
rect 508498 223292 508504 223304
rect 493100 223264 508504 223292
rect 493100 223252 493106 223264
rect 508498 223252 508504 223264
rect 508556 223252 508562 223304
rect 514662 223252 514668 223304
rect 514720 223292 514726 223304
rect 535454 223292 535460 223304
rect 514720 223264 535460 223292
rect 514720 223252 514726 223264
rect 535454 223252 535460 223264
rect 535512 223252 535518 223304
rect 154942 223156 154948 223168
rect 146720 223128 152136 223156
rect 152200 223128 154948 223156
rect 146720 223116 146726 223128
rect 75822 222980 75828 223032
rect 75880 223020 75886 223032
rect 152200 223020 152228 223128
rect 154942 223116 154948 223128
rect 155000 223116 155006 223168
rect 156414 223116 156420 223168
rect 156472 223156 156478 223168
rect 176102 223156 176108 223168
rect 156472 223128 176108 223156
rect 156472 223116 156478 223128
rect 176102 223116 176108 223128
rect 176160 223116 176166 223168
rect 181990 223116 181996 223168
rect 182048 223156 182054 223168
rect 240318 223156 240324 223168
rect 182048 223128 240324 223156
rect 182048 223116 182054 223128
rect 240318 223116 240324 223128
rect 240376 223116 240382 223168
rect 241330 223116 241336 223168
rect 241388 223156 241394 223168
rect 283466 223156 283472 223168
rect 241388 223128 283472 223156
rect 241388 223116 241394 223128
rect 283466 223116 283472 223128
rect 283524 223116 283530 223168
rect 288250 223116 288256 223168
rect 288308 223156 288314 223168
rect 321462 223156 321468 223168
rect 288308 223128 321468 223156
rect 288308 223116 288314 223128
rect 321462 223116 321468 223128
rect 321520 223116 321526 223168
rect 323946 223116 323952 223168
rect 324004 223156 324010 223168
rect 348510 223156 348516 223168
rect 324004 223128 348516 223156
rect 324004 223116 324010 223128
rect 348510 223116 348516 223128
rect 348568 223116 348574 223168
rect 358538 223116 358544 223168
rect 358596 223156 358602 223168
rect 374638 223156 374644 223168
rect 358596 223128 374644 223156
rect 358596 223116 358602 223128
rect 374638 223116 374644 223128
rect 374696 223116 374702 223168
rect 483106 223116 483112 223168
rect 483164 223156 483170 223168
rect 496078 223156 496084 223168
rect 483164 223128 496084 223156
rect 483164 223116 483170 223128
rect 496078 223116 496084 223128
rect 496136 223116 496142 223168
rect 503346 223116 503352 223168
rect 503404 223156 503410 223168
rect 521746 223156 521752 223168
rect 503404 223128 521752 223156
rect 503404 223116 503410 223128
rect 521746 223116 521752 223128
rect 521804 223116 521810 223168
rect 529474 223116 529480 223168
rect 529532 223156 529538 223168
rect 555694 223156 555700 223168
rect 529532 223128 555700 223156
rect 529532 223116 529538 223128
rect 555694 223116 555700 223128
rect 555752 223116 555758 223168
rect 75880 222992 152228 223020
rect 75880 222980 75886 222992
rect 152366 222980 152372 223032
rect 152424 223020 152430 223032
rect 152424 222992 156920 223020
rect 152424 222980 152430 222992
rect 71406 222844 71412 222896
rect 71464 222884 71470 222896
rect 151630 222884 151636 222896
rect 71464 222856 151636 222884
rect 71464 222844 71470 222856
rect 151630 222844 151636 222856
rect 151688 222844 151694 222896
rect 151768 222844 151774 222896
rect 151826 222884 151832 222896
rect 156414 222884 156420 222896
rect 151826 222856 156420 222884
rect 151826 222844 151832 222856
rect 156414 222844 156420 222856
rect 156472 222844 156478 222896
rect 156892 222884 156920 222992
rect 158070 222980 158076 223032
rect 158128 223020 158134 223032
rect 219066 223020 219072 223032
rect 158128 222992 219072 223020
rect 158128 222980 158134 222992
rect 219066 222980 219072 222992
rect 219124 222980 219130 223032
rect 245286 222980 245292 223032
rect 245344 223020 245350 223032
rect 289262 223020 289268 223032
rect 245344 222992 289268 223020
rect 245344 222980 245350 222992
rect 289262 222980 289268 222992
rect 289320 222980 289326 223032
rect 291654 222980 291660 223032
rect 291712 223020 291718 223032
rect 300210 223020 300216 223032
rect 291712 222992 300216 223020
rect 291712 222980 291718 222992
rect 300210 222980 300216 222992
rect 300268 222980 300274 223032
rect 315666 222980 315672 223032
rect 315724 223020 315730 223032
rect 344646 223020 344652 223032
rect 315724 222992 344652 223020
rect 315724 222980 315730 222992
rect 344646 222980 344652 222992
rect 344704 222980 344710 223032
rect 346578 223020 346584 223032
rect 344986 222992 346584 223020
rect 171778 222884 171784 222896
rect 156892 222856 171784 222884
rect 171778 222844 171784 222856
rect 171836 222844 171842 222896
rect 172882 222844 172888 222896
rect 172940 222884 172946 222896
rect 212626 222884 212632 222896
rect 172940 222856 212632 222884
rect 172940 222844 172946 222856
rect 212626 222844 212632 222856
rect 212684 222844 212690 222896
rect 213178 222844 213184 222896
rect 213236 222884 213242 222896
rect 233326 222884 233332 222896
rect 213236 222856 233332 222884
rect 213236 222844 213242 222856
rect 233326 222844 233332 222856
rect 233384 222844 233390 222896
rect 234522 222844 234528 222896
rect 234580 222884 234586 222896
rect 281534 222884 281540 222896
rect 234580 222856 281540 222884
rect 234580 222844 234586 222856
rect 281534 222844 281540 222856
rect 281592 222844 281598 222896
rect 282730 222844 282736 222896
rect 282788 222884 282794 222896
rect 316310 222884 316316 222896
rect 282788 222856 316316 222884
rect 282788 222844 282794 222856
rect 316310 222844 316316 222856
rect 316368 222844 316374 222896
rect 321462 222844 321468 222896
rect 321520 222884 321526 222896
rect 344986 222884 345014 222992
rect 346578 222980 346584 222992
rect 346636 222980 346642 223032
rect 349062 222980 349068 223032
rect 349120 223020 349126 223032
rect 367186 223020 367192 223032
rect 349120 222992 367192 223020
rect 349120 222980 349126 222992
rect 367186 222980 367192 222992
rect 367244 222980 367250 223032
rect 368382 222980 368388 223032
rect 368440 223020 368446 223032
rect 382642 223020 382648 223032
rect 368440 222992 382648 223020
rect 368440 222980 368446 222992
rect 382642 222980 382648 222992
rect 382700 222980 382706 223032
rect 383562 222980 383568 223032
rect 383620 223020 383626 223032
rect 394878 223020 394884 223032
rect 383620 222992 394884 223020
rect 383620 222980 383626 222992
rect 394878 222980 394884 222992
rect 394936 222980 394942 223032
rect 486602 222980 486608 223032
rect 486660 223020 486666 223032
rect 500034 223020 500040 223032
rect 486660 222992 500040 223020
rect 486660 222980 486666 222992
rect 500034 222980 500040 222992
rect 500092 222980 500098 223032
rect 508222 222980 508228 223032
rect 508280 223020 508286 223032
rect 527726 223020 527732 223032
rect 508280 222992 527732 223020
rect 508280 222980 508286 222992
rect 527726 222980 527732 222992
rect 527784 222980 527790 223032
rect 532050 222980 532056 223032
rect 532108 223020 532114 223032
rect 559006 223020 559012 223032
rect 532108 222992 559012 223020
rect 532108 222980 532114 222992
rect 559006 222980 559012 222992
rect 559064 222980 559070 223032
rect 670620 223020 670648 223332
rect 670786 223116 670792 223168
rect 670844 223156 670850 223168
rect 670844 223128 670956 223156
rect 670844 223116 670850 223128
rect 670620 222992 670832 223020
rect 321520 222856 345014 222884
rect 321520 222844 321526 222856
rect 345290 222844 345296 222896
rect 345348 222884 345354 222896
rect 347866 222884 347872 222896
rect 345348 222856 347872 222884
rect 345348 222844 345354 222856
rect 347866 222844 347872 222856
rect 347924 222844 347930 222896
rect 367830 222884 367836 222896
rect 354646 222856 367836 222884
rect 78582 222708 78588 222760
rect 78640 222748 78646 222760
rect 127618 222748 127624 222760
rect 78640 222720 127624 222748
rect 78640 222708 78646 222720
rect 127618 222708 127624 222720
rect 127676 222708 127682 222760
rect 127802 222708 127808 222760
rect 127860 222748 127866 222760
rect 191374 222748 191380 222760
rect 127860 222720 191380 222748
rect 127860 222708 127866 222720
rect 191374 222708 191380 222720
rect 191432 222708 191438 222760
rect 197170 222708 197176 222760
rect 197228 222748 197234 222760
rect 249978 222748 249984 222760
rect 197228 222720 249984 222748
rect 197228 222708 197234 222720
rect 249978 222708 249984 222720
rect 250036 222708 250042 222760
rect 284202 222708 284208 222760
rect 284260 222748 284266 222760
rect 316954 222748 316960 222760
rect 284260 222720 316960 222748
rect 284260 222708 284266 222720
rect 316954 222708 316960 222720
rect 317012 222708 317018 222760
rect 347222 222708 347228 222760
rect 347280 222748 347286 222760
rect 354646 222748 354674 222856
rect 367830 222844 367836 222856
rect 367888 222844 367894 222896
rect 375190 222844 375196 222896
rect 375248 222884 375254 222896
rect 391014 222884 391020 222896
rect 375248 222856 391020 222884
rect 375248 222844 375254 222856
rect 391014 222844 391020 222856
rect 391072 222844 391078 222896
rect 395798 222844 395804 222896
rect 395856 222884 395862 222896
rect 406470 222884 406476 222896
rect 395856 222856 406476 222884
rect 395856 222844 395862 222856
rect 406470 222844 406476 222856
rect 406528 222844 406534 222896
rect 420822 222844 420828 222896
rect 420880 222884 420886 222896
rect 425146 222884 425152 222896
rect 420880 222856 425152 222884
rect 420880 222844 420886 222856
rect 425146 222844 425152 222856
rect 425204 222844 425210 222896
rect 459922 222844 459928 222896
rect 459980 222884 459986 222896
rect 467098 222884 467104 222896
rect 459980 222856 467104 222884
rect 459980 222844 459986 222856
rect 467098 222844 467104 222856
rect 467156 222844 467162 222896
rect 467466 222844 467472 222896
rect 467524 222884 467530 222896
rect 473722 222884 473728 222896
rect 467524 222856 473728 222884
rect 467524 222844 467530 222856
rect 473722 222844 473728 222856
rect 473780 222844 473786 222896
rect 479886 222844 479892 222896
rect 479944 222884 479950 222896
rect 492030 222884 492036 222896
rect 479944 222856 492036 222884
rect 479944 222844 479950 222856
rect 492030 222844 492036 222856
rect 492088 222844 492094 222896
rect 500770 222844 500776 222896
rect 500828 222884 500834 222896
rect 517514 222884 517520 222896
rect 500828 222856 517520 222884
rect 500828 222844 500834 222856
rect 517514 222844 517520 222856
rect 517572 222844 517578 222896
rect 519814 222844 519820 222896
rect 519872 222884 519878 222896
rect 543366 222884 543372 222896
rect 519872 222856 543372 222884
rect 519872 222844 519878 222856
rect 543366 222844 543372 222856
rect 543424 222844 543430 222896
rect 554038 222844 554044 222896
rect 554096 222884 554102 222896
rect 632698 222884 632704 222896
rect 554096 222856 632704 222884
rect 554096 222844 554102 222856
rect 632698 222844 632704 222856
rect 632756 222844 632762 222896
rect 651282 222844 651288 222896
rect 651340 222884 651346 222896
rect 666462 222884 666468 222896
rect 651340 222856 666468 222884
rect 651340 222844 651346 222856
rect 666462 222844 666468 222856
rect 666520 222844 666526 222896
rect 347280 222720 354674 222748
rect 347280 222708 347286 222720
rect 532510 222708 532516 222760
rect 532568 222748 532574 222760
rect 542998 222748 543004 222760
rect 532568 222720 543004 222748
rect 532568 222708 532574 222720
rect 542998 222708 543004 222720
rect 543056 222708 543062 222760
rect 558178 222708 558184 222760
rect 558236 222748 558242 222760
rect 558236 222720 596174 222748
rect 558236 222708 558242 222720
rect 426434 222640 426440 222692
rect 426492 222680 426498 222692
rect 426986 222680 426992 222692
rect 426492 222652 426992 222680
rect 426492 222640 426498 222652
rect 426986 222640 426992 222652
rect 427044 222640 427050 222692
rect 85298 222572 85304 222624
rect 85356 222612 85362 222624
rect 156598 222612 156604 222624
rect 85356 222584 156604 222612
rect 85356 222572 85362 222584
rect 156598 222572 156604 222584
rect 156656 222572 156662 222624
rect 166350 222572 166356 222624
rect 166408 222612 166414 222624
rect 192018 222612 192024 222624
rect 166408 222584 192024 222612
rect 166408 222572 166414 222584
rect 192018 222572 192024 222584
rect 192076 222572 192082 222624
rect 194502 222572 194508 222624
rect 194560 222612 194566 222624
rect 247402 222612 247408 222624
rect 194560 222584 247408 222612
rect 194560 222572 194566 222584
rect 247402 222572 247408 222584
rect 247460 222572 247466 222624
rect 482738 222572 482744 222624
rect 482796 222612 482802 222624
rect 593966 222612 593972 222624
rect 482796 222584 593972 222612
rect 482796 222572 482802 222584
rect 593966 222572 593972 222584
rect 594024 222572 594030 222624
rect 596146 222612 596174 222720
rect 630674 222612 630680 222624
rect 596146 222584 630680 222612
rect 630674 222572 630680 222584
rect 630732 222572 630738 222624
rect 118418 222436 118424 222488
rect 118476 222476 118482 222488
rect 118476 222448 122834 222476
rect 118476 222436 118482 222448
rect 122806 222340 122834 222448
rect 127618 222436 127624 222488
rect 127676 222476 127682 222488
rect 146662 222476 146668 222488
rect 127676 222448 146668 222476
rect 127676 222436 127682 222448
rect 146662 222436 146668 222448
rect 146720 222436 146726 222488
rect 206830 222476 206836 222488
rect 146956 222448 206836 222476
rect 127802 222340 127808 222352
rect 122806 222312 127808 222340
rect 127802 222300 127808 222312
rect 127860 222300 127866 222352
rect 139118 222300 139124 222352
rect 139176 222340 139182 222352
rect 146956 222340 146984 222448
rect 206830 222436 206836 222448
rect 206888 222436 206894 222488
rect 207842 222436 207848 222488
rect 207900 222476 207906 222488
rect 258350 222476 258356 222488
rect 207900 222448 258356 222476
rect 207900 222436 207906 222448
rect 258350 222436 258356 222448
rect 258408 222436 258414 222488
rect 500218 222436 500224 222488
rect 500276 222476 500282 222488
rect 542814 222476 542820 222488
rect 500276 222448 542820 222476
rect 500276 222436 500282 222448
rect 542814 222436 542820 222448
rect 542872 222436 542878 222488
rect 542998 222436 543004 222488
rect 543056 222476 543062 222488
rect 621198 222476 621204 222488
rect 543056 222448 621204 222476
rect 543056 222436 543062 222448
rect 621198 222436 621204 222448
rect 621256 222436 621262 222488
rect 490006 222368 490012 222420
rect 490064 222408 490070 222420
rect 490064 222380 495434 222408
rect 490064 222368 490070 222380
rect 139176 222312 146984 222340
rect 139176 222300 139182 222312
rect 147122 222300 147128 222352
rect 147180 222340 147186 222352
rect 211982 222340 211988 222352
rect 147180 222312 211988 222340
rect 147180 222300 147186 222312
rect 211982 222300 211988 222312
rect 212040 222300 212046 222352
rect 237006 222300 237012 222352
rect 237064 222340 237070 222352
rect 280890 222340 280896 222352
rect 237064 222312 280896 222340
rect 237064 222300 237070 222312
rect 280890 222300 280896 222312
rect 280948 222300 280954 222352
rect 484578 222300 484584 222352
rect 484636 222340 484642 222352
rect 495406 222340 495434 222380
rect 629846 222340 629852 222352
rect 484636 222312 489914 222340
rect 495406 222312 629852 222340
rect 484636 222300 484642 222312
rect 489886 222204 489914 222312
rect 629846 222300 629852 222312
rect 629904 222300 629910 222352
rect 500218 222204 500224 222216
rect 489886 222176 500224 222204
rect 500218 222164 500224 222176
rect 500276 222164 500282 222216
rect 542814 222164 542820 222216
rect 542872 222204 542878 222216
rect 558178 222204 558184 222216
rect 542872 222176 558184 222204
rect 542872 222164 542878 222176
rect 558178 222164 558184 222176
rect 558236 222164 558242 222216
rect 558546 222164 558552 222216
rect 558604 222204 558610 222216
rect 559926 222204 559932 222216
rect 558604 222176 559932 222204
rect 558604 222164 558610 222176
rect 559926 222164 559932 222176
rect 559984 222204 559990 222216
rect 627086 222204 627092 222216
rect 559984 222176 627092 222204
rect 559984 222164 559990 222176
rect 627086 222164 627092 222176
rect 627144 222164 627150 222216
rect 670804 222148 670832 222992
rect 111978 222096 111984 222148
rect 112036 222136 112042 222148
rect 185946 222136 185952 222148
rect 112036 222108 185952 222136
rect 112036 222096 112042 222108
rect 185946 222096 185952 222108
rect 186004 222096 186010 222148
rect 200390 222096 200396 222148
rect 200448 222136 200454 222148
rect 252922 222136 252928 222148
rect 200448 222108 252928 222136
rect 200448 222096 200454 222108
rect 252922 222096 252928 222108
rect 252980 222096 252986 222148
rect 258074 222096 258080 222148
rect 258132 222136 258138 222148
rect 263870 222136 263876 222148
rect 258132 222108 263876 222136
rect 258132 222096 258138 222108
rect 263870 222096 263876 222108
rect 263928 222096 263934 222148
rect 270034 222096 270040 222148
rect 270092 222136 270098 222148
rect 306374 222136 306380 222148
rect 270092 222108 306380 222136
rect 270092 222096 270098 222108
rect 306374 222096 306380 222108
rect 306432 222096 306438 222148
rect 310698 222096 310704 222148
rect 310756 222136 310762 222148
rect 312630 222136 312636 222148
rect 310756 222108 312636 222136
rect 310756 222096 310762 222108
rect 312630 222096 312636 222108
rect 312688 222096 312694 222148
rect 331398 222096 331404 222148
rect 331456 222136 331462 222148
rect 353938 222136 353944 222148
rect 331456 222108 353944 222136
rect 331456 222096 331462 222108
rect 353938 222096 353944 222108
rect 353996 222096 354002 222148
rect 424962 222096 424968 222148
rect 425020 222136 425026 222148
rect 429286 222136 429292 222148
rect 425020 222108 429292 222136
rect 425020 222096 425026 222108
rect 429286 222096 429292 222108
rect 429344 222096 429350 222148
rect 452562 222096 452568 222148
rect 452620 222136 452626 222148
rect 455598 222136 455604 222148
rect 452620 222108 455604 222136
rect 452620 222096 452626 222108
rect 455598 222096 455604 222108
rect 455656 222096 455662 222148
rect 462130 222096 462136 222148
rect 462188 222136 462194 222148
rect 468754 222136 468760 222148
rect 462188 222108 468760 222136
rect 462188 222096 462194 222108
rect 468754 222096 468760 222108
rect 468812 222096 468818 222148
rect 471882 222096 471888 222148
rect 471940 222136 471946 222148
rect 477862 222136 477868 222148
rect 471940 222108 477868 222136
rect 471940 222096 471946 222108
rect 477862 222096 477868 222108
rect 477920 222096 477926 222148
rect 533154 222096 533160 222148
rect 533212 222136 533218 222148
rect 538674 222136 538680 222148
rect 533212 222108 538680 222136
rect 533212 222096 533218 222108
rect 538674 222096 538680 222108
rect 538732 222096 538738 222148
rect 539502 222096 539508 222148
rect 539560 222136 539566 222148
rect 542262 222136 542268 222148
rect 539560 222108 542268 222136
rect 539560 222096 539566 222108
rect 542262 222096 542268 222108
rect 542320 222096 542326 222148
rect 670786 222096 670792 222148
rect 670844 222096 670850 222148
rect 543826 222028 543832 222080
rect 543884 222068 543890 222080
rect 605006 222068 605012 222080
rect 543884 222040 605012 222068
rect 543884 222028 543890 222040
rect 605006 222028 605012 222040
rect 605064 222028 605070 222080
rect 91278 221960 91284 222012
rect 91336 222000 91342 222012
rect 167178 222000 167184 222012
rect 91336 221972 167184 222000
rect 91336 221960 91342 221972
rect 167178 221960 167184 221972
rect 167236 221960 167242 222012
rect 167454 221960 167460 222012
rect 167512 222000 167518 222012
rect 172698 222000 172704 222012
rect 167512 221972 172704 222000
rect 167512 221960 167518 221972
rect 172698 221960 172704 221972
rect 172756 221960 172762 222012
rect 226518 222000 226524 222012
rect 172900 221972 226524 222000
rect 94590 221824 94596 221876
rect 94648 221864 94654 221876
rect 161428 221864 161434 221876
rect 94648 221836 161434 221864
rect 94648 221824 94654 221836
rect 161428 221824 161434 221836
rect 161486 221824 161492 221876
rect 161566 221824 161572 221876
rect 161624 221864 161630 221876
rect 164326 221864 164332 221876
rect 161624 221836 164332 221864
rect 161624 221824 161630 221836
rect 164326 221824 164332 221836
rect 164384 221824 164390 221876
rect 164510 221824 164516 221876
rect 164568 221864 164574 221876
rect 169846 221864 169852 221876
rect 164568 221836 169852 221864
rect 164568 221824 164574 221836
rect 169846 221824 169852 221836
rect 169904 221824 169910 221876
rect 97718 221688 97724 221740
rect 97776 221728 97782 221740
rect 167454 221728 167460 221740
rect 97776 221700 167460 221728
rect 97776 221688 97782 221700
rect 167454 221688 167460 221700
rect 167512 221688 167518 221740
rect 167638 221688 167644 221740
rect 167696 221728 167702 221740
rect 167696 221700 168052 221728
rect 167696 221688 167702 221700
rect 73890 221552 73896 221604
rect 73948 221592 73954 221604
rect 82078 221592 82084 221604
rect 73948 221564 82084 221592
rect 73948 221552 73954 221564
rect 82078 221552 82084 221564
rect 82136 221552 82142 221604
rect 86310 221552 86316 221604
rect 86368 221592 86374 221604
rect 161474 221592 161480 221604
rect 86368 221564 161480 221592
rect 86368 221552 86374 221564
rect 161474 221552 161480 221564
rect 161532 221552 161538 221604
rect 161658 221552 161664 221604
rect 161716 221592 161722 221604
rect 167822 221592 167828 221604
rect 161716 221564 167828 221592
rect 161716 221552 161722 221564
rect 167822 221552 167828 221564
rect 167880 221552 167886 221604
rect 168024 221592 168052 221700
rect 168190 221688 168196 221740
rect 168248 221728 168254 221740
rect 172900 221728 172928 221972
rect 226518 221960 226524 221972
rect 226576 221960 226582 222012
rect 232130 221960 232136 222012
rect 232188 222000 232194 222012
rect 234706 222000 234712 222012
rect 232188 221972 234712 222000
rect 232188 221960 232194 221972
rect 234706 221960 234712 221972
rect 234764 221960 234770 222012
rect 261018 221960 261024 222012
rect 261076 222000 261082 222012
rect 301682 222000 301688 222012
rect 261076 221972 301688 222000
rect 261076 221960 261082 221972
rect 301682 221960 301688 221972
rect 301740 221960 301746 222012
rect 313182 221960 313188 222012
rect 313240 222000 313246 222012
rect 340414 222000 340420 222012
rect 313240 221972 340420 222000
rect 313240 221960 313246 221972
rect 340414 221960 340420 221972
rect 340472 221960 340478 222012
rect 516778 221960 516784 222012
rect 516836 222000 516842 222012
rect 527542 222000 527548 222012
rect 516836 221972 527548 222000
rect 516836 221960 516842 221972
rect 527542 221960 527548 221972
rect 527600 221960 527606 222012
rect 527726 221960 527732 222012
rect 527784 222000 527790 222012
rect 528186 222000 528192 222012
rect 527784 221972 528192 222000
rect 527784 221960 527790 221972
rect 528186 221960 528192 221972
rect 528244 222000 528250 222012
rect 533522 222000 533528 222012
rect 528244 221972 533528 222000
rect 528244 221960 528250 221972
rect 533522 221960 533528 221972
rect 533580 221960 533586 222012
rect 533982 221960 533988 222012
rect 534040 222000 534046 222012
rect 542998 222000 543004 222012
rect 534040 221972 543004 222000
rect 534040 221960 534046 221972
rect 542998 221960 543004 221972
rect 543056 221960 543062 222012
rect 543366 221960 543372 222012
rect 543424 222000 543430 222012
rect 543688 222000 543694 222012
rect 543424 221972 543694 222000
rect 543424 221960 543430 221972
rect 543688 221960 543694 221972
rect 543746 221960 543752 222012
rect 174078 221824 174084 221876
rect 174136 221864 174142 221876
rect 231946 221864 231952 221876
rect 174136 221836 231952 221864
rect 174136 221824 174142 221836
rect 231946 221824 231952 221836
rect 232004 221824 232010 221876
rect 233694 221824 233700 221876
rect 233752 221864 233758 221876
rect 277946 221864 277952 221876
rect 233752 221836 277952 221864
rect 233752 221824 233758 221836
rect 277946 221824 277952 221836
rect 278004 221824 278010 221876
rect 280062 221824 280068 221876
rect 280120 221864 280126 221876
rect 313734 221864 313740 221876
rect 280120 221836 313740 221864
rect 280120 221824 280126 221836
rect 313734 221824 313740 221836
rect 313792 221824 313798 221876
rect 318242 221824 318248 221876
rect 318300 221864 318306 221876
rect 343634 221864 343640 221876
rect 318300 221836 343640 221864
rect 318300 221824 318306 221836
rect 343634 221824 343640 221836
rect 343692 221824 343698 221876
rect 353294 221824 353300 221876
rect 353352 221864 353358 221876
rect 372706 221864 372712 221876
rect 353352 221836 372712 221864
rect 353352 221824 353358 221836
rect 372706 221824 372712 221836
rect 372764 221824 372770 221876
rect 380342 221864 380348 221876
rect 373966 221836 380348 221864
rect 168248 221700 172928 221728
rect 168248 221688 168254 221700
rect 174906 221688 174912 221740
rect 174964 221728 174970 221740
rect 174964 221700 185348 221728
rect 174964 221688 174970 221700
rect 185320 221660 185348 221700
rect 185762 221688 185768 221740
rect 185820 221728 185826 221740
rect 243078 221728 243084 221740
rect 185820 221700 243084 221728
rect 185820 221688 185826 221700
rect 243078 221688 243084 221700
rect 243136 221688 243142 221740
rect 263134 221728 263140 221740
rect 243556 221700 263140 221728
rect 185320 221632 185440 221660
rect 182634 221592 182640 221604
rect 168024 221564 182640 221592
rect 182634 221552 182640 221564
rect 182692 221552 182698 221604
rect 185412 221592 185440 221632
rect 232130 221592 232136 221604
rect 185412 221564 232136 221592
rect 232130 221552 232136 221564
rect 232188 221552 232194 221604
rect 243556 221592 243584 221700
rect 263134 221688 263140 221700
rect 263192 221688 263198 221740
rect 263502 221688 263508 221740
rect 263560 221728 263566 221740
rect 301038 221728 301044 221740
rect 263560 221700 301044 221728
rect 263560 221688 263566 221700
rect 301038 221688 301044 221700
rect 301096 221688 301102 221740
rect 303246 221688 303252 221740
rect 303304 221728 303310 221740
rect 332778 221728 332784 221740
rect 303304 221700 332784 221728
rect 303304 221688 303310 221700
rect 332778 221688 332784 221700
rect 332836 221688 332842 221740
rect 344646 221688 344652 221740
rect 344704 221728 344710 221740
rect 364518 221728 364524 221740
rect 344704 221700 364524 221728
rect 344704 221688 344710 221700
rect 364518 221688 364524 221700
rect 364576 221688 364582 221740
rect 370958 221688 370964 221740
rect 371016 221728 371022 221740
rect 373966 221728 373994 221836
rect 380342 221824 380348 221836
rect 380400 221824 380406 221876
rect 492490 221824 492496 221876
rect 492548 221864 492554 221876
rect 506842 221864 506848 221876
rect 492548 221836 506848 221864
rect 492548 221824 492554 221836
rect 506842 221824 506848 221836
rect 506900 221824 506906 221876
rect 515766 221824 515772 221876
rect 515824 221864 515830 221876
rect 600314 221864 600320 221876
rect 515824 221836 600320 221864
rect 515824 221824 515830 221836
rect 600314 221824 600320 221836
rect 600372 221824 600378 221876
rect 371016 221700 373994 221728
rect 371016 221688 371022 221700
rect 380066 221688 380072 221740
rect 380124 221728 380130 221740
rect 386506 221728 386512 221740
rect 380124 221700 386512 221728
rect 380124 221688 380130 221700
rect 386506 221688 386512 221700
rect 386564 221688 386570 221740
rect 484762 221688 484768 221740
rect 484820 221728 484826 221740
rect 497734 221728 497740 221740
rect 484820 221700 497740 221728
rect 484820 221688 484826 221700
rect 497734 221688 497740 221700
rect 497792 221688 497798 221740
rect 501322 221688 501328 221740
rect 501380 221728 501386 221740
rect 519630 221728 519636 221740
rect 501380 221700 519636 221728
rect 501380 221688 501386 221700
rect 519630 221688 519636 221700
rect 519688 221688 519694 221740
rect 522666 221688 522672 221740
rect 522724 221728 522730 221740
rect 542354 221728 542360 221740
rect 522724 221700 542360 221728
rect 522724 221688 522730 221700
rect 542354 221688 542360 221700
rect 542412 221688 542418 221740
rect 542998 221688 543004 221740
rect 543056 221728 543062 221740
rect 543688 221728 543694 221740
rect 543056 221700 543694 221728
rect 543056 221688 543062 221700
rect 543688 221688 543694 221700
rect 543746 221688 543752 221740
rect 543826 221688 543832 221740
rect 543884 221728 543890 221740
rect 601142 221728 601148 221740
rect 543884 221700 601148 221728
rect 543884 221688 543890 221700
rect 601142 221688 601148 221700
rect 601200 221688 601206 221740
rect 233896 221564 243584 221592
rect 59354 221416 59360 221468
rect 59412 221456 59418 221468
rect 141326 221456 141332 221468
rect 59412 221428 141332 221456
rect 59412 221416 59418 221428
rect 141326 221416 141332 221428
rect 141384 221416 141390 221468
rect 147582 221416 147588 221468
rect 147640 221456 147646 221468
rect 204898 221456 204904 221468
rect 147640 221428 204904 221456
rect 147640 221416 147646 221428
rect 204898 221416 204904 221428
rect 204956 221416 204962 221468
rect 205082 221416 205088 221468
rect 205140 221456 205146 221468
rect 220170 221456 220176 221468
rect 205140 221428 220176 221456
rect 205140 221416 205146 221428
rect 220170 221416 220176 221428
rect 220228 221416 220234 221468
rect 220998 221416 221004 221468
rect 221056 221456 221062 221468
rect 233896 221456 233924 221564
rect 243722 221552 243728 221604
rect 243780 221592 243786 221604
rect 283742 221592 283748 221604
rect 243780 221564 283748 221592
rect 243780 221552 243786 221564
rect 283742 221552 283748 221564
rect 283800 221552 283806 221604
rect 302418 221552 302424 221604
rect 302476 221592 302482 221604
rect 334066 221592 334072 221604
rect 302476 221564 334072 221592
rect 302476 221552 302482 221564
rect 334066 221552 334072 221564
rect 334124 221552 334130 221604
rect 348786 221552 348792 221604
rect 348844 221592 348850 221604
rect 370038 221592 370044 221604
rect 348844 221564 370044 221592
rect 348844 221552 348850 221564
rect 370038 221552 370044 221564
rect 370096 221552 370102 221604
rect 373718 221552 373724 221604
rect 373776 221592 373782 221604
rect 384298 221592 384304 221604
rect 373776 221564 384304 221592
rect 373776 221552 373782 221564
rect 384298 221552 384304 221564
rect 384356 221552 384362 221604
rect 391014 221552 391020 221604
rect 391072 221592 391078 221604
rect 400306 221592 400312 221604
rect 391072 221564 400312 221592
rect 391072 221552 391078 221564
rect 400306 221552 400312 221564
rect 400364 221552 400370 221604
rect 401226 221552 401232 221604
rect 401284 221592 401290 221604
rect 405826 221592 405832 221604
rect 401284 221564 405832 221592
rect 401284 221552 401290 221564
rect 405826 221552 405832 221564
rect 405884 221552 405890 221604
rect 475838 221552 475844 221604
rect 475896 221592 475902 221604
rect 486142 221592 486148 221604
rect 475896 221564 486148 221592
rect 475896 221552 475902 221564
rect 486142 221552 486148 221564
rect 486200 221552 486206 221604
rect 496262 221552 496268 221604
rect 496320 221592 496326 221604
rect 513558 221592 513564 221604
rect 496320 221564 513564 221592
rect 496320 221552 496326 221564
rect 513558 221552 513564 221564
rect 513616 221552 513622 221604
rect 524230 221552 524236 221604
rect 524288 221592 524294 221604
rect 524288 221564 533384 221592
rect 524288 221552 524294 221564
rect 221056 221428 233924 221456
rect 221056 221416 221062 221428
rect 234062 221416 234068 221468
rect 234120 221456 234126 221468
rect 276106 221456 276112 221468
rect 234120 221428 276112 221456
rect 234120 221416 234126 221428
rect 276106 221416 276112 221428
rect 276164 221416 276170 221468
rect 284018 221416 284024 221468
rect 284076 221456 284082 221468
rect 320358 221456 320364 221468
rect 284076 221428 320364 221456
rect 284076 221416 284082 221428
rect 320358 221416 320364 221428
rect 320416 221416 320422 221468
rect 333606 221416 333612 221468
rect 333664 221456 333670 221468
rect 357526 221456 357532 221468
rect 333664 221428 357532 221456
rect 333664 221416 333670 221428
rect 357526 221416 357532 221428
rect 357584 221416 357590 221468
rect 369486 221416 369492 221468
rect 369544 221456 369550 221468
rect 384114 221456 384120 221468
rect 369544 221428 384120 221456
rect 369544 221416 369550 221428
rect 384114 221416 384120 221428
rect 384172 221416 384178 221468
rect 384390 221416 384396 221468
rect 384448 221456 384454 221468
rect 395154 221456 395160 221468
rect 384448 221428 395160 221456
rect 384448 221416 384454 221428
rect 395154 221416 395160 221428
rect 395212 221416 395218 221468
rect 396810 221416 396816 221468
rect 396868 221456 396874 221468
rect 407298 221456 407304 221468
rect 396868 221428 407304 221456
rect 396868 221416 396874 221428
rect 407298 221416 407304 221428
rect 407356 221416 407362 221468
rect 408402 221416 408408 221468
rect 408460 221456 408466 221468
rect 416866 221456 416872 221468
rect 408460 221428 416872 221456
rect 408460 221416 408466 221428
rect 416866 221416 416872 221428
rect 416924 221416 416930 221468
rect 468938 221416 468944 221468
rect 468996 221456 469002 221468
rect 476206 221456 476212 221468
rect 468996 221428 476212 221456
rect 468996 221416 469002 221428
rect 476206 221416 476212 221428
rect 476264 221416 476270 221468
rect 483750 221416 483756 221468
rect 483808 221456 483814 221468
rect 533154 221456 533160 221468
rect 483808 221428 533160 221456
rect 483808 221416 483814 221428
rect 533154 221416 533160 221428
rect 533212 221416 533218 221468
rect 533356 221456 533384 221564
rect 533522 221552 533528 221604
rect 533580 221592 533586 221604
rect 600682 221592 600688 221604
rect 533580 221564 600688 221592
rect 533580 221552 533586 221564
rect 600682 221552 600688 221564
rect 600740 221552 600746 221604
rect 606110 221592 606116 221604
rect 600976 221564 606116 221592
rect 543734 221456 543740 221468
rect 533356 221428 543740 221456
rect 543734 221416 543740 221428
rect 543792 221416 543798 221468
rect 544746 221416 544752 221468
rect 544804 221456 544810 221468
rect 600976 221456 601004 221564
rect 606110 221552 606116 221564
rect 606168 221552 606174 221604
rect 544804 221428 601004 221456
rect 544804 221416 544810 221428
rect 601142 221416 601148 221468
rect 601200 221456 601206 221468
rect 605926 221456 605932 221468
rect 601200 221428 605932 221456
rect 601200 221416 601206 221428
rect 605926 221416 605932 221428
rect 605984 221416 605990 221468
rect 104526 221280 104532 221332
rect 104584 221320 104590 221332
rect 176470 221320 176476 221332
rect 104584 221292 176476 221320
rect 104584 221280 104590 221292
rect 176470 221280 176476 221292
rect 176528 221280 176534 221332
rect 176626 221292 185532 221320
rect 111150 221144 111156 221196
rect 111208 221184 111214 221196
rect 167638 221184 167644 221196
rect 111208 221156 167644 221184
rect 111208 221144 111214 221156
rect 167638 221144 167644 221156
rect 167696 221144 167702 221196
rect 167822 221144 167828 221196
rect 167880 221184 167886 221196
rect 176626 221184 176654 221292
rect 185504 221252 185532 221292
rect 185854 221280 185860 221332
rect 185912 221320 185918 221332
rect 234246 221320 234252 221332
rect 185912 221292 234252 221320
rect 185912 221280 185918 221292
rect 234246 221280 234252 221292
rect 234304 221280 234310 221332
rect 237834 221280 237840 221332
rect 237892 221320 237898 221332
rect 243722 221320 243728 221332
rect 237892 221292 243728 221320
rect 237892 221280 237898 221292
rect 243722 221280 243728 221292
rect 243780 221280 243786 221332
rect 266814 221280 266820 221332
rect 266872 221320 266878 221332
rect 303798 221320 303804 221332
rect 266872 221292 303804 221320
rect 266872 221280 266878 221292
rect 303798 221280 303804 221292
rect 303856 221280 303862 221332
rect 600682 221280 600688 221332
rect 600740 221320 600746 221332
rect 603166 221320 603172 221332
rect 600740 221292 603172 221320
rect 600740 221280 600746 221292
rect 603166 221280 603172 221292
rect 603224 221280 603230 221332
rect 185504 221224 185716 221252
rect 167880 221156 176654 221184
rect 167880 221144 167886 221156
rect 177298 221144 177304 221196
rect 177356 221184 177362 221196
rect 185302 221184 185308 221196
rect 177356 221156 185308 221184
rect 177356 221144 177362 221156
rect 185302 221144 185308 221156
rect 185360 221144 185366 221196
rect 185688 221184 185716 221224
rect 520918 221212 520924 221264
rect 520976 221252 520982 221264
rect 600498 221252 600504 221264
rect 520976 221224 600504 221252
rect 520976 221212 520982 221224
rect 600498 221212 600504 221224
rect 600556 221212 600562 221264
rect 185688 221156 200114 221184
rect 124398 221008 124404 221060
rect 124456 221048 124462 221060
rect 193306 221048 193312 221060
rect 124456 221020 193312 221048
rect 124456 221008 124462 221020
rect 193306 221008 193312 221020
rect 193364 221008 193370 221060
rect 200086 221048 200114 221156
rect 204898 221144 204904 221196
rect 204956 221184 204962 221196
rect 211154 221184 211160 221196
rect 204956 221156 211160 221184
rect 204956 221144 204962 221156
rect 211154 221144 211160 221156
rect 211212 221144 211218 221196
rect 211522 221144 211528 221196
rect 211580 221184 211586 221196
rect 260834 221184 260840 221196
rect 211580 221156 260840 221184
rect 211580 221144 211586 221156
rect 260834 221144 260840 221156
rect 260892 221144 260898 221196
rect 517514 221076 517520 221128
rect 517572 221116 517578 221128
rect 518434 221116 518440 221128
rect 517572 221088 518440 221116
rect 517572 221076 517578 221088
rect 518434 221076 518440 221088
rect 518492 221116 518498 221128
rect 600682 221116 600688 221128
rect 518492 221088 600688 221116
rect 518492 221076 518498 221088
rect 600682 221076 600688 221088
rect 600740 221076 600746 221128
rect 205082 221048 205088 221060
rect 200086 221020 205088 221048
rect 205082 221008 205088 221020
rect 205140 221008 205146 221060
rect 218054 221008 218060 221060
rect 218112 221048 218118 221060
rect 220998 221048 221004 221060
rect 218112 221020 221004 221048
rect 218112 221008 218118 221020
rect 220998 221008 221004 221020
rect 221056 221008 221062 221060
rect 227898 221008 227904 221060
rect 227956 221048 227962 221060
rect 234062 221048 234068 221060
rect 227956 221020 234068 221048
rect 227956 221008 227962 221020
rect 234062 221008 234068 221020
rect 234120 221008 234126 221060
rect 268194 221048 268200 221060
rect 238726 221020 268200 221048
rect 82998 220940 83004 220992
rect 83056 220980 83062 220992
rect 83056 220952 93854 220980
rect 83056 220940 83062 220952
rect 93826 220912 93854 220952
rect 151078 220912 151084 220924
rect 93826 220884 151084 220912
rect 151078 220872 151084 220884
rect 151136 220872 151142 220924
rect 155034 220872 155040 220924
rect 155092 220912 155098 220924
rect 158254 220912 158260 220924
rect 155092 220884 158260 220912
rect 155092 220872 155098 220884
rect 158254 220872 158260 220884
rect 158312 220872 158318 220924
rect 158438 220872 158444 220924
rect 158496 220912 158502 220924
rect 222286 220912 222292 220924
rect 158496 220884 222292 220912
rect 158496 220872 158502 220884
rect 222286 220872 222292 220884
rect 222344 220872 222350 220924
rect 223482 220872 223488 220924
rect 223540 220912 223546 220924
rect 238726 220912 238754 221020
rect 268194 221008 268200 221020
rect 268252 221008 268258 221060
rect 523494 220940 523500 220992
rect 523552 220980 523558 220992
rect 601694 220980 601700 220992
rect 523552 220952 601700 220980
rect 523552 220940 523558 220952
rect 601694 220940 601700 220952
rect 601752 220940 601758 220992
rect 223540 220884 238754 220912
rect 223540 220872 223546 220884
rect 253382 220872 253388 220924
rect 253440 220912 253446 220924
rect 258626 220912 258632 220924
rect 253440 220884 258632 220912
rect 253440 220872 253446 220884
rect 258626 220872 258632 220884
rect 258684 220872 258690 220924
rect 80514 220804 80520 220856
rect 80572 220844 80578 220856
rect 86126 220844 86132 220856
rect 80572 220816 86132 220844
rect 80572 220804 80578 220816
rect 86126 220804 86132 220816
rect 86184 220804 86190 220856
rect 418338 220804 418344 220856
rect 418396 220844 418402 220856
rect 424042 220844 424048 220856
rect 418396 220816 424048 220844
rect 418396 220804 418402 220816
rect 424042 220804 424048 220816
rect 424100 220804 424106 220856
rect 456702 220804 456708 220856
rect 456760 220844 456766 220856
rect 462130 220844 462136 220856
rect 456760 220816 462136 220844
rect 456760 220804 456766 220816
rect 462130 220804 462136 220816
rect 462188 220804 462194 220856
rect 466086 220804 466092 220856
rect 466144 220844 466150 220856
rect 471330 220844 471336 220856
rect 466144 220816 471336 220844
rect 466144 220804 466150 220816
rect 471330 220804 471336 220816
rect 471388 220804 471394 220856
rect 538490 220804 538496 220856
rect 538548 220844 538554 220856
rect 539502 220844 539508 220856
rect 538548 220816 539508 220844
rect 538548 220804 538554 220816
rect 539502 220804 539508 220816
rect 539560 220804 539566 220856
rect 542354 220804 542360 220856
rect 542412 220844 542418 220856
rect 542412 220816 543872 220844
rect 542412 220804 542418 220816
rect 107838 220736 107844 220788
rect 107896 220776 107902 220788
rect 176470 220776 176476 220788
rect 107896 220748 176476 220776
rect 107896 220736 107902 220748
rect 176470 220736 176476 220748
rect 176528 220736 176534 220788
rect 176608 220736 176614 220788
rect 176666 220776 176672 220788
rect 180518 220776 180524 220788
rect 176666 220748 180524 220776
rect 176666 220736 176672 220748
rect 180518 220736 180524 220748
rect 180576 220736 180582 220788
rect 180702 220736 180708 220788
rect 180760 220776 180766 220788
rect 236730 220776 236736 220788
rect 180760 220748 236736 220776
rect 180760 220736 180766 220748
rect 236730 220736 236736 220748
rect 236788 220736 236794 220788
rect 246942 220736 246948 220788
rect 247000 220776 247006 220788
rect 288618 220776 288624 220788
rect 247000 220748 288624 220776
rect 247000 220736 247006 220748
rect 288618 220736 288624 220748
rect 288676 220736 288682 220788
rect 340046 220736 340052 220788
rect 340104 220776 340110 220788
rect 342346 220776 342352 220788
rect 340104 220748 342352 220776
rect 340104 220736 340110 220748
rect 342346 220736 342352 220748
rect 342404 220736 342410 220788
rect 414198 220736 414204 220788
rect 414256 220776 414262 220788
rect 418154 220776 418160 220788
rect 414256 220748 418160 220776
rect 414256 220736 414262 220748
rect 418154 220736 418160 220748
rect 418212 220736 418218 220788
rect 473998 220736 474004 220788
rect 474056 220776 474062 220788
rect 475378 220776 475384 220788
rect 474056 220748 475384 220776
rect 474056 220736 474062 220748
rect 475378 220736 475384 220748
rect 475436 220736 475442 220788
rect 476758 220736 476764 220788
rect 476816 220776 476822 220788
rect 478690 220776 478696 220788
rect 476816 220748 478696 220776
rect 476816 220736 476822 220748
rect 478690 220736 478696 220748
rect 478748 220736 478754 220788
rect 500402 220736 500408 220788
rect 500460 220776 500466 220788
rect 511810 220776 511816 220788
rect 500460 220748 511816 220776
rect 500460 220736 500466 220748
rect 511810 220736 511816 220748
rect 511868 220736 511874 220788
rect 543844 220776 543872 220816
rect 544378 220804 544384 220856
rect 544436 220844 544442 220856
rect 553394 220844 553400 220856
rect 544436 220816 553400 220844
rect 544436 220804 544442 220816
rect 553394 220804 553400 220816
rect 553452 220804 553458 220856
rect 559558 220804 559564 220856
rect 559616 220844 559622 220856
rect 563054 220844 563060 220856
rect 559616 220816 563060 220844
rect 559616 220804 559622 220816
rect 563054 220804 563060 220816
rect 563112 220804 563118 220856
rect 563238 220804 563244 220856
rect 563296 220844 563302 220856
rect 609422 220844 609428 220856
rect 563296 220816 609428 220844
rect 563296 220804 563302 220816
rect 609422 220804 609428 220816
rect 609480 220804 609486 220856
rect 543844 220748 543964 220776
rect 455322 220668 455328 220720
rect 455380 220708 455386 220720
rect 458818 220708 458824 220720
rect 455380 220680 458824 220708
rect 455380 220668 455386 220680
rect 458818 220668 458824 220680
rect 458876 220668 458882 220720
rect 465718 220668 465724 220720
rect 465776 220708 465782 220720
rect 469582 220708 469588 220720
rect 465776 220680 469588 220708
rect 465776 220668 465782 220680
rect 469582 220668 469588 220680
rect 469640 220668 469646 220720
rect 543936 220708 543964 220748
rect 546586 220708 546592 220720
rect 543936 220680 546592 220708
rect 546586 220668 546592 220680
rect 546644 220668 546650 220720
rect 79686 220600 79692 220652
rect 79744 220640 79750 220652
rect 154022 220640 154028 220652
rect 79744 220612 154028 220640
rect 79744 220600 79750 220612
rect 154022 220600 154028 220612
rect 154080 220600 154086 220652
rect 154206 220600 154212 220652
rect 154264 220640 154270 220652
rect 156782 220640 156788 220652
rect 154264 220612 156788 220640
rect 154264 220600 154270 220612
rect 156782 220600 156788 220612
rect 156840 220600 156846 220652
rect 156966 220600 156972 220652
rect 157024 220640 157030 220652
rect 158898 220640 158904 220652
rect 157024 220612 158904 220640
rect 157024 220600 157030 220612
rect 158898 220600 158904 220612
rect 158956 220600 158962 220652
rect 160830 220600 160836 220652
rect 160888 220640 160894 220652
rect 221274 220640 221280 220652
rect 160888 220612 221280 220640
rect 160888 220600 160894 220612
rect 221274 220600 221280 220612
rect 221332 220600 221338 220652
rect 223758 220640 223764 220652
rect 221568 220612 223764 220640
rect 76374 220464 76380 220516
rect 76432 220504 76438 220516
rect 156138 220504 156144 220516
rect 76432 220476 156144 220504
rect 76432 220464 76438 220476
rect 156138 220464 156144 220476
rect 156196 220464 156202 220516
rect 156598 220464 156604 220516
rect 156656 220504 156662 220516
rect 166948 220504 166954 220516
rect 156656 220476 166954 220504
rect 156656 220464 156662 220476
rect 166948 220464 166954 220476
rect 167006 220464 167012 220516
rect 167086 220464 167092 220516
rect 167144 220504 167150 220516
rect 221568 220504 221596 220612
rect 223758 220600 223764 220612
rect 223816 220600 223822 220652
rect 236178 220600 236184 220652
rect 236236 220640 236242 220652
rect 246482 220640 246488 220652
rect 236236 220612 246488 220640
rect 236236 220600 236242 220612
rect 246482 220600 246488 220612
rect 246540 220600 246546 220652
rect 254394 220600 254400 220652
rect 254452 220640 254458 220652
rect 296806 220640 296812 220652
rect 254452 220612 296812 220640
rect 254452 220600 254458 220612
rect 296806 220600 296812 220612
rect 296864 220600 296870 220652
rect 304902 220600 304908 220652
rect 304960 220640 304966 220652
rect 333422 220640 333428 220652
rect 304960 220612 333428 220640
rect 304960 220600 304966 220612
rect 333422 220600 333428 220612
rect 333480 220600 333486 220652
rect 509878 220600 509884 220652
rect 509936 220640 509942 220652
rect 522574 220640 522580 220652
rect 509936 220612 522580 220640
rect 509936 220600 509942 220612
rect 522574 220600 522580 220612
rect 522632 220600 522638 220652
rect 529014 220600 529020 220652
rect 529072 220640 529078 220652
rect 529072 220612 543780 220640
rect 529072 220600 529078 220612
rect 167144 220476 221596 220504
rect 167144 220464 167150 220476
rect 223758 220464 223764 220516
rect 223816 220504 223822 220516
rect 270586 220504 270592 220516
rect 223816 220476 270592 220504
rect 223816 220464 223822 220476
rect 270586 220464 270592 220476
rect 270644 220464 270650 220516
rect 292482 220464 292488 220516
rect 292540 220504 292546 220516
rect 326154 220504 326160 220516
rect 292540 220476 326160 220504
rect 292540 220464 292546 220476
rect 326154 220464 326160 220476
rect 326212 220464 326218 220516
rect 328086 220464 328092 220516
rect 328144 220504 328150 220516
rect 351270 220504 351276 220516
rect 328144 220476 351276 220504
rect 328144 220464 328150 220476
rect 351270 220464 351276 220476
rect 351328 220464 351334 220516
rect 364518 220464 364524 220516
rect 364576 220504 364582 220516
rect 379698 220504 379704 220516
rect 364576 220476 379704 220504
rect 364576 220464 364582 220476
rect 379698 220464 379704 220476
rect 379756 220464 379762 220516
rect 469122 220464 469128 220516
rect 469180 220504 469186 220516
rect 474550 220504 474556 220516
rect 469180 220476 474556 220504
rect 469180 220464 469186 220476
rect 474550 220464 474556 220476
rect 474608 220464 474614 220516
rect 488442 220464 488448 220516
rect 488500 220504 488506 220516
rect 501874 220504 501880 220516
rect 488500 220476 501880 220504
rect 488500 220464 488506 220476
rect 501874 220464 501880 220476
rect 501932 220464 501938 220516
rect 511626 220464 511632 220516
rect 511684 220504 511690 220516
rect 531682 220504 531688 220516
rect 511684 220476 531688 220504
rect 511684 220464 511690 220476
rect 531682 220464 531688 220476
rect 531740 220464 531746 220516
rect 540790 220464 540796 220516
rect 540848 220504 540854 220516
rect 543550 220504 543556 220516
rect 540848 220476 543556 220504
rect 540848 220464 540854 220476
rect 543550 220464 543556 220476
rect 543608 220464 543614 220516
rect 543752 220504 543780 220612
rect 557994 220600 558000 220652
rect 558052 220640 558058 220652
rect 566458 220640 566464 220652
rect 558052 220612 566464 220640
rect 558052 220600 558058 220612
rect 566458 220600 566464 220612
rect 566516 220600 566522 220652
rect 566642 220600 566648 220652
rect 566700 220640 566706 220652
rect 567286 220640 567292 220652
rect 566700 220612 567292 220640
rect 566700 220600 566706 220612
rect 567286 220600 567292 220612
rect 567344 220600 567350 220652
rect 568574 220600 568580 220652
rect 568632 220640 568638 220652
rect 569770 220640 569776 220652
rect 568632 220612 569776 220640
rect 568632 220600 568638 220612
rect 569770 220600 569776 220612
rect 569828 220600 569834 220652
rect 569954 220600 569960 220652
rect 570012 220640 570018 220652
rect 610526 220640 610532 220652
rect 570012 220612 610532 220640
rect 570012 220600 570018 220612
rect 610526 220600 610532 220612
rect 610584 220600 610590 220652
rect 544930 220504 544936 220516
rect 543752 220476 544936 220504
rect 544930 220464 544936 220476
rect 544988 220464 544994 220516
rect 553026 220504 553032 220516
rect 548444 220476 553032 220504
rect 64598 220328 64604 220380
rect 64656 220368 64662 220380
rect 141970 220368 141976 220380
rect 64656 220340 141976 220368
rect 64656 220328 64662 220340
rect 141970 220328 141976 220340
rect 142028 220328 142034 220380
rect 151630 220368 151636 220380
rect 142126 220340 151636 220368
rect 73062 220192 73068 220244
rect 73120 220232 73126 220244
rect 142126 220232 142154 220340
rect 151630 220328 151636 220340
rect 151688 220328 151694 220380
rect 151768 220328 151774 220380
rect 151826 220368 151832 220380
rect 208578 220368 208584 220380
rect 151826 220340 208584 220368
rect 151826 220328 151832 220340
rect 208578 220328 208584 220340
rect 208636 220328 208642 220380
rect 213822 220328 213828 220380
rect 213880 220368 213886 220380
rect 262398 220368 262404 220380
rect 213880 220340 262404 220368
rect 213880 220328 213886 220340
rect 262398 220328 262404 220340
rect 262456 220328 262462 220380
rect 262674 220328 262680 220380
rect 262732 220368 262738 220380
rect 264238 220368 264244 220380
rect 262732 220340 264244 220368
rect 262732 220328 262738 220340
rect 264238 220328 264244 220340
rect 264296 220328 264302 220380
rect 264606 220328 264612 220380
rect 264664 220368 264670 220380
rect 269298 220368 269304 220380
rect 264664 220340 269304 220368
rect 264664 220328 264670 220340
rect 269298 220328 269304 220340
rect 269356 220328 269362 220380
rect 273438 220328 273444 220380
rect 273496 220368 273502 220380
rect 309226 220368 309232 220380
rect 273496 220340 309232 220368
rect 273496 220328 273502 220340
rect 309226 220328 309232 220340
rect 309284 220328 309290 220380
rect 316494 220328 316500 220380
rect 316552 220368 316558 220380
rect 342898 220368 342904 220380
rect 316552 220340 342904 220368
rect 316552 220328 316558 220340
rect 342898 220328 342904 220340
rect 342956 220328 342962 220380
rect 351270 220328 351276 220380
rect 351328 220368 351334 220380
rect 369302 220368 369308 220380
rect 351328 220340 369308 220368
rect 351328 220328 351334 220340
rect 369302 220328 369308 220340
rect 369360 220328 369366 220380
rect 376938 220328 376944 220380
rect 376996 220368 377002 220380
rect 388438 220368 388444 220380
rect 376996 220340 388444 220368
rect 376996 220328 377002 220340
rect 388438 220328 388444 220340
rect 388496 220328 388502 220380
rect 436278 220328 436284 220380
rect 436336 220368 436342 220380
rect 437014 220368 437020 220380
rect 436336 220340 437020 220368
rect 436336 220328 436342 220340
rect 437014 220328 437020 220340
rect 437072 220328 437078 220380
rect 473170 220328 473176 220380
rect 473228 220368 473234 220380
rect 481174 220368 481180 220380
rect 473228 220340 481180 220368
rect 473228 220328 473234 220340
rect 481174 220328 481180 220340
rect 481232 220328 481238 220380
rect 496446 220328 496452 220380
rect 496504 220368 496510 220380
rect 509326 220368 509332 220380
rect 496504 220340 509332 220368
rect 496504 220328 496510 220340
rect 509326 220328 509332 220340
rect 509384 220328 509390 220380
rect 515398 220328 515404 220380
rect 515456 220368 515462 220380
rect 530026 220368 530032 220380
rect 515456 220340 530032 220368
rect 515456 220328 515462 220340
rect 530026 220328 530032 220340
rect 530084 220328 530090 220380
rect 531130 220328 531136 220380
rect 531188 220368 531194 220380
rect 548444 220368 548472 220476
rect 553026 220464 553032 220476
rect 553084 220464 553090 220516
rect 553854 220464 553860 220516
rect 553912 220504 553918 220516
rect 608594 220504 608600 220516
rect 553912 220476 608600 220504
rect 553912 220464 553918 220476
rect 608594 220464 608600 220476
rect 608652 220464 608658 220516
rect 647234 220464 647240 220516
rect 647292 220504 647298 220516
rect 651466 220504 651472 220516
rect 647292 220476 651472 220504
rect 647292 220464 647298 220476
rect 651466 220464 651472 220476
rect 651524 220464 651530 220516
rect 554038 220368 554044 220380
rect 531188 220340 548472 220368
rect 548536 220340 554044 220368
rect 531188 220328 531194 220340
rect 73120 220204 142154 220232
rect 73120 220192 73126 220204
rect 144270 220192 144276 220244
rect 144328 220232 144334 220244
rect 146754 220232 146760 220244
rect 144328 220204 146760 220232
rect 144328 220192 144334 220204
rect 146754 220192 146760 220204
rect 146812 220192 146818 220244
rect 146938 220192 146944 220244
rect 146996 220232 147002 220244
rect 156598 220232 156604 220244
rect 146996 220204 156604 220232
rect 146996 220192 147002 220204
rect 156598 220192 156604 220204
rect 156656 220192 156662 220244
rect 156782 220192 156788 220244
rect 156840 220232 156846 220244
rect 215938 220232 215944 220244
rect 156840 220204 215944 220232
rect 156840 220192 156846 220204
rect 215938 220192 215944 220204
rect 215996 220192 216002 220244
rect 217134 220192 217140 220244
rect 217192 220232 217198 220244
rect 265158 220232 265164 220244
rect 217192 220204 265164 220232
rect 217192 220192 217198 220204
rect 265158 220192 265164 220204
rect 265216 220192 265222 220244
rect 267642 220192 267648 220244
rect 267700 220232 267706 220244
rect 306834 220232 306840 220244
rect 267700 220204 306840 220232
rect 267700 220192 267706 220204
rect 306834 220192 306840 220204
rect 306892 220192 306898 220244
rect 309042 220192 309048 220244
rect 309100 220232 309106 220244
rect 339678 220232 339684 220244
rect 309100 220204 339684 220232
rect 309100 220192 309106 220204
rect 339678 220192 339684 220204
rect 339736 220192 339742 220244
rect 342990 220192 342996 220244
rect 343048 220232 343054 220244
rect 363322 220232 363328 220244
rect 343048 220204 363328 220232
rect 343048 220192 343054 220204
rect 363322 220192 363328 220204
rect 363380 220192 363386 220244
rect 363690 220192 363696 220244
rect 363748 220232 363754 220244
rect 381078 220232 381084 220244
rect 363748 220204 381084 220232
rect 363748 220192 363754 220204
rect 381078 220192 381084 220204
rect 381136 220192 381142 220244
rect 388438 220192 388444 220244
rect 388496 220232 388502 220244
rect 400950 220232 400956 220244
rect 388496 220204 400956 220232
rect 388496 220192 388502 220204
rect 400950 220192 400956 220204
rect 401008 220192 401014 220244
rect 430114 220192 430120 220244
rect 430172 220232 430178 220244
rect 432046 220232 432052 220244
rect 430172 220204 432052 220232
rect 430172 220192 430178 220204
rect 432046 220192 432052 220204
rect 432104 220192 432110 220244
rect 459462 220192 459468 220244
rect 459520 220232 459526 220244
rect 465442 220232 465448 220244
rect 459520 220204 465448 220232
rect 459520 220192 459526 220204
rect 465442 220192 465448 220204
rect 465500 220192 465506 220244
rect 472986 220192 472992 220244
rect 473044 220232 473050 220244
rect 482002 220232 482008 220244
rect 473044 220204 482008 220232
rect 473044 220192 473050 220204
rect 482002 220192 482008 220204
rect 482060 220192 482066 220244
rect 482922 220192 482928 220244
rect 482980 220232 482986 220244
rect 495342 220232 495348 220244
rect 482980 220204 495348 220232
rect 482980 220192 482986 220204
rect 495342 220192 495348 220204
rect 495400 220192 495406 220244
rect 497458 220192 497464 220244
rect 497516 220232 497522 220244
rect 515214 220232 515220 220244
rect 497516 220204 515220 220232
rect 497516 220192 497522 220204
rect 515214 220192 515220 220204
rect 515272 220192 515278 220244
rect 528370 220192 528376 220244
rect 528428 220232 528434 220244
rect 548536 220232 548564 220340
rect 554038 220328 554044 220340
rect 554096 220328 554102 220380
rect 563054 220328 563060 220380
rect 563112 220368 563118 220380
rect 610066 220368 610072 220380
rect 563112 220340 610072 220368
rect 563112 220328 563118 220340
rect 610066 220328 610072 220340
rect 610124 220328 610130 220380
rect 560754 220260 560760 220312
rect 560812 220300 560818 220312
rect 562870 220300 562876 220312
rect 560812 220272 562876 220300
rect 560812 220260 560818 220272
rect 562870 220260 562876 220272
rect 562928 220260 562934 220312
rect 528428 220204 548564 220232
rect 528428 220192 528434 220204
rect 548702 220192 548708 220244
rect 548760 220232 548766 220244
rect 548760 220204 558224 220232
rect 548760 220192 548766 220204
rect 101214 220056 101220 220108
rect 101272 220096 101278 220108
rect 166948 220096 166954 220108
rect 101272 220068 166954 220096
rect 101272 220056 101278 220068
rect 166948 220056 166954 220068
rect 167006 220056 167012 220108
rect 167086 220056 167092 220108
rect 167144 220096 167150 220108
rect 167144 220068 181392 220096
rect 167144 220056 167150 220068
rect 114462 219920 114468 219972
rect 114520 219960 114526 219972
rect 180886 219960 180892 219972
rect 114520 219932 180892 219960
rect 114520 219920 114526 219932
rect 180886 219920 180892 219932
rect 180944 219920 180950 219972
rect 181364 219960 181392 220068
rect 181530 220056 181536 220108
rect 181588 220096 181594 220108
rect 229278 220096 229284 220108
rect 181588 220068 229284 220096
rect 181588 220056 181594 220068
rect 229278 220056 229284 220068
rect 229336 220056 229342 220108
rect 230198 220056 230204 220108
rect 230256 220096 230262 220108
rect 275278 220096 275284 220108
rect 230256 220068 275284 220096
rect 230256 220056 230262 220068
rect 275278 220056 275284 220068
rect 275336 220056 275342 220108
rect 276750 220056 276756 220108
rect 276808 220096 276814 220108
rect 311342 220096 311348 220108
rect 276808 220068 311348 220096
rect 276808 220056 276814 220068
rect 311342 220056 311348 220068
rect 311400 220056 311406 220108
rect 328914 220056 328920 220108
rect 328972 220096 328978 220108
rect 354766 220096 354772 220108
rect 328972 220068 354772 220096
rect 328972 220056 328978 220068
rect 354766 220056 354772 220068
rect 354824 220056 354830 220108
rect 355410 220056 355416 220108
rect 355468 220096 355474 220108
rect 375558 220096 375564 220108
rect 355468 220068 375564 220096
rect 355468 220056 355474 220068
rect 375558 220056 375564 220068
rect 375616 220056 375622 220108
rect 379422 220056 379428 220108
rect 379480 220096 379486 220108
rect 392118 220096 392124 220108
rect 379480 220068 392124 220096
rect 379480 220056 379486 220068
rect 392118 220056 392124 220068
rect 392176 220056 392182 220108
rect 395982 220056 395988 220108
rect 396040 220096 396046 220108
rect 404722 220096 404728 220108
rect 396040 220068 404728 220096
rect 396040 220056 396046 220068
rect 404722 220056 404728 220068
rect 404780 220056 404786 220108
rect 421650 220056 421656 220108
rect 421708 220096 421714 220108
rect 426710 220096 426716 220108
rect 421708 220068 426716 220096
rect 421708 220056 421714 220068
rect 426710 220056 426716 220068
rect 426768 220056 426774 220108
rect 431954 220056 431960 220108
rect 432012 220096 432018 220108
rect 434806 220096 434812 220108
rect 432012 220068 434812 220096
rect 432012 220056 432018 220068
rect 434806 220056 434812 220068
rect 434864 220056 434870 220108
rect 478322 220056 478328 220108
rect 478380 220096 478386 220108
rect 489454 220096 489460 220108
rect 478380 220068 489460 220096
rect 478380 220056 478386 220068
rect 489454 220056 489460 220068
rect 489512 220056 489518 220108
rect 489638 220056 489644 220108
rect 489696 220096 489702 220108
rect 504358 220096 504364 220108
rect 489696 220068 504364 220096
rect 489696 220056 489702 220068
rect 504358 220056 504364 220068
rect 504416 220056 504422 220108
rect 513098 220056 513104 220108
rect 513156 220096 513162 220108
rect 534166 220096 534172 220108
rect 513156 220068 534172 220096
rect 513156 220056 513162 220068
rect 534166 220056 534172 220068
rect 534224 220056 534230 220108
rect 538122 220056 538128 220108
rect 538180 220096 538186 220108
rect 557994 220096 558000 220108
rect 538180 220068 558000 220096
rect 538180 220056 538186 220068
rect 557994 220056 558000 220068
rect 558052 220056 558058 220108
rect 558196 220028 558224 220204
rect 576762 220192 576768 220244
rect 576820 220232 576826 220244
rect 611630 220232 611636 220244
rect 576820 220204 611636 220232
rect 576820 220192 576826 220204
rect 611630 220192 611636 220204
rect 611688 220192 611694 220244
rect 668946 220192 668952 220244
rect 669004 220232 669010 220244
rect 669004 220204 669176 220232
rect 669004 220192 669010 220204
rect 558362 220124 558368 220176
rect 558420 220164 558426 220176
rect 576578 220164 576584 220176
rect 558420 220136 576584 220164
rect 558420 220124 558426 220136
rect 576578 220124 576584 220136
rect 576636 220124 576642 220176
rect 582466 220056 582472 220108
rect 582524 220096 582530 220108
rect 633434 220096 633440 220108
rect 582524 220068 633440 220096
rect 582524 220056 582530 220068
rect 633434 220056 633440 220068
rect 633492 220056 633498 220108
rect 669148 220040 669176 220204
rect 576762 220028 576768 220040
rect 558196 220000 576768 220028
rect 576762 219988 576768 220000
rect 576820 219988 576826 220040
rect 576946 219988 576952 220040
rect 577004 220028 577010 220040
rect 581638 220028 581644 220040
rect 577004 220000 581644 220028
rect 577004 219988 577010 220000
rect 581638 219988 581644 220000
rect 581696 219988 581702 220040
rect 581822 219988 581828 220040
rect 581880 220028 581886 220040
rect 582328 220028 582334 220040
rect 581880 220000 582334 220028
rect 581880 219988 581886 220000
rect 582328 219988 582334 220000
rect 582386 219988 582392 220040
rect 669130 219988 669136 220040
rect 669188 219988 669194 220040
rect 190454 219960 190460 219972
rect 181364 219932 190460 219960
rect 190454 219920 190460 219932
rect 190512 219920 190518 219972
rect 190638 219920 190644 219972
rect 190696 219960 190702 219972
rect 244458 219960 244464 219972
rect 190696 219932 244464 219960
rect 190696 219920 190702 219932
rect 244458 219920 244464 219932
rect 244516 219920 244522 219972
rect 253566 219920 253572 219972
rect 253624 219960 253630 219972
rect 293310 219960 293316 219972
rect 253624 219932 293316 219960
rect 253624 219920 253630 219932
rect 293310 219920 293316 219932
rect 293368 219920 293374 219972
rect 530026 219852 530032 219904
rect 530084 219892 530090 219904
rect 558362 219892 558368 219904
rect 530084 219864 558368 219892
rect 530084 219852 530090 219864
rect 558362 219852 558368 219864
rect 558420 219852 558426 219904
rect 558730 219852 558736 219904
rect 558788 219892 558794 219904
rect 600958 219892 600964 219904
rect 558788 219864 600964 219892
rect 558788 219852 558794 219864
rect 600958 219852 600964 219864
rect 601016 219852 601022 219904
rect 601142 219852 601148 219904
rect 601200 219892 601206 219904
rect 619818 219892 619824 219904
rect 601200 219864 619824 219892
rect 601200 219852 601206 219864
rect 619818 219852 619824 219864
rect 619876 219852 619882 219904
rect 121086 219784 121092 219836
rect 121144 219824 121150 219836
rect 121144 219796 122834 219824
rect 121144 219784 121150 219796
rect 122806 219688 122834 219796
rect 134334 219784 134340 219836
rect 134392 219824 134398 219836
rect 140774 219824 140780 219836
rect 134392 219796 140780 219824
rect 134392 219784 134398 219796
rect 140774 219784 140780 219796
rect 140832 219784 140838 219836
rect 140958 219784 140964 219836
rect 141016 219824 141022 219836
rect 141970 219824 141976 219836
rect 141016 219796 141976 219824
rect 141016 219784 141022 219796
rect 141970 219784 141976 219796
rect 142028 219784 142034 219836
rect 142154 219784 142160 219836
rect 142212 219824 142218 219836
rect 200206 219824 200212 219836
rect 142212 219796 200212 219824
rect 142212 219784 142218 219796
rect 200206 219784 200212 219796
rect 200264 219784 200270 219836
rect 200574 219784 200580 219836
rect 200632 219824 200638 219836
rect 252738 219824 252744 219836
rect 200632 219796 252744 219824
rect 200632 219784 200638 219796
rect 252738 219784 252744 219796
rect 252796 219784 252802 219836
rect 286686 219784 286692 219836
rect 286744 219824 286750 219836
rect 319070 219824 319076 219836
rect 286744 219796 319076 219824
rect 286744 219784 286750 219796
rect 319070 219784 319076 219796
rect 319128 219784 319134 219836
rect 527542 219716 527548 219768
rect 527600 219756 527606 219768
rect 548702 219756 548708 219768
rect 527600 219728 548708 219756
rect 527600 219716 527606 219728
rect 548702 219716 548708 219728
rect 548760 219716 548766 219768
rect 548886 219716 548892 219768
rect 548944 219756 548950 219768
rect 548944 219728 601372 219756
rect 548944 219716 548950 219728
rect 146938 219688 146944 219700
rect 122806 219660 146944 219688
rect 146938 219648 146944 219660
rect 146996 219648 147002 219700
rect 205818 219688 205824 219700
rect 147140 219660 205824 219688
rect 69750 219512 69756 219564
rect 69808 219552 69814 219564
rect 142154 219552 142160 219564
rect 69808 219524 142160 219552
rect 69808 219512 69814 219524
rect 142154 219512 142160 219524
rect 142212 219512 142218 219564
rect 142338 219512 142344 219564
rect 142396 219552 142402 219564
rect 147140 219552 147168 219660
rect 205818 219648 205824 219660
rect 205876 219648 205882 219700
rect 207198 219648 207204 219700
rect 207256 219688 207262 219700
rect 257246 219688 257252 219700
rect 207256 219660 257252 219688
rect 207256 219648 207262 219660
rect 257246 219648 257252 219660
rect 257304 219648 257310 219700
rect 464982 219580 464988 219632
rect 465040 219620 465046 219632
rect 472066 219620 472072 219632
rect 465040 219592 472072 219620
rect 465040 219580 465046 219592
rect 472066 219580 472072 219592
rect 472124 219580 472130 219632
rect 506014 219580 506020 219632
rect 506072 219620 506078 219632
rect 576762 219620 576768 219632
rect 506072 219592 576768 219620
rect 506072 219580 506078 219592
rect 576762 219580 576768 219592
rect 576820 219580 576826 219632
rect 581638 219580 581644 219632
rect 581696 219620 581702 219632
rect 582374 219620 582380 219632
rect 581696 219592 582380 219620
rect 581696 219580 581702 219592
rect 582374 219580 582380 219592
rect 582432 219580 582438 219632
rect 582650 219580 582656 219632
rect 582708 219620 582714 219632
rect 601142 219620 601148 219632
rect 582708 219592 601148 219620
rect 582708 219580 582714 219592
rect 601142 219580 601148 219592
rect 601200 219580 601206 219632
rect 601344 219620 601372 219728
rect 601510 219716 601516 219768
rect 601568 219756 601574 219768
rect 620002 219756 620008 219768
rect 601568 219728 620008 219756
rect 601568 219716 601574 219728
rect 620002 219716 620008 219728
rect 620060 219716 620066 219768
rect 607490 219620 607496 219632
rect 601344 219592 607496 219620
rect 607490 219580 607496 219592
rect 607548 219580 607554 219632
rect 142396 219524 147168 219552
rect 142396 219512 142402 219524
rect 147766 219512 147772 219564
rect 147824 219552 147830 219564
rect 150710 219552 150716 219564
rect 147824 219524 150716 219552
rect 147824 219512 147830 219524
rect 150710 219512 150716 219524
rect 150768 219512 150774 219564
rect 150894 219512 150900 219564
rect 150952 219552 150958 219564
rect 214006 219552 214012 219564
rect 150952 219524 214012 219552
rect 150952 219512 150958 219524
rect 214006 219512 214012 219524
rect 214064 219512 214070 219564
rect 270770 219512 270776 219564
rect 270828 219552 270834 219564
rect 279142 219552 279148 219564
rect 270828 219524 279148 219552
rect 270828 219512 270834 219524
rect 279142 219512 279148 219524
rect 279200 219512 279206 219564
rect 289814 219512 289820 219564
rect 289872 219552 289878 219564
rect 289872 219524 290136 219552
rect 289872 219512 289878 219524
rect 63954 219376 63960 219428
rect 64012 219416 64018 219428
rect 64874 219416 64880 219428
rect 64012 219388 64880 219416
rect 64012 219376 64018 219388
rect 64874 219376 64880 219388
rect 64932 219376 64938 219428
rect 105814 219394 105820 219446
rect 105872 219434 105878 219446
rect 105872 219416 106182 219434
rect 147122 219416 147128 219428
rect 105872 219406 147128 219416
rect 105872 219394 105878 219406
rect 106154 219388 147128 219406
rect 147122 219376 147128 219388
rect 147180 219376 147186 219428
rect 159818 219376 159824 219428
rect 159876 219416 159882 219428
rect 204530 219416 204536 219428
rect 159876 219388 204536 219416
rect 159876 219376 159882 219388
rect 204530 219376 204536 219388
rect 204588 219376 204594 219428
rect 209682 219376 209688 219428
rect 209740 219416 209746 219428
rect 210418 219416 210424 219428
rect 209740 219388 210424 219416
rect 209740 219376 209746 219388
rect 210418 219376 210424 219388
rect 210476 219376 210482 219428
rect 212994 219376 213000 219428
rect 213052 219416 213058 219428
rect 258074 219416 258080 219428
rect 213052 219388 258080 219416
rect 213052 219376 213058 219388
rect 258074 219376 258080 219388
rect 258132 219376 258138 219428
rect 272886 219376 272892 219428
rect 272944 219416 272950 219428
rect 290108 219416 290136 219524
rect 366726 219512 366732 219564
rect 366784 219552 366790 219564
rect 366784 219524 367048 219552
rect 366784 219512 366790 219524
rect 367020 219434 367048 219524
rect 576964 219524 579752 219552
rect 405918 219444 405924 219496
rect 405976 219484 405982 219496
rect 412726 219484 412732 219496
rect 405976 219456 412732 219484
rect 405976 219444 405982 219456
rect 412726 219444 412732 219456
rect 412784 219444 412790 219496
rect 421006 219484 421012 219496
rect 418172 219456 421012 219484
rect 297542 219416 297548 219428
rect 272944 219388 290044 219416
rect 290108 219388 297548 219416
rect 272944 219376 272950 219388
rect 106918 219280 106924 219292
rect 64846 219252 106924 219280
rect 63126 219104 63132 219156
rect 63184 219144 63190 219156
rect 64846 219144 64874 219252
rect 106918 219240 106924 219252
rect 106976 219240 106982 219292
rect 113634 219240 113640 219292
rect 113692 219280 113698 219292
rect 156230 219280 156236 219292
rect 113692 219252 156236 219280
rect 113692 219240 113698 219252
rect 156230 219240 156236 219252
rect 156288 219240 156294 219292
rect 162486 219240 162492 219292
rect 162544 219280 162550 219292
rect 166534 219280 166540 219292
rect 162544 219252 166540 219280
rect 162544 219240 162550 219252
rect 166534 219240 166540 219252
rect 166592 219240 166598 219292
rect 167454 219240 167460 219292
rect 167512 219280 167518 219292
rect 168190 219280 168196 219292
rect 167512 219252 168196 219280
rect 167512 219240 167518 219252
rect 168190 219240 168196 219252
rect 168248 219240 168254 219292
rect 169110 219240 169116 219292
rect 169168 219280 169174 219292
rect 169662 219280 169668 219292
rect 169168 219252 169668 219280
rect 169168 219240 169174 219252
rect 169662 219240 169668 219252
rect 169720 219240 169726 219292
rect 169938 219240 169944 219292
rect 169996 219280 170002 219292
rect 171042 219280 171048 219292
rect 169996 219252 171048 219280
rect 169996 219240 170002 219252
rect 171042 219240 171048 219252
rect 171100 219240 171106 219292
rect 171594 219240 171600 219292
rect 171652 219280 171658 219292
rect 172146 219280 172152 219292
rect 171652 219252 172152 219280
rect 171652 219240 171658 219252
rect 172146 219240 172152 219252
rect 172204 219240 172210 219292
rect 172422 219240 172428 219292
rect 172480 219280 172486 219292
rect 173158 219280 173164 219292
rect 172480 219252 173164 219280
rect 172480 219240 172486 219252
rect 173158 219240 173164 219252
rect 173216 219240 173222 219292
rect 182358 219240 182364 219292
rect 182416 219280 182422 219292
rect 189718 219280 189724 219292
rect 182416 219252 189724 219280
rect 182416 219240 182422 219252
rect 189718 219240 189724 219252
rect 189776 219240 189782 219292
rect 192846 219240 192852 219292
rect 192904 219280 192910 219292
rect 198182 219280 198188 219292
rect 192904 219252 198188 219280
rect 192904 219240 192910 219252
rect 198182 219240 198188 219252
rect 198240 219240 198246 219292
rect 198918 219240 198924 219292
rect 198976 219280 198982 219292
rect 200022 219280 200028 219292
rect 198976 219252 200028 219280
rect 198976 219240 198982 219252
rect 200022 219240 200028 219252
rect 200080 219240 200086 219292
rect 202598 219240 202604 219292
rect 202656 219280 202662 219292
rect 207658 219280 207664 219292
rect 202656 219252 207664 219280
rect 202656 219240 202662 219252
rect 207658 219240 207664 219252
rect 207716 219240 207722 219292
rect 211338 219240 211344 219292
rect 211396 219280 211402 219292
rect 218054 219280 218060 219292
rect 211396 219252 218060 219280
rect 211396 219240 211402 219252
rect 218054 219240 218060 219252
rect 218112 219240 218118 219292
rect 239490 219240 239496 219292
rect 239548 219280 239554 219292
rect 272702 219280 272708 219292
rect 239548 219252 272708 219280
rect 239548 219240 239554 219252
rect 272702 219240 272708 219252
rect 272760 219240 272766 219292
rect 289814 219280 289820 219292
rect 277366 219252 289820 219280
rect 63184 219116 64874 219144
rect 63184 219104 63190 219116
rect 70578 219104 70584 219156
rect 70636 219144 70642 219156
rect 117958 219144 117964 219156
rect 70636 219116 117964 219144
rect 70636 219104 70642 219116
rect 117958 219104 117964 219116
rect 118016 219104 118022 219156
rect 132586 219104 132592 219156
rect 132644 219144 132650 219156
rect 177482 219144 177488 219156
rect 132644 219116 177488 219144
rect 132644 219104 132650 219116
rect 177482 219104 177488 219116
rect 177540 219104 177546 219156
rect 179046 219104 179052 219156
rect 179104 219144 179110 219156
rect 196618 219144 196624 219156
rect 179104 219116 196624 219144
rect 179104 219104 179110 219116
rect 196618 219104 196624 219116
rect 196676 219104 196682 219156
rect 199746 219104 199752 219156
rect 199804 219144 199810 219156
rect 243538 219144 243544 219156
rect 199804 219116 243544 219144
rect 199804 219104 199810 219116
rect 243538 219104 243544 219116
rect 243596 219104 243602 219156
rect 272334 219104 272340 219156
rect 272392 219144 272398 219156
rect 277366 219144 277394 219252
rect 289814 219240 289820 219252
rect 289872 219240 289878 219292
rect 290016 219280 290044 219388
rect 297542 219376 297548 219388
rect 297600 219376 297606 219428
rect 304074 219376 304080 219428
rect 304132 219416 304138 219428
rect 308398 219416 308404 219428
rect 304132 219388 308404 219416
rect 304132 219376 304138 219388
rect 308398 219376 308404 219388
rect 308456 219376 308462 219428
rect 320634 219376 320640 219428
rect 320692 219416 320698 219428
rect 320692 219388 335354 219416
rect 320692 219376 320698 219388
rect 290016 219252 291884 219280
rect 272392 219116 277394 219144
rect 272392 219104 272398 219116
rect 279050 219104 279056 219156
rect 279108 219144 279114 219156
rect 286318 219144 286324 219156
rect 279108 219116 286324 219144
rect 279108 219104 279114 219116
rect 286318 219104 286324 219116
rect 286376 219104 286382 219156
rect 291856 219144 291884 219252
rect 292022 219240 292028 219292
rect 292080 219280 292086 219292
rect 313918 219280 313924 219292
rect 292080 219252 313924 219280
rect 292080 219240 292086 219252
rect 313918 219240 313924 219252
rect 313976 219240 313982 219292
rect 335326 219280 335354 219388
rect 341334 219376 341340 219428
rect 341392 219416 341398 219428
rect 342254 219416 342260 219428
rect 341392 219388 342260 219416
rect 341392 219376 341398 219388
rect 342254 219376 342260 219388
rect 342312 219376 342318 219428
rect 343818 219376 343824 219428
rect 343876 219416 343882 219428
rect 347038 219416 347044 219428
rect 343876 219388 347044 219416
rect 343876 219376 343882 219388
rect 347038 219376 347044 219388
rect 347096 219376 347102 219428
rect 366174 219376 366180 219428
rect 366232 219416 366238 219428
rect 366928 219416 367048 219434
rect 366232 219406 367048 219416
rect 366232 219388 366956 219406
rect 366232 219376 366238 219388
rect 399294 219376 399300 219428
rect 399352 219416 399358 219428
rect 400214 219416 400220 219428
rect 399352 219388 400220 219416
rect 399352 219376 399358 219388
rect 400214 219376 400220 219388
rect 400272 219376 400278 219428
rect 415854 219376 415860 219428
rect 415912 219416 415918 219428
rect 416774 219416 416780 219428
rect 415912 219388 416780 219416
rect 415912 219376 415918 219388
rect 416774 219376 416780 219388
rect 416832 219376 416838 219428
rect 417510 219376 417516 219428
rect 417568 219416 417574 219428
rect 418172 219416 418200 219456
rect 421006 219444 421012 219456
rect 421064 219444 421070 219496
rect 501046 219444 501052 219496
rect 501104 219484 501110 219496
rect 576964 219484 576992 219524
rect 501104 219456 576992 219484
rect 579724 219484 579752 219524
rect 579724 219456 591712 219484
rect 501104 219444 501110 219456
rect 417568 219388 418200 219416
rect 577130 219394 577136 219446
rect 577188 219434 577194 219446
rect 577188 219406 579614 219434
rect 577188 219394 577194 219406
rect 417568 219376 417574 219388
rect 579586 219348 579614 219406
rect 582650 219348 582656 219360
rect 579586 219320 582656 219348
rect 582650 219308 582656 219320
rect 582708 219308 582714 219360
rect 591684 219348 591712 219456
rect 591942 219444 591948 219496
rect 592000 219484 592006 219496
rect 600130 219484 600136 219496
rect 592000 219456 600136 219484
rect 592000 219444 592006 219456
rect 600130 219444 600136 219456
rect 600188 219444 600194 219496
rect 600958 219444 600964 219496
rect 601016 219484 601022 219496
rect 607306 219484 607312 219496
rect 601016 219456 607312 219484
rect 601016 219444 601022 219456
rect 607306 219444 607312 219456
rect 607364 219444 607370 219496
rect 596818 219348 596824 219360
rect 591684 219320 596824 219348
rect 596818 219308 596824 219320
rect 596876 219308 596882 219360
rect 345290 219280 345296 219292
rect 335326 219252 345296 219280
rect 345290 219240 345296 219252
rect 345348 219240 345354 219292
rect 419166 219240 419172 219292
rect 419224 219280 419230 219292
rect 422662 219280 422668 219292
rect 419224 219252 422668 219280
rect 419224 219240 419230 219252
rect 422662 219240 422668 219252
rect 422720 219240 422726 219292
rect 552474 219240 552480 219292
rect 552532 219280 552538 219292
rect 574738 219280 574744 219292
rect 552532 219252 574744 219280
rect 552532 219240 552538 219252
rect 574738 219240 574744 219252
rect 574796 219240 574802 219292
rect 582466 219172 582472 219224
rect 582524 219212 582530 219224
rect 597922 219212 597928 219224
rect 582524 219184 597928 219212
rect 582524 219172 582530 219184
rect 597922 219172 597928 219184
rect 597980 219172 597986 219224
rect 291856 219116 291976 219144
rect 62298 218968 62304 219020
rect 62356 219008 62362 219020
rect 72418 219008 72424 219020
rect 62356 218980 72424 219008
rect 62356 218968 62362 218980
rect 72418 218968 72424 218980
rect 72476 218968 72482 219020
rect 77202 218968 77208 219020
rect 77260 219008 77266 219020
rect 140038 219008 140044 219020
rect 77260 218980 140044 219008
rect 77260 218968 77266 218980
rect 140038 218968 140044 218980
rect 140096 218968 140102 219020
rect 142430 218968 142436 219020
rect 142488 219008 142494 219020
rect 143718 219008 143724 219020
rect 142488 218980 143724 219008
rect 142488 218968 142494 218980
rect 143718 218968 143724 218980
rect 143776 218968 143782 219020
rect 146754 218968 146760 219020
rect 146812 219008 146818 219020
rect 150434 219008 150440 219020
rect 146812 218980 150440 219008
rect 146812 218968 146818 218980
rect 150434 218968 150440 218980
rect 150492 218968 150498 219020
rect 153378 218968 153384 219020
rect 153436 219008 153442 219020
rect 203518 219008 203524 219020
rect 153436 218980 203524 219008
rect 153436 218968 153442 218980
rect 203518 218968 203524 218980
rect 203576 218968 203582 219020
rect 206370 218968 206376 219020
rect 206428 219008 206434 219020
rect 253382 219008 253388 219020
rect 206428 218980 253388 219008
rect 206428 218968 206434 218980
rect 253382 218968 253388 218980
rect 253440 218968 253446 219020
rect 259178 218968 259184 219020
rect 259236 219008 259242 219020
rect 291654 219008 291660 219020
rect 259236 218980 291660 219008
rect 259236 218968 259242 218980
rect 291654 218968 291660 218980
rect 291712 218968 291718 219020
rect 291948 219008 291976 219116
rect 295794 219104 295800 219156
rect 295852 219144 295858 219156
rect 296714 219144 296720 219156
rect 295852 219116 296720 219144
rect 295852 219104 295858 219116
rect 296714 219104 296720 219116
rect 296772 219104 296778 219156
rect 300486 219104 300492 219156
rect 300544 219144 300550 219156
rect 322106 219144 322112 219156
rect 300544 219116 322112 219144
rect 300544 219104 300550 219116
rect 322106 219104 322112 219116
rect 322164 219104 322170 219156
rect 325326 219104 325332 219156
rect 325384 219144 325390 219156
rect 327718 219144 327724 219156
rect 325384 219116 327724 219144
rect 325384 219104 325390 219116
rect 327718 219104 327724 219116
rect 327776 219104 327782 219156
rect 340506 219104 340512 219156
rect 340564 219144 340570 219156
rect 352558 219144 352564 219156
rect 340564 219116 352564 219144
rect 340564 219104 340570 219116
rect 352558 219104 352564 219116
rect 352616 219104 352622 219156
rect 362034 219104 362040 219156
rect 362092 219144 362098 219156
rect 370958 219144 370964 219156
rect 362092 219116 370964 219144
rect 362092 219104 362098 219116
rect 370958 219104 370964 219116
rect 371016 219104 371022 219156
rect 543734 219104 543740 219156
rect 543792 219144 543798 219156
rect 549070 219144 549076 219156
rect 543792 219116 549076 219144
rect 543792 219104 543798 219116
rect 549070 219104 549076 219116
rect 549128 219104 549134 219156
rect 553026 219104 553032 219156
rect 553084 219144 553090 219156
rect 556614 219144 556620 219156
rect 553084 219116 556620 219144
rect 553084 219104 553090 219116
rect 556614 219104 556620 219116
rect 556672 219104 556678 219156
rect 561674 219104 561680 219156
rect 561732 219144 561738 219156
rect 562410 219144 562416 219156
rect 561732 219116 562416 219144
rect 561732 219104 561738 219116
rect 562410 219104 562416 219116
rect 562468 219144 562474 219156
rect 571334 219144 571340 219156
rect 562468 219116 571340 219144
rect 562468 219104 562474 219116
rect 571334 219104 571340 219116
rect 571392 219104 571398 219156
rect 571518 219104 571524 219156
rect 571576 219144 571582 219156
rect 571576 219116 576854 219144
rect 571576 219104 571582 219116
rect 297358 219008 297364 219020
rect 291948 218980 297364 219008
rect 297358 218968 297364 218980
rect 297416 218968 297422 219020
rect 307386 218968 307392 219020
rect 307444 219008 307450 219020
rect 331858 219008 331864 219020
rect 307444 218980 331864 219008
rect 307444 218968 307450 218980
rect 331858 218968 331864 218980
rect 331916 218968 331922 219020
rect 333422 218968 333428 219020
rect 333480 219008 333486 219020
rect 355226 219008 355232 219020
rect 333480 218980 355232 219008
rect 333480 218968 333486 218980
rect 355226 218968 355232 218980
rect 355284 218968 355290 219020
rect 357066 218968 357072 219020
rect 357124 219008 357130 219020
rect 369118 219008 369124 219020
rect 357124 218980 369124 219008
rect 357124 218968 357130 218980
rect 369118 218968 369124 218980
rect 369176 218968 369182 219020
rect 370314 218968 370320 219020
rect 370372 219008 370378 219020
rect 380066 219008 380072 219020
rect 370372 218980 380072 219008
rect 370372 218968 370378 218980
rect 380066 218968 380072 218980
rect 380124 218968 380130 219020
rect 380250 218968 380256 219020
rect 380308 219008 380314 219020
rect 388622 219008 388628 219020
rect 380308 218980 388628 219008
rect 380308 218968 380314 218980
rect 388622 218968 388628 218980
rect 388680 218968 388686 219020
rect 572070 219008 572076 219020
rect 543706 218980 572076 219008
rect 50706 218832 50712 218884
rect 50764 218872 50770 218884
rect 62666 218872 62672 218884
rect 50764 218844 62672 218872
rect 50764 218832 50770 218844
rect 62666 218832 62672 218844
rect 62724 218832 62730 218884
rect 83826 218832 83832 218884
rect 83884 218872 83890 218884
rect 153838 218872 153844 218884
rect 83884 218844 153844 218872
rect 83884 218832 83890 218844
rect 153838 218832 153844 218844
rect 153896 218832 153902 218884
rect 156230 218832 156236 218884
rect 156288 218872 156294 218884
rect 162118 218872 162124 218884
rect 156288 218844 162124 218872
rect 156288 218832 156294 218844
rect 162118 218832 162124 218844
rect 162176 218832 162182 218884
rect 165798 218832 165804 218884
rect 165856 218872 165862 218884
rect 165856 218844 166396 218872
rect 165856 218832 165862 218844
rect 59814 218696 59820 218748
rect 59872 218736 59878 218748
rect 142430 218736 142436 218748
rect 59872 218708 142436 218736
rect 59872 218696 59878 218708
rect 142430 218696 142436 218708
rect 142488 218696 142494 218748
rect 142614 218696 142620 218748
rect 142672 218736 142678 218748
rect 143258 218736 143264 218748
rect 142672 218708 143264 218736
rect 142672 218696 142678 218708
rect 143258 218696 143264 218708
rect 143316 218696 143322 218748
rect 145098 218696 145104 218748
rect 145156 218736 145162 218748
rect 145926 218736 145932 218748
rect 145156 218708 145932 218736
rect 145156 218696 145162 218708
rect 145926 218696 145932 218708
rect 145984 218696 145990 218748
rect 148410 218696 148416 218748
rect 148468 218736 148474 218748
rect 148962 218736 148968 218748
rect 148468 218708 148968 218736
rect 148468 218696 148474 218708
rect 148962 218696 148968 218708
rect 149020 218696 149026 218748
rect 149238 218696 149244 218748
rect 149296 218736 149302 218748
rect 150066 218736 150072 218748
rect 149296 218708 150072 218736
rect 149296 218696 149302 218708
rect 150066 218696 150072 218708
rect 150124 218696 150130 218748
rect 150434 218696 150440 218748
rect 150492 218736 150498 218748
rect 166368 218736 166396 218844
rect 166534 218832 166540 218884
rect 166592 218872 166598 218884
rect 171134 218872 171140 218884
rect 166592 218844 171140 218872
rect 166592 218832 166598 218844
rect 171134 218832 171140 218844
rect 171192 218832 171198 218884
rect 180058 218872 180064 218884
rect 171796 218844 180064 218872
rect 171796 218736 171824 218844
rect 180058 218832 180064 218844
rect 180116 218832 180122 218884
rect 180766 218844 184612 218872
rect 150492 218708 166304 218736
rect 166368 218708 171824 218736
rect 150492 218696 150498 218708
rect 100386 218560 100392 218612
rect 100444 218600 100450 218612
rect 105814 218600 105820 218612
rect 100444 218572 105820 218600
rect 100444 218560 100450 218572
rect 105814 218560 105820 218572
rect 105872 218560 105878 218612
rect 107010 218560 107016 218612
rect 107068 218600 107074 218612
rect 152366 218600 152372 218612
rect 107068 218572 152372 218600
rect 107068 218560 107074 218572
rect 152366 218560 152372 218572
rect 152424 218560 152430 218612
rect 152550 218560 152556 218612
rect 152608 218600 152614 218612
rect 153102 218600 153108 218612
rect 152608 218572 153108 218600
rect 152608 218560 152614 218572
rect 153102 218560 153108 218572
rect 153160 218560 153166 218612
rect 156690 218560 156696 218612
rect 156748 218600 156754 218612
rect 157242 218600 157248 218612
rect 156748 218572 157248 218600
rect 156748 218560 156754 218572
rect 157242 218560 157248 218572
rect 157300 218560 157306 218612
rect 157518 218560 157524 218612
rect 157576 218600 157582 218612
rect 158254 218600 158260 218612
rect 157576 218572 158260 218600
rect 157576 218560 157582 218572
rect 158254 218560 158260 218572
rect 158312 218560 158318 218612
rect 159174 218560 159180 218612
rect 159232 218600 159238 218612
rect 160002 218600 160008 218612
rect 159232 218572 160008 218600
rect 159232 218560 159238 218572
rect 160002 218560 160008 218572
rect 160060 218560 160066 218612
rect 161474 218560 161480 218612
rect 161532 218600 161538 218612
rect 166074 218600 166080 218612
rect 161532 218572 166080 218600
rect 161532 218560 161538 218572
rect 166074 218560 166080 218572
rect 166132 218560 166138 218612
rect 120258 218424 120264 218476
rect 120316 218464 120322 218476
rect 166074 218464 166080 218476
rect 120316 218436 166080 218464
rect 120316 218424 120322 218436
rect 166074 218424 166080 218436
rect 166132 218424 166138 218476
rect 166276 218464 166304 218708
rect 175734 218696 175740 218748
rect 175792 218736 175798 218748
rect 180766 218736 180794 218844
rect 175792 218708 180794 218736
rect 175792 218696 175798 218708
rect 181162 218696 181168 218748
rect 181220 218736 181226 218748
rect 184382 218736 184388 218748
rect 181220 218708 184388 218736
rect 181220 218696 181226 218708
rect 184382 218696 184388 218708
rect 184440 218696 184446 218748
rect 184584 218736 184612 218844
rect 186498 218832 186504 218884
rect 186556 218872 186562 218884
rect 239306 218872 239312 218884
rect 186556 218844 239312 218872
rect 186556 218832 186562 218844
rect 239306 218832 239312 218844
rect 239364 218832 239370 218884
rect 246114 218832 246120 218884
rect 246172 218872 246178 218884
rect 279050 218872 279056 218884
rect 246172 218844 279056 218872
rect 246172 218832 246178 218844
rect 279050 218832 279056 218844
rect 279108 218832 279114 218884
rect 279234 218832 279240 218884
rect 279292 218872 279298 218884
rect 279292 218844 282316 218872
rect 279292 218832 279298 218844
rect 189902 218736 189908 218748
rect 184584 218708 189908 218736
rect 189902 218696 189908 218708
rect 189960 218696 189966 218748
rect 191926 218696 191932 218748
rect 191984 218736 191990 218748
rect 195238 218736 195244 218748
rect 191984 218708 195244 218736
rect 191984 218696 191990 218708
rect 195238 218696 195244 218708
rect 195296 218696 195302 218748
rect 195606 218696 195612 218748
rect 195664 218736 195670 218748
rect 197998 218736 198004 218748
rect 195664 218708 198004 218736
rect 195664 218696 195670 218708
rect 197998 218696 198004 218708
rect 198056 218696 198062 218748
rect 198182 218696 198188 218748
rect 198240 218736 198246 218748
rect 246298 218736 246304 218748
rect 198240 218708 246304 218736
rect 198240 218696 198246 218708
rect 246298 218696 246304 218708
rect 246356 218696 246362 218748
rect 252738 218696 252744 218748
rect 252796 218736 252802 218748
rect 252796 218708 282224 218736
rect 252796 218696 252802 218708
rect 166626 218560 166632 218612
rect 166684 218600 166690 218612
rect 202598 218600 202604 218612
rect 166684 218572 202604 218600
rect 166684 218560 166690 218572
rect 202598 218560 202604 218572
rect 202656 218560 202662 218612
rect 203058 218560 203064 218612
rect 203116 218600 203122 218612
rect 206186 218600 206192 218612
rect 203116 218572 206192 218600
rect 203116 218560 203122 218572
rect 206186 218560 206192 218572
rect 206244 218560 206250 218612
rect 208026 218560 208032 218612
rect 208084 218600 208090 218612
rect 208084 218572 209774 218600
rect 208084 218560 208090 218572
rect 170950 218464 170956 218476
rect 166276 218436 170956 218464
rect 170950 218424 170956 218436
rect 171008 218424 171014 218476
rect 171134 218424 171140 218476
rect 171192 218464 171198 218476
rect 181346 218464 181352 218476
rect 171192 218436 181352 218464
rect 171192 218424 171198 218436
rect 181346 218424 181352 218436
rect 181404 218424 181410 218476
rect 189810 218424 189816 218476
rect 189868 218464 189874 218476
rect 191926 218464 191932 218476
rect 189868 218436 191932 218464
rect 189868 218424 189874 218436
rect 191926 218424 191932 218436
rect 191984 218424 191990 218476
rect 193766 218464 193772 218476
rect 192128 218436 193772 218464
rect 117958 218288 117964 218340
rect 118016 218328 118022 218340
rect 123478 218328 123484 218340
rect 118016 218300 123484 218328
rect 118016 218288 118022 218300
rect 123478 218288 123484 218300
rect 123536 218288 123542 218340
rect 131850 218288 131856 218340
rect 131908 218328 131914 218340
rect 132402 218328 132408 218340
rect 131908 218300 132408 218328
rect 131908 218288 131914 218300
rect 132402 218288 132408 218300
rect 132460 218288 132466 218340
rect 136818 218288 136824 218340
rect 136876 218328 136882 218340
rect 139486 218328 139492 218340
rect 136876 218300 139492 218328
rect 136876 218288 136882 218300
rect 139486 218288 139492 218300
rect 139544 218288 139550 218340
rect 140130 218288 140136 218340
rect 140188 218328 140194 218340
rect 181162 218328 181168 218340
rect 140188 218300 181168 218328
rect 140188 218288 140194 218300
rect 181162 218288 181168 218300
rect 181220 218288 181226 218340
rect 181530 218288 181536 218340
rect 181588 218328 181594 218340
rect 181990 218328 181996 218340
rect 181588 218300 181996 218328
rect 181588 218288 181594 218300
rect 181990 218288 181996 218300
rect 182048 218288 182054 218340
rect 184014 218288 184020 218340
rect 184072 218328 184078 218340
rect 184934 218328 184940 218340
rect 184072 218300 184940 218328
rect 184072 218288 184078 218300
rect 184934 218288 184940 218300
rect 184992 218288 184998 218340
rect 185670 218288 185676 218340
rect 185728 218328 185734 218340
rect 186130 218328 186136 218340
rect 185728 218300 186136 218328
rect 185728 218288 185734 218300
rect 186130 218288 186136 218300
rect 186188 218288 186194 218340
rect 188154 218288 188160 218340
rect 188212 218328 188218 218340
rect 188890 218328 188896 218340
rect 188212 218300 188896 218328
rect 188212 218288 188218 218300
rect 188890 218288 188896 218300
rect 188948 218288 188954 218340
rect 189074 218288 189080 218340
rect 189132 218328 189138 218340
rect 192128 218328 192156 218436
rect 193766 218424 193772 218436
rect 193824 218424 193830 218476
rect 198090 218424 198096 218476
rect 198148 218464 198154 218476
rect 200390 218464 200396 218476
rect 198148 218436 200396 218464
rect 198148 218424 198154 218436
rect 200390 218424 200396 218436
rect 200448 218424 200454 218476
rect 202230 218424 202236 218476
rect 202288 218464 202294 218476
rect 202782 218464 202788 218476
rect 202288 218436 202788 218464
rect 202288 218424 202294 218436
rect 202782 218424 202788 218436
rect 202840 218424 202846 218476
rect 204714 218424 204720 218476
rect 204772 218464 204778 218476
rect 207842 218464 207848 218476
rect 204772 218436 207848 218464
rect 204772 218424 204778 218436
rect 207842 218424 207848 218436
rect 207900 218424 207906 218476
rect 208854 218424 208860 218476
rect 208912 218464 208918 218476
rect 209498 218464 209504 218476
rect 208912 218436 209504 218464
rect 208912 218424 208918 218436
rect 209498 218424 209504 218436
rect 209556 218424 209562 218476
rect 209746 218464 209774 218572
rect 210142 218560 210148 218612
rect 210200 218600 210206 218612
rect 217318 218600 217324 218612
rect 210200 218572 217324 218600
rect 210200 218560 210206 218572
rect 217318 218560 217324 218572
rect 217376 218560 217382 218612
rect 219618 218560 219624 218612
rect 219676 218600 219682 218612
rect 264606 218600 264612 218612
rect 219676 218572 264612 218600
rect 219676 218560 219682 218572
rect 264606 218560 264612 218572
rect 264664 218560 264670 218612
rect 265986 218560 265992 218612
rect 266044 218600 266050 218612
rect 272334 218600 272340 218612
rect 266044 218572 272340 218600
rect 266044 218560 266050 218572
rect 272334 218560 272340 218572
rect 272392 218560 272398 218612
rect 272702 218560 272708 218612
rect 272760 218600 272766 218612
rect 279418 218600 279424 218612
rect 272760 218572 279424 218600
rect 272760 218560 272766 218572
rect 279418 218560 279424 218572
rect 279476 218560 279482 218612
rect 211522 218464 211528 218476
rect 209746 218436 211528 218464
rect 211522 218424 211528 218436
rect 211580 218424 211586 218476
rect 217962 218424 217968 218476
rect 218020 218464 218026 218476
rect 223482 218464 223488 218476
rect 218020 218436 223488 218464
rect 218020 218424 218026 218436
rect 223482 218424 223488 218436
rect 223540 218424 223546 218476
rect 225966 218424 225972 218476
rect 226024 218464 226030 218476
rect 266998 218464 267004 218476
rect 226024 218436 267004 218464
rect 226024 218424 226030 218436
rect 266998 218424 267004 218436
rect 267056 218424 267062 218476
rect 282196 218464 282224 218708
rect 282288 218600 282316 218844
rect 285858 218832 285864 218884
rect 285916 218872 285922 218884
rect 292022 218872 292028 218884
rect 285916 218844 292028 218872
rect 285916 218832 285922 218844
rect 292022 218832 292028 218844
rect 292080 218832 292086 218884
rect 314010 218832 314016 218884
rect 314068 218872 314074 218884
rect 340046 218872 340052 218884
rect 314068 218844 340052 218872
rect 314068 218832 314074 218844
rect 340046 218832 340052 218844
rect 340104 218832 340110 218884
rect 347038 218832 347044 218884
rect 347096 218872 347102 218884
rect 363506 218872 363512 218884
rect 347096 218844 363512 218872
rect 347096 218832 347102 218844
rect 363506 218832 363512 218844
rect 363564 218832 363570 218884
rect 368658 218832 368664 218884
rect 368716 218872 368722 218884
rect 378778 218872 378784 218884
rect 368716 218844 378784 218872
rect 368716 218832 368722 218844
rect 378778 218832 378784 218844
rect 378836 218832 378842 218884
rect 382734 218832 382740 218884
rect 382792 218872 382798 218884
rect 383562 218872 383568 218884
rect 382792 218844 383568 218872
rect 382792 218832 382798 218844
rect 383562 218832 383568 218844
rect 383620 218832 383626 218884
rect 386874 218832 386880 218884
rect 386932 218872 386938 218884
rect 398098 218872 398104 218884
rect 386932 218844 398104 218872
rect 386932 218832 386938 218844
rect 398098 218832 398104 218844
rect 398156 218832 398162 218884
rect 402606 218832 402612 218884
rect 402664 218872 402670 218884
rect 409046 218872 409052 218884
rect 402664 218844 409052 218872
rect 402664 218832 402670 218844
rect 409046 218832 409052 218844
rect 409104 218832 409110 218884
rect 411714 218832 411720 218884
rect 411772 218872 411778 218884
rect 412542 218872 412548 218884
rect 411772 218844 412548 218872
rect 411772 218832 411778 218844
rect 412542 218832 412548 218844
rect 412600 218832 412606 218884
rect 291654 218696 291660 218748
rect 291712 218736 291718 218748
rect 324590 218736 324596 218748
rect 291712 218708 324596 218736
rect 291712 218696 291718 218708
rect 324590 218696 324596 218708
rect 324648 218696 324654 218748
rect 327258 218696 327264 218748
rect 327316 218736 327322 218748
rect 351086 218736 351092 218748
rect 327316 218708 351092 218736
rect 327316 218696 327322 218708
rect 351086 218696 351092 218708
rect 351144 218696 351150 218748
rect 353754 218696 353760 218748
rect 353812 218736 353818 218748
rect 371786 218736 371792 218748
rect 353812 218708 371792 218736
rect 353812 218696 353818 218708
rect 371786 218696 371792 218708
rect 371844 218696 371850 218748
rect 383562 218696 383568 218748
rect 383620 218736 383626 218748
rect 396258 218736 396264 218748
rect 383620 218708 396264 218736
rect 383620 218696 383626 218708
rect 396258 218696 396264 218708
rect 396316 218696 396322 218748
rect 412542 218696 412548 218748
rect 412600 218736 412606 218748
rect 417142 218736 417148 218748
rect 412600 218708 417148 218736
rect 412600 218696 412606 218708
rect 417142 218696 417148 218708
rect 417200 218696 417206 218748
rect 429930 218696 429936 218748
rect 429988 218736 429994 218748
rect 432690 218736 432696 218748
rect 429988 218708 432696 218736
rect 429988 218696 429994 218708
rect 432690 218696 432696 218708
rect 432748 218696 432754 218748
rect 471330 218696 471336 218748
rect 471388 218736 471394 218748
rect 472894 218736 472900 218748
rect 471388 218708 472900 218736
rect 471388 218696 471394 218708
rect 472894 218696 472900 218708
rect 472952 218696 472958 218748
rect 482738 218696 482744 218748
rect 482796 218736 482802 218748
rect 485314 218736 485320 218748
rect 482796 218708 485320 218736
rect 482796 218696 482802 218708
rect 485314 218696 485320 218708
rect 485372 218696 485378 218748
rect 542814 218696 542820 218748
rect 542872 218736 542878 218748
rect 542872 218708 543228 218736
rect 542872 218696 542878 218708
rect 304258 218600 304264 218612
rect 282288 218572 304264 218600
rect 304258 218560 304264 218572
rect 304316 218560 304322 218612
rect 398466 218560 398472 218612
rect 398524 218600 398530 218612
rect 407758 218600 407764 218612
rect 398524 218572 407764 218600
rect 398524 218560 398530 218572
rect 407758 218560 407764 218572
rect 407816 218560 407822 218612
rect 469858 218560 469864 218612
rect 469916 218600 469922 218612
rect 471238 218600 471244 218612
rect 469916 218572 471244 218600
rect 469916 218560 469922 218572
rect 471238 218560 471244 218572
rect 471296 218560 471302 218612
rect 475562 218560 475568 218612
rect 475620 218600 475626 218612
rect 482830 218600 482836 218612
rect 475620 218572 482836 218600
rect 475620 218560 475626 218572
rect 482830 218560 482836 218572
rect 482888 218560 482894 218612
rect 537478 218560 537484 218612
rect 537536 218600 537542 218612
rect 542998 218600 543004 218612
rect 537536 218572 543004 218600
rect 537536 218560 537542 218572
rect 542998 218560 543004 218572
rect 543056 218560 543062 218612
rect 543200 218600 543228 218708
rect 543706 218600 543734 218980
rect 572070 218968 572076 218980
rect 572128 218968 572134 219020
rect 575474 219008 575480 219020
rect 572686 218980 575480 219008
rect 544930 218832 544936 218884
rect 544988 218872 544994 218884
rect 555970 218872 555976 218884
rect 544988 218844 555976 218872
rect 544988 218832 544994 218844
rect 555970 218832 555976 218844
rect 556028 218832 556034 218884
rect 567654 218872 567660 218884
rect 556172 218844 567660 218872
rect 547414 218696 547420 218748
rect 547472 218736 547478 218748
rect 556172 218736 556200 218844
rect 567654 218832 567660 218844
rect 567712 218832 567718 218884
rect 568206 218832 568212 218884
rect 568264 218872 568270 218884
rect 572686 218872 572714 218980
rect 575474 218968 575480 218980
rect 575532 218968 575538 219020
rect 568264 218844 572714 218872
rect 576826 218872 576854 219116
rect 626350 218872 626356 218884
rect 576826 218844 626356 218872
rect 568264 218832 568270 218844
rect 626350 218832 626356 218844
rect 626408 218832 626414 218884
rect 547472 218708 556200 218736
rect 547472 218696 547478 218708
rect 556430 218696 556436 218748
rect 556488 218736 556494 218748
rect 567838 218736 567844 218748
rect 556488 218708 567844 218736
rect 556488 218696 556494 218708
rect 567838 218696 567844 218708
rect 567896 218696 567902 218748
rect 568022 218696 568028 218748
rect 568080 218736 568086 218748
rect 570966 218736 570972 218748
rect 568080 218708 570972 218736
rect 568080 218696 568086 218708
rect 570966 218696 570972 218708
rect 571024 218696 571030 218748
rect 572530 218696 572536 218748
rect 572588 218736 572594 218748
rect 601878 218736 601884 218748
rect 572588 218708 601884 218736
rect 572588 218696 572594 218708
rect 601878 218696 601884 218708
rect 601936 218696 601942 218748
rect 644934 218696 644940 218748
rect 644992 218736 644998 218748
rect 656158 218736 656164 218748
rect 644992 218708 656164 218736
rect 644992 218696 644998 218708
rect 656158 218696 656164 218708
rect 656216 218696 656222 218748
rect 543200 218572 543734 218600
rect 555970 218560 555976 218612
rect 556028 218600 556034 218612
rect 598842 218600 598848 218612
rect 556028 218572 598848 218600
rect 556028 218560 556034 218572
rect 598842 218560 598848 218572
rect 598900 218560 598906 218612
rect 288986 218464 288992 218476
rect 282196 218436 288992 218464
rect 288986 218424 288992 218436
rect 289044 218424 289050 218476
rect 294138 218424 294144 218476
rect 294196 218464 294202 218476
rect 316678 218464 316684 218476
rect 294196 218436 316684 218464
rect 294196 218424 294202 218436
rect 316678 218424 316684 218436
rect 316736 218424 316742 218476
rect 500034 218424 500040 218476
rect 500092 218464 500098 218476
rect 609882 218464 609888 218476
rect 500092 218436 609888 218464
rect 500092 218424 500098 218436
rect 609882 218424 609888 218436
rect 609940 218424 609946 218476
rect 458174 218356 458180 218408
rect 458232 218396 458238 218408
rect 458232 218368 460934 218396
rect 458232 218356 458238 218368
rect 189132 218300 192156 218328
rect 189132 218288 189138 218300
rect 192294 218288 192300 218340
rect 192352 218328 192358 218340
rect 193030 218328 193036 218340
rect 192352 218300 193036 218328
rect 192352 218288 192358 218300
rect 193030 218288 193036 218300
rect 193088 218288 193094 218340
rect 193950 218288 193956 218340
rect 194008 218328 194014 218340
rect 194502 218328 194508 218340
rect 194008 218300 194508 218328
rect 194008 218288 194014 218300
rect 194502 218288 194508 218300
rect 194560 218288 194566 218340
rect 194778 218288 194784 218340
rect 194836 218328 194842 218340
rect 195882 218328 195888 218340
rect 194836 218300 195888 218328
rect 194836 218288 194842 218300
rect 195882 218288 195888 218300
rect 195940 218288 195946 218340
rect 196434 218288 196440 218340
rect 196492 218328 196498 218340
rect 210142 218328 210148 218340
rect 196492 218300 210148 218328
rect 196492 218288 196498 218300
rect 210142 218288 210148 218300
rect 210200 218288 210206 218340
rect 210326 218288 210332 218340
rect 210384 218328 210390 218340
rect 213178 218328 213184 218340
rect 210384 218300 213184 218328
rect 210384 218288 210390 218300
rect 213178 218288 213184 218300
rect 213236 218288 213242 218340
rect 222930 218288 222936 218340
rect 222988 218328 222994 218340
rect 231026 218328 231032 218340
rect 222988 218300 231032 218328
rect 222988 218288 222994 218300
rect 231026 218288 231032 218300
rect 231084 218288 231090 218340
rect 232866 218288 232872 218340
rect 232924 218328 232930 218340
rect 270770 218328 270776 218340
rect 232924 218300 270776 218328
rect 232924 218288 232930 218300
rect 270770 218288 270776 218300
rect 270828 218288 270834 218340
rect 426618 218288 426624 218340
rect 426676 218328 426682 218340
rect 429562 218328 429568 218340
rect 426676 218300 429568 218328
rect 426676 218288 426682 218300
rect 429562 218288 429568 218300
rect 429620 218288 429626 218340
rect 450722 218288 450728 218340
rect 450780 218328 450786 218340
rect 453850 218328 453856 218340
rect 450780 218300 453856 218328
rect 450780 218288 450786 218300
rect 453850 218288 453856 218300
rect 453908 218288 453914 218340
rect 460906 218328 460934 218368
rect 461302 218328 461308 218340
rect 460906 218300 461308 218328
rect 461302 218288 461308 218300
rect 461360 218288 461366 218340
rect 503162 218288 503168 218340
rect 503220 218328 503226 218340
rect 503220 218300 558224 218328
rect 503220 218288 503226 218300
rect 55674 218152 55680 218204
rect 55732 218192 55738 218204
rect 56502 218192 56508 218204
rect 55732 218164 56508 218192
rect 55732 218152 55738 218164
rect 56502 218152 56508 218164
rect 56560 218152 56566 218204
rect 57422 218152 57428 218204
rect 57480 218192 57486 218204
rect 61654 218192 61660 218204
rect 57480 218164 61660 218192
rect 57480 218152 57486 218164
rect 61654 218152 61660 218164
rect 61712 218152 61718 218204
rect 67266 218152 67272 218204
rect 67324 218192 67330 218204
rect 68278 218192 68284 218204
rect 67324 218164 68284 218192
rect 67324 218152 67330 218164
rect 68278 218152 68284 218164
rect 68336 218152 68342 218204
rect 75546 218152 75552 218204
rect 75604 218192 75610 218204
rect 76558 218192 76564 218204
rect 75604 218164 76564 218192
rect 75604 218152 75610 218164
rect 76558 218152 76564 218164
rect 76616 218152 76622 218204
rect 123570 218152 123576 218204
rect 123628 218192 123634 218204
rect 161474 218192 161480 218204
rect 123628 218164 161480 218192
rect 123628 218152 123634 218164
rect 161474 218152 161480 218164
rect 161532 218152 161538 218204
rect 161658 218152 161664 218204
rect 161716 218192 161722 218204
rect 162762 218192 162768 218204
rect 161716 218164 162768 218192
rect 161716 218152 161722 218164
rect 162762 218152 162768 218164
rect 162820 218152 162826 218204
rect 163314 218152 163320 218204
rect 163372 218192 163378 218204
rect 163958 218192 163964 218204
rect 163372 218164 163964 218192
rect 163372 218152 163378 218164
rect 163958 218152 163964 218164
rect 164016 218152 164022 218204
rect 164970 218152 164976 218204
rect 165028 218192 165034 218204
rect 165522 218192 165528 218204
rect 165028 218164 165528 218192
rect 165028 218152 165034 218164
rect 165522 218152 165528 218164
rect 165580 218152 165586 218204
rect 171410 218192 171416 218204
rect 166966 218164 171416 218192
rect 56502 218016 56508 218068
rect 56560 218056 56566 218068
rect 57238 218056 57244 218068
rect 56560 218028 57244 218056
rect 56560 218016 56566 218028
rect 57238 218016 57244 218028
rect 57296 218016 57302 218068
rect 58158 218016 58164 218068
rect 58216 218056 58222 218068
rect 59354 218056 59360 218068
rect 58216 218028 59360 218056
rect 58216 218016 58222 218028
rect 59354 218016 59360 218028
rect 59412 218016 59418 218068
rect 61470 218016 61476 218068
rect 61528 218056 61534 218068
rect 62022 218056 62028 218068
rect 61528 218028 62028 218056
rect 61528 218016 61534 218028
rect 62022 218016 62028 218028
rect 62080 218016 62086 218068
rect 65610 218016 65616 218068
rect 65668 218056 65674 218068
rect 66162 218056 66168 218068
rect 65668 218028 66168 218056
rect 65668 218016 65674 218028
rect 66162 218016 66168 218028
rect 66220 218016 66226 218068
rect 66438 218016 66444 218068
rect 66496 218056 66502 218068
rect 67542 218056 67548 218068
rect 66496 218028 67548 218056
rect 66496 218016 66502 218028
rect 67542 218016 67548 218028
rect 67600 218016 67606 218068
rect 68094 218016 68100 218068
rect 68152 218056 68158 218068
rect 68738 218056 68744 218068
rect 68152 218028 68744 218056
rect 68152 218016 68158 218028
rect 68738 218016 68744 218028
rect 68796 218016 68802 218068
rect 72234 218016 72240 218068
rect 72292 218056 72298 218068
rect 73706 218056 73712 218068
rect 72292 218028 73712 218056
rect 72292 218016 72298 218028
rect 73706 218016 73712 218028
rect 73764 218016 73770 218068
rect 74718 218016 74724 218068
rect 74776 218056 74782 218068
rect 75822 218056 75828 218068
rect 74776 218028 75828 218056
rect 74776 218016 74782 218028
rect 75822 218016 75828 218028
rect 75880 218016 75886 218068
rect 78030 218016 78036 218068
rect 78088 218056 78094 218068
rect 78582 218056 78588 218068
rect 78088 218028 78588 218056
rect 78088 218016 78094 218028
rect 78582 218016 78588 218028
rect 78640 218016 78646 218068
rect 78858 218016 78864 218068
rect 78916 218056 78922 218068
rect 79962 218056 79968 218068
rect 78916 218028 79968 218056
rect 78916 218016 78922 218028
rect 79962 218016 79968 218028
rect 80020 218016 80026 218068
rect 82170 218016 82176 218068
rect 82228 218056 82234 218068
rect 83458 218056 83464 218068
rect 82228 218028 83464 218056
rect 82228 218016 82234 218028
rect 83458 218016 83464 218028
rect 83516 218016 83522 218068
rect 84654 218016 84660 218068
rect 84712 218056 84718 218068
rect 85298 218056 85304 218068
rect 84712 218028 85304 218056
rect 84712 218016 84718 218028
rect 85298 218016 85304 218028
rect 85356 218016 85362 218068
rect 87138 218016 87144 218068
rect 87196 218056 87202 218068
rect 88242 218056 88248 218068
rect 87196 218028 88248 218056
rect 87196 218016 87202 218028
rect 88242 218016 88248 218028
rect 88300 218016 88306 218068
rect 88794 218016 88800 218068
rect 88852 218056 88858 218068
rect 89438 218056 89444 218068
rect 88852 218028 89444 218056
rect 88852 218016 88858 218028
rect 89438 218016 89444 218028
rect 89496 218016 89502 218068
rect 90450 218016 90456 218068
rect 90508 218056 90514 218068
rect 91738 218056 91744 218068
rect 90508 218028 91744 218056
rect 90508 218016 90514 218028
rect 91738 218016 91744 218028
rect 91796 218016 91802 218068
rect 92934 218016 92940 218068
rect 92992 218056 92998 218068
rect 93762 218056 93768 218068
rect 92992 218028 93768 218056
rect 92992 218016 92998 218028
rect 93762 218016 93768 218028
rect 93820 218016 93826 218068
rect 95418 218016 95424 218068
rect 95476 218056 95482 218068
rect 96246 218056 96252 218068
rect 95476 218028 96252 218056
rect 95476 218016 95482 218028
rect 96246 218016 96252 218028
rect 96304 218016 96310 218068
rect 97074 218016 97080 218068
rect 97132 218056 97138 218068
rect 97994 218056 98000 218068
rect 97132 218028 98000 218056
rect 97132 218016 97138 218028
rect 97994 218016 98000 218028
rect 98052 218016 98058 218068
rect 98730 218016 98736 218068
rect 98788 218056 98794 218068
rect 99282 218056 99288 218068
rect 98788 218028 99288 218056
rect 98788 218016 98794 218028
rect 99282 218016 99288 218028
rect 99340 218016 99346 218068
rect 99558 218016 99564 218068
rect 99616 218056 99622 218068
rect 100662 218056 100668 218068
rect 99616 218028 100668 218056
rect 99616 218016 99622 218028
rect 100662 218016 100668 218028
rect 100720 218016 100726 218068
rect 102870 218016 102876 218068
rect 102928 218056 102934 218068
rect 103422 218056 103428 218068
rect 102928 218028 103428 218056
rect 102928 218016 102934 218028
rect 103422 218016 103428 218028
rect 103480 218016 103486 218068
rect 105354 218016 105360 218068
rect 105412 218056 105418 218068
rect 105998 218056 106004 218068
rect 105412 218028 106004 218056
rect 105412 218016 105418 218028
rect 105998 218016 106004 218028
rect 106056 218016 106062 218068
rect 109494 218016 109500 218068
rect 109552 218056 109558 218068
rect 110138 218056 110144 218068
rect 109552 218028 110144 218056
rect 109552 218016 109558 218028
rect 110138 218016 110144 218028
rect 110196 218016 110202 218068
rect 116118 218016 116124 218068
rect 116176 218056 116182 218068
rect 117222 218056 117228 218068
rect 116176 218028 117228 218056
rect 116176 218016 116182 218028
rect 117222 218016 117228 218028
rect 117280 218016 117286 218068
rect 117774 218016 117780 218068
rect 117832 218056 117838 218068
rect 118694 218056 118700 218068
rect 117832 218028 118700 218056
rect 117832 218016 117838 218028
rect 118694 218016 118700 218028
rect 118752 218016 118758 218068
rect 119430 218016 119436 218068
rect 119488 218056 119494 218068
rect 119982 218056 119988 218068
rect 119488 218028 119988 218056
rect 119488 218016 119494 218028
rect 119982 218016 119988 218028
rect 120040 218016 120046 218068
rect 121914 218016 121920 218068
rect 121972 218056 121978 218068
rect 122558 218056 122564 218068
rect 121972 218028 122564 218056
rect 121972 218016 121978 218028
rect 122558 218016 122564 218028
rect 122616 218016 122622 218068
rect 126054 218016 126060 218068
rect 126112 218056 126118 218068
rect 126698 218056 126704 218068
rect 126112 218028 126704 218056
rect 126112 218016 126118 218028
rect 126698 218016 126704 218028
rect 126756 218016 126762 218068
rect 127710 218016 127716 218068
rect 127768 218056 127774 218068
rect 128262 218056 128268 218068
rect 127768 218028 128268 218056
rect 127768 218016 127774 218028
rect 128262 218016 128268 218028
rect 128320 218016 128326 218068
rect 128538 218016 128544 218068
rect 128596 218056 128602 218068
rect 129366 218056 129372 218068
rect 128596 218028 129372 218056
rect 128596 218016 128602 218028
rect 129366 218016 129372 218028
rect 129424 218016 129430 218068
rect 130194 218016 130200 218068
rect 130252 218056 130258 218068
rect 132494 218056 132500 218068
rect 130252 218028 132500 218056
rect 130252 218016 130258 218028
rect 132494 218016 132500 218028
rect 132552 218016 132558 218068
rect 132678 218016 132684 218068
rect 132736 218056 132742 218068
rect 133506 218056 133512 218068
rect 132736 218028 133512 218056
rect 132736 218016 132742 218028
rect 133506 218016 133512 218028
rect 133564 218016 133570 218068
rect 135990 218016 135996 218068
rect 136048 218056 136054 218068
rect 136542 218056 136548 218068
rect 136048 218028 136548 218056
rect 136048 218016 136054 218028
rect 136542 218016 136548 218028
rect 136600 218016 136606 218068
rect 138474 218016 138480 218068
rect 138532 218056 138538 218068
rect 139118 218056 139124 218068
rect 138532 218028 139124 218056
rect 138532 218016 138538 218028
rect 139118 218016 139124 218028
rect 139176 218016 139182 218068
rect 139486 218016 139492 218068
rect 139544 218056 139550 218068
rect 166966 218056 166994 218164
rect 171410 218152 171416 218164
rect 171468 218152 171474 218204
rect 173250 218152 173256 218204
rect 173308 218192 173314 218204
rect 173308 218164 179552 218192
rect 173308 218152 173314 218164
rect 139544 218028 166994 218056
rect 139544 218016 139550 218028
rect 170766 218016 170772 218068
rect 170824 218056 170830 218068
rect 176470 218056 176476 218068
rect 170824 218028 176476 218056
rect 170824 218016 170830 218028
rect 176470 218016 176476 218028
rect 176528 218016 176534 218068
rect 178218 218016 178224 218068
rect 178276 218056 178282 218068
rect 179322 218056 179328 218068
rect 178276 218028 179328 218056
rect 178276 218016 178282 218028
rect 179322 218016 179328 218028
rect 179380 218016 179386 218068
rect 179524 218056 179552 218164
rect 179874 218152 179880 218204
rect 179932 218192 179938 218204
rect 225598 218192 225604 218204
rect 179932 218164 225604 218192
rect 179932 218152 179938 218164
rect 225598 218152 225604 218164
rect 225656 218152 225662 218204
rect 241974 218152 241980 218204
rect 242032 218192 242038 218204
rect 242894 218192 242900 218204
rect 242032 218164 242900 218192
rect 242032 218152 242038 218164
rect 242894 218152 242900 218164
rect 242952 218152 242958 218204
rect 243538 218152 243544 218204
rect 243596 218192 243602 218204
rect 249058 218192 249064 218204
rect 243596 218164 249064 218192
rect 243596 218152 243602 218164
rect 249058 218152 249064 218164
rect 249116 218152 249122 218204
rect 297450 218152 297456 218204
rect 297508 218192 297514 218204
rect 302878 218192 302884 218204
rect 297508 218164 302884 218192
rect 297508 218152 297514 218164
rect 302878 218152 302884 218164
rect 302936 218152 302942 218204
rect 333054 218152 333060 218204
rect 333112 218192 333118 218204
rect 333882 218192 333888 218204
rect 333112 218164 333888 218192
rect 333112 218152 333118 218164
rect 333882 218152 333888 218164
rect 333940 218152 333946 218204
rect 335538 218152 335544 218204
rect 335596 218192 335602 218204
rect 338666 218192 338672 218204
rect 335596 218164 338672 218192
rect 335596 218152 335602 218164
rect 338666 218152 338672 218164
rect 338724 218152 338730 218204
rect 358722 218152 358728 218204
rect 358780 218192 358786 218204
rect 359458 218192 359464 218204
rect 358780 218164 359464 218192
rect 358780 218152 358786 218164
rect 359458 218152 359464 218164
rect 359516 218152 359522 218204
rect 381906 218152 381912 218204
rect 381964 218192 381970 218204
rect 382918 218192 382924 218204
rect 381964 218164 382924 218192
rect 381964 218152 381970 218164
rect 382918 218152 382924 218164
rect 382976 218152 382982 218204
rect 400950 218152 400956 218204
rect 401008 218192 401014 218204
rect 402238 218192 402244 218204
rect 401008 218164 402244 218192
rect 401008 218152 401014 218164
rect 402238 218152 402244 218164
rect 402296 218152 402302 218204
rect 407574 218152 407580 218204
rect 407632 218192 407638 218204
rect 411898 218192 411904 218204
rect 407632 218164 411904 218192
rect 407632 218152 407638 218164
rect 411898 218152 411904 218164
rect 411956 218152 411962 218204
rect 422478 218152 422484 218204
rect 422536 218192 422542 218204
rect 425422 218192 425428 218204
rect 422536 218164 425428 218192
rect 422536 218152 422542 218164
rect 425422 218152 425428 218164
rect 425480 218152 425486 218204
rect 425790 218152 425796 218204
rect 425848 218192 425854 218204
rect 427906 218192 427912 218204
rect 425848 218164 427912 218192
rect 425848 218152 425854 218164
rect 427906 218152 427912 218164
rect 427964 218152 427970 218204
rect 428458 218152 428464 218204
rect 428516 218192 428522 218204
rect 430114 218192 430120 218204
rect 428516 218164 430120 218192
rect 428516 218152 428522 218164
rect 430114 218152 430120 218164
rect 430172 218152 430178 218204
rect 433242 218152 433248 218204
rect 433300 218192 433306 218204
rect 435266 218192 435272 218204
rect 433300 218164 435272 218192
rect 433300 218152 433306 218164
rect 435266 218152 435272 218164
rect 435324 218152 435330 218204
rect 435726 218152 435732 218204
rect 435784 218192 435790 218204
rect 436646 218192 436652 218204
rect 435784 218164 436652 218192
rect 435784 218152 435790 218164
rect 436646 218152 436652 218164
rect 436704 218152 436710 218204
rect 461946 218152 461952 218204
rect 462004 218192 462010 218204
rect 466270 218192 466276 218204
rect 462004 218164 466276 218192
rect 462004 218152 462010 218164
rect 466270 218152 466276 218164
rect 466328 218152 466334 218204
rect 507670 218152 507676 218204
rect 507728 218192 507734 218204
rect 542814 218192 542820 218204
rect 507728 218164 542820 218192
rect 507728 218152 507734 218164
rect 542814 218152 542820 218164
rect 542872 218152 542878 218204
rect 542998 218152 543004 218204
rect 543056 218192 543062 218204
rect 556430 218192 556436 218204
rect 543056 218164 556436 218192
rect 543056 218152 543062 218164
rect 556430 218152 556436 218164
rect 556488 218152 556494 218204
rect 558196 218192 558224 218300
rect 562226 218288 562232 218340
rect 562284 218328 562290 218340
rect 562870 218328 562876 218340
rect 562284 218300 562876 218328
rect 562284 218288 562290 218300
rect 562870 218288 562876 218300
rect 562928 218288 562934 218340
rect 614482 218328 614488 218340
rect 563026 218300 614488 218328
rect 563026 218192 563054 218300
rect 614482 218288 614488 218300
rect 614540 218288 614546 218340
rect 558196 218164 563054 218192
rect 572668 218152 572674 218204
rect 572726 218192 572732 218204
rect 615678 218192 615684 218204
rect 572726 218164 615684 218192
rect 572726 218152 572732 218164
rect 615678 218152 615684 218164
rect 615736 218152 615742 218204
rect 572438 218124 572444 218136
rect 563210 218096 572444 218124
rect 210326 218056 210332 218068
rect 179524 218028 210332 218056
rect 210326 218016 210332 218028
rect 210384 218016 210390 218068
rect 210510 218016 210516 218068
rect 210568 218056 210574 218068
rect 210970 218056 210976 218068
rect 210568 218028 210976 218056
rect 210568 218016 210574 218028
rect 210970 218016 210976 218028
rect 211028 218016 211034 218068
rect 214650 218016 214656 218068
rect 214708 218056 214714 218068
rect 215202 218056 215208 218068
rect 214708 218028 215208 218056
rect 214708 218016 214714 218028
rect 215202 218016 215208 218028
rect 215260 218016 215266 218068
rect 215478 218016 215484 218068
rect 215536 218056 215542 218068
rect 216122 218056 216128 218068
rect 215536 218028 216128 218056
rect 215536 218016 215542 218028
rect 216122 218016 216128 218028
rect 216180 218016 216186 218068
rect 218790 218016 218796 218068
rect 218848 218056 218854 218068
rect 219342 218056 219348 218068
rect 218848 218028 219348 218056
rect 218848 218016 218854 218028
rect 219342 218016 219348 218028
rect 219400 218016 219406 218068
rect 221274 218016 221280 218068
rect 221332 218056 221338 218068
rect 221826 218056 221832 218068
rect 221332 218028 221832 218056
rect 221332 218016 221338 218028
rect 221826 218016 221832 218028
rect 221884 218016 221890 218068
rect 225414 218016 225420 218068
rect 225472 218056 225478 218068
rect 226150 218056 226156 218068
rect 225472 218028 226156 218056
rect 225472 218016 225478 218028
rect 226150 218016 226156 218028
rect 226208 218016 226214 218068
rect 227070 218016 227076 218068
rect 227128 218056 227134 218068
rect 227530 218056 227536 218068
rect 227128 218028 227536 218056
rect 227128 218016 227134 218028
rect 227530 218016 227536 218028
rect 227588 218016 227594 218068
rect 229554 218016 229560 218068
rect 229612 218056 229618 218068
rect 230474 218056 230480 218068
rect 229612 218028 230480 218056
rect 229612 218016 229618 218028
rect 230474 218016 230480 218028
rect 230532 218016 230538 218068
rect 231210 218016 231216 218068
rect 231268 218056 231274 218068
rect 231670 218056 231676 218068
rect 231268 218028 231676 218056
rect 231268 218016 231274 218028
rect 231670 218016 231676 218028
rect 231728 218016 231734 218068
rect 232038 218016 232044 218068
rect 232096 218056 232102 218068
rect 233142 218056 233148 218068
rect 232096 218028 233148 218056
rect 232096 218016 232102 218028
rect 233142 218016 233148 218028
rect 233200 218016 233206 218068
rect 235350 218016 235356 218068
rect 235408 218056 235414 218068
rect 235810 218056 235816 218068
rect 235408 218028 235816 218056
rect 235408 218016 235414 218028
rect 235810 218016 235816 218028
rect 235868 218016 235874 218068
rect 240318 218016 240324 218068
rect 240376 218056 240382 218068
rect 241330 218056 241336 218068
rect 240376 218028 241336 218056
rect 240376 218016 240382 218028
rect 241330 218016 241336 218028
rect 241388 218016 241394 218068
rect 243630 218016 243636 218068
rect 243688 218056 243694 218068
rect 244090 218056 244096 218068
rect 243688 218028 244096 218056
rect 243688 218016 243694 218028
rect 244090 218016 244096 218028
rect 244148 218016 244154 218068
rect 244458 218016 244464 218068
rect 244516 218056 244522 218068
rect 245286 218056 245292 218068
rect 244516 218028 245292 218056
rect 244516 218016 244522 218028
rect 245286 218016 245292 218028
rect 245344 218016 245350 218068
rect 247770 218016 247776 218068
rect 247828 218056 247834 218068
rect 248322 218056 248328 218068
rect 247828 218028 248328 218056
rect 247828 218016 247834 218028
rect 248322 218016 248328 218028
rect 248380 218016 248386 218068
rect 248598 218016 248604 218068
rect 248656 218056 248662 218068
rect 249242 218056 249248 218068
rect 248656 218028 249248 218056
rect 248656 218016 248662 218028
rect 249242 218016 249248 218028
rect 249300 218016 249306 218068
rect 250254 218016 250260 218068
rect 250312 218056 250318 218068
rect 250898 218056 250904 218068
rect 250312 218028 250904 218056
rect 250312 218016 250318 218028
rect 250898 218016 250904 218028
rect 250956 218016 250962 218068
rect 251910 218016 251916 218068
rect 251968 218056 251974 218068
rect 252462 218056 252468 218068
rect 251968 218028 252468 218056
rect 251968 218016 251974 218028
rect 252462 218016 252468 218028
rect 252520 218016 252526 218068
rect 256050 218016 256056 218068
rect 256108 218056 256114 218068
rect 256510 218056 256516 218068
rect 256108 218028 256516 218056
rect 256108 218016 256114 218028
rect 256510 218016 256516 218028
rect 256568 218016 256574 218068
rect 256878 218016 256884 218068
rect 256936 218056 256942 218068
rect 257522 218056 257528 218068
rect 256936 218028 257528 218056
rect 256936 218016 256942 218028
rect 257522 218016 257528 218028
rect 257580 218016 257586 218068
rect 258534 218016 258540 218068
rect 258592 218056 258598 218068
rect 259362 218056 259368 218068
rect 258592 218028 259368 218056
rect 258592 218016 258598 218028
rect 259362 218016 259368 218028
rect 259420 218016 259426 218068
rect 260190 218016 260196 218068
rect 260248 218056 260254 218068
rect 260742 218056 260748 218068
rect 260248 218028 260748 218056
rect 260248 218016 260254 218028
rect 260742 218016 260748 218028
rect 260800 218016 260806 218068
rect 264330 218016 264336 218068
rect 264388 218056 264394 218068
rect 264790 218056 264796 218068
rect 264388 218028 264796 218056
rect 264388 218016 264394 218028
rect 264790 218016 264796 218028
rect 264848 218016 264854 218068
rect 265158 218016 265164 218068
rect 265216 218056 265222 218068
rect 266262 218056 266268 218068
rect 265216 218028 266268 218056
rect 265216 218016 265222 218028
rect 266262 218016 266268 218028
rect 266320 218016 266326 218068
rect 268470 218016 268476 218068
rect 268528 218056 268534 218068
rect 268930 218056 268936 218068
rect 268528 218028 268936 218056
rect 268528 218016 268534 218028
rect 268930 218016 268936 218028
rect 268988 218016 268994 218068
rect 269298 218016 269304 218068
rect 269356 218056 269362 218068
rect 270218 218056 270224 218068
rect 269356 218028 270224 218056
rect 269356 218016 269362 218028
rect 270218 218016 270224 218028
rect 270276 218016 270282 218068
rect 270954 218016 270960 218068
rect 271012 218056 271018 218068
rect 272518 218056 272524 218068
rect 271012 218028 272524 218056
rect 271012 218016 271018 218028
rect 272518 218016 272524 218028
rect 272576 218016 272582 218068
rect 277578 218016 277584 218068
rect 277636 218056 277642 218068
rect 278590 218056 278596 218068
rect 277636 218028 278596 218056
rect 277636 218016 277642 218028
rect 278590 218016 278596 218028
rect 278648 218016 278654 218068
rect 280890 218016 280896 218068
rect 280948 218056 280954 218068
rect 281442 218056 281448 218068
rect 280948 218028 281448 218056
rect 280948 218016 280954 218028
rect 281442 218016 281448 218028
rect 281500 218016 281506 218068
rect 281718 218016 281724 218068
rect 281776 218056 281782 218068
rect 282730 218056 282736 218068
rect 281776 218028 282736 218056
rect 281776 218016 281782 218028
rect 282730 218016 282736 218028
rect 282788 218016 282794 218068
rect 283374 218016 283380 218068
rect 283432 218056 283438 218068
rect 284294 218056 284300 218068
rect 283432 218028 284300 218056
rect 283432 218016 283438 218028
rect 284294 218016 284300 218028
rect 284352 218016 284358 218068
rect 285030 218016 285036 218068
rect 285088 218056 285094 218068
rect 285490 218056 285496 218068
rect 285088 218028 285496 218056
rect 285088 218016 285094 218028
rect 285490 218016 285496 218028
rect 285548 218016 285554 218068
rect 287514 218016 287520 218068
rect 287572 218056 287578 218068
rect 288066 218056 288072 218068
rect 287572 218028 288072 218056
rect 287572 218016 287578 218028
rect 288066 218016 288072 218028
rect 288124 218016 288130 218068
rect 289170 218016 289176 218068
rect 289228 218056 289234 218068
rect 289630 218056 289636 218068
rect 289228 218028 289636 218056
rect 289228 218016 289234 218028
rect 289630 218016 289636 218028
rect 289688 218016 289694 218068
rect 289998 218016 290004 218068
rect 290056 218056 290062 218068
rect 291102 218056 291108 218068
rect 290056 218028 291108 218056
rect 290056 218016 290062 218028
rect 291102 218016 291108 218028
rect 291160 218016 291166 218068
rect 293310 218016 293316 218068
rect 293368 218056 293374 218068
rect 293770 218056 293776 218068
rect 293368 218028 293776 218056
rect 293368 218016 293374 218028
rect 293770 218016 293776 218028
rect 293828 218016 293834 218068
rect 298278 218016 298284 218068
rect 298336 218056 298342 218068
rect 299382 218056 299388 218068
rect 298336 218028 299388 218056
rect 298336 218016 298342 218028
rect 299382 218016 299388 218028
rect 299440 218016 299446 218068
rect 299934 218016 299940 218068
rect 299992 218056 299998 218068
rect 300670 218056 300676 218068
rect 299992 218028 300676 218056
rect 299992 218016 299998 218028
rect 300670 218016 300676 218028
rect 300728 218016 300734 218068
rect 301590 218016 301596 218068
rect 301648 218056 301654 218068
rect 302142 218056 302148 218068
rect 301648 218028 302148 218056
rect 301648 218016 301654 218028
rect 302142 218016 302148 218028
rect 302200 218016 302206 218068
rect 305730 218016 305736 218068
rect 305788 218056 305794 218068
rect 306190 218056 306196 218068
rect 305788 218028 306196 218056
rect 305788 218016 305794 218028
rect 306190 218016 306196 218028
rect 306248 218016 306254 218068
rect 306558 218016 306564 218068
rect 306616 218056 306622 218068
rect 307662 218056 307668 218068
rect 306616 218028 307668 218056
rect 306616 218016 306622 218028
rect 307662 218016 307668 218028
rect 307720 218016 307726 218068
rect 308214 218016 308220 218068
rect 308272 218056 308278 218068
rect 308858 218056 308864 218068
rect 308272 218028 308864 218056
rect 308272 218016 308278 218028
rect 308858 218016 308864 218028
rect 308916 218016 308922 218068
rect 309870 218016 309876 218068
rect 309928 218056 309934 218068
rect 310330 218056 310336 218068
rect 309928 218028 310336 218056
rect 309928 218016 309934 218028
rect 310330 218016 310336 218028
rect 310388 218016 310394 218068
rect 312354 218016 312360 218068
rect 312412 218056 312418 218068
rect 312906 218056 312912 218068
rect 312412 218028 312912 218056
rect 312412 218016 312418 218028
rect 312906 218016 312912 218028
rect 312964 218016 312970 218068
rect 314838 218016 314844 218068
rect 314896 218056 314902 218068
rect 315482 218056 315488 218068
rect 314896 218028 315488 218056
rect 314896 218016 314902 218028
rect 315482 218016 315488 218028
rect 315540 218016 315546 218068
rect 317322 218016 317328 218068
rect 317380 218056 317386 218068
rect 317966 218056 317972 218068
rect 317380 218028 317972 218056
rect 317380 218016 317386 218028
rect 317966 218016 317972 218028
rect 318024 218016 318030 218068
rect 318978 218016 318984 218068
rect 319036 218056 319042 218068
rect 320082 218056 320088 218068
rect 319036 218028 320088 218056
rect 319036 218016 319042 218028
rect 320082 218016 320088 218028
rect 320140 218016 320146 218068
rect 322290 218016 322296 218068
rect 322348 218056 322354 218068
rect 322842 218056 322848 218068
rect 322348 218028 322848 218056
rect 322348 218016 322354 218028
rect 322842 218016 322848 218028
rect 322900 218016 322906 218068
rect 323118 218016 323124 218068
rect 323176 218056 323182 218068
rect 323946 218056 323952 218068
rect 323176 218028 323952 218056
rect 323176 218016 323182 218028
rect 323946 218016 323952 218028
rect 324004 218016 324010 218068
rect 324774 218016 324780 218068
rect 324832 218056 324838 218068
rect 325510 218056 325516 218068
rect 324832 218028 325516 218056
rect 324832 218016 324838 218028
rect 325510 218016 325516 218028
rect 325568 218016 325574 218068
rect 326430 218016 326436 218068
rect 326488 218056 326494 218068
rect 326890 218056 326896 218068
rect 326488 218028 326896 218056
rect 326488 218016 326494 218028
rect 326890 218016 326896 218028
rect 326948 218016 326954 218068
rect 330570 218016 330576 218068
rect 330628 218056 330634 218068
rect 331030 218056 331036 218068
rect 330628 218028 331036 218056
rect 330628 218016 330634 218028
rect 331030 218016 331036 218028
rect 331088 218016 331094 218068
rect 332226 218016 332232 218068
rect 332284 218056 332290 218068
rect 333606 218056 333612 218068
rect 332284 218028 333612 218056
rect 332284 218016 332290 218028
rect 333606 218016 333612 218028
rect 333664 218016 333670 218068
rect 334710 218016 334716 218068
rect 334768 218056 334774 218068
rect 335170 218056 335176 218068
rect 334768 218028 335176 218056
rect 334768 218016 334774 218028
rect 335170 218016 335176 218028
rect 335228 218016 335234 218068
rect 337194 218016 337200 218068
rect 337252 218056 337258 218068
rect 337746 218056 337752 218068
rect 337252 218028 337752 218056
rect 337252 218016 337258 218028
rect 337746 218016 337752 218028
rect 337804 218016 337810 218068
rect 338850 218016 338856 218068
rect 338908 218056 338914 218068
rect 339402 218056 339408 218068
rect 338908 218028 339408 218056
rect 338908 218016 338914 218028
rect 339402 218016 339408 218028
rect 339460 218016 339466 218068
rect 339678 218016 339684 218068
rect 339736 218056 339742 218068
rect 340690 218056 340696 218068
rect 339736 218028 340696 218056
rect 339736 218016 339742 218028
rect 340690 218016 340696 218028
rect 340748 218016 340754 218068
rect 345474 218016 345480 218068
rect 345532 218056 345538 218068
rect 347222 218056 347228 218068
rect 345532 218028 347228 218056
rect 345532 218016 345538 218028
rect 347222 218016 347228 218028
rect 347280 218016 347286 218068
rect 347958 218016 347964 218068
rect 348016 218056 348022 218068
rect 349062 218056 349068 218068
rect 348016 218028 349068 218056
rect 348016 218016 348022 218028
rect 349062 218016 349068 218028
rect 349120 218016 349126 218068
rect 349614 218016 349620 218068
rect 349672 218056 349678 218068
rect 350166 218056 350172 218068
rect 349672 218028 350172 218056
rect 349672 218016 349678 218028
rect 350166 218016 350172 218028
rect 350224 218016 350230 218068
rect 352098 218016 352104 218068
rect 352156 218056 352162 218068
rect 353294 218056 353300 218068
rect 352156 218028 353300 218056
rect 352156 218016 352162 218028
rect 353294 218016 353300 218028
rect 353352 218016 353358 218068
rect 356238 218016 356244 218068
rect 356296 218056 356302 218068
rect 357250 218056 357256 218068
rect 356296 218028 357256 218056
rect 356296 218016 356302 218028
rect 357250 218016 357256 218028
rect 357308 218016 357314 218068
rect 357894 218016 357900 218068
rect 357952 218056 357958 218068
rect 358538 218056 358544 218068
rect 357952 218028 358544 218056
rect 357952 218016 357958 218028
rect 358538 218016 358544 218028
rect 358596 218016 358602 218068
rect 359550 218016 359556 218068
rect 359608 218056 359614 218068
rect 360102 218056 360108 218068
rect 359608 218028 360108 218056
rect 359608 218016 359614 218028
rect 360102 218016 360108 218028
rect 360160 218016 360166 218068
rect 360378 218016 360384 218068
rect 360436 218056 360442 218068
rect 361022 218056 361028 218068
rect 360436 218028 361028 218056
rect 360436 218016 360442 218028
rect 361022 218016 361028 218028
rect 361080 218016 361086 218068
rect 367830 218016 367836 218068
rect 367888 218056 367894 218068
rect 368382 218056 368388 218068
rect 367888 218028 368388 218056
rect 367888 218016 367894 218028
rect 368382 218016 368388 218028
rect 368440 218016 368446 218068
rect 371970 218016 371976 218068
rect 372028 218056 372034 218068
rect 372522 218056 372528 218068
rect 372028 218028 372528 218056
rect 372028 218016 372034 218028
rect 372522 218016 372528 218028
rect 372580 218016 372586 218068
rect 372798 218016 372804 218068
rect 372856 218056 372862 218068
rect 373534 218056 373540 218068
rect 372856 218028 373540 218056
rect 372856 218016 372862 218028
rect 373534 218016 373540 218028
rect 373592 218016 373598 218068
rect 374454 218016 374460 218068
rect 374512 218056 374518 218068
rect 375006 218056 375012 218068
rect 374512 218028 375012 218056
rect 374512 218016 374518 218028
rect 375006 218016 375012 218028
rect 375064 218016 375070 218068
rect 376110 218016 376116 218068
rect 376168 218056 376174 218068
rect 376662 218056 376668 218068
rect 376168 218028 376668 218056
rect 376168 218016 376174 218028
rect 376662 218016 376668 218028
rect 376720 218016 376726 218068
rect 378594 218016 378600 218068
rect 378652 218056 378658 218068
rect 379238 218056 379244 218068
rect 378652 218028 379244 218056
rect 378652 218016 378658 218028
rect 379238 218016 379244 218028
rect 379296 218016 379302 218068
rect 381078 218016 381084 218068
rect 381136 218056 381142 218068
rect 382090 218056 382096 218068
rect 381136 218028 382096 218056
rect 381136 218016 381142 218028
rect 382090 218016 382096 218028
rect 382148 218016 382154 218068
rect 385218 218016 385224 218068
rect 385276 218056 385282 218068
rect 386046 218056 386052 218068
rect 385276 218028 386052 218056
rect 385276 218016 385282 218028
rect 386046 218016 386052 218028
rect 386104 218016 386110 218068
rect 389358 218016 389364 218068
rect 389416 218056 389422 218068
rect 390462 218056 390468 218068
rect 389416 218028 390468 218056
rect 389416 218016 389422 218028
rect 390462 218016 390468 218028
rect 390520 218016 390526 218068
rect 392670 218016 392676 218068
rect 392728 218056 392734 218068
rect 393130 218056 393136 218068
rect 392728 218028 393136 218056
rect 392728 218016 392734 218028
rect 393130 218016 393136 218028
rect 393188 218016 393194 218068
rect 393498 218016 393504 218068
rect 393556 218056 393562 218068
rect 394510 218056 394516 218068
rect 393556 218028 394516 218056
rect 393556 218016 393562 218028
rect 394510 218016 394516 218028
rect 394568 218016 394574 218068
rect 395154 218016 395160 218068
rect 395212 218056 395218 218068
rect 395798 218056 395804 218068
rect 395212 218028 395804 218056
rect 395212 218016 395218 218028
rect 395798 218016 395804 218028
rect 395856 218016 395862 218068
rect 397638 218016 397644 218068
rect 397696 218056 397702 218068
rect 401226 218056 401232 218068
rect 397696 218028 401232 218056
rect 397696 218016 397702 218028
rect 401226 218016 401232 218028
rect 401284 218016 401290 218068
rect 401778 218016 401784 218068
rect 401836 218056 401842 218068
rect 402790 218056 402796 218068
rect 401836 218028 402796 218056
rect 401836 218016 401842 218028
rect 402790 218016 402796 218028
rect 402848 218016 402854 218068
rect 403434 218016 403440 218068
rect 403492 218056 403498 218068
rect 403986 218056 403992 218068
rect 403492 218028 403992 218056
rect 403492 218016 403498 218028
rect 403986 218016 403992 218028
rect 404044 218016 404050 218068
rect 405090 218016 405096 218068
rect 405148 218056 405154 218068
rect 405550 218056 405556 218068
rect 405148 218028 405556 218056
rect 405148 218016 405154 218028
rect 405550 218016 405556 218028
rect 405608 218016 405614 218068
rect 409230 218016 409236 218068
rect 409288 218056 409294 218068
rect 409782 218056 409788 218068
rect 409288 218028 409788 218056
rect 409288 218016 409294 218028
rect 409782 218016 409788 218028
rect 409840 218016 409846 218068
rect 410058 218016 410064 218068
rect 410116 218056 410122 218068
rect 410702 218056 410708 218068
rect 410116 218028 410708 218056
rect 410116 218016 410122 218028
rect 410702 218016 410708 218028
rect 410760 218016 410766 218068
rect 413370 218016 413376 218068
rect 413428 218056 413434 218068
rect 413830 218056 413836 218068
rect 413428 218028 413836 218056
rect 413428 218016 413434 218028
rect 413830 218016 413836 218028
rect 413888 218016 413894 218068
rect 419994 218016 420000 218068
rect 420052 218056 420058 218068
rect 420914 218056 420920 218068
rect 420052 218028 420920 218056
rect 420052 218016 420058 218028
rect 420914 218016 420920 218028
rect 420972 218016 420978 218068
rect 424134 218016 424140 218068
rect 424192 218056 424198 218068
rect 426986 218056 426992 218068
rect 424192 218028 426992 218056
rect 424192 218016 424198 218028
rect 426986 218016 426992 218028
rect 427044 218016 427050 218068
rect 427446 218016 427452 218068
rect 427504 218056 427510 218068
rect 428274 218056 428280 218068
rect 427504 218028 428280 218056
rect 427504 218016 427510 218028
rect 428274 218016 428280 218028
rect 428332 218016 428338 218068
rect 429102 218016 429108 218068
rect 429160 218056 429166 218068
rect 430574 218056 430580 218068
rect 429160 218028 430580 218056
rect 429160 218016 429166 218028
rect 430574 218016 430580 218028
rect 430632 218016 430638 218068
rect 432414 218016 432420 218068
rect 432472 218056 432478 218068
rect 433794 218056 433800 218068
rect 432472 218028 433800 218056
rect 432472 218016 432478 218028
rect 433794 218016 433800 218028
rect 433852 218016 433858 218068
rect 434898 218016 434904 218068
rect 434956 218056 434962 218068
rect 436278 218056 436284 218068
rect 434956 218028 436284 218056
rect 434956 218016 434962 218028
rect 436278 218016 436284 218028
rect 436336 218016 436342 218068
rect 436554 218016 436560 218068
rect 436612 218056 436618 218068
rect 437474 218056 437480 218068
rect 436612 218028 437480 218056
rect 436612 218016 436618 218028
rect 437474 218016 437480 218028
rect 437532 218016 437538 218068
rect 438210 218016 438216 218068
rect 438268 218056 438274 218068
rect 438854 218056 438860 218068
rect 438268 218028 438860 218056
rect 438268 218016 438274 218028
rect 438854 218016 438860 218028
rect 438912 218016 438918 218068
rect 439866 218016 439872 218068
rect 439924 218056 439930 218068
rect 440326 218056 440332 218068
rect 439924 218028 440332 218056
rect 439924 218016 439930 218028
rect 440326 218016 440332 218028
rect 440384 218016 440390 218068
rect 453298 218016 453304 218068
rect 453356 218056 453362 218068
rect 455414 218056 455420 218068
rect 453356 218028 455420 218056
rect 453356 218016 453362 218028
rect 455414 218016 455420 218028
rect 455472 218016 455478 218068
rect 455598 218016 455604 218068
rect 455656 218056 455662 218068
rect 457162 218056 457168 218068
rect 455656 218028 457168 218056
rect 455656 218016 455662 218028
rect 457162 218016 457168 218028
rect 457220 218016 457226 218068
rect 463142 218016 463148 218068
rect 463200 218056 463206 218068
rect 464614 218056 464620 218068
rect 463200 218028 464620 218056
rect 463200 218016 463206 218028
rect 464614 218016 464620 218028
rect 464672 218016 464678 218068
rect 467282 218016 467288 218068
rect 467340 218056 467346 218068
rect 467926 218056 467932 218068
rect 467340 218028 467932 218056
rect 467340 218016 467346 218028
rect 467926 218016 467932 218028
rect 467984 218016 467990 218068
rect 492030 218016 492036 218068
rect 492088 218056 492094 218068
rect 505646 218056 505652 218068
rect 492088 218028 505652 218056
rect 492088 218016 492094 218028
rect 505646 218016 505652 218028
rect 505704 218016 505710 218068
rect 512730 218016 512736 218068
rect 512788 218056 512794 218068
rect 512788 218028 563100 218056
rect 512788 218016 512794 218028
rect 563072 217988 563100 218028
rect 563210 217988 563238 218096
rect 572438 218084 572444 218096
rect 572496 218084 572502 218136
rect 572622 218016 572628 218068
rect 572680 218056 572686 218068
rect 604638 218056 604644 218068
rect 572680 218028 604644 218056
rect 572680 218016 572686 218028
rect 604638 218016 604644 218028
rect 604696 218016 604702 218068
rect 563072 217960 563238 217988
rect 563606 217948 563612 218000
rect 563664 217988 563670 218000
rect 572438 217988 572444 218000
rect 563664 217960 572444 217988
rect 563664 217948 563670 217960
rect 572438 217948 572444 217960
rect 572496 217948 572502 218000
rect 675846 217948 675852 218000
rect 675904 217988 675910 218000
rect 676674 217988 676680 218000
rect 675904 217960 676680 217988
rect 675904 217948 675910 217960
rect 676674 217948 676680 217960
rect 676732 217948 676738 218000
rect 131022 217812 131028 217864
rect 131080 217852 131086 217864
rect 197722 217852 197728 217864
rect 131080 217824 197728 217852
rect 131080 217812 131086 217824
rect 197722 217812 197728 217824
rect 197780 217812 197786 217864
rect 523034 217812 523040 217864
rect 523092 217852 523098 217864
rect 524230 217852 524236 217864
rect 523092 217824 524236 217852
rect 523092 217812 523098 217824
rect 524230 217812 524236 217824
rect 524288 217812 524294 217864
rect 535454 217812 535460 217864
rect 535512 217852 535518 217864
rect 536650 217852 536656 217864
rect 535512 217824 536656 217852
rect 535512 217812 535518 217824
rect 536650 217812 536656 217824
rect 536708 217812 536714 217864
rect 598290 217852 598296 217864
rect 536852 217824 598296 217852
rect 116946 217676 116952 217728
rect 117004 217716 117010 217728
rect 189258 217716 189264 217728
rect 117004 217688 189264 217716
rect 117004 217676 117010 217688
rect 189258 217676 189264 217688
rect 189316 217676 189322 217728
rect 525978 217676 525984 217728
rect 526036 217716 526042 217728
rect 526530 217716 526536 217728
rect 526036 217688 526536 217716
rect 526036 217676 526042 217688
rect 526530 217676 526536 217688
rect 526588 217676 526594 217728
rect 533430 217676 533436 217728
rect 533488 217716 533494 217728
rect 536852 217716 536880 217824
rect 598290 217812 598296 217824
rect 598348 217812 598354 217864
rect 602982 217852 602988 217864
rect 598492 217824 602988 217852
rect 598492 217716 598520 217824
rect 602982 217812 602988 217824
rect 603040 217812 603046 217864
rect 603350 217812 603356 217864
rect 603408 217852 603414 217864
rect 613378 217852 613384 217864
rect 603408 217824 613384 217852
rect 603408 217812 603414 217824
rect 613378 217812 613384 217824
rect 613436 217812 613442 217864
rect 533488 217688 536880 217716
rect 536944 217688 598520 217716
rect 533488 217676 533494 217688
rect 103698 217540 103704 217592
rect 103756 217580 103762 217592
rect 178402 217580 178408 217592
rect 103756 217552 178408 217580
rect 103756 217540 103762 217552
rect 178402 217540 178408 217552
rect 178460 217540 178466 217592
rect 530946 217540 530952 217592
rect 531004 217580 531010 217592
rect 536944 217580 536972 217688
rect 598658 217676 598664 217728
rect 598716 217716 598722 217728
rect 604270 217716 604276 217728
rect 598716 217688 604276 217716
rect 598716 217676 598722 217688
rect 604270 217676 604276 217688
rect 604328 217676 604334 217728
rect 604638 217676 604644 217728
rect 604696 217716 604702 217728
rect 616874 217716 616880 217728
rect 604696 217688 616880 217716
rect 604696 217676 604702 217688
rect 616874 217676 616880 217688
rect 616932 217676 616938 217728
rect 531004 217552 536972 217580
rect 531004 217540 531010 217552
rect 538214 217540 538220 217592
rect 538272 217580 538278 217592
rect 539134 217580 539140 217592
rect 538272 217552 539140 217580
rect 538272 217540 538278 217552
rect 539134 217540 539140 217552
rect 539192 217540 539198 217592
rect 545758 217540 545764 217592
rect 545816 217580 545822 217592
rect 606754 217580 606760 217592
rect 545816 217552 606760 217580
rect 545816 217540 545822 217552
rect 606754 217540 606760 217552
rect 606812 217540 606818 217592
rect 92106 217404 92112 217456
rect 92164 217444 92170 217456
rect 170306 217444 170312 217456
rect 92164 217416 170312 217444
rect 92164 217404 92170 217416
rect 170306 217404 170312 217416
rect 170364 217404 170370 217456
rect 526530 217404 526536 217456
rect 526588 217444 526594 217456
rect 526588 217416 601602 217444
rect 526588 217404 526594 217416
rect 93762 217268 93768 217320
rect 93820 217308 93826 217320
rect 171226 217308 171232 217320
rect 93820 217280 171232 217308
rect 93820 217268 93826 217280
rect 171226 217268 171232 217280
rect 171284 217268 171290 217320
rect 535822 217268 535828 217320
rect 535880 217308 535886 217320
rect 598658 217308 598664 217320
rect 535880 217280 598664 217308
rect 535880 217268 535886 217280
rect 598658 217268 598664 217280
rect 598716 217268 598722 217320
rect 598842 217268 598848 217320
rect 598900 217308 598906 217320
rect 601142 217308 601148 217320
rect 598900 217280 601148 217308
rect 598900 217268 598906 217280
rect 601142 217268 601148 217280
rect 601200 217268 601206 217320
rect 601574 217308 601602 217416
rect 601878 217404 601884 217456
rect 601936 217444 601942 217456
rect 628282 217444 628288 217456
rect 601936 217416 628288 217444
rect 601936 217404 601942 217416
rect 628282 217404 628288 217416
rect 628340 217404 628346 217456
rect 602338 217308 602344 217320
rect 601574 217280 602344 217308
rect 602338 217268 602344 217280
rect 602396 217268 602402 217320
rect 602982 217268 602988 217320
rect 603040 217308 603046 217320
rect 603442 217308 603448 217320
rect 603040 217280 603448 217308
rect 603040 217268 603046 217280
rect 603442 217268 603448 217280
rect 603500 217268 603506 217320
rect 436094 217200 436100 217252
rect 436152 217240 436158 217252
rect 437336 217240 437342 217252
rect 436152 217212 437342 217240
rect 436152 217200 436158 217212
rect 437336 217200 437342 217212
rect 437394 217200 437400 217252
rect 447134 217200 447140 217252
rect 447192 217240 447198 217252
rect 448100 217240 448106 217252
rect 447192 217212 448106 217240
rect 447192 217200 447198 217212
rect 448100 217200 448106 217212
rect 448158 217200 448164 217252
rect 448606 217200 448612 217252
rect 448664 217240 448670 217252
rect 449756 217240 449762 217252
rect 448664 217212 449762 217240
rect 448664 217200 448670 217212
rect 449756 217200 449762 217212
rect 449814 217200 449820 217252
rect 469306 217200 469312 217252
rect 469364 217240 469370 217252
rect 470456 217240 470462 217252
rect 469364 217212 470462 217240
rect 469364 217200 469370 217212
rect 470456 217200 470462 217212
rect 470514 217200 470520 217252
rect 489914 217200 489920 217252
rect 489972 217240 489978 217252
rect 491156 217240 491162 217252
rect 489972 217212 491162 217240
rect 489972 217200 489978 217212
rect 491156 217200 491162 217212
rect 491214 217200 491220 217252
rect 498286 217200 498292 217252
rect 498344 217240 498350 217252
rect 499436 217240 499442 217252
rect 498344 217212 499442 217240
rect 498344 217200 498350 217212
rect 499436 217200 499442 217212
rect 499494 217200 499500 217252
rect 502978 217200 502984 217252
rect 503036 217240 503042 217252
rect 503576 217240 503582 217252
rect 503036 217212 503582 217240
rect 503036 217200 503042 217212
rect 503576 217200 503582 217212
rect 503634 217200 503640 217252
rect 511028 217132 511034 217184
rect 511086 217172 511092 217184
rect 562226 217172 562232 217184
rect 511086 217144 562232 217172
rect 511086 217132 511092 217144
rect 562226 217132 562232 217144
rect 562284 217132 562290 217184
rect 562502 217132 562508 217184
rect 562560 217132 562566 217184
rect 562686 217132 562692 217184
rect 562744 217132 562750 217184
rect 563054 217132 563060 217184
rect 563112 217172 563118 217184
rect 599026 217172 599032 217184
rect 563112 217144 599032 217172
rect 563112 217132 563118 217144
rect 599026 217132 599032 217144
rect 599084 217132 599090 217184
rect 600130 217132 600136 217184
rect 600188 217172 600194 217184
rect 603994 217172 604000 217184
rect 600188 217144 604000 217172
rect 600188 217132 600194 217144
rect 603994 217132 604000 217144
rect 604052 217132 604058 217184
rect 503576 217064 503582 217116
rect 503634 217104 503640 217116
rect 503634 217076 505094 217104
rect 503634 217064 503640 217076
rect 505066 217036 505094 217076
rect 562520 217036 562548 217132
rect 505066 217008 562548 217036
rect 562704 217036 562732 217132
rect 608962 217036 608968 217048
rect 562704 217008 608968 217036
rect 608962 216996 608968 217008
rect 609020 216996 609026 217048
rect 609882 216996 609888 217048
rect 609940 217036 609946 217048
rect 614114 217036 614120 217048
rect 609940 217008 614120 217036
rect 609940 216996 609946 217008
rect 614114 216996 614120 217008
rect 614172 216996 614178 217048
rect 574094 216860 574100 216912
rect 574152 216900 574158 216912
rect 597554 216900 597560 216912
rect 574152 216872 597560 216900
rect 574152 216860 574158 216872
rect 597554 216860 597560 216872
rect 597612 216860 597618 216912
rect 598290 216860 598296 216912
rect 598348 216900 598354 216912
rect 600130 216900 600136 216912
rect 598348 216872 600136 216900
rect 598348 216860 598354 216872
rect 600130 216860 600136 216872
rect 600188 216860 600194 216912
rect 612274 216900 612280 216912
rect 600976 216872 612280 216900
rect 594794 216724 594800 216776
rect 594852 216764 594858 216776
rect 600976 216764 601004 216872
rect 612274 216860 612280 216872
rect 612332 216860 612338 216912
rect 594852 216736 601004 216764
rect 594852 216724 594858 216736
rect 601142 216724 601148 216776
rect 601200 216764 601206 216776
rect 623866 216764 623872 216776
rect 601200 216736 623872 216764
rect 601200 216724 601206 216736
rect 623866 216724 623872 216736
rect 623924 216724 623930 216776
rect 675846 216452 675852 216504
rect 675904 216492 675910 216504
rect 676950 216492 676956 216504
rect 675904 216464 676956 216492
rect 675904 216452 675910 216464
rect 676950 216452 676956 216464
rect 677008 216452 677014 216504
rect 649902 215908 649908 215960
rect 649960 215948 649966 215960
rect 663058 215948 663064 215960
rect 649960 215920 663064 215948
rect 649960 215908 649966 215920
rect 663058 215908 663064 215920
rect 663116 215908 663122 215960
rect 676030 215296 676036 215348
rect 676088 215336 676094 215348
rect 676582 215336 676588 215348
rect 676088 215308 676588 215336
rect 676088 215296 676094 215308
rect 676582 215296 676588 215308
rect 676640 215296 676646 215348
rect 575474 214820 575480 214872
rect 575532 214860 575538 214872
rect 622302 214860 622308 214872
rect 575532 214832 622308 214860
rect 575532 214820 575538 214832
rect 622302 214820 622308 214832
rect 622360 214820 622366 214872
rect 574922 214684 574928 214736
rect 574980 214724 574986 214736
rect 616690 214724 616696 214736
rect 574980 214696 616696 214724
rect 574980 214684 574986 214696
rect 616690 214684 616696 214696
rect 616748 214684 616754 214736
rect 617058 214684 617064 214736
rect 617116 214724 617122 214736
rect 617794 214724 617800 214736
rect 617116 214696 617800 214724
rect 617116 214684 617122 214696
rect 617794 214684 617800 214696
rect 617852 214684 617858 214736
rect 619818 214684 619824 214736
rect 619876 214724 619882 214736
rect 620554 214724 620560 214736
rect 619876 214696 620560 214724
rect 619876 214684 619882 214696
rect 620554 214684 620560 214696
rect 620612 214684 620618 214736
rect 621014 214684 621020 214736
rect 621072 214724 621078 214736
rect 621658 214724 621664 214736
rect 621072 214696 621664 214724
rect 621072 214684 621078 214696
rect 621658 214684 621664 214696
rect 621716 214684 621722 214736
rect 622486 214684 622492 214736
rect 622544 214724 622550 214736
rect 623314 214724 623320 214736
rect 622544 214696 623320 214724
rect 622544 214684 622550 214696
rect 623314 214684 623320 214696
rect 623372 214684 623378 214736
rect 630030 214684 630036 214736
rect 630088 214724 630094 214736
rect 632882 214724 632888 214736
rect 630088 214696 632888 214724
rect 630088 214684 630094 214696
rect 632882 214684 632888 214696
rect 632940 214684 632946 214736
rect 574738 214548 574744 214600
rect 574796 214588 574802 214600
rect 625522 214588 625528 214600
rect 574796 214560 625528 214588
rect 574796 214548 574802 214560
rect 625522 214548 625528 214560
rect 625580 214548 625586 214600
rect 600498 214412 600504 214464
rect 600556 214452 600562 214464
rect 601234 214452 601240 214464
rect 600556 214424 601240 214452
rect 600556 214412 600562 214424
rect 601234 214412 601240 214424
rect 601292 214412 601298 214464
rect 605926 214412 605932 214464
rect 605984 214452 605990 214464
rect 606294 214452 606300 214464
rect 605984 214424 606300 214452
rect 605984 214412 605990 214424
rect 606294 214412 606300 214424
rect 606352 214412 606358 214464
rect 607306 214412 607312 214464
rect 607364 214452 607370 214464
rect 607858 214452 607864 214464
rect 607364 214424 607864 214452
rect 607364 214412 607370 214424
rect 607858 214412 607864 214424
rect 607916 214412 607922 214464
rect 611446 214412 611452 214464
rect 611504 214452 611510 214464
rect 611814 214452 611820 214464
rect 611504 214424 611820 214452
rect 611504 214412 611510 214424
rect 611814 214412 611820 214424
rect 611872 214412 611878 214464
rect 616690 214412 616696 214464
rect 616748 214452 616754 214464
rect 624418 214452 624424 214464
rect 616748 214424 624424 214452
rect 616748 214412 616754 214424
rect 624418 214412 624424 214424
rect 624476 214412 624482 214464
rect 653214 214412 653220 214464
rect 653272 214452 653278 214464
rect 660206 214452 660212 214464
rect 653272 214424 660212 214452
rect 653272 214412 653278 214424
rect 660206 214412 660212 214424
rect 660264 214412 660270 214464
rect 663426 214412 663432 214464
rect 663484 214452 663490 214464
rect 665818 214452 665824 214464
rect 663484 214424 665824 214452
rect 663484 214412 663490 214424
rect 665818 214412 665824 214424
rect 665876 214412 665882 214464
rect 626350 214276 626356 214328
rect 626408 214316 626414 214328
rect 628834 214316 628840 214328
rect 626408 214288 628840 214316
rect 626408 214276 626414 214288
rect 628834 214276 628840 214288
rect 628892 214276 628898 214328
rect 35802 214208 35808 214260
rect 35860 214248 35866 214260
rect 39666 214248 39672 214260
rect 35860 214220 39672 214248
rect 35860 214208 35866 214220
rect 39666 214208 39672 214220
rect 39724 214208 39730 214260
rect 646314 214208 646320 214260
rect 646372 214248 646378 214260
rect 653398 214248 653404 214260
rect 646372 214220 653404 214248
rect 646372 214208 646378 214220
rect 653398 214208 653404 214220
rect 653456 214208 653462 214260
rect 627454 213936 627460 213988
rect 627512 213976 627518 213988
rect 629386 213976 629392 213988
rect 627512 213948 629392 213976
rect 627512 213936 627518 213948
rect 629386 213936 629392 213948
rect 629444 213936 629450 213988
rect 663150 213868 663156 213920
rect 663208 213908 663214 213920
rect 663610 213908 663616 213920
rect 663208 213880 663616 213908
rect 663208 213868 663214 213880
rect 663610 213868 663616 213880
rect 663668 213868 663674 213920
rect 646038 213528 646044 213580
rect 646096 213568 646102 213580
rect 646498 213568 646504 213580
rect 646096 213540 646504 213568
rect 646096 213528 646102 213540
rect 646498 213528 646504 213540
rect 646556 213528 646562 213580
rect 652110 213528 652116 213580
rect 652168 213568 652174 213580
rect 654318 213568 654324 213580
rect 652168 213540 654324 213568
rect 652168 213528 652174 213540
rect 654318 213528 654324 213540
rect 654376 213528 654382 213580
rect 574094 213460 574100 213512
rect 574152 213500 574158 213512
rect 594794 213500 594800 213512
rect 574152 213472 594800 213500
rect 574152 213460 574158 213472
rect 594794 213460 594800 213472
rect 594852 213460 594858 213512
rect 574370 213324 574376 213376
rect 574428 213364 574434 213376
rect 612826 213364 612832 213376
rect 574428 213336 612832 213364
rect 574428 213324 574434 213336
rect 612826 213324 612832 213336
rect 612884 213324 612890 213376
rect 666002 213364 666008 213376
rect 644446 213336 666008 213364
rect 574554 213188 574560 213240
rect 574612 213228 574618 213240
rect 616138 213228 616144 213240
rect 574612 213200 616144 213228
rect 574612 213188 574618 213200
rect 616138 213188 616144 213200
rect 616196 213188 616202 213240
rect 643830 213188 643836 213240
rect 643888 213228 643894 213240
rect 644446 213228 644474 213336
rect 666002 213324 666008 213336
rect 666060 213324 666066 213376
rect 643888 213200 644474 213228
rect 643888 213188 643894 213200
rect 654594 213120 654600 213172
rect 654652 213160 654658 213172
rect 657538 213160 657544 213172
rect 654652 213132 657544 213160
rect 654652 213120 654658 213132
rect 657538 213120 657544 213132
rect 657596 213120 657602 213172
rect 654134 212984 654140 213036
rect 654192 213024 654198 213036
rect 654778 213024 654784 213036
rect 654192 212996 654784 213024
rect 654192 212984 654198 212996
rect 654778 212984 654784 212996
rect 654836 212984 654842 213036
rect 662046 212984 662052 213036
rect 662104 213024 662110 213036
rect 664714 213024 664720 213036
rect 662104 212996 664720 213024
rect 662104 212984 662110 212996
rect 664714 212984 664720 212996
rect 664772 212984 664778 213036
rect 645486 212848 645492 212900
rect 645544 212888 645550 212900
rect 651926 212888 651932 212900
rect 645544 212860 651932 212888
rect 645544 212848 645550 212860
rect 651926 212848 651932 212860
rect 651984 212848 651990 212900
rect 650454 212712 650460 212764
rect 650512 212752 650518 212764
rect 651282 212752 651288 212764
rect 650512 212724 651288 212752
rect 650512 212712 650518 212724
rect 651282 212712 651288 212724
rect 651340 212712 651346 212764
rect 658734 212712 658740 212764
rect 658792 212752 658798 212764
rect 659562 212752 659568 212764
rect 658792 212724 659568 212752
rect 658792 212712 658798 212724
rect 659562 212712 659568 212724
rect 659620 212712 659626 212764
rect 664254 212712 664260 212764
rect 664312 212752 664318 212764
rect 665082 212752 665088 212764
rect 664312 212724 665088 212752
rect 664312 212712 664318 212724
rect 665082 212712 665088 212724
rect 665140 212712 665146 212764
rect 632698 212508 632704 212560
rect 632756 212548 632762 212560
rect 634354 212548 634360 212560
rect 632756 212520 634360 212548
rect 632756 212508 632762 212520
rect 634354 212508 634360 212520
rect 634412 212508 634418 212560
rect 630674 212372 630680 212424
rect 630732 212412 630738 212424
rect 631594 212412 631600 212424
rect 630732 212384 631600 212412
rect 630732 212372 630738 212384
rect 631594 212372 631600 212384
rect 631652 212372 631658 212424
rect 35802 211556 35808 211608
rect 35860 211596 35866 211608
rect 35860 211556 35894 211596
rect 35866 211460 35894 211556
rect 41506 211460 41512 211472
rect 35866 211432 41512 211460
rect 41506 211420 41512 211432
rect 41564 211420 41570 211472
rect 35618 211284 35624 211336
rect 35676 211324 35682 211336
rect 41690 211324 41696 211336
rect 35676 211296 41696 211324
rect 35676 211284 35682 211296
rect 41690 211284 41696 211296
rect 41748 211284 41754 211336
rect 35802 211148 35808 211200
rect 35860 211188 35866 211200
rect 40126 211188 40132 211200
rect 35860 211160 40132 211188
rect 35860 211148 35866 211160
rect 40126 211148 40132 211160
rect 40184 211148 40190 211200
rect 578326 211148 578332 211200
rect 578384 211188 578390 211200
rect 580902 211188 580908 211200
rect 578384 211160 580908 211188
rect 578384 211148 578390 211160
rect 580902 211148 580908 211160
rect 580960 211148 580966 211200
rect 633434 211012 633440 211064
rect 633492 211052 633498 211064
rect 633802 211052 633808 211064
rect 633492 211024 633808 211052
rect 633492 211012 633498 211024
rect 633802 211012 633808 211024
rect 633860 211012 633866 211064
rect 35802 209924 35808 209976
rect 35860 209964 35866 209976
rect 40126 209964 40132 209976
rect 35860 209936 40132 209964
rect 35860 209924 35866 209936
rect 40126 209924 40132 209936
rect 40184 209924 40190 209976
rect 35526 209788 35532 209840
rect 35584 209828 35590 209840
rect 40770 209828 40776 209840
rect 35584 209800 40776 209828
rect 35584 209788 35590 209800
rect 40770 209788 40776 209800
rect 40828 209788 40834 209840
rect 579522 209788 579528 209840
rect 579580 209828 579586 209840
rect 582282 209828 582288 209840
rect 579580 209800 582288 209828
rect 579580 209788 579586 209800
rect 582282 209788 582288 209800
rect 582340 209788 582346 209840
rect 632146 209556 632152 209568
rect 625126 209528 632152 209556
rect 35802 208564 35808 208616
rect 35860 208604 35866 208616
rect 40954 208604 40960 208616
rect 35860 208576 40960 208604
rect 35860 208564 35866 208576
rect 40954 208564 40960 208576
rect 41012 208564 41018 208616
rect 581638 208564 581644 208616
rect 581696 208604 581702 208616
rect 625126 208604 625154 209528
rect 632146 209516 632152 209528
rect 632204 209516 632210 209568
rect 581696 208576 625154 208604
rect 581696 208564 581702 208576
rect 578878 208292 578884 208344
rect 578936 208332 578942 208344
rect 589458 208332 589464 208344
rect 578936 208304 589464 208332
rect 578936 208292 578942 208304
rect 589458 208292 589464 208304
rect 589516 208292 589522 208344
rect 35802 207204 35808 207256
rect 35860 207244 35866 207256
rect 40770 207244 40776 207256
rect 35860 207216 40776 207244
rect 35860 207204 35866 207216
rect 40770 207204 40776 207216
rect 40828 207204 40834 207256
rect 580902 206864 580908 206916
rect 580960 206904 580966 206916
rect 589458 206904 589464 206916
rect 580960 206876 589464 206904
rect 580960 206864 580966 206876
rect 589458 206864 589464 206876
rect 589516 206864 589522 206916
rect 579522 205776 579528 205828
rect 579580 205816 579586 205828
rect 580994 205816 581000 205828
rect 579580 205788 581000 205816
rect 579580 205776 579586 205788
rect 580994 205776 581000 205788
rect 581052 205776 581058 205828
rect 582282 205504 582288 205556
rect 582340 205544 582346 205556
rect 589458 205544 589464 205556
rect 582340 205516 589464 205544
rect 582340 205504 582346 205516
rect 589458 205504 589464 205516
rect 589516 205504 589522 205556
rect 35802 204416 35808 204468
rect 35860 204456 35866 204468
rect 41690 204456 41696 204468
rect 35860 204428 41696 204456
rect 35860 204416 35866 204428
rect 41690 204416 41696 204428
rect 41748 204416 41754 204468
rect 35618 204280 35624 204332
rect 35676 204320 35682 204332
rect 41690 204320 41696 204332
rect 35676 204292 41696 204320
rect 35676 204280 35682 204292
rect 41690 204280 41696 204292
rect 41748 204280 41754 204332
rect 579706 204212 579712 204264
rect 579764 204252 579770 204264
rect 589458 204252 589464 204264
rect 579764 204224 589464 204252
rect 579764 204212 579770 204224
rect 589458 204212 589464 204224
rect 589516 204212 589522 204264
rect 578326 202852 578332 202904
rect 578384 202892 578390 202904
rect 580258 202892 580264 202904
rect 578384 202864 580264 202892
rect 578384 202852 578390 202864
rect 580258 202852 580264 202864
rect 580316 202852 580322 202904
rect 580994 202784 581000 202836
rect 581052 202824 581058 202836
rect 589458 202824 589464 202836
rect 581052 202796 589464 202824
rect 581052 202784 581058 202796
rect 589458 202784 589464 202796
rect 589516 202784 589522 202836
rect 578786 200132 578792 200184
rect 578844 200172 578850 200184
rect 590378 200172 590384 200184
rect 578844 200144 590384 200172
rect 578844 200132 578850 200144
rect 590378 200132 590384 200144
rect 590436 200132 590442 200184
rect 580258 199996 580264 200048
rect 580316 200036 580322 200048
rect 589458 200036 589464 200048
rect 580316 200008 589464 200036
rect 580316 199996 580322 200008
rect 589458 199996 589464 200008
rect 589516 199996 589522 200048
rect 579522 198704 579528 198756
rect 579580 198744 579586 198756
rect 589458 198744 589464 198756
rect 579580 198716 589464 198744
rect 579580 198704 579586 198716
rect 589458 198704 589464 198716
rect 589516 198704 589522 198756
rect 578510 195984 578516 196036
rect 578568 196024 578574 196036
rect 589274 196024 589280 196036
rect 578568 195996 589280 196024
rect 578568 195984 578574 195996
rect 589274 195984 589280 195996
rect 589332 195984 589338 196036
rect 579522 194556 579528 194608
rect 579580 194596 579586 194608
rect 589458 194596 589464 194608
rect 579580 194568 589464 194596
rect 579580 194556 579586 194568
rect 589458 194556 589464 194568
rect 589516 194556 589522 194608
rect 579522 191836 579528 191888
rect 579580 191876 579586 191888
rect 589458 191876 589464 191888
rect 579580 191848 589464 191876
rect 579580 191836 579586 191848
rect 589458 191836 589464 191848
rect 589516 191836 589522 191888
rect 579522 190476 579528 190528
rect 579580 190516 579586 190528
rect 590562 190516 590568 190528
rect 579580 190488 590568 190516
rect 579580 190476 579586 190488
rect 590562 190476 590568 190488
rect 590620 190476 590626 190528
rect 579522 187688 579528 187740
rect 579580 187728 579586 187740
rect 589458 187728 589464 187740
rect 579580 187700 589464 187728
rect 579580 187688 579586 187700
rect 589458 187688 589464 187700
rect 589516 187688 589522 187740
rect 579522 186260 579528 186312
rect 579580 186300 579586 186312
rect 589642 186300 589648 186312
rect 579580 186272 589648 186300
rect 579580 186260 579586 186272
rect 589642 186260 589648 186272
rect 589700 186260 589706 186312
rect 579522 184832 579528 184884
rect 579580 184872 579586 184884
rect 589458 184872 589464 184884
rect 579580 184844 589464 184872
rect 579580 184832 579586 184844
rect 589458 184832 589464 184844
rect 589516 184832 589522 184884
rect 42150 183472 42156 183524
rect 42208 183512 42214 183524
rect 42978 183512 42984 183524
rect 42208 183484 42984 183512
rect 42208 183472 42214 183484
rect 42978 183472 42984 183484
rect 43036 183472 43042 183524
rect 42426 182112 42432 182164
rect 42484 182152 42490 182164
rect 43162 182152 43168 182164
rect 42484 182124 43168 182152
rect 42484 182112 42490 182124
rect 43162 182112 43168 182124
rect 43220 182112 43226 182164
rect 579522 182112 579528 182164
rect 579580 182152 579586 182164
rect 589458 182152 589464 182164
rect 579580 182124 589464 182152
rect 579580 182112 579586 182124
rect 589458 182112 589464 182124
rect 589516 182112 589522 182164
rect 578786 180752 578792 180804
rect 578844 180792 578850 180804
rect 590562 180792 590568 180804
rect 578844 180764 590568 180792
rect 578844 180752 578850 180764
rect 590562 180752 590568 180764
rect 590620 180752 590626 180804
rect 578786 178032 578792 178084
rect 578844 178072 578850 178084
rect 589458 178072 589464 178084
rect 578844 178044 589464 178072
rect 578844 178032 578850 178044
rect 589458 178032 589464 178044
rect 589516 178032 589522 178084
rect 579522 177896 579528 177948
rect 579580 177936 579586 177948
rect 589642 177936 589648 177948
rect 579580 177908 589648 177936
rect 579580 177896 579586 177908
rect 589642 177896 589648 177908
rect 589700 177896 589706 177948
rect 589458 175352 589464 175364
rect 586486 175324 589464 175352
rect 579982 175244 579988 175296
rect 580040 175284 580046 175296
rect 586486 175284 586514 175324
rect 589458 175312 589464 175324
rect 589516 175312 589522 175364
rect 580040 175256 586514 175284
rect 580040 175244 580046 175256
rect 668026 174700 668032 174752
rect 668084 174740 668090 174752
rect 670326 174740 670332 174752
rect 668084 174712 670332 174740
rect 668084 174700 668090 174712
rect 670326 174700 670332 174712
rect 670384 174700 670390 174752
rect 578418 174496 578424 174548
rect 578476 174536 578482 174548
rect 589642 174536 589648 174548
rect 578476 174508 589648 174536
rect 578476 174496 578482 174508
rect 589642 174496 589648 174508
rect 589700 174496 589706 174548
rect 667934 173068 667940 173120
rect 667992 173108 667998 173120
rect 669590 173108 669596 173120
rect 667992 173080 669596 173108
rect 667992 173068 667998 173080
rect 669590 173068 669596 173080
rect 669648 173068 669654 173120
rect 578234 172864 578240 172916
rect 578292 172904 578298 172916
rect 579982 172904 579988 172916
rect 578292 172876 579988 172904
rect 578292 172864 578298 172876
rect 579982 172864 579988 172876
rect 580040 172864 580046 172916
rect 580902 172524 580908 172576
rect 580960 172564 580966 172576
rect 589458 172564 589464 172576
rect 580960 172536 589464 172564
rect 580960 172524 580966 172536
rect 589458 172524 589464 172536
rect 589516 172524 589522 172576
rect 580258 171096 580264 171148
rect 580316 171136 580322 171148
rect 589458 171136 589464 171148
rect 580316 171108 589464 171136
rect 580316 171096 580322 171108
rect 589458 171096 589464 171108
rect 589516 171096 589522 171148
rect 578694 169736 578700 169788
rect 578752 169776 578758 169788
rect 580902 169776 580908 169788
rect 578752 169748 580908 169776
rect 578752 169736 578758 169748
rect 580902 169736 580908 169748
rect 580960 169736 580966 169788
rect 582374 168376 582380 168428
rect 582432 168416 582438 168428
rect 589458 168416 589464 168428
rect 582432 168388 589464 168416
rect 582432 168376 582438 168388
rect 589458 168376 589464 168388
rect 589516 168376 589522 168428
rect 668210 168172 668216 168224
rect 668268 168212 668274 168224
rect 670786 168212 670792 168224
rect 668268 168184 670792 168212
rect 668268 168172 668274 168184
rect 670786 168172 670792 168184
rect 670844 168172 670850 168224
rect 578234 167288 578240 167340
rect 578292 167328 578298 167340
rect 580258 167328 580264 167340
rect 578292 167300 580264 167328
rect 578292 167288 578298 167300
rect 580258 167288 580264 167300
rect 580316 167288 580322 167340
rect 579982 167016 579988 167068
rect 580040 167056 580046 167068
rect 589458 167056 589464 167068
rect 580040 167028 589464 167056
rect 580040 167016 580046 167028
rect 589458 167016 589464 167028
rect 589516 167016 589522 167068
rect 579522 166268 579528 166320
rect 579580 166308 579586 166320
rect 589642 166308 589648 166320
rect 579580 166280 589648 166308
rect 579580 166268 579586 166280
rect 589642 166268 589648 166280
rect 589700 166268 589706 166320
rect 579338 165180 579344 165232
rect 579396 165220 579402 165232
rect 582374 165220 582380 165232
rect 579396 165192 582380 165220
rect 579396 165180 579402 165192
rect 582374 165180 582380 165192
rect 582432 165180 582438 165232
rect 667934 164908 667940 164960
rect 667992 164948 667998 164960
rect 669774 164948 669780 164960
rect 667992 164920 669780 164948
rect 667992 164908 667998 164920
rect 669774 164908 669780 164920
rect 669832 164908 669838 164960
rect 582466 164228 582472 164280
rect 582524 164268 582530 164280
rect 589458 164268 589464 164280
rect 582524 164240 589464 164268
rect 582524 164228 582530 164240
rect 589458 164228 589464 164240
rect 589516 164228 589522 164280
rect 578234 163616 578240 163668
rect 578292 163656 578298 163668
rect 579982 163656 579988 163668
rect 578292 163628 579988 163656
rect 578292 163616 578298 163628
rect 579982 163616 579988 163628
rect 580040 163616 580046 163668
rect 580902 162868 580908 162920
rect 580960 162908 580966 162920
rect 589458 162908 589464 162920
rect 580960 162880 589464 162908
rect 580960 162868 580966 162880
rect 589458 162868 589464 162880
rect 589516 162868 589522 162920
rect 578418 162664 578424 162716
rect 578476 162704 578482 162716
rect 582466 162704 582472 162716
rect 578476 162676 582472 162704
rect 578476 162664 578482 162676
rect 582466 162664 582472 162676
rect 582524 162664 582530 162716
rect 675938 161712 675944 161764
rect 675996 161752 676002 161764
rect 679618 161752 679624 161764
rect 675996 161724 679624 161752
rect 675996 161712 676002 161724
rect 679618 161712 679624 161724
rect 679676 161712 679682 161764
rect 580534 161440 580540 161492
rect 580592 161480 580598 161492
rect 589458 161480 589464 161492
rect 580592 161452 589464 161480
rect 580592 161440 580598 161452
rect 589458 161440 589464 161452
rect 589516 161440 589522 161492
rect 580718 160080 580724 160132
rect 580776 160120 580782 160132
rect 589458 160120 589464 160132
rect 580776 160092 589464 160120
rect 580776 160080 580782 160092
rect 589458 160080 589464 160092
rect 589516 160080 589522 160132
rect 578878 158720 578884 158772
rect 578936 158760 578942 158772
rect 580902 158760 580908 158772
rect 578936 158732 580908 158760
rect 578936 158720 578942 158732
rect 580902 158720 580908 158732
rect 580960 158720 580966 158772
rect 585778 158720 585784 158772
rect 585836 158760 585842 158772
rect 589458 158760 589464 158772
rect 585836 158732 589464 158760
rect 585836 158720 585842 158732
rect 589458 158720 589464 158732
rect 589516 158720 589522 158772
rect 587158 157360 587164 157412
rect 587216 157400 587222 157412
rect 589274 157400 589280 157412
rect 587216 157372 589280 157400
rect 587216 157360 587222 157372
rect 589274 157360 589280 157372
rect 589332 157360 589338 157412
rect 578326 154776 578332 154828
rect 578384 154816 578390 154828
rect 580534 154816 580540 154828
rect 578384 154788 580540 154816
rect 578384 154776 578390 154788
rect 580534 154776 580540 154788
rect 580592 154776 580598 154828
rect 584398 154572 584404 154624
rect 584456 154612 584462 154624
rect 589458 154612 589464 154624
rect 584456 154584 589464 154612
rect 584456 154572 584462 154584
rect 589458 154572 589464 154584
rect 589516 154572 589522 154624
rect 583018 153212 583024 153264
rect 583076 153252 583082 153264
rect 589458 153252 589464 153264
rect 583076 153224 589464 153252
rect 583076 153212 583082 153224
rect 589458 153212 589464 153224
rect 589516 153212 589522 153264
rect 578234 152736 578240 152788
rect 578292 152776 578298 152788
rect 580718 152776 580724 152788
rect 578292 152748 580724 152776
rect 578292 152736 578298 152748
rect 580718 152736 580724 152748
rect 580776 152736 580782 152788
rect 580258 151784 580264 151836
rect 580316 151824 580322 151836
rect 589458 151824 589464 151836
rect 580316 151796 589464 151824
rect 580316 151784 580322 151796
rect 589458 151784 589464 151796
rect 589516 151784 589522 151836
rect 578878 150560 578884 150612
rect 578936 150600 578942 150612
rect 585778 150600 585784 150612
rect 578936 150572 585784 150600
rect 578936 150560 578942 150572
rect 585778 150560 585784 150572
rect 585836 150560 585842 150612
rect 585134 149064 585140 149116
rect 585192 149104 585198 149116
rect 589458 149104 589464 149116
rect 585192 149076 589464 149104
rect 585192 149064 585198 149076
rect 589458 149064 589464 149076
rect 589516 149064 589522 149116
rect 668394 149064 668400 149116
rect 668452 149104 668458 149116
rect 670786 149104 670792 149116
rect 668452 149076 670792 149104
rect 668452 149064 668458 149076
rect 670786 149064 670792 149076
rect 670844 149064 670850 149116
rect 579522 148316 579528 148368
rect 579580 148356 579586 148368
rect 587158 148356 587164 148368
rect 579580 148328 587164 148356
rect 579580 148316 579586 148328
rect 587158 148316 587164 148328
rect 587216 148316 587222 148368
rect 578878 146276 578884 146328
rect 578936 146316 578942 146328
rect 585134 146316 585140 146328
rect 578936 146288 585140 146316
rect 578936 146276 578942 146288
rect 585134 146276 585140 146288
rect 585192 146276 585198 146328
rect 584766 144916 584772 144968
rect 584824 144956 584830 144968
rect 589458 144956 589464 144968
rect 584824 144928 589464 144956
rect 584824 144916 584830 144928
rect 589458 144916 589464 144928
rect 589516 144916 589522 144968
rect 579246 144644 579252 144696
rect 579304 144684 579310 144696
rect 584398 144684 584404 144696
rect 579304 144656 584404 144684
rect 579304 144644 579310 144656
rect 584398 144644 584404 144656
rect 584456 144644 584462 144696
rect 585778 143556 585784 143608
rect 585836 143596 585842 143608
rect 589458 143596 589464 143608
rect 585836 143568 589464 143596
rect 585836 143556 585842 143568
rect 589458 143556 589464 143568
rect 589516 143556 589522 143608
rect 579522 143420 579528 143472
rect 579580 143460 579586 143472
rect 583018 143460 583024 143472
rect 579580 143432 583024 143460
rect 579580 143420 579586 143432
rect 583018 143420 583024 143432
rect 583076 143420 583082 143472
rect 587158 142400 587164 142452
rect 587216 142440 587222 142452
rect 589826 142440 589832 142452
rect 587216 142412 589832 142440
rect 587216 142400 587222 142412
rect 589826 142400 589832 142412
rect 589884 142400 589890 142452
rect 580442 140768 580448 140820
rect 580500 140808 580506 140820
rect 589458 140808 589464 140820
rect 580500 140780 589464 140808
rect 580500 140768 580506 140780
rect 589458 140768 589464 140780
rect 589516 140768 589522 140820
rect 578602 140700 578608 140752
rect 578660 140740 578666 140752
rect 580258 140740 580264 140752
rect 578660 140712 580264 140740
rect 578660 140700 578666 140712
rect 580258 140700 580264 140712
rect 580316 140700 580322 140752
rect 668210 140632 668216 140684
rect 668268 140672 668274 140684
rect 670786 140672 670792 140684
rect 668268 140644 670792 140672
rect 668268 140632 668274 140644
rect 670786 140632 670792 140644
rect 670844 140632 670850 140684
rect 583018 139408 583024 139460
rect 583076 139448 583082 139460
rect 589458 139448 589464 139460
rect 583076 139420 589464 139448
rect 583076 139408 583082 139420
rect 589458 139408 589464 139420
rect 589516 139408 589522 139460
rect 578602 139272 578608 139324
rect 578660 139312 578666 139324
rect 589918 139312 589924 139324
rect 578660 139284 589924 139312
rect 578660 139272 578666 139284
rect 589918 139272 589924 139284
rect 589976 139272 589982 139324
rect 579522 138660 579528 138712
rect 579580 138700 579586 138712
rect 588538 138700 588544 138712
rect 579580 138672 588544 138700
rect 579580 138660 579586 138672
rect 588538 138660 588544 138672
rect 588596 138660 588602 138712
rect 668578 137980 668584 138032
rect 668636 138020 668642 138032
rect 670142 138020 670148 138032
rect 668636 137992 670148 138020
rect 668636 137980 668642 137992
rect 670142 137980 670148 137992
rect 670200 137980 670206 138032
rect 579062 137300 579068 137352
rect 579120 137340 579126 137352
rect 584766 137340 584772 137352
rect 579120 137312 584772 137340
rect 579120 137300 579126 137312
rect 584766 137300 584772 137312
rect 584824 137300 584830 137352
rect 584582 136620 584588 136672
rect 584640 136660 584646 136672
rect 589458 136660 589464 136672
rect 584640 136632 589464 136660
rect 584640 136620 584646 136632
rect 589458 136620 589464 136632
rect 589516 136620 589522 136672
rect 580258 134512 580264 134564
rect 580316 134552 580322 134564
rect 589458 134552 589464 134564
rect 580316 134524 589464 134552
rect 580316 134512 580322 134524
rect 589458 134512 589464 134524
rect 589516 134512 589522 134564
rect 585962 132472 585968 132524
rect 586020 132512 586026 132524
rect 589458 132512 589464 132524
rect 586020 132484 589464 132512
rect 586020 132472 586026 132484
rect 589458 132472 589464 132484
rect 589516 132472 589522 132524
rect 581822 131248 581828 131300
rect 581880 131288 581886 131300
rect 589458 131288 589464 131300
rect 581880 131260 589464 131288
rect 581880 131248 581886 131260
rect 589458 131248 589464 131260
rect 589516 131248 589522 131300
rect 578878 131112 578884 131164
rect 578936 131152 578942 131164
rect 585778 131152 585784 131164
rect 578936 131124 585784 131152
rect 578936 131112 578942 131124
rect 585778 131112 585784 131124
rect 585836 131112 585842 131164
rect 667934 130636 667940 130688
rect 667992 130676 667998 130688
rect 669958 130676 669964 130688
rect 667992 130648 669964 130676
rect 667992 130636 667998 130648
rect 669958 130636 669964 130648
rect 670016 130636 670022 130688
rect 583386 129140 583392 129192
rect 583444 129180 583450 129192
rect 590378 129180 590384 129192
rect 583444 129152 590384 129180
rect 583444 129140 583450 129152
rect 590378 129140 590384 129152
rect 590436 129140 590442 129192
rect 579522 129004 579528 129056
rect 579580 129044 579586 129056
rect 587158 129044 587164 129056
rect 579580 129016 587164 129044
rect 579580 129004 579586 129016
rect 587158 129004 587164 129016
rect 587216 129004 587222 129056
rect 668762 128596 668768 128648
rect 668820 128636 668826 128648
rect 670786 128636 670792 128648
rect 668820 128608 670792 128636
rect 668820 128596 668826 128608
rect 670786 128596 670792 128608
rect 670844 128596 670850 128648
rect 587802 126964 587808 127016
rect 587860 127004 587866 127016
rect 589458 127004 589464 127016
rect 587860 126976 589464 127004
rect 587860 126964 587866 126976
rect 589458 126964 589464 126976
rect 589516 126964 589522 127016
rect 578326 125604 578332 125656
rect 578384 125644 578390 125656
rect 580442 125644 580448 125656
rect 578384 125616 580448 125644
rect 578384 125604 578390 125616
rect 580442 125604 580448 125616
rect 580500 125604 580506 125656
rect 676030 125400 676036 125452
rect 676088 125440 676094 125452
rect 676398 125440 676404 125452
rect 676088 125412 676404 125440
rect 676088 125400 676094 125412
rect 676398 125400 676404 125412
rect 676456 125400 676462 125452
rect 579062 124856 579068 124908
rect 579120 124896 579126 124908
rect 587802 124896 587808 124908
rect 579120 124868 587808 124896
rect 579120 124856 579126 124868
rect 587802 124856 587808 124868
rect 587860 124856 587866 124908
rect 578694 124108 578700 124160
rect 578752 124148 578758 124160
rect 583018 124148 583024 124160
rect 578752 124120 583024 124148
rect 578752 124108 578758 124120
rect 583018 124108 583024 124120
rect 583076 124108 583082 124160
rect 584398 122816 584404 122868
rect 584456 122856 584462 122868
rect 589458 122856 589464 122868
rect 584456 122828 589464 122856
rect 584456 122816 584462 122828
rect 589458 122816 589464 122828
rect 589516 122816 589522 122868
rect 578878 122136 578884 122188
rect 578936 122176 578942 122188
rect 584582 122176 584588 122188
rect 578936 122148 584588 122176
rect 578936 122136 578942 122148
rect 584582 122136 584588 122148
rect 584640 122136 584646 122188
rect 580626 122000 580632 122052
rect 580684 122040 580690 122052
rect 590102 122040 590108 122052
rect 580684 122012 590108 122040
rect 580684 122000 580690 122012
rect 590102 122000 590108 122012
rect 590160 122000 590166 122052
rect 587342 121456 587348 121508
rect 587400 121496 587406 121508
rect 589274 121496 589280 121508
rect 587400 121468 589280 121496
rect 587400 121456 587406 121468
rect 589274 121456 589280 121468
rect 589332 121456 589338 121508
rect 583202 120708 583208 120760
rect 583260 120748 583266 120760
rect 590562 120748 590568 120760
rect 583260 120720 590568 120748
rect 583260 120708 583266 120720
rect 590562 120708 590568 120720
rect 590620 120708 590626 120760
rect 578510 118532 578516 118584
rect 578568 118572 578574 118584
rect 580258 118572 580264 118584
rect 578568 118544 580264 118572
rect 578568 118532 578574 118544
rect 580258 118532 580264 118544
rect 580316 118532 580322 118584
rect 579522 116900 579528 116952
rect 579580 116940 579586 116952
rect 583386 116940 583392 116952
rect 579580 116912 583392 116940
rect 579580 116900 579586 116912
rect 583386 116900 583392 116912
rect 583444 116900 583450 116952
rect 675846 116628 675852 116680
rect 675904 116668 675910 116680
rect 678238 116668 678244 116680
rect 675904 116640 678244 116668
rect 675904 116628 675910 116640
rect 678238 116628 678244 116640
rect 678296 116628 678302 116680
rect 585778 115948 585784 116000
rect 585836 115988 585842 116000
rect 589458 115988 589464 116000
rect 585836 115960 589464 115988
rect 585836 115948 585842 115960
rect 589458 115948 589464 115960
rect 589516 115948 589522 116000
rect 584582 115200 584588 115252
rect 584640 115240 584646 115252
rect 589642 115240 589648 115252
rect 584640 115212 589648 115240
rect 584640 115200 584646 115212
rect 589642 115200 589648 115212
rect 589700 115200 589706 115252
rect 579246 114452 579252 114504
rect 579304 114492 579310 114504
rect 581638 114492 581644 114504
rect 579304 114464 581644 114492
rect 579304 114452 579310 114464
rect 581638 114452 581644 114464
rect 581696 114452 581702 114504
rect 583018 113160 583024 113212
rect 583076 113200 583082 113212
rect 589458 113200 589464 113212
rect 583076 113172 589464 113200
rect 583076 113160 583082 113172
rect 589458 113160 589464 113172
rect 589516 113160 589522 113212
rect 579522 112820 579528 112872
rect 579580 112860 579586 112872
rect 585962 112860 585968 112872
rect 579580 112832 585968 112860
rect 579580 112820 579586 112832
rect 585962 112820 585968 112832
rect 586020 112820 586026 112872
rect 586146 112412 586152 112464
rect 586204 112452 586210 112464
rect 590102 112452 590108 112464
rect 586204 112424 590108 112452
rect 586204 112412 586210 112424
rect 590102 112412 590108 112424
rect 590160 112412 590166 112464
rect 581638 110440 581644 110492
rect 581696 110480 581702 110492
rect 589458 110480 589464 110492
rect 581696 110452 589464 110480
rect 581696 110440 581702 110452
rect 589458 110440 589464 110452
rect 589516 110440 589522 110492
rect 579338 110236 579344 110288
rect 579396 110276 579402 110288
rect 581822 110276 581828 110288
rect 579396 110248 581828 110276
rect 579396 110236 579402 110248
rect 581822 110236 581828 110248
rect 581880 110236 581886 110288
rect 580442 109080 580448 109132
rect 580500 109120 580506 109132
rect 589458 109120 589464 109132
rect 580500 109092 589464 109120
rect 580500 109080 580506 109092
rect 589458 109080 589464 109092
rect 589516 109080 589522 109132
rect 578326 108944 578332 108996
rect 578384 108984 578390 108996
rect 580626 108984 580632 108996
rect 578384 108956 580632 108984
rect 578384 108944 578390 108956
rect 580626 108944 580632 108956
rect 580684 108944 580690 108996
rect 667934 107992 667940 108044
rect 667992 108032 667998 108044
rect 670142 108032 670148 108044
rect 667992 108004 670148 108032
rect 667992 107992 667998 108004
rect 670142 107992 670148 108004
rect 670200 107992 670206 108044
rect 582282 107652 582288 107704
rect 582340 107692 582346 107704
rect 589458 107692 589464 107704
rect 582340 107664 589464 107692
rect 582340 107652 582346 107664
rect 589458 107652 589464 107664
rect 589516 107652 589522 107704
rect 580258 106292 580264 106344
rect 580316 106332 580322 106344
rect 589458 106332 589464 106344
rect 580316 106304 589464 106332
rect 580316 106292 580322 106304
rect 589458 106292 589464 106304
rect 589516 106292 589522 106344
rect 668394 106156 668400 106208
rect 668452 106196 668458 106208
rect 670786 106196 670792 106208
rect 668452 106168 670792 106196
rect 668452 106156 668458 106168
rect 670786 106156 670792 106168
rect 670844 106156 670850 106208
rect 579338 105612 579344 105664
rect 579396 105652 579402 105664
rect 582282 105652 582288 105664
rect 579396 105624 582288 105652
rect 579396 105612 579402 105624
rect 582282 105612 582288 105624
rect 582340 105612 582346 105664
rect 587158 104864 587164 104916
rect 587216 104904 587222 104916
rect 589826 104904 589832 104916
rect 587216 104876 589832 104904
rect 587216 104864 587222 104876
rect 589826 104864 589832 104876
rect 589884 104864 589890 104916
rect 668302 104796 668308 104848
rect 668360 104836 668366 104848
rect 670786 104836 670792 104848
rect 668360 104808 670792 104836
rect 668360 104796 668366 104808
rect 670786 104796 670792 104808
rect 670844 104796 670850 104848
rect 578510 103368 578516 103420
rect 578568 103408 578574 103420
rect 588722 103408 588728 103420
rect 578568 103380 588728 103408
rect 578568 103368 578574 103380
rect 588722 103368 588728 103380
rect 588780 103368 588786 103420
rect 579154 102076 579160 102128
rect 579212 102116 579218 102128
rect 584398 102116 584404 102128
rect 579212 102088 584404 102116
rect 579212 102076 579218 102088
rect 584398 102076 584404 102088
rect 584456 102076 584462 102128
rect 584398 100104 584404 100156
rect 584456 100144 584462 100156
rect 589458 100144 589464 100156
rect 584456 100116 589464 100144
rect 584456 100104 584462 100116
rect 589458 100104 589464 100116
rect 589516 100104 589522 100156
rect 578602 99968 578608 100020
rect 578660 100008 578666 100020
rect 587342 100008 587348 100020
rect 578660 99980 587348 100008
rect 578660 99968 578666 99980
rect 587342 99968 587348 99980
rect 587400 99968 587406 100020
rect 592678 99968 592684 100020
rect 592736 100008 592742 100020
rect 667934 100008 667940 100020
rect 592736 99980 667940 100008
rect 592736 99968 592742 99980
rect 667934 99968 667940 99980
rect 667992 99968 667998 100020
rect 622302 99288 622308 99340
rect 622360 99328 622366 99340
rect 630766 99328 630772 99340
rect 622360 99300 630772 99328
rect 622360 99288 622366 99300
rect 630766 99288 630772 99300
rect 630824 99288 630830 99340
rect 579522 99220 579528 99272
rect 579580 99260 579586 99272
rect 583202 99260 583208 99272
rect 579580 99232 583208 99260
rect 579580 99220 579586 99232
rect 583202 99220 583208 99232
rect 583260 99220 583266 99272
rect 623682 99152 623688 99204
rect 623740 99192 623746 99204
rect 633434 99192 633440 99204
rect 623740 99164 633440 99192
rect 623740 99152 623746 99164
rect 633434 99152 633440 99164
rect 633492 99152 633498 99204
rect 577498 99084 577504 99136
rect 577556 99124 577562 99136
rect 595254 99124 595260 99136
rect 577556 99096 595260 99124
rect 577556 99084 577562 99096
rect 595254 99084 595260 99096
rect 595312 99084 595318 99136
rect 624602 99016 624608 99068
rect 624660 99056 624666 99068
rect 634998 99056 635004 99068
rect 624660 99028 635004 99056
rect 624660 99016 624666 99028
rect 634998 99016 635004 99028
rect 635056 99016 635062 99068
rect 625062 98880 625068 98932
rect 625120 98920 625126 98932
rect 636286 98920 636292 98932
rect 625120 98892 636292 98920
rect 625120 98880 625126 98892
rect 636286 98880 636292 98892
rect 636344 98880 636350 98932
rect 629018 98744 629024 98796
rect 629076 98784 629082 98796
rect 643646 98784 643652 98796
rect 629076 98756 643652 98784
rect 629076 98744 629082 98756
rect 643646 98744 643652 98756
rect 643704 98744 643710 98796
rect 647142 98744 647148 98796
rect 647200 98784 647206 98796
rect 661954 98784 661960 98796
rect 647200 98756 661960 98784
rect 647200 98744 647206 98756
rect 661954 98744 661960 98756
rect 662012 98744 662018 98796
rect 630490 98608 630496 98660
rect 630548 98648 630554 98660
rect 646590 98648 646596 98660
rect 630548 98620 646596 98648
rect 630548 98608 630554 98620
rect 646590 98608 646596 98620
rect 646648 98608 646654 98660
rect 631410 98268 631416 98320
rect 631468 98308 631474 98320
rect 642174 98308 642180 98320
rect 631468 98280 642180 98308
rect 631468 98268 631474 98280
rect 642174 98268 642180 98280
rect 642232 98268 642238 98320
rect 633618 98132 633624 98184
rect 633676 98172 633682 98184
rect 640702 98172 640708 98184
rect 633676 98144 640708 98172
rect 633676 98132 633682 98144
rect 640702 98132 640708 98144
rect 640760 98132 640766 98184
rect 631980 98076 632192 98104
rect 618714 97928 618720 97980
rect 618772 97968 618778 97980
rect 625798 97968 625804 97980
rect 618772 97940 625804 97968
rect 618772 97928 618778 97940
rect 625798 97928 625804 97940
rect 625856 97928 625862 97980
rect 629754 97928 629760 97980
rect 629812 97968 629818 97980
rect 631980 97968 632008 98076
rect 632164 98036 632192 98076
rect 645302 98036 645308 98048
rect 632164 98008 645308 98036
rect 645302 97996 645308 98008
rect 645360 97996 645366 98048
rect 629812 97940 632008 97968
rect 629812 97928 629818 97940
rect 659194 97928 659200 97980
rect 659252 97968 659258 97980
rect 664162 97968 664168 97980
rect 659252 97940 664168 97968
rect 659252 97928 659258 97940
rect 664162 97928 664168 97940
rect 664220 97928 664226 97980
rect 628282 97792 628288 97844
rect 628340 97832 628346 97844
rect 631410 97832 631416 97844
rect 628340 97804 631416 97832
rect 628340 97792 628346 97804
rect 631410 97792 631416 97804
rect 631468 97792 631474 97844
rect 632698 97792 632704 97844
rect 632756 97832 632762 97844
rect 647510 97832 647516 97844
rect 632756 97804 647516 97832
rect 632756 97792 632762 97804
rect 647510 97792 647516 97804
rect 647568 97792 647574 97844
rect 655238 97792 655244 97844
rect 655296 97832 655302 97844
rect 659746 97832 659752 97844
rect 655296 97804 659752 97832
rect 655296 97792 655302 97804
rect 659746 97792 659752 97804
rect 659804 97792 659810 97844
rect 659930 97792 659936 97844
rect 659988 97832 659994 97844
rect 665358 97832 665364 97844
rect 659988 97804 665364 97832
rect 659988 97792 659994 97804
rect 665358 97792 665364 97804
rect 665416 97792 665422 97844
rect 631226 97656 631232 97708
rect 631284 97696 631290 97708
rect 647326 97696 647332 97708
rect 631284 97668 647332 97696
rect 631284 97656 631290 97668
rect 647326 97656 647332 97668
rect 647384 97656 647390 97708
rect 651834 97656 651840 97708
rect 651892 97696 651898 97708
rect 659562 97696 659568 97708
rect 651892 97668 659568 97696
rect 651892 97656 651898 97668
rect 659562 97656 659568 97668
rect 659620 97656 659626 97708
rect 627546 97520 627552 97572
rect 627604 97560 627610 97572
rect 633618 97560 633624 97572
rect 627604 97532 633624 97560
rect 627604 97520 627610 97532
rect 633618 97520 633624 97532
rect 633676 97520 633682 97572
rect 633802 97520 633808 97572
rect 633860 97560 633866 97572
rect 637758 97560 637764 97572
rect 633860 97532 637764 97560
rect 633860 97520 633866 97532
rect 637758 97520 637764 97532
rect 637816 97520 637822 97572
rect 643002 97520 643008 97572
rect 643060 97560 643066 97572
rect 655238 97560 655244 97572
rect 643060 97532 655244 97560
rect 643060 97520 643066 97532
rect 655238 97520 655244 97532
rect 655296 97520 655302 97572
rect 655422 97520 655428 97572
rect 655480 97560 655486 97572
rect 662506 97560 662512 97572
rect 655480 97532 662512 97560
rect 655480 97520 655486 97532
rect 662506 97520 662512 97532
rect 662564 97520 662570 97572
rect 605466 97384 605472 97436
rect 605524 97424 605530 97436
rect 611906 97424 611912 97436
rect 605524 97396 611912 97424
rect 605524 97384 605530 97396
rect 611906 97384 611912 97396
rect 611964 97384 611970 97436
rect 612642 97384 612648 97436
rect 612700 97424 612706 97436
rect 620278 97424 620284 97436
rect 612700 97396 620284 97424
rect 612700 97384 612706 97396
rect 620278 97384 620284 97396
rect 620336 97384 620342 97436
rect 621658 97384 621664 97436
rect 621716 97424 621722 97436
rect 629294 97424 629300 97436
rect 621716 97396 629300 97424
rect 621716 97384 621722 97396
rect 629294 97384 629300 97396
rect 629352 97384 629358 97436
rect 631962 97384 631968 97436
rect 632020 97424 632026 97436
rect 648614 97424 648620 97436
rect 632020 97396 648620 97424
rect 632020 97384 632026 97396
rect 648614 97384 648620 97396
rect 648672 97384 648678 97436
rect 653950 97384 653956 97436
rect 654008 97424 654014 97436
rect 655238 97424 655244 97436
rect 654008 97396 655244 97424
rect 654008 97384 654014 97396
rect 655238 97384 655244 97396
rect 655296 97384 655302 97436
rect 658182 97384 658188 97436
rect 658240 97424 658246 97436
rect 663058 97424 663064 97436
rect 658240 97396 663064 97424
rect 658240 97384 658246 97396
rect 663058 97384 663064 97396
rect 663116 97384 663122 97436
rect 623130 97248 623136 97300
rect 623188 97288 623194 97300
rect 632054 97288 632060 97300
rect 623188 97260 632060 97288
rect 623188 97248 623194 97260
rect 632054 97248 632060 97260
rect 632112 97248 632118 97300
rect 633250 97248 633256 97300
rect 633308 97288 633314 97300
rect 633308 97260 649994 97288
rect 633308 97248 633314 97260
rect 620094 97112 620100 97164
rect 620152 97152 620158 97164
rect 626442 97152 626448 97164
rect 620152 97124 626448 97152
rect 620152 97112 620158 97124
rect 626442 97112 626448 97124
rect 626500 97112 626506 97164
rect 634170 97112 634176 97164
rect 634228 97152 634234 97164
rect 649074 97152 649080 97164
rect 634228 97124 649080 97152
rect 634228 97112 634234 97124
rect 649074 97112 649080 97124
rect 649132 97112 649138 97164
rect 649966 97152 649994 97260
rect 650362 97248 650368 97300
rect 650420 97288 650426 97300
rect 658274 97288 658280 97300
rect 650420 97260 658280 97288
rect 650420 97248 650426 97260
rect 658274 97248 658280 97260
rect 658332 97248 658338 97300
rect 650546 97152 650552 97164
rect 649966 97124 650552 97152
rect 650546 97112 650552 97124
rect 650604 97112 650610 97164
rect 656802 97112 656808 97164
rect 656860 97152 656866 97164
rect 661402 97152 661408 97164
rect 656860 97124 661408 97152
rect 656860 97112 656866 97124
rect 661402 97112 661408 97124
rect 661460 97112 661466 97164
rect 626074 96976 626080 97028
rect 626132 97016 626138 97028
rect 633802 97016 633808 97028
rect 626132 96988 633808 97016
rect 626132 96976 626138 96988
rect 633802 96976 633808 96988
rect 633860 96976 633866 97028
rect 634722 96976 634728 97028
rect 634780 97016 634786 97028
rect 647050 97016 647056 97028
rect 634780 96988 647056 97016
rect 634780 96976 634786 96988
rect 647050 96976 647056 96988
rect 647108 96976 647114 97028
rect 597646 96908 597652 96960
rect 597704 96948 597710 96960
rect 598198 96948 598204 96960
rect 597704 96920 598204 96948
rect 597704 96908 597710 96920
rect 598198 96908 598204 96920
rect 598256 96908 598262 96960
rect 600314 96908 600320 96960
rect 600372 96948 600378 96960
rect 601142 96948 601148 96960
rect 600372 96920 601148 96948
rect 600372 96908 600378 96920
rect 601142 96908 601148 96920
rect 601200 96908 601206 96960
rect 606202 96908 606208 96960
rect 606260 96948 606266 96960
rect 607122 96948 607128 96960
rect 606260 96920 607128 96948
rect 606260 96908 606266 96920
rect 607122 96908 607128 96920
rect 607180 96908 607186 96960
rect 615770 96908 615776 96960
rect 615828 96948 615834 96960
rect 616782 96948 616788 96960
rect 615828 96920 616788 96948
rect 615828 96908 615834 96920
rect 616782 96908 616788 96920
rect 616840 96908 616846 96960
rect 656710 96908 656716 96960
rect 656768 96948 656774 96960
rect 660114 96948 660120 96960
rect 656768 96920 660120 96948
rect 656768 96908 656774 96920
rect 660114 96908 660120 96920
rect 660172 96908 660178 96960
rect 612090 96840 612096 96892
rect 612148 96880 612154 96892
rect 612642 96880 612648 96892
rect 612148 96852 612648 96880
rect 612148 96840 612154 96852
rect 612642 96840 612648 96852
rect 612700 96840 612706 96892
rect 617242 96840 617248 96892
rect 617300 96880 617306 96892
rect 618162 96880 618168 96892
rect 617300 96852 618168 96880
rect 617300 96840 617306 96852
rect 618162 96840 618168 96852
rect 618220 96840 618226 96892
rect 626810 96840 626816 96892
rect 626868 96880 626874 96892
rect 639230 96880 639236 96892
rect 626868 96852 639236 96880
rect 626868 96840 626874 96852
rect 639230 96840 639236 96852
rect 639288 96840 639294 96892
rect 644290 96840 644296 96892
rect 644348 96880 644354 96892
rect 644348 96852 656572 96880
rect 644348 96840 644354 96852
rect 656544 96812 656572 96852
rect 658826 96812 658832 96824
rect 656544 96784 658832 96812
rect 658826 96772 658832 96784
rect 658884 96772 658890 96824
rect 609146 96704 609152 96756
rect 609204 96744 609210 96756
rect 609698 96744 609704 96756
rect 609204 96716 609704 96744
rect 609204 96704 609210 96716
rect 609698 96704 609704 96716
rect 609756 96704 609762 96756
rect 654778 96704 654784 96756
rect 654836 96744 654842 96756
rect 655422 96744 655428 96756
rect 654836 96716 655428 96744
rect 654836 96704 654842 96716
rect 655422 96704 655428 96716
rect 655480 96704 655486 96756
rect 640058 96568 640064 96620
rect 640116 96608 640122 96620
rect 645118 96608 645124 96620
rect 640116 96580 645124 96608
rect 640116 96568 640122 96580
rect 645118 96568 645124 96580
rect 645176 96568 645182 96620
rect 646406 96568 646412 96620
rect 646464 96608 646470 96620
rect 652202 96608 652208 96620
rect 646464 96580 652208 96608
rect 646464 96568 646470 96580
rect 652202 96568 652208 96580
rect 652260 96568 652266 96620
rect 652570 96568 652576 96620
rect 652628 96608 652634 96620
rect 664346 96608 664352 96620
rect 652628 96580 664352 96608
rect 652628 96568 652634 96580
rect 664346 96568 664352 96580
rect 664404 96568 664410 96620
rect 638586 96432 638592 96484
rect 638644 96472 638650 96484
rect 641346 96472 641352 96484
rect 638644 96444 641352 96472
rect 638644 96432 638650 96444
rect 641346 96432 641352 96444
rect 641404 96432 641410 96484
rect 641530 96432 641536 96484
rect 641588 96472 641594 96484
rect 648062 96472 648068 96484
rect 641588 96444 648068 96472
rect 641588 96432 641594 96444
rect 648062 96432 648068 96444
rect 648120 96432 648126 96484
rect 648890 96432 648896 96484
rect 648948 96472 648954 96484
rect 664530 96472 664536 96484
rect 648948 96444 664536 96472
rect 648948 96432 648954 96444
rect 664530 96432 664536 96444
rect 664588 96432 664594 96484
rect 648264 96376 648568 96404
rect 637574 96296 637580 96348
rect 637632 96336 637638 96348
rect 648264 96336 648292 96376
rect 637632 96308 648292 96336
rect 648540 96336 648568 96376
rect 660666 96336 660672 96348
rect 648540 96308 660672 96336
rect 637632 96296 637638 96308
rect 660666 96296 660672 96308
rect 660724 96296 660730 96348
rect 645486 96160 645492 96212
rect 645544 96200 645550 96212
rect 647878 96200 647884 96212
rect 645544 96172 647884 96200
rect 645544 96160 645550 96172
rect 647878 96160 647884 96172
rect 647936 96160 647942 96212
rect 649258 96160 649264 96212
rect 649316 96200 649322 96212
rect 663794 96200 663800 96212
rect 649316 96172 663800 96200
rect 649316 96160 649322 96172
rect 663794 96160 663800 96172
rect 663852 96160 663858 96212
rect 640518 96092 640524 96144
rect 640576 96132 640582 96144
rect 644934 96132 644940 96144
rect 640576 96104 644940 96132
rect 640576 96092 640582 96104
rect 644934 96092 644940 96104
rect 644992 96092 644998 96144
rect 591298 96024 591304 96076
rect 591356 96064 591362 96076
rect 602614 96064 602620 96076
rect 591356 96036 602620 96064
rect 591356 96024 591362 96036
rect 602614 96024 602620 96036
rect 602672 96024 602678 96076
rect 610618 96024 610624 96076
rect 610676 96064 610682 96076
rect 621658 96064 621664 96076
rect 610676 96036 621664 96064
rect 610676 96024 610682 96036
rect 621658 96024 621664 96036
rect 621716 96024 621722 96076
rect 645762 96024 645768 96076
rect 645820 96064 645826 96076
rect 648062 96064 648068 96076
rect 645820 96036 648068 96064
rect 645820 96024 645826 96036
rect 648062 96024 648068 96036
rect 648120 96024 648126 96076
rect 648614 96024 648620 96076
rect 648672 96064 648678 96076
rect 663978 96064 663984 96076
rect 648672 96036 663984 96064
rect 648672 96024 648678 96036
rect 663978 96024 663984 96036
rect 664036 96024 664042 96076
rect 594058 95888 594064 95940
rect 594116 95928 594122 95940
rect 668118 95928 668124 95940
rect 594116 95900 668124 95928
rect 594116 95888 594122 95900
rect 668118 95888 668124 95900
rect 668176 95888 668182 95940
rect 598934 95752 598940 95804
rect 598992 95792 598998 95804
rect 599670 95792 599676 95804
rect 598992 95764 599676 95792
rect 598992 95752 598998 95764
rect 599670 95752 599676 95764
rect 599728 95752 599734 95804
rect 639046 95752 639052 95804
rect 639104 95792 639110 95804
rect 648614 95792 648620 95804
rect 639104 95764 648620 95792
rect 639104 95752 639110 95764
rect 648614 95752 648620 95764
rect 648672 95752 648678 95804
rect 653306 95752 653312 95804
rect 653364 95792 653370 95804
rect 665174 95792 665180 95804
rect 653364 95764 665180 95792
rect 653364 95752 653370 95764
rect 665174 95752 665180 95764
rect 665232 95752 665238 95804
rect 645118 95616 645124 95668
rect 645176 95656 645182 95668
rect 652018 95656 652024 95668
rect 645176 95628 652024 95656
rect 645176 95616 645182 95628
rect 652018 95616 652024 95628
rect 652076 95616 652082 95668
rect 656158 95520 656164 95532
rect 654106 95492 656164 95520
rect 641346 95412 641352 95464
rect 641404 95412 641410 95464
rect 643462 95412 643468 95464
rect 643520 95452 643526 95464
rect 647878 95452 647884 95464
rect 643520 95424 647884 95452
rect 643520 95412 643526 95424
rect 647878 95412 647884 95424
rect 647936 95412 647942 95464
rect 641364 95316 641392 95412
rect 648062 95344 648068 95396
rect 648120 95384 648126 95396
rect 654106 95384 654134 95492
rect 656158 95480 656164 95492
rect 656216 95480 656222 95532
rect 648120 95356 654134 95384
rect 648120 95344 648126 95356
rect 647694 95316 647700 95328
rect 641364 95288 647700 95316
rect 647694 95276 647700 95288
rect 647752 95276 647758 95328
rect 578326 95140 578332 95192
rect 578384 95180 578390 95192
rect 584582 95180 584588 95192
rect 578384 95152 584588 95180
rect 578384 95140 578390 95152
rect 584582 95140 584588 95152
rect 584640 95140 584646 95192
rect 620922 95140 620928 95192
rect 620980 95180 620986 95192
rect 625430 95180 625436 95192
rect 620980 95152 625436 95180
rect 620980 95140 620986 95152
rect 625430 95140 625436 95152
rect 625488 95140 625494 95192
rect 647050 95140 647056 95192
rect 647108 95180 647114 95192
rect 650270 95180 650276 95192
rect 647108 95152 650276 95180
rect 647108 95140 647114 95152
rect 650270 95140 650276 95152
rect 650328 95140 650334 95192
rect 616506 94936 616512 94988
rect 616564 94976 616570 94988
rect 624970 94976 624976 94988
rect 616564 94948 624976 94976
rect 616564 94936 616570 94948
rect 624970 94936 624976 94948
rect 625028 94936 625034 94988
rect 607674 94460 607680 94512
rect 607732 94500 607738 94512
rect 620646 94500 620652 94512
rect 607732 94472 620652 94500
rect 607732 94460 607738 94472
rect 620646 94460 620652 94472
rect 620704 94460 620710 94512
rect 619542 93780 619548 93832
rect 619600 93820 619606 93832
rect 626258 93820 626264 93832
rect 619600 93792 626264 93820
rect 619600 93780 619606 93792
rect 626258 93780 626264 93792
rect 626316 93780 626322 93832
rect 647510 93712 647516 93764
rect 647568 93752 647574 93764
rect 648246 93752 648252 93764
rect 647568 93724 648252 93752
rect 647568 93712 647574 93724
rect 648246 93712 648252 93724
rect 648304 93712 648310 93764
rect 651282 93576 651288 93628
rect 651340 93616 651346 93628
rect 654686 93616 654692 93628
rect 651340 93588 654692 93616
rect 651340 93576 651346 93588
rect 654686 93576 654692 93588
rect 654744 93576 654750 93628
rect 579246 93372 579252 93424
rect 579304 93412 579310 93424
rect 586146 93412 586152 93424
rect 579304 93384 586152 93412
rect 579304 93372 579310 93384
rect 586146 93372 586152 93384
rect 586204 93372 586210 93424
rect 609698 93100 609704 93152
rect 609756 93140 609762 93152
rect 618622 93140 618628 93152
rect 609756 93112 618628 93140
rect 609756 93100 609762 93112
rect 618622 93100 618628 93112
rect 618680 93100 618686 93152
rect 617978 92420 617984 92472
rect 618036 92460 618042 92472
rect 626442 92460 626448 92472
rect 618036 92432 626448 92460
rect 618036 92420 618042 92432
rect 626442 92420 626448 92432
rect 626500 92420 626506 92472
rect 647694 92420 647700 92472
rect 647752 92460 647758 92472
rect 655422 92460 655428 92472
rect 647752 92432 655428 92460
rect 647752 92420 647758 92432
rect 655422 92420 655428 92432
rect 655480 92420 655486 92472
rect 606938 91740 606944 91792
rect 606996 91780 607002 91792
rect 622394 91780 622400 91792
rect 606996 91752 622400 91780
rect 606996 91740 607002 91752
rect 622394 91740 622400 91752
rect 622452 91740 622458 91792
rect 578602 91128 578608 91180
rect 578660 91168 578666 91180
rect 585778 91168 585784 91180
rect 578660 91140 585784 91168
rect 578660 91128 578666 91140
rect 585778 91128 585784 91140
rect 585836 91128 585842 91180
rect 618162 91128 618168 91180
rect 618220 91168 618226 91180
rect 618220 91140 618392 91168
rect 618220 91128 618226 91140
rect 611262 90992 611268 91044
rect 611320 91032 611326 91044
rect 618162 91032 618168 91044
rect 611320 91004 618168 91032
rect 611320 90992 611326 91004
rect 618162 90992 618168 91004
rect 618220 90992 618226 91044
rect 618364 91032 618392 91140
rect 626442 91032 626448 91044
rect 618364 91004 626448 91032
rect 626442 90992 626448 91004
rect 626500 90992 626506 91044
rect 648614 90788 648620 90840
rect 648672 90828 648678 90840
rect 655422 90828 655428 90840
rect 648672 90800 655428 90828
rect 648672 90788 648678 90800
rect 655422 90788 655428 90800
rect 655480 90788 655486 90840
rect 620646 89632 620652 89684
rect 620704 89672 620710 89684
rect 625430 89672 625436 89684
rect 620704 89644 625436 89672
rect 620704 89632 620710 89644
rect 625430 89632 625436 89644
rect 625488 89632 625494 89684
rect 649718 88748 649724 88800
rect 649776 88788 649782 88800
rect 658550 88788 658556 88800
rect 649776 88760 658556 88788
rect 649776 88748 649782 88760
rect 658550 88748 658556 88760
rect 658608 88748 658614 88800
rect 662322 88748 662328 88800
rect 662380 88788 662386 88800
rect 664162 88788 664168 88800
rect 662380 88760 664168 88788
rect 662380 88748 662386 88760
rect 664162 88748 664168 88760
rect 664220 88748 664226 88800
rect 656158 88612 656164 88664
rect 656216 88652 656222 88664
rect 657446 88652 657452 88664
rect 656216 88624 657452 88652
rect 656216 88612 656222 88624
rect 657446 88612 657452 88624
rect 657504 88612 657510 88664
rect 579246 88272 579252 88324
rect 579304 88312 579310 88324
rect 589918 88312 589924 88324
rect 579304 88284 589924 88312
rect 579304 88272 579310 88284
rect 589918 88272 589924 88284
rect 589976 88272 589982 88324
rect 622394 88272 622400 88324
rect 622452 88312 622458 88324
rect 626442 88312 626448 88324
rect 622452 88284 626448 88312
rect 622452 88272 622458 88284
rect 626442 88272 626448 88284
rect 626500 88272 626506 88324
rect 655238 88272 655244 88324
rect 655296 88312 655302 88324
rect 658458 88312 658464 88324
rect 655296 88284 658464 88312
rect 655296 88272 655302 88284
rect 658458 88272 658464 88284
rect 658516 88272 658522 88324
rect 618162 88136 618168 88188
rect 618220 88176 618226 88188
rect 626258 88176 626264 88188
rect 618220 88148 626264 88176
rect 618220 88136 618226 88148
rect 626258 88136 626264 88148
rect 626316 88136 626322 88188
rect 648430 86980 648436 87032
rect 648488 87020 648494 87032
rect 662506 87020 662512 87032
rect 648488 86992 662512 87020
rect 648488 86980 648494 86992
rect 662506 86980 662512 86992
rect 662564 86980 662570 87032
rect 578326 86912 578332 86964
rect 578384 86952 578390 86964
rect 580442 86952 580448 86964
rect 578384 86924 580448 86952
rect 578384 86912 578390 86924
rect 580442 86912 580448 86924
rect 580500 86912 580506 86964
rect 656710 86844 656716 86896
rect 656768 86884 656774 86896
rect 659562 86884 659568 86896
rect 656768 86856 659568 86884
rect 656768 86844 656774 86856
rect 659562 86844 659568 86856
rect 659620 86844 659626 86896
rect 652018 86708 652024 86760
rect 652076 86748 652082 86760
rect 660114 86748 660120 86760
rect 652076 86720 660120 86748
rect 652076 86708 652082 86720
rect 660114 86708 660120 86720
rect 660172 86708 660178 86760
rect 647878 86572 647884 86624
rect 647936 86612 647942 86624
rect 661402 86612 661408 86624
rect 647936 86584 661408 86612
rect 647936 86572 647942 86584
rect 661402 86572 661408 86584
rect 661460 86572 661466 86624
rect 652202 86436 652208 86488
rect 652260 86476 652266 86488
rect 657170 86476 657176 86488
rect 652260 86448 657176 86476
rect 652260 86436 652266 86448
rect 657170 86436 657176 86448
rect 657228 86436 657234 86488
rect 621658 86300 621664 86352
rect 621716 86340 621722 86352
rect 626442 86340 626448 86352
rect 621716 86312 626448 86340
rect 621716 86300 621722 86312
rect 626442 86300 626448 86312
rect 626500 86300 626506 86352
rect 656342 86300 656348 86352
rect 656400 86340 656406 86352
rect 660666 86340 660672 86352
rect 656400 86312 660672 86340
rect 656400 86300 656406 86312
rect 660666 86300 660672 86312
rect 660724 86300 660730 86352
rect 609882 85484 609888 85536
rect 609940 85524 609946 85536
rect 626442 85524 626448 85536
rect 609940 85496 626448 85524
rect 609940 85484 609946 85496
rect 626442 85484 626448 85496
rect 626500 85484 626506 85536
rect 618622 85348 618628 85400
rect 618680 85388 618686 85400
rect 625246 85388 625252 85400
rect 618680 85360 625252 85388
rect 618680 85348 618686 85360
rect 625246 85348 625252 85360
rect 625304 85348 625310 85400
rect 608502 84124 608508 84176
rect 608560 84164 608566 84176
rect 626442 84164 626448 84176
rect 608560 84136 626448 84164
rect 608560 84124 608566 84136
rect 626442 84124 626448 84136
rect 626500 84124 626506 84176
rect 579246 83988 579252 84040
rect 579304 84028 579310 84040
rect 581638 84028 581644 84040
rect 579304 84000 581644 84028
rect 579304 83988 579310 84000
rect 581638 83988 581644 84000
rect 581696 83988 581702 84040
rect 578878 82764 578884 82816
rect 578936 82804 578942 82816
rect 583018 82804 583024 82816
rect 578936 82776 583024 82804
rect 578936 82764 578942 82776
rect 583018 82764 583024 82776
rect 583076 82764 583082 82816
rect 579246 82084 579252 82136
rect 579304 82124 579310 82136
rect 587158 82124 587164 82136
rect 579304 82096 587164 82124
rect 579304 82084 579310 82096
rect 587158 82084 587164 82096
rect 587216 82084 587222 82136
rect 628742 81064 628748 81116
rect 628800 81104 628806 81116
rect 642450 81104 642456 81116
rect 628800 81076 642456 81104
rect 628800 81064 628806 81076
rect 642450 81064 642456 81076
rect 642508 81064 642514 81116
rect 615402 80928 615408 80980
rect 615460 80968 615466 80980
rect 646314 80968 646320 80980
rect 615460 80940 646320 80968
rect 615460 80928 615466 80940
rect 646314 80928 646320 80940
rect 646372 80928 646378 80980
rect 613838 80792 613844 80844
rect 613896 80832 613902 80844
rect 647326 80832 647332 80844
rect 613896 80804 647332 80832
rect 613896 80792 613902 80804
rect 647326 80792 647332 80804
rect 647384 80792 647390 80844
rect 595438 80656 595444 80708
rect 595496 80696 595502 80708
rect 636746 80696 636752 80708
rect 595496 80668 636752 80696
rect 595496 80656 595502 80668
rect 636746 80656 636752 80668
rect 636804 80656 636810 80708
rect 629202 79976 629208 80028
rect 629260 80016 629266 80028
rect 633434 80016 633440 80028
rect 629260 79988 633440 80016
rect 629260 79976 629266 79988
rect 633434 79976 633440 79988
rect 633492 79976 633498 80028
rect 614022 79432 614028 79484
rect 614080 79472 614086 79484
rect 646038 79472 646044 79484
rect 614080 79444 646044 79472
rect 614080 79432 614086 79444
rect 646038 79432 646044 79444
rect 646096 79432 646102 79484
rect 583018 79296 583024 79348
rect 583076 79336 583082 79348
rect 600314 79336 600320 79348
rect 583076 79308 600320 79336
rect 583076 79296 583082 79308
rect 600314 79296 600320 79308
rect 600372 79296 600378 79348
rect 612642 79296 612648 79348
rect 612700 79336 612706 79348
rect 648614 79336 648620 79348
rect 612700 79308 648620 79336
rect 612700 79296 612706 79308
rect 648614 79296 648620 79308
rect 648672 79296 648678 79348
rect 578234 78072 578240 78124
rect 578292 78112 578298 78124
rect 580258 78112 580264 78124
rect 578292 78084 580264 78112
rect 578292 78072 578298 78084
rect 580258 78072 580264 78084
rect 580316 78072 580322 78124
rect 633434 78072 633440 78124
rect 633492 78112 633498 78124
rect 645302 78112 645308 78124
rect 633492 78084 645308 78112
rect 633492 78072 633498 78084
rect 645302 78072 645308 78084
rect 645360 78072 645366 78124
rect 631042 77936 631048 77988
rect 631100 77976 631106 77988
rect 643094 77976 643100 77988
rect 631100 77948 643100 77976
rect 631100 77936 631106 77948
rect 643094 77936 643100 77948
rect 643152 77936 643158 77988
rect 628466 77596 628472 77648
rect 628524 77636 628530 77648
rect 632790 77636 632796 77648
rect 628524 77608 632796 77636
rect 628524 77596 628530 77608
rect 632790 77596 632796 77608
rect 632848 77596 632854 77648
rect 628466 77432 628472 77444
rect 625126 77404 628472 77432
rect 624418 77256 624424 77308
rect 624476 77296 624482 77308
rect 625126 77296 625154 77404
rect 628466 77392 628472 77404
rect 628524 77392 628530 77444
rect 624476 77268 625154 77296
rect 624476 77256 624482 77268
rect 625798 77256 625804 77308
rect 625856 77296 625862 77308
rect 631042 77296 631048 77308
rect 625856 77268 631048 77296
rect 625856 77256 625862 77268
rect 631042 77256 631048 77268
rect 631100 77256 631106 77308
rect 620278 76780 620284 76832
rect 620336 76820 620342 76832
rect 648982 76820 648988 76832
rect 620336 76792 648988 76820
rect 620336 76780 620342 76792
rect 648982 76780 648988 76792
rect 649040 76780 649046 76832
rect 611998 76644 612004 76696
rect 612056 76684 612062 76696
rect 662414 76684 662420 76696
rect 612056 76656 662420 76684
rect 612056 76644 612062 76656
rect 662414 76644 662420 76656
rect 662472 76644 662478 76696
rect 587158 76508 587164 76560
rect 587216 76548 587222 76560
rect 668210 76548 668216 76560
rect 587216 76520 668216 76548
rect 587216 76508 587222 76520
rect 668210 76508 668216 76520
rect 668268 76508 668274 76560
rect 616782 75420 616788 75472
rect 616840 75460 616846 75472
rect 646682 75460 646688 75472
rect 616840 75432 646688 75460
rect 616840 75420 616846 75432
rect 646682 75420 646688 75432
rect 646740 75420 646746 75472
rect 607122 75284 607128 75336
rect 607180 75324 607186 75336
rect 646498 75324 646504 75336
rect 607180 75296 646504 75324
rect 607180 75284 607186 75296
rect 646498 75284 646504 75296
rect 646556 75284 646562 75336
rect 578878 75148 578884 75200
rect 578936 75188 578942 75200
rect 666554 75188 666560 75200
rect 578936 75160 666560 75188
rect 578936 75148 578942 75160
rect 666554 75148 666560 75160
rect 666612 75148 666618 75200
rect 579522 73108 579528 73160
rect 579580 73148 579586 73160
rect 588538 73148 588544 73160
rect 579580 73120 588544 73148
rect 579580 73108 579586 73120
rect 588538 73108 588544 73120
rect 588596 73108 588602 73160
rect 578510 71544 578516 71596
rect 578568 71584 578574 71596
rect 584398 71584 584404 71596
rect 578568 71556 584404 71584
rect 578568 71544 578574 71556
rect 584398 71544 584404 71556
rect 584456 71544 584462 71596
rect 579522 66852 579528 66904
rect 579580 66892 579586 66904
rect 625982 66892 625988 66904
rect 579580 66864 625988 66892
rect 579580 66852 579586 66864
rect 625982 66852 625988 66864
rect 626040 66852 626046 66904
rect 579522 64812 579528 64864
rect 579580 64852 579586 64864
rect 592678 64852 592684 64864
rect 579580 64824 592684 64852
rect 579580 64812 579586 64824
rect 592678 64812 592684 64824
rect 592736 64812 592742 64864
rect 579522 62024 579528 62076
rect 579580 62064 579586 62076
rect 587158 62064 587164 62076
rect 579580 62036 587164 62064
rect 579580 62024 579586 62036
rect 587158 62024 587164 62036
rect 587216 62024 587222 62076
rect 578326 59984 578332 60036
rect 578384 60024 578390 60036
rect 624418 60024 624424 60036
rect 578384 59996 624424 60024
rect 578384 59984 578390 59996
rect 624418 59984 624424 59996
rect 624476 59984 624482 60036
rect 576118 58760 576124 58812
rect 576176 58800 576182 58812
rect 603074 58800 603080 58812
rect 576176 58772 603080 58800
rect 576176 58760 576182 58772
rect 603074 58760 603080 58772
rect 603132 58760 603138 58812
rect 577498 58624 577504 58676
rect 577556 58664 577562 58676
rect 604454 58664 604460 58676
rect 577556 58636 604460 58664
rect 577556 58624 577562 58636
rect 604454 58624 604460 58636
rect 604512 58624 604518 58676
rect 579522 57876 579528 57928
rect 579580 57916 579586 57928
rect 594058 57916 594064 57928
rect 579580 57888 594064 57916
rect 579580 57876 579586 57888
rect 594058 57876 594064 57888
rect 594116 57876 594122 57928
rect 574922 57196 574928 57248
rect 574980 57236 574986 57248
rect 600498 57236 600504 57248
rect 574980 57208 600504 57236
rect 574980 57196 574986 57208
rect 600498 57196 600504 57208
rect 600556 57196 600562 57248
rect 574738 55972 574744 56024
rect 574796 56012 574802 56024
rect 598934 56012 598940 56024
rect 574796 55984 598940 56012
rect 574796 55972 574802 55984
rect 598934 55972 598940 55984
rect 598992 55972 598998 56024
rect 574462 55836 574468 55888
rect 574520 55876 574526 55888
rect 601878 55876 601884 55888
rect 574520 55848 601884 55876
rect 574520 55836 574526 55848
rect 601878 55836 601884 55848
rect 601936 55836 601942 55888
rect 471946 55236 473354 55264
rect 471946 55196 471974 55236
rect 464908 55168 471974 55196
rect 473326 55196 473354 55236
rect 596450 55196 596456 55208
rect 473326 55168 596456 55196
rect 464908 54652 464936 55168
rect 596450 55156 596456 55168
rect 596508 55156 596514 55208
rect 597830 55060 597836 55072
rect 463988 54624 464936 54652
rect 465046 55032 597836 55060
rect 463988 53836 464016 54624
rect 465046 54380 465074 55032
rect 597830 55020 597836 55032
rect 597888 55020 597894 55072
rect 597646 54924 597652 54936
rect 463896 53808 464016 53836
rect 464540 54352 465074 54380
rect 473326 54896 597652 54924
rect 463896 53644 463924 53808
rect 464540 53644 464568 54352
rect 473326 54312 473354 54896
rect 597646 54884 597652 54896
rect 597704 54884 597710 54936
rect 599118 54788 599124 54800
rect 474706 54760 599124 54788
rect 474706 54720 474734 54760
rect 599118 54748 599124 54760
rect 599176 54748 599182 54800
rect 465184 54284 473354 54312
rect 474200 54692 474734 54720
rect 465184 53768 465212 54284
rect 474200 54176 474228 54692
rect 623038 54652 623044 54664
rect 477466 54624 623044 54652
rect 477466 54584 477494 54624
rect 623038 54612 623044 54624
rect 623096 54612 623102 54664
rect 464678 53740 465212 53768
rect 473326 54148 474228 54176
rect 474292 54556 477494 54584
rect 463878 53592 463884 53644
rect 463936 53592 463942 53644
rect 464522 53592 464528 53644
rect 464580 53592 464586 53644
rect 463602 53456 463608 53508
rect 463660 53496 463666 53508
rect 464678 53496 464706 53740
rect 464798 53592 464804 53644
rect 464856 53632 464862 53644
rect 473326 53632 473354 54148
rect 474292 53644 474320 54556
rect 625798 54516 625804 54528
rect 478846 54488 625804 54516
rect 478846 54448 478874 54488
rect 625798 54476 625804 54488
rect 625856 54476 625862 54528
rect 474476 54420 478874 54448
rect 474476 53644 474504 54420
rect 596174 54380 596180 54392
rect 479812 54352 596180 54380
rect 479812 54312 479840 54352
rect 596174 54340 596180 54352
rect 596232 54340 596238 54392
rect 474936 54284 479840 54312
rect 464856 53604 473354 53632
rect 464856 53592 464862 53604
rect 474274 53592 474280 53644
rect 474332 53592 474338 53644
rect 474458 53592 474464 53644
rect 474516 53592 474522 53644
rect 463660 53468 464706 53496
rect 463660 53456 463666 53468
rect 464982 53456 464988 53508
rect 465040 53496 465046 53508
rect 474936 53496 474964 54284
rect 583018 54244 583024 54256
rect 479904 54216 583024 54244
rect 479904 54176 479932 54216
rect 583018 54204 583024 54216
rect 583076 54204 583082 54256
rect 479812 54148 479932 54176
rect 479812 53904 479840 54148
rect 580442 54108 580448 54120
rect 479996 54080 580448 54108
rect 479996 54040 480024 54080
rect 580442 54068 580448 54080
rect 580500 54068 580506 54120
rect 475212 53876 479840 53904
rect 479904 54012 480024 54040
rect 475212 53644 475240 53876
rect 479904 53768 479932 54012
rect 574738 53972 574744 53984
rect 475396 53740 479932 53768
rect 480088 53944 574744 53972
rect 475396 53644 475424 53740
rect 480088 53644 480116 53944
rect 574738 53932 574744 53944
rect 574796 53932 574802 53984
rect 574922 53836 574928 53848
rect 480226 53808 574928 53836
rect 475194 53592 475200 53644
rect 475252 53592 475258 53644
rect 475378 53592 475384 53644
rect 475436 53592 475442 53644
rect 480070 53592 480076 53644
rect 480128 53592 480134 53644
rect 465040 53468 474964 53496
rect 465040 53456 465046 53468
rect 462222 53320 462228 53372
rect 462280 53360 462286 53372
rect 480226 53360 480254 53808
rect 574922 53796 574928 53808
rect 574980 53796 574986 53848
rect 462280 53332 480254 53360
rect 462280 53320 462286 53332
rect 48958 53184 48964 53236
rect 49016 53224 49022 53236
rect 128998 53224 129004 53236
rect 49016 53196 129004 53224
rect 49016 53184 49022 53196
rect 128998 53184 129004 53196
rect 129056 53184 129062 53236
rect 463142 53184 463148 53236
rect 463200 53224 463206 53236
rect 468294 53224 468300 53236
rect 463200 53196 468300 53224
rect 463200 53184 463206 53196
rect 468294 53184 468300 53196
rect 468352 53184 468358 53236
rect 312354 53116 312360 53168
rect 312412 53156 312418 53168
rect 313734 53156 313740 53168
rect 312412 53128 313740 53156
rect 312412 53116 312418 53128
rect 313734 53116 313740 53128
rect 313792 53116 313798 53168
rect 316310 53116 316316 53168
rect 316368 53156 316374 53168
rect 317690 53156 317696 53168
rect 316368 53128 317696 53156
rect 316368 53116 316374 53128
rect 317690 53116 317696 53128
rect 317748 53116 317754 53168
rect 46198 53048 46204 53100
rect 46256 53088 46262 53100
rect 130378 53088 130384 53100
rect 46256 53060 130384 53088
rect 46256 53048 46262 53060
rect 130378 53048 130384 53060
rect 130436 53048 130442 53100
rect 461302 53048 461308 53100
rect 461360 53088 461366 53100
rect 480070 53088 480076 53100
rect 461360 53060 480076 53088
rect 461360 53048 461366 53060
rect 480070 53048 480076 53060
rect 480128 53048 480134 53100
rect 460382 52912 460388 52964
rect 460440 52952 460446 52964
rect 474458 52952 474464 52964
rect 460440 52924 474464 52952
rect 460440 52912 460446 52924
rect 474458 52912 474464 52924
rect 474516 52912 474522 52964
rect 459140 52776 459146 52828
rect 459198 52816 459204 52828
rect 464798 52816 464804 52828
rect 459198 52788 464804 52816
rect 459198 52776 459204 52788
rect 464798 52776 464804 52788
rect 464856 52776 464862 52828
rect 465120 52776 465126 52828
rect 465178 52816 465184 52828
rect 475378 52816 475384 52828
rect 465178 52788 475384 52816
rect 465178 52776 465184 52788
rect 475378 52776 475384 52788
rect 475436 52776 475442 52828
rect 465902 52640 465908 52692
rect 465960 52680 465966 52692
rect 474274 52680 474280 52692
rect 465960 52652 474280 52680
rect 465960 52640 465966 52652
rect 474274 52640 474280 52652
rect 474332 52640 474338 52692
rect 51718 51960 51724 52012
rect 51776 52000 51782 52012
rect 129366 52000 129372 52012
rect 51776 51972 129372 52000
rect 51776 51960 51782 51972
rect 129366 51960 129372 51972
rect 129424 51960 129430 52012
rect 50522 51824 50528 51876
rect 50580 51864 50586 51876
rect 130562 51864 130568 51876
rect 50580 51836 130568 51864
rect 50580 51824 50586 51836
rect 130562 51824 130568 51836
rect 130620 51824 130626 51876
rect 47578 51688 47584 51740
rect 47636 51728 47642 51740
rect 129182 51728 129188 51740
rect 47636 51700 129188 51728
rect 47636 51688 47642 51700
rect 129182 51688 129188 51700
rect 129240 51688 129246 51740
rect 145374 51688 145380 51740
rect 145432 51728 145438 51740
rect 306006 51728 306012 51740
rect 145432 51700 306012 51728
rect 145432 51688 145438 51700
rect 306006 51688 306012 51700
rect 306064 51688 306070 51740
rect 318334 50464 318340 50516
rect 318392 50504 318398 50516
rect 458358 50504 458364 50516
rect 318392 50476 458364 50504
rect 318392 50464 318398 50476
rect 458358 50464 458364 50476
rect 458416 50464 458422 50516
rect 45462 50328 45468 50380
rect 45520 50368 45526 50380
rect 129642 50368 129648 50380
rect 45520 50340 129648 50368
rect 45520 50328 45526 50340
rect 129642 50328 129648 50340
rect 129700 50328 129706 50380
rect 314010 50328 314016 50380
rect 314068 50368 314074 50380
rect 458174 50368 458180 50380
rect 314068 50340 458180 50368
rect 314068 50328 314074 50340
rect 458174 50328 458180 50340
rect 458232 50328 458238 50380
rect 522942 50328 522948 50380
rect 523000 50368 523006 50380
rect 544010 50368 544016 50380
rect 523000 50340 544016 50368
rect 523000 50328 523006 50340
rect 544010 50328 544016 50340
rect 544068 50328 544074 50380
rect 49142 48968 49148 49020
rect 49200 49008 49206 49020
rect 131022 49008 131028 49020
rect 49200 48980 131028 49008
rect 49200 48968 49206 48980
rect 131022 48968 131028 48980
rect 131080 48968 131086 49020
rect 129182 47812 129188 47864
rect 129240 47852 129246 47864
rect 131574 47852 131580 47864
rect 129240 47824 131580 47852
rect 129240 47812 129246 47824
rect 131574 47812 131580 47824
rect 131632 47812 131638 47864
rect 625982 46452 625988 46504
rect 626040 46492 626046 46504
rect 661770 46492 661776 46504
rect 626040 46464 661776 46492
rect 626040 46452 626046 46464
rect 661770 46452 661776 46464
rect 661828 46452 661834 46504
rect 129642 46044 129648 46096
rect 129700 46084 129706 46096
rect 132034 46084 132040 46096
rect 129700 46056 132040 46084
rect 129700 46044 129706 46056
rect 132034 46044 132040 46056
rect 132092 46044 132098 46096
rect 130378 45500 130384 45552
rect 130436 45540 130442 45552
rect 132218 45540 132224 45552
rect 130436 45512 132224 45540
rect 130436 45500 130442 45512
rect 132218 45500 132224 45512
rect 132276 45500 132282 45552
rect 131298 45364 131304 45416
rect 131356 45404 131362 45416
rect 132954 45404 132960 45416
rect 131356 45376 132960 45404
rect 131356 45364 131362 45376
rect 132954 45364 132960 45376
rect 133012 45364 133018 45416
rect 129366 45296 129372 45348
rect 129424 45336 129430 45348
rect 130930 45336 130936 45348
rect 129424 45308 130936 45336
rect 129424 45296 129430 45308
rect 130930 45296 130936 45308
rect 130988 45296 130994 45348
rect 43806 45160 43812 45212
rect 43864 45200 43870 45212
rect 43864 45172 122834 45200
rect 43864 45160 43870 45172
rect 122806 44996 122834 45172
rect 130930 45064 130936 45116
rect 130988 45104 130994 45116
rect 130988 45076 131192 45104
rect 130988 45064 130994 45076
rect 129366 44996 129372 45008
rect 122806 44968 129372 44996
rect 129366 44956 129372 44968
rect 129424 44956 129430 45008
rect 131178 44992 131330 45020
rect 131178 44928 131206 44992
rect 131500 44928 131606 44936
rect 131040 44900 131206 44928
rect 131408 44908 131606 44928
rect 131408 44900 131528 44908
rect 128354 44820 128360 44872
rect 128412 44860 128418 44872
rect 131040 44860 131068 44900
rect 131408 44860 131436 44900
rect 128412 44832 131068 44860
rect 131362 44832 131436 44860
rect 128412 44820 128418 44832
rect 131362 44736 131390 44832
rect 131362 44696 131396 44736
rect 131390 44684 131396 44696
rect 131448 44684 131454 44736
rect 128998 44616 129004 44668
rect 129056 44656 129062 44668
rect 131776 44656 131804 44838
rect 129056 44628 131252 44656
rect 129056 44616 129062 44628
rect 131224 44588 131252 44628
rect 131684 44628 131804 44656
rect 131868 44740 131974 44768
rect 131684 44588 131712 44628
rect 131224 44560 131712 44588
rect 131868 44516 131896 44740
rect 132144 44516 132172 44670
rect 131776 44488 131896 44516
rect 131960 44488 132172 44516
rect 50338 44412 50344 44464
rect 50396 44452 50402 44464
rect 128354 44452 128360 44464
rect 50396 44424 128360 44452
rect 50396 44412 50402 44424
rect 128354 44412 128360 44424
rect 128412 44412 128418 44464
rect 131776 44452 131804 44488
rect 131270 44424 131804 44452
rect 43622 44276 43628 44328
rect 43680 44316 43686 44328
rect 131270 44316 131298 44424
rect 131960 44384 131988 44488
rect 132374 44384 132402 44586
rect 131868 44356 131988 44384
rect 132052 44356 132402 44384
rect 132466 44488 132526 44516
rect 43680 44288 131298 44316
rect 43680 44276 43686 44288
rect 131574 44276 131580 44328
rect 131632 44316 131638 44328
rect 131868 44316 131896 44356
rect 131632 44288 131896 44316
rect 131632 44276 131638 44288
rect 132052 44260 132080 44356
rect 132034 44208 132040 44260
rect 132092 44208 132098 44260
rect 132218 44208 132224 44260
rect 132276 44248 132282 44260
rect 132466 44248 132494 44488
rect 132586 44364 132592 44416
rect 132644 44404 132650 44416
rect 132644 44376 132756 44404
rect 132644 44364 132650 44376
rect 132954 44252 132960 44304
rect 133012 44252 133018 44304
rect 132276 44220 132494 44248
rect 132276 44208 132282 44220
rect 43438 44140 43444 44192
rect 43496 44180 43502 44192
rect 131390 44180 131396 44192
rect 43496 44152 131396 44180
rect 43496 44140 43502 44152
rect 131390 44140 131396 44152
rect 131448 44140 131454 44192
rect 129366 44004 129372 44056
rect 129424 44044 129430 44056
rect 133156 44044 133184 44166
rect 129424 44016 133184 44044
rect 129424 44004 129430 44016
rect 440234 43800 440240 43852
rect 440292 43840 440298 43852
rect 441062 43840 441068 43852
rect 440292 43812 441068 43840
rect 440292 43800 440298 43812
rect 441062 43800 441068 43812
rect 441120 43800 441126 43852
rect 410886 42848 410892 42900
rect 410944 42888 410950 42900
rect 415578 42888 415584 42900
rect 410944 42860 415584 42888
rect 410944 42848 410950 42860
rect 415578 42848 415584 42860
rect 415636 42848 415642 42900
rect 187326 42780 187332 42832
rect 187384 42820 187390 42832
rect 255866 42820 255872 42832
rect 187384 42792 255872 42820
rect 187384 42780 187390 42792
rect 255866 42780 255872 42792
rect 255924 42780 255930 42832
rect 310422 42712 310428 42764
rect 310480 42752 310486 42764
rect 364518 42752 364524 42764
rect 310480 42724 364524 42752
rect 310480 42712 310486 42724
rect 364518 42712 364524 42724
rect 364576 42712 364582 42764
rect 431218 42752 431224 42764
rect 364720 42724 431224 42752
rect 361758 42440 361764 42492
rect 361816 42480 361822 42492
rect 364720 42480 364748 42724
rect 431218 42712 431224 42724
rect 431276 42712 431282 42764
rect 441062 42712 441068 42764
rect 441120 42752 441126 42764
rect 449158 42752 449164 42764
rect 441120 42724 449164 42752
rect 441120 42712 441126 42724
rect 449158 42712 449164 42724
rect 449216 42712 449222 42764
rect 453574 42712 453580 42764
rect 453632 42752 453638 42764
rect 464338 42752 464344 42764
rect 453632 42724 464344 42752
rect 453632 42712 453638 42724
rect 464338 42712 464344 42724
rect 464396 42712 464402 42764
rect 364886 42576 364892 42628
rect 364944 42616 364950 42628
rect 427078 42616 427084 42628
rect 364944 42588 427084 42616
rect 364944 42576 364950 42588
rect 427078 42576 427084 42588
rect 427136 42576 427142 42628
rect 441246 42576 441252 42628
rect 441304 42616 441310 42628
rect 446398 42616 446404 42628
rect 441304 42588 446404 42616
rect 441304 42576 441310 42588
rect 446398 42576 446404 42588
rect 446456 42576 446462 42628
rect 454678 42576 454684 42628
rect 454736 42616 454742 42628
rect 462958 42616 462964 42628
rect 454736 42588 462964 42616
rect 454736 42576 454742 42588
rect 462958 42576 462964 42588
rect 463016 42576 463022 42628
rect 410886 42480 410892 42492
rect 361816 42452 364748 42480
rect 373966 42452 410892 42480
rect 361816 42440 361822 42452
rect 364518 42304 364524 42356
rect 364576 42344 364582 42356
rect 373966 42344 373994 42452
rect 410886 42440 410892 42452
rect 410944 42440 410950 42492
rect 429102 42480 429108 42492
rect 422266 42452 429108 42480
rect 364576 42316 373994 42344
rect 364576 42304 364582 42316
rect 415578 42304 415584 42356
rect 415636 42344 415642 42356
rect 422266 42344 422294 42452
rect 429102 42440 429108 42452
rect 429160 42440 429166 42492
rect 454494 42440 454500 42492
rect 454552 42480 454558 42492
rect 463694 42480 463700 42492
rect 454552 42452 463700 42480
rect 454552 42440 454558 42452
rect 463694 42440 463700 42452
rect 463752 42440 463758 42492
rect 415636 42316 422294 42344
rect 415636 42304 415642 42316
rect 661402 42129 661408 42181
rect 661460 42129 661466 42181
rect 427078 41964 427084 42016
rect 427136 42004 427142 42016
rect 427136 41976 427814 42004
rect 427136 41964 427142 41976
rect 427786 41868 427814 41976
rect 431218 41964 431224 42016
rect 431276 42004 431282 42016
rect 441062 42004 441068 42016
rect 431276 41976 441068 42004
rect 431276 41964 431282 41976
rect 441062 41964 441068 41976
rect 441120 41964 441126 42016
rect 446398 41964 446404 42016
rect 446456 42004 446462 42016
rect 454494 42004 454500 42016
rect 446456 41976 454500 42004
rect 446456 41964 446462 41976
rect 454494 41964 454500 41976
rect 454552 41964 454558 42016
rect 441246 41868 441252 41880
rect 427786 41840 441252 41868
rect 441246 41828 441252 41840
rect 441304 41828 441310 41880
rect 454678 41868 454684 41880
rect 441586 41840 454684 41868
rect 429102 41692 429108 41744
rect 429160 41732 429166 41744
rect 441586 41732 441614 41840
rect 454678 41828 454684 41840
rect 454736 41828 454742 41880
rect 429160 41704 441614 41732
rect 429160 41692 429166 41704
rect 449158 41692 449164 41744
rect 449216 41732 449222 41744
rect 453574 41732 453580 41744
rect 449216 41704 453580 41732
rect 449216 41692 449222 41704
rect 453574 41692 453580 41704
rect 453632 41692 453638 41744
<< via1 >>
rect 652024 896996 652076 897048
rect 676036 897064 676088 897116
rect 654784 895772 654836 895824
rect 675852 895772 675904 895824
rect 672724 895636 672776 895688
rect 676036 895636 676088 895688
rect 672172 894412 672224 894464
rect 675852 894412 675904 894464
rect 673368 894276 673420 894328
rect 676036 894276 676088 894328
rect 671988 892984 672040 893036
rect 676036 892984 676088 893036
rect 670976 892848 671028 892900
rect 675852 892848 675904 892900
rect 676220 891488 676272 891540
rect 676864 891488 676916 891540
rect 674840 890740 674892 890792
rect 676036 890740 676088 890792
rect 676036 889992 676088 890044
rect 677048 889992 677100 890044
rect 674656 888904 674708 888956
rect 676036 888904 676088 888956
rect 675024 888768 675076 888820
rect 675852 888768 675904 888820
rect 674288 888496 674340 888548
rect 676036 888496 676088 888548
rect 673184 886864 673236 886916
rect 676036 886864 676088 886916
rect 671804 885640 671856 885692
rect 676036 885640 676088 885692
rect 675208 881016 675260 881068
rect 683304 881016 683356 881068
rect 653404 880472 653456 880524
rect 675576 880540 675628 880592
rect 675760 880404 675812 880456
rect 679624 880404 679676 880456
rect 675392 879316 675444 879368
rect 677048 879316 677100 879368
rect 674840 879180 674892 879232
rect 675300 879180 675352 879232
rect 674840 879044 674892 879096
rect 678244 879044 678296 879096
rect 676864 878500 676916 878552
rect 675484 876528 675536 876580
rect 674472 876188 674524 876240
rect 674840 876188 674892 876240
rect 674840 872856 674892 872908
rect 675392 872856 675444 872908
rect 674288 870272 674340 870324
rect 674932 870272 674984 870324
rect 657544 869388 657596 869440
rect 675208 869320 675260 869372
rect 675208 869116 675260 869168
rect 675024 868980 675076 869032
rect 651472 868844 651524 868896
rect 654784 868844 654836 868896
rect 654140 868028 654192 868080
rect 674840 868028 674892 868080
rect 651472 866600 651524 866652
rect 672724 866600 672776 866652
rect 651380 865172 651432 865224
rect 653404 865172 653456 865224
rect 651472 863812 651524 863864
rect 657544 863812 657596 863864
rect 651472 862452 651524 862504
rect 654140 862452 654192 862504
rect 35624 817096 35676 817148
rect 35808 817096 35860 817148
rect 44824 817096 44876 817148
rect 61384 816960 61436 817012
rect 35624 815736 35676 815788
rect 43444 815736 43496 815788
rect 35808 815600 35860 815652
rect 44180 815600 44232 815652
rect 35808 814376 35860 814428
rect 44364 814376 44416 814428
rect 35624 814240 35676 814292
rect 44548 814240 44600 814292
rect 41328 812812 41380 812864
rect 43260 812812 43312 812864
rect 41328 811452 41380 811504
rect 41788 811452 41840 811504
rect 31668 809344 31720 809396
rect 42432 809344 42484 809396
rect 41328 808664 41380 808716
rect 43076 808664 43128 808716
rect 43444 807916 43496 807968
rect 62764 807916 62816 807968
rect 41328 807440 41380 807492
rect 42892 807440 42944 807492
rect 41144 807304 41196 807356
rect 43444 807304 43496 807356
rect 41328 806080 41380 806132
rect 43812 806080 43864 806132
rect 41144 805944 41196 805996
rect 64144 805944 64196 805996
rect 30288 805196 30340 805248
rect 42708 805196 42760 805248
rect 32220 802408 32272 802460
rect 41788 802408 41840 802460
rect 33784 801184 33836 801236
rect 42616 801184 42668 801236
rect 31024 801048 31076 801100
rect 40500 801048 40552 801100
rect 43628 799076 43680 799128
rect 53104 799076 53156 799128
rect 45008 797648 45060 797700
rect 57244 797648 57296 797700
rect 42248 796832 42300 796884
rect 42616 796832 42668 796884
rect 42708 794724 42760 794776
rect 43444 794724 43496 794776
rect 653404 790780 653456 790832
rect 675392 790780 675444 790832
rect 53104 790712 53156 790764
rect 62212 790712 62264 790764
rect 42248 789692 42300 789744
rect 42248 789488 42300 789540
rect 670608 789352 670660 789404
rect 675116 789352 675168 789404
rect 57244 789148 57296 789200
rect 62120 789148 62172 789200
rect 42616 786632 42668 786684
rect 62120 786632 62172 786684
rect 44824 785136 44876 785188
rect 62120 785136 62172 785188
rect 674472 783844 674524 783896
rect 675116 783844 675168 783896
rect 674748 782620 674800 782672
rect 675208 782620 675260 782672
rect 655520 781056 655572 781108
rect 675208 781056 675260 781108
rect 655060 778336 655112 778388
rect 675208 778336 675260 778388
rect 651472 777588 651524 777640
rect 660304 777588 660356 777640
rect 674288 776976 674340 777028
rect 675300 776976 675352 777028
rect 651472 775548 651524 775600
rect 669964 775548 670016 775600
rect 670792 775548 670844 775600
rect 674840 775548 674892 775600
rect 651380 775276 651432 775328
rect 653404 775276 653456 775328
rect 35808 774188 35860 774240
rect 41696 774188 41748 774240
rect 42064 774188 42116 774240
rect 60004 774188 60056 774240
rect 651472 774120 651524 774172
rect 655520 774120 655572 774172
rect 651472 773780 651524 773832
rect 655060 773780 655112 773832
rect 35440 773372 35492 773424
rect 41512 773372 41564 773424
rect 35808 773100 35860 773152
rect 41696 773168 41748 773220
rect 42064 773168 42116 773220
rect 44180 773168 44232 773220
rect 35624 772964 35676 773016
rect 41696 773032 41748 773084
rect 42064 773032 42116 773084
rect 46204 773032 46256 773084
rect 35256 772828 35308 772880
rect 41696 772828 41748 772880
rect 42064 772828 42116 772880
rect 61384 772828 61436 772880
rect 35808 771808 35860 771860
rect 39488 771808 39540 771860
rect 42064 771604 42116 771656
rect 44548 771604 44600 771656
rect 35624 771536 35676 771588
rect 41696 771536 41748 771588
rect 35808 771400 35860 771452
rect 41696 771400 41748 771452
rect 42064 771400 42116 771452
rect 44364 771400 44416 771452
rect 35808 770448 35860 770500
rect 39120 770448 39172 770500
rect 35808 770176 35860 770228
rect 39856 770176 39908 770228
rect 35624 770040 35676 770092
rect 41696 770040 41748 770092
rect 42064 770040 42116 770092
rect 45376 770040 45428 770092
rect 35808 768952 35860 769004
rect 41696 768952 41748 769004
rect 35808 768816 35860 768868
rect 39764 768816 39816 768868
rect 35624 768680 35676 768732
rect 40040 768680 40092 768732
rect 35808 767320 35860 767372
rect 36544 767320 36596 767372
rect 35808 766096 35860 766148
rect 39580 766096 39632 766148
rect 35808 764804 35860 764856
rect 40132 764804 40184 764856
rect 35808 764532 35860 764584
rect 41696 764532 41748 764584
rect 42064 764532 42116 764584
rect 44180 764532 44232 764584
rect 35624 763376 35676 763428
rect 40500 763308 40552 763360
rect 42064 763308 42116 763360
rect 35808 763172 35860 763224
rect 41696 763172 41748 763224
rect 58624 763172 58676 763224
rect 35808 761880 35860 761932
rect 39948 761880 40000 761932
rect 35164 759772 35216 759824
rect 41696 759772 41748 759824
rect 32404 759636 32456 759688
rect 41604 759636 41656 759688
rect 33784 758276 33836 758328
rect 39856 758276 39908 758328
rect 44732 755488 44784 755540
rect 62764 755488 62816 755540
rect 42248 754264 42300 754316
rect 44732 754264 44784 754316
rect 42432 754128 42484 754180
rect 42800 754128 42852 754180
rect 42248 751476 42300 751528
rect 42248 751136 42300 751188
rect 61384 747124 61436 747176
rect 63040 747124 63092 747176
rect 45100 746512 45152 746564
rect 62120 746512 62172 746564
rect 671344 743996 671396 744048
rect 675392 743996 675444 744048
rect 42524 743860 42576 743912
rect 62120 743860 62172 743912
rect 46204 743724 46256 743776
rect 62120 743724 62172 743776
rect 671160 743180 671212 743232
rect 675300 743180 675352 743232
rect 672356 742772 672408 742824
rect 675484 742772 675536 742824
rect 60004 742364 60056 742416
rect 62120 742364 62172 742416
rect 669228 741072 669280 741124
rect 674840 741072 674892 741124
rect 674840 740596 674892 740648
rect 675392 740596 675444 740648
rect 652024 736176 652076 736228
rect 653404 736176 653456 736228
rect 657544 735564 657596 735616
rect 675208 735700 675260 735752
rect 654784 734136 654836 734188
rect 675116 734204 675168 734256
rect 668676 733864 668728 733916
rect 651472 733388 651524 733440
rect 668032 733388 668084 733440
rect 675300 733320 675352 733372
rect 651472 732776 651524 732828
rect 661684 732776 661736 732828
rect 651472 731416 651524 731468
rect 658924 731416 658976 731468
rect 651472 731280 651524 731332
rect 671344 731280 671396 731332
rect 41144 730192 41196 730244
rect 41696 730260 41748 730312
rect 42064 730260 42116 730312
rect 46204 730260 46256 730312
rect 43444 730124 43496 730176
rect 61384 730056 61436 730108
rect 651472 729988 651524 730040
rect 657544 729988 657596 730040
rect 43628 729308 43680 729360
rect 62764 729308 62816 729360
rect 41328 729036 41380 729088
rect 41696 729036 41748 729088
rect 42064 728628 42116 728680
rect 43076 728628 43128 728680
rect 651472 728492 651524 728544
rect 654784 728492 654836 728544
rect 671804 728288 671856 728340
rect 673184 728084 673236 728136
rect 674472 727880 674524 727932
rect 683488 727880 683540 727932
rect 674840 727472 674892 727524
rect 675116 727472 675168 727524
rect 675484 727472 675536 727524
rect 41052 727404 41104 727456
rect 41696 727404 41748 727456
rect 42064 727404 42116 727456
rect 45008 727404 45060 727456
rect 40776 727268 40828 727320
rect 41696 727268 41748 727320
rect 42064 727268 42116 727320
rect 45376 727268 45428 727320
rect 678244 727200 678296 727252
rect 674656 726656 674708 726708
rect 683304 726656 683356 726708
rect 674288 726520 674340 726572
rect 684132 726520 684184 726572
rect 41328 726180 41380 726232
rect 41696 726180 41748 726232
rect 41144 725908 41196 725960
rect 41604 725908 41656 725960
rect 42064 725908 42116 725960
rect 42708 725908 42760 725960
rect 673736 722168 673788 722220
rect 673920 722168 673972 722220
rect 675116 721692 675168 721744
rect 675300 721692 675352 721744
rect 675116 721216 675168 721268
rect 675300 721216 675352 721268
rect 675116 720808 675168 720860
rect 675300 720808 675352 720860
rect 675116 720468 675168 720520
rect 675300 720468 675352 720520
rect 42064 718972 42116 719024
rect 57244 718972 57296 719024
rect 42248 717204 42300 717256
rect 42708 717204 42760 717256
rect 653404 716252 653456 716304
rect 673828 716252 673880 716304
rect 672172 716116 672224 716168
rect 673368 716116 673420 716168
rect 669964 715708 670016 715760
rect 672816 715708 672868 715760
rect 35164 715640 35216 715692
rect 33784 715504 33836 715556
rect 40776 715504 40828 715556
rect 41512 715164 41564 715216
rect 660304 714960 660356 715012
rect 673828 714960 673880 715012
rect 670148 714824 670200 714876
rect 673368 714824 673420 714876
rect 671804 714008 671856 714060
rect 673828 714008 673880 714060
rect 670976 713668 671028 713720
rect 673828 713668 673880 713720
rect 671344 713192 671396 713244
rect 673828 713192 673880 713244
rect 671988 712852 672040 712904
rect 673828 712852 673880 712904
rect 671988 712376 672040 712428
rect 673828 712376 673880 712428
rect 43628 712104 43680 712156
rect 50344 712104 50396 712156
rect 669780 711628 669832 711680
rect 673828 711628 673880 711680
rect 670792 709996 670844 710048
rect 673828 709996 673880 710048
rect 670608 709588 670660 709640
rect 673828 709588 673880 709640
rect 43628 709316 43680 709368
rect 44456 709316 44508 709368
rect 674288 707956 674340 708008
rect 676036 707956 676088 708008
rect 674472 705576 674524 705628
rect 676036 705576 676088 705628
rect 42248 705508 42300 705560
rect 43444 705508 43496 705560
rect 668400 705508 668452 705560
rect 673368 705508 673420 705560
rect 674288 705304 674340 705356
rect 683120 705304 683172 705356
rect 50344 705100 50396 705152
rect 62120 705100 62172 705152
rect 674288 703876 674340 703928
rect 676036 703876 676088 703928
rect 667848 703808 667900 703860
rect 673184 703808 673236 703860
rect 44456 703740 44508 703792
rect 62120 703740 62172 703792
rect 42248 702176 42300 702228
rect 42248 701904 42300 701956
rect 654784 701156 654836 701208
rect 673184 701156 673236 701208
rect 42708 701088 42760 701140
rect 62212 701020 62264 701072
rect 666468 701020 666520 701072
rect 673000 701020 673052 701072
rect 46204 698164 46256 698216
rect 62120 698164 62172 698216
rect 656808 690004 656860 690056
rect 673184 690004 673236 690056
rect 652760 688780 652812 688832
rect 673184 688780 673236 688832
rect 651472 688644 651524 688696
rect 657544 688644 657596 688696
rect 42708 687284 42760 687336
rect 61384 687216 61436 687268
rect 651472 687216 651524 687268
rect 669964 687216 670016 687268
rect 675116 687216 675168 687268
rect 674472 687080 674524 687132
rect 651472 687012 651524 687064
rect 654784 687012 654836 687064
rect 43444 686468 43496 686520
rect 62764 686468 62816 686520
rect 651656 686468 651708 686520
rect 667204 686468 667256 686520
rect 41144 685992 41196 686044
rect 41696 685992 41748 686044
rect 42064 685992 42116 686044
rect 45376 685992 45428 686044
rect 668216 685924 668268 685976
rect 673644 685924 673696 685976
rect 40868 685856 40920 685908
rect 41696 685856 41748 685908
rect 42064 685856 42116 685908
rect 45192 685856 45244 685908
rect 651472 685516 651524 685568
rect 656808 685516 656860 685568
rect 41328 683408 41380 683460
rect 41696 683408 41748 683460
rect 41052 682932 41104 682984
rect 41696 682932 41748 682984
rect 674656 682388 674708 682440
rect 683212 682388 683264 682440
rect 41144 676200 41196 676252
rect 41696 676200 41748 676252
rect 42064 676200 42116 676252
rect 55864 676200 55916 676252
rect 31668 674092 31720 674144
rect 41512 674092 41564 674144
rect 35164 672732 35216 672784
rect 41696 672732 41748 672784
rect 42064 672664 42116 672716
rect 42524 672664 42576 672716
rect 33784 671304 33836 671356
rect 41696 671304 41748 671356
rect 673736 671304 673788 671356
rect 668032 671100 668084 671152
rect 673736 671100 673788 671152
rect 661684 670692 661736 670744
rect 670148 670148 670200 670200
rect 672172 670148 672224 670200
rect 670148 669672 670200 669724
rect 672172 669672 672224 669724
rect 658924 669468 658976 669520
rect 673552 669536 673604 669588
rect 42340 669332 42392 669384
rect 53104 669332 53156 669384
rect 671804 669332 671856 669384
rect 673552 669196 673604 669248
rect 669780 668652 669832 668704
rect 673552 668652 673604 668704
rect 671344 668244 671396 668296
rect 673552 668244 673604 668296
rect 60004 667904 60056 667956
rect 671436 667904 671488 667956
rect 673552 667904 673604 667956
rect 675208 667836 675260 667888
rect 676036 667836 676088 667888
rect 42248 667224 42300 667276
rect 671988 666884 672040 666936
rect 673552 666884 673604 666936
rect 671804 666680 671856 666732
rect 673552 666680 673604 666732
rect 671160 665660 671212 665712
rect 673552 665660 673604 665712
rect 42340 665388 42392 665440
rect 43628 665388 43680 665440
rect 671252 665320 671304 665372
rect 671804 665320 671856 665372
rect 669596 665184 669648 665236
rect 673552 665184 673604 665236
rect 670332 664300 670384 664352
rect 673552 664300 673604 664352
rect 674840 663892 674892 663944
rect 676220 663892 676272 663944
rect 42432 663824 42484 663876
rect 669228 663756 669280 663808
rect 673552 663756 673604 663808
rect 673552 663348 673604 663400
rect 673920 663348 673972 663400
rect 42432 663008 42484 663060
rect 674656 662940 674708 662992
rect 676220 662940 676272 662992
rect 668676 662736 668728 662788
rect 673920 662736 673972 662788
rect 671620 661512 671672 661564
rect 673920 661512 673972 661564
rect 669228 661104 669280 661156
rect 673920 661104 673972 661156
rect 53104 660900 53156 660952
rect 62120 660900 62172 660952
rect 42156 660492 42208 660544
rect 43076 660492 43128 660544
rect 668952 660084 669004 660136
rect 673920 660084 673972 660136
rect 674656 659812 674708 659864
rect 683120 659812 683172 659864
rect 60004 659540 60056 659592
rect 62120 659540 62172 659592
rect 42524 657364 42576 657416
rect 62120 657500 62172 657552
rect 653404 655528 653456 655580
rect 673920 655528 673972 655580
rect 44824 655460 44876 655512
rect 62120 655460 62172 655512
rect 667020 647300 667072 647352
rect 674012 647300 674064 647352
rect 655520 645872 655572 645924
rect 674012 645872 674064 645924
rect 35808 644444 35860 644496
rect 41696 644444 41748 644496
rect 42064 644444 42116 644496
rect 54484 644444 54536 644496
rect 35808 643492 35860 643544
rect 40500 643492 40552 643544
rect 35532 643220 35584 643272
rect 41696 643288 41748 643340
rect 42064 643288 42116 643340
rect 45376 643288 45428 643340
rect 35348 643084 35400 643136
rect 41696 643084 41748 643136
rect 42064 643084 42116 643136
rect 61384 643084 61436 643136
rect 655336 643084 655388 643136
rect 674012 643084 674064 643136
rect 38568 642472 38620 642524
rect 41696 642472 41748 642524
rect 42064 642336 42116 642388
rect 62948 642336 63000 642388
rect 651472 642336 651524 642388
rect 660304 642336 660356 642388
rect 35624 641996 35676 642048
rect 39488 641996 39540 642048
rect 35808 641724 35860 641776
rect 41696 641724 41748 641776
rect 42064 641724 42116 641776
rect 44640 641724 44692 641776
rect 35808 640772 35860 640824
rect 39580 640704 39632 640756
rect 35808 640432 35860 640484
rect 39948 640432 40000 640484
rect 35624 640296 35676 640348
rect 41696 640296 41748 640348
rect 42064 640296 42116 640348
rect 45376 640296 45428 640348
rect 651472 640296 651524 640348
rect 668584 640296 668636 640348
rect 651380 640092 651432 640144
rect 653404 640092 653456 640144
rect 35808 639072 35860 639124
rect 41696 639072 41748 639124
rect 35532 638936 35584 638988
rect 37924 638936 37976 638988
rect 651656 638868 651708 638920
rect 655336 638868 655388 638920
rect 651472 638732 651524 638784
rect 655520 638732 655572 638784
rect 35348 638188 35400 638240
rect 41696 638188 41748 638240
rect 35808 637576 35860 637628
rect 36544 637576 36596 637628
rect 672356 637372 672408 637424
rect 672816 637372 672868 637424
rect 35624 637168 35676 637220
rect 675484 636964 675536 637016
rect 683304 636964 683356 637016
rect 40408 636896 40460 636948
rect 674380 636828 674432 636880
rect 683948 636828 684000 636880
rect 674288 636692 674340 636744
rect 675484 636692 675536 636744
rect 35624 636488 35676 636540
rect 39856 636488 39908 636540
rect 35808 636216 35860 636268
rect 39028 636148 39080 636200
rect 675116 635468 675168 635520
rect 675484 635468 675536 635520
rect 35808 634924 35860 634976
rect 39488 634924 39540 634976
rect 35808 633836 35860 633888
rect 40132 633836 40184 633888
rect 35808 633564 35860 633616
rect 39764 633632 39816 633684
rect 35624 633428 35676 633480
rect 41604 633428 41656 633480
rect 42064 633428 42116 633480
rect 63408 633428 63460 633480
rect 672356 632680 672408 632732
rect 672724 632680 672776 632732
rect 36544 630572 36596 630624
rect 41604 630572 41656 630624
rect 35164 628668 35216 628720
rect 40500 628668 40552 628720
rect 673552 627648 673604 627700
rect 673920 627648 673972 627700
rect 674288 626220 674340 626272
rect 674840 626220 674892 626272
rect 674288 626016 674340 626068
rect 676220 626016 676272 626068
rect 44456 625812 44508 625864
rect 63132 625812 63184 625864
rect 667204 625608 667256 625660
rect 674012 625608 674064 625660
rect 674288 625608 674340 625660
rect 676220 625608 676272 625660
rect 657544 625268 657596 625320
rect 674012 625336 674064 625388
rect 669964 625200 670016 625252
rect 674012 625200 674064 625252
rect 674288 625200 674340 625252
rect 676220 625200 676272 625252
rect 670240 625064 670292 625116
rect 674012 625064 674064 625116
rect 674288 625064 674340 625116
rect 676496 625064 676548 625116
rect 669780 624588 669832 624640
rect 674012 624588 674064 624640
rect 674288 624452 674340 624504
rect 676220 624452 676272 624504
rect 674288 624316 674340 624368
rect 676036 624316 676088 624368
rect 669872 624248 669924 624300
rect 674012 624248 674064 624300
rect 670240 623840 670292 623892
rect 674012 623840 674064 623892
rect 671436 623636 671488 623688
rect 674012 623636 674064 623688
rect 674288 623568 674340 623620
rect 676220 623568 676272 623620
rect 670056 623024 670108 623076
rect 674012 623024 674064 623076
rect 671252 622820 671304 622872
rect 674012 622820 674064 622872
rect 674288 622820 674340 622872
rect 676220 622820 676272 622872
rect 671436 622208 671488 622260
rect 674012 622208 674064 622260
rect 42248 621664 42300 621716
rect 44548 621664 44600 621716
rect 674288 621188 674340 621240
rect 676220 621188 676272 621240
rect 666468 621120 666520 621172
rect 674012 621120 674064 621172
rect 670608 620780 670660 620832
rect 674012 620780 674064 620832
rect 674288 620780 674340 620832
rect 676220 620780 676272 620832
rect 42248 620372 42300 620424
rect 42708 620372 42760 620424
rect 674840 620168 674892 620220
rect 683120 620168 683172 620220
rect 674288 619760 674340 619812
rect 676036 619760 676088 619812
rect 668216 619692 668268 619744
rect 674012 619692 674064 619744
rect 42248 619624 42300 619676
rect 44272 619624 44324 619676
rect 673184 619284 673236 619336
rect 674012 619284 674064 619336
rect 674288 619148 674340 619200
rect 676496 619148 676548 619200
rect 674288 618332 674340 618384
rect 676220 618332 676272 618384
rect 668400 618264 668452 618316
rect 674012 618264 674064 618316
rect 674472 618196 674524 618248
rect 676036 618196 676088 618248
rect 670976 618060 671028 618112
rect 674012 618060 674064 618112
rect 674288 617924 674340 617976
rect 676220 617924 676272 617976
rect 42248 617312 42300 617364
rect 43076 617312 43128 617364
rect 44732 616768 44784 616820
rect 62120 616768 62172 616820
rect 669412 616700 669464 616752
rect 674012 616700 674064 616752
rect 674288 616632 674340 616684
rect 676220 616632 676272 616684
rect 43076 616496 43128 616548
rect 43812 616496 43864 616548
rect 672816 615612 672868 615664
rect 674012 615612 674064 615664
rect 674288 615476 674340 615528
rect 683120 615476 683172 615528
rect 670608 614864 670660 614916
rect 674012 614864 674064 614916
rect 43536 614660 43588 614712
rect 44364 614660 44416 614712
rect 42708 614116 42760 614168
rect 62120 614116 62172 614168
rect 673552 613504 673604 613556
rect 673736 613300 673788 613352
rect 42892 612756 42944 612808
rect 54484 612620 54536 612672
rect 62120 612620 62172 612672
rect 43076 612484 43128 612536
rect 43904 612212 43956 612264
rect 44548 612212 44600 612264
rect 43766 612144 43818 612196
rect 43875 611872 43927 611924
rect 47032 612008 47084 612060
rect 47216 611872 47268 611924
rect 44364 611600 44416 611652
rect 653404 611328 653456 611380
rect 674012 611328 674064 611380
rect 674288 611328 674340 611380
rect 675392 611328 675444 611380
rect 44318 611124 44370 611176
rect 44824 611192 44876 611244
rect 44548 611056 44600 611108
rect 657544 600312 657596 600364
rect 670884 600312 670936 600364
rect 670792 599088 670844 599140
rect 654784 598952 654836 599004
rect 674656 598884 674708 598936
rect 674656 598612 674708 598664
rect 651472 597524 651524 597576
rect 667388 597524 667440 597576
rect 42892 597388 42944 597440
rect 42892 596980 42944 597032
rect 672356 596232 672408 596284
rect 672724 596232 672776 596284
rect 651472 596164 651524 596216
rect 661684 596164 661736 596216
rect 39948 595756 40000 595808
rect 41696 595756 41748 595808
rect 651656 595484 651708 595536
rect 653404 595484 653456 595536
rect 651472 594804 651524 594856
rect 658924 594804 658976 594856
rect 651472 594668 651524 594720
rect 657544 594668 657596 594720
rect 38568 594124 38620 594176
rect 41696 594124 41748 594176
rect 651472 593036 651524 593088
rect 654784 593036 654836 593088
rect 674840 592492 674892 592544
rect 683396 592492 683448 592544
rect 675576 588548 675628 588600
rect 684040 588548 684092 588600
rect 35440 587120 35492 587172
rect 41512 587120 41564 587172
rect 36544 586100 36596 586152
rect 39672 586100 39724 586152
rect 32404 585896 32456 585948
rect 41696 585896 41748 585948
rect 31024 585760 31076 585812
rect 39764 585760 39816 585812
rect 652024 581000 652076 581052
rect 673920 581000 673972 581052
rect 668584 580252 668636 580304
rect 673920 580252 673972 580304
rect 669872 579844 669924 579896
rect 673920 579844 673972 579896
rect 660304 579640 660356 579692
rect 673552 579640 673604 579692
rect 669596 579368 669648 579420
rect 673920 579368 673972 579420
rect 670240 579028 670292 579080
rect 673920 579028 673972 579080
rect 670240 578552 670292 578604
rect 673920 578552 673972 578604
rect 670056 578144 670108 578196
rect 673920 578144 673972 578196
rect 669412 577736 669464 577788
rect 673920 577736 673972 577788
rect 42432 577600 42484 577652
rect 42616 577532 42668 577584
rect 42616 577396 42668 577448
rect 42340 577260 42392 577312
rect 671436 577396 671488 577448
rect 673920 577396 673972 577448
rect 671344 576920 671396 576972
rect 673920 576920 673972 576972
rect 45100 575424 45152 575476
rect 62396 575424 62448 575476
rect 671804 575356 671856 575408
rect 673920 575356 673972 575408
rect 670424 574540 670476 574592
rect 673552 574540 673604 574592
rect 671988 574268 672040 574320
rect 673552 574268 673604 574320
rect 667020 574064 667072 574116
rect 673920 574064 673972 574116
rect 45560 573996 45612 574048
rect 62396 573996 62448 574048
rect 672540 573724 672592 573776
rect 673920 573724 673972 573776
rect 671620 572092 671672 572144
rect 673920 572092 673972 572144
rect 674656 571548 674708 571600
rect 676220 571548 676272 571600
rect 671988 570800 672040 570852
rect 673920 570800 673972 570852
rect 667204 570528 667256 570580
rect 667664 570528 667716 570580
rect 667664 570188 667716 570240
rect 673920 570188 673972 570240
rect 674656 569916 674708 569968
rect 683120 569916 683172 569968
rect 669780 569576 669832 569628
rect 673552 569576 673604 569628
rect 42432 569372 42484 569424
rect 42432 569168 42484 569220
rect 653404 565836 653456 565888
rect 673552 565836 673604 565888
rect 674656 558016 674708 558068
rect 675300 558016 675352 558068
rect 657820 554752 657872 554804
rect 674012 554752 674064 554804
rect 655152 553392 655204 553444
rect 674012 553392 674064 553444
rect 40040 553324 40092 553376
rect 41696 553324 41748 553376
rect 651472 552644 651524 552696
rect 665824 552644 665876 552696
rect 41328 552100 41380 552152
rect 41696 552100 41748 552152
rect 651472 550604 651524 550656
rect 669964 550604 670016 550656
rect 41144 550536 41196 550588
rect 41696 550536 41748 550588
rect 651380 550332 651432 550384
rect 653404 550332 653456 550384
rect 675300 550060 675352 550112
rect 674748 549924 674800 549976
rect 674840 549788 674892 549840
rect 674748 549244 674800 549296
rect 651472 549176 651524 549228
rect 657820 549176 657872 549228
rect 651472 548836 651524 548888
rect 655152 548836 655204 548888
rect 674380 547272 674432 547324
rect 683212 547272 683264 547324
rect 675300 546864 675352 546916
rect 682384 546864 682436 546916
rect 672632 544552 672684 544604
rect 675024 544552 675076 544604
rect 675392 544552 675444 544604
rect 29644 544348 29696 544400
rect 41696 544348 41748 544400
rect 672816 544348 672868 544400
rect 674288 537140 674340 537192
rect 675484 537140 675536 537192
rect 673920 536392 673972 536444
rect 673920 536120 673972 536172
rect 673736 535984 673788 536036
rect 667388 535780 667440 535832
rect 673736 535780 673788 535832
rect 661684 535440 661736 535492
rect 669596 534964 669648 535016
rect 672632 534964 672684 535016
rect 670240 534284 670292 534336
rect 672632 534284 672684 534336
rect 674288 534216 674340 534268
rect 676220 534216 676272 534268
rect 658924 534080 658976 534132
rect 673736 534080 673788 534132
rect 42248 533400 42300 533452
rect 42984 533400 43036 533452
rect 669412 533332 669464 533384
rect 672632 533332 672684 533384
rect 675484 533332 675536 533384
rect 683580 533332 683632 533384
rect 674288 532788 674340 532840
rect 676036 532788 676088 532840
rect 44732 531224 44784 531276
rect 62304 531224 62356 531276
rect 53104 531088 53156 531140
rect 62120 531088 62172 531140
rect 673184 530068 673236 530120
rect 673736 530068 673788 530120
rect 668952 529932 669004 529984
rect 673736 529932 673788 529984
rect 670976 529456 671028 529508
rect 673736 529456 673788 529508
rect 671160 529184 671212 529236
rect 673736 529184 673788 529236
rect 673000 528844 673052 528896
rect 673736 528776 673788 528828
rect 45100 528572 45152 528624
rect 62120 528572 62172 528624
rect 674380 527552 674432 527604
rect 676220 527552 676272 527604
rect 54484 527076 54536 527128
rect 62120 527076 62172 527128
rect 674288 526736 674340 526788
rect 676036 526736 676088 526788
rect 674472 526328 674524 526380
rect 676036 526328 676088 526380
rect 674288 524560 674340 524612
rect 683120 524560 683172 524612
rect 668768 524356 668820 524408
rect 674012 524424 674064 524476
rect 652208 520888 652260 520940
rect 668768 520888 668820 520940
rect 675668 520208 675720 520260
rect 680360 520208 680412 520260
rect 675484 520072 675536 520124
rect 678980 520072 679032 520124
rect 674932 503820 674984 503872
rect 678244 503820 678296 503872
rect 675116 503616 675168 503668
rect 679624 503616 679676 503668
rect 675300 503480 675352 503532
rect 681004 503480 681056 503532
rect 652024 493280 652076 493332
rect 673184 493280 673236 493332
rect 669964 491444 670016 491496
rect 673828 491444 673880 491496
rect 674288 491444 674340 491496
rect 676036 491444 676088 491496
rect 665824 491308 665876 491360
rect 674012 491308 674064 491360
rect 670792 490900 670844 490952
rect 674012 490900 674064 490952
rect 672632 490084 672684 490136
rect 674012 490084 674064 490136
rect 672632 489880 672684 489932
rect 673184 489880 673236 489932
rect 672448 489608 672500 489660
rect 674012 489608 674064 489660
rect 671528 489268 671580 489320
rect 674012 489268 674064 489320
rect 671344 488452 671396 488504
rect 674012 488452 674064 488504
rect 671804 486820 671856 486872
rect 674012 486820 674064 486872
rect 672264 486004 672316 486056
rect 674012 486004 674064 486056
rect 676036 485324 676088 485376
rect 677140 485324 677192 485376
rect 674288 485120 674340 485172
rect 676036 485120 676088 485172
rect 667020 484372 667072 484424
rect 674012 484372 674064 484424
rect 674472 484372 674524 484424
rect 675852 484372 675904 484424
rect 676220 484304 676272 484356
rect 677416 484304 677468 484356
rect 674288 482468 674340 482520
rect 676036 482468 676088 482520
rect 668400 481924 668452 481976
rect 674012 482128 674064 482180
rect 674288 482060 674340 482112
rect 676036 482060 676088 482112
rect 667572 481788 667624 481840
rect 674012 481788 674064 481840
rect 658924 480904 658976 480956
rect 670424 480904 670476 480956
rect 674012 480904 674064 480956
rect 674288 480360 674340 480412
rect 683120 480360 683172 480412
rect 650644 476076 650696 476128
rect 652208 476076 652260 476128
rect 673368 475464 673420 475516
rect 674012 475464 674064 475516
rect 674288 475464 674340 475516
rect 676220 475464 676272 475516
rect 676036 475124 676088 475176
rect 680360 475124 680412 475176
rect 656164 466420 656216 466472
rect 658924 466420 658976 466472
rect 651380 458396 651432 458448
rect 656164 458396 656216 458448
rect 667848 456560 667900 456612
rect 674288 456084 674340 456136
rect 676220 456084 676272 456136
rect 673828 456016 673880 456068
rect 672816 455744 672868 455796
rect 669228 455608 669280 455660
rect 673276 455336 673328 455388
rect 672080 455064 672132 455116
rect 673388 455200 673440 455252
rect 673506 455200 673558 455252
rect 673046 454724 673098 454776
rect 674288 454724 674340 454776
rect 675668 454724 675720 454776
rect 650828 454520 650880 454572
rect 651380 454520 651432 454572
rect 674288 454452 674340 454504
rect 675484 454452 675536 454504
rect 672954 454384 673006 454436
rect 672816 454180 672868 454232
rect 674288 454180 674340 454232
rect 675852 454180 675904 454232
rect 672264 453908 672316 453960
rect 674288 453908 674340 453960
rect 676036 453908 676088 453960
rect 35808 429156 35860 429208
rect 41328 429156 41380 429208
rect 41144 425348 41196 425400
rect 41696 425348 41748 425400
rect 40960 420928 41012 420980
rect 41696 420928 41748 420980
rect 33048 415896 33100 415948
rect 40592 415896 40644 415948
rect 42248 406036 42300 406088
rect 42248 405628 42300 405680
rect 45100 404268 45152 404320
rect 62120 404268 62172 404320
rect 674564 403248 674616 403300
rect 676220 403248 676272 403300
rect 46112 402908 46164 402960
rect 62120 402908 62172 402960
rect 51080 400188 51132 400240
rect 62120 400188 62172 400240
rect 47952 400052 48004 400104
rect 62120 400052 62172 400104
rect 674932 398828 674984 398880
rect 676036 398828 676088 398880
rect 54484 398760 54536 398812
rect 62120 398760 62172 398812
rect 47584 397400 47636 397452
rect 50712 397400 50764 397452
rect 674380 396040 674432 396092
rect 676036 396040 676088 396092
rect 675024 395700 675076 395752
rect 676220 395700 676272 395752
rect 674472 394272 674524 394324
rect 676220 394272 676272 394324
rect 679624 386724 679676 386776
rect 674840 386112 674892 386164
rect 675300 386112 675352 386164
rect 675484 385976 675536 386028
rect 41328 382372 41380 382424
rect 41696 382372 41748 382424
rect 674380 382168 674432 382220
rect 675116 382168 675168 382220
rect 674564 378088 674616 378140
rect 675116 378088 675168 378140
rect 674380 375300 674432 375352
rect 675116 375300 675168 375352
rect 651472 373940 651524 373992
rect 657544 373940 657596 373992
rect 32404 373260 32456 373312
rect 41696 373260 41748 373312
rect 42064 373192 42116 373244
rect 42616 373192 42668 373244
rect 674748 372512 674800 372564
rect 675300 372512 675352 372564
rect 37924 372308 37976 372360
rect 41696 372308 41748 372360
rect 651472 370948 651524 371000
rect 654784 370948 654836 371000
rect 45376 361496 45428 361548
rect 62120 361496 62172 361548
rect 46756 360136 46808 360188
rect 62120 360136 62172 360188
rect 42156 359932 42208 359984
rect 42800 359932 42852 359984
rect 44640 359048 44692 359100
rect 45376 359048 45428 359100
rect 51724 357416 51776 357468
rect 62120 357416 62172 357468
rect 47952 355988 48004 356040
rect 62120 355988 62172 356040
rect 44640 354968 44692 355020
rect 44640 354628 44692 354680
rect 44732 354424 44784 354476
rect 45284 354356 45336 354408
rect 45284 353880 45336 353932
rect 45303 353676 45355 353728
rect 45836 353472 45888 353524
rect 45422 353200 45474 353252
rect 35808 344564 35860 344616
rect 40040 344564 40092 344616
rect 35532 343748 35584 343800
rect 39856 343748 39908 343800
rect 35808 342184 35860 342236
rect 40224 342184 40276 342236
rect 45468 342184 45520 342236
rect 62304 342184 62356 342236
rect 35808 341164 35860 341216
rect 40224 341164 40276 341216
rect 35624 341028 35676 341080
rect 39672 341028 39724 341080
rect 35532 339600 35584 339652
rect 36544 339600 36596 339652
rect 35808 339464 35860 339516
rect 38568 339464 38620 339516
rect 660304 338716 660356 338768
rect 669320 338716 669372 338768
rect 674380 336676 674432 336728
rect 675116 336676 675168 336728
rect 674380 336472 674432 336524
rect 675300 336472 675352 336524
rect 35808 336200 35860 336252
rect 40040 336200 40092 336252
rect 35532 335316 35584 335368
rect 40224 335316 40276 335368
rect 35808 334092 35860 334144
rect 39764 334092 39816 334144
rect 674472 331100 674524 331152
rect 675300 331100 675352 331152
rect 651472 328380 651524 328432
rect 667388 328380 667440 328432
rect 651380 325592 651432 325644
rect 653404 325592 653456 325644
rect 42248 319880 42300 319932
rect 43352 319880 43404 319932
rect 53840 317364 53892 317416
rect 62120 317364 62172 317416
rect 53104 315936 53156 315988
rect 62120 315936 62172 315988
rect 53840 314712 53892 314764
rect 62120 314712 62172 314764
rect 652024 313896 652076 313948
rect 660304 313896 660356 313948
rect 674564 311992 674616 312044
rect 675484 311992 675536 312044
rect 674840 306348 674892 306400
rect 675484 306348 675536 306400
rect 676220 306348 676272 306400
rect 676864 306348 676916 306400
rect 675852 304852 675904 304904
rect 676404 304852 676456 304904
rect 651472 302132 651524 302184
rect 667388 302132 667440 302184
rect 47584 301724 47636 301776
rect 51908 301724 51960 301776
rect 651472 300772 651524 300824
rect 660304 300772 660356 300824
rect 35624 298732 35676 298784
rect 41604 298732 41656 298784
rect 35808 298256 35860 298308
rect 41604 298256 41656 298308
rect 676128 298052 676180 298104
rect 678244 298052 678296 298104
rect 678980 298052 679032 298104
rect 675944 297916 675996 297968
rect 675024 297304 675076 297356
rect 675208 297100 675260 297152
rect 675024 296964 675076 297016
rect 674840 296828 674892 296880
rect 651748 296760 651800 296812
rect 35808 296692 35860 296744
rect 41604 296692 41656 296744
rect 665824 296692 665876 296744
rect 674472 295672 674524 295724
rect 675484 295672 675536 295724
rect 35624 295468 35676 295520
rect 39304 295468 39356 295520
rect 35808 295332 35860 295384
rect 41328 295332 41380 295384
rect 51908 295060 51960 295112
rect 56508 295060 56560 295112
rect 35440 294584 35492 294636
rect 41696 294584 41748 294636
rect 35808 293972 35860 294024
rect 40040 293972 40092 294024
rect 53104 293972 53156 294024
rect 62212 293972 62264 294024
rect 651472 293972 651524 294024
rect 664444 293972 664496 294024
rect 35808 292884 35860 292936
rect 39856 292816 39908 292868
rect 35808 292544 35860 292596
rect 54484 292544 54536 292596
rect 62304 292544 62356 292596
rect 46204 292408 46256 292460
rect 62120 292408 62172 292460
rect 41604 292340 41656 292392
rect 40776 292068 40828 292120
rect 41604 292068 41656 292120
rect 649264 291864 649316 291916
rect 652024 291864 652076 291916
rect 40040 291320 40092 291372
rect 41696 291320 41748 291372
rect 42156 291320 42208 291372
rect 43352 291320 43404 291372
rect 42064 291184 42116 291236
rect 42616 291184 42668 291236
rect 39856 291116 39908 291168
rect 41604 291116 41656 291168
rect 60004 291116 60056 291168
rect 62304 291116 62356 291168
rect 651472 289824 651524 289876
rect 663064 289824 663116 289876
rect 56508 289756 56560 289808
rect 58808 289756 58860 289808
rect 60004 288464 60056 288516
rect 62120 288464 62172 288516
rect 651472 288396 651524 288448
rect 672080 288396 672132 288448
rect 651656 287648 651708 287700
rect 672448 287648 672500 287700
rect 31024 286288 31076 286340
rect 41512 286288 41564 286340
rect 46204 285676 46256 285728
rect 62120 285676 62172 285728
rect 651472 285676 651524 285728
rect 672264 285676 672316 285728
rect 674656 285132 674708 285184
rect 35808 284928 35860 284980
rect 41696 284928 41748 284980
rect 674656 284928 674708 284980
rect 47584 284316 47636 284368
rect 62948 284316 63000 284368
rect 651472 284316 651524 284368
rect 672264 284316 672316 284368
rect 651472 282888 651524 282940
rect 667388 282888 667440 282940
rect 651472 281528 651524 281580
rect 667756 281528 667808 281580
rect 47952 280168 48004 280220
rect 62120 280168 62172 280220
rect 651472 280168 651524 280220
rect 667572 280168 667624 280220
rect 47768 278672 47820 278724
rect 650828 278672 650880 278724
rect 62856 278536 62908 278588
rect 672632 278536 672684 278588
rect 58808 278400 58860 278452
rect 650644 278400 650696 278452
rect 50712 278264 50764 278316
rect 649264 278264 649316 278316
rect 63224 278128 63276 278180
rect 667204 278128 667256 278180
rect 503536 277380 503588 277432
rect 587072 277380 587124 277432
rect 484032 277176 484084 277228
rect 561128 277176 561180 277228
rect 485504 277040 485556 277092
rect 562324 277040 562376 277092
rect 495072 276904 495124 276956
rect 576492 276904 576544 276956
rect 514484 276768 514536 276820
rect 603632 276768 603684 276820
rect 521108 276632 521160 276684
rect 613108 276632 613160 276684
rect 479984 276496 480036 276548
rect 554044 276496 554096 276548
rect 478512 276360 478564 276412
rect 551652 276360 551704 276412
rect 470416 276224 470468 276276
rect 539876 276224 539928 276276
rect 107200 275952 107252 276004
rect 163504 275952 163556 276004
rect 167552 275952 167604 276004
rect 178684 275952 178736 276004
rect 185216 275952 185268 276004
rect 221280 275952 221332 276004
rect 410800 275952 410852 276004
rect 455880 275952 455932 276004
rect 456432 275952 456484 276004
rect 509056 275952 509108 276004
rect 513196 275952 513248 276004
rect 601332 275952 601384 276004
rect 139124 275816 139176 275868
rect 174268 275816 174320 275868
rect 178132 275816 178184 275868
rect 216680 275816 216732 275868
rect 224224 275816 224276 275868
rect 233056 275816 233108 275868
rect 236092 275816 236144 275868
rect 250444 275816 250496 275868
rect 284576 275816 284628 275868
rect 290096 275816 290148 275868
rect 430212 275816 430264 275868
rect 484308 275816 484360 275868
rect 485044 275816 485096 275868
rect 491392 275816 491444 275868
rect 522764 275816 522816 275868
rect 615500 275816 615552 275868
rect 260932 275748 260984 275800
rect 266360 275748 266412 275800
rect 93032 275680 93084 275732
rect 152832 275680 152884 275732
rect 160468 275680 160520 275732
rect 199384 275680 199436 275732
rect 217140 275680 217192 275732
rect 224224 275680 224276 275732
rect 229008 275680 229060 275732
rect 243728 275680 243780 275732
rect 250260 275680 250312 275732
rect 259368 275680 259420 275732
rect 286876 275680 286928 275732
rect 291844 275680 291896 275732
rect 416412 275680 416464 275732
rect 462964 275680 463016 275732
rect 463148 275680 463200 275732
rect 516232 275680 516284 275732
rect 528192 275680 528244 275732
rect 622584 275680 622636 275732
rect 76472 275544 76524 275596
rect 86224 275544 86276 275596
rect 90732 275544 90784 275596
rect 154764 275544 154816 275596
rect 171048 275544 171100 275596
rect 211436 275544 211488 275596
rect 218336 275544 218388 275596
rect 233884 275544 233936 275596
rect 239588 275544 239640 275596
rect 255964 275544 256016 275596
rect 257344 275544 257396 275596
rect 262312 275544 262364 275596
rect 266820 275544 266872 275596
rect 276480 275544 276532 275596
rect 363880 275544 363932 275596
rect 388536 275544 388588 275596
rect 445024 275544 445076 275596
rect 498476 275544 498528 275596
rect 498844 275544 498896 275596
rect 505560 275544 505612 275596
rect 505744 275544 505796 275596
rect 512644 275544 512696 275596
rect 516784 275544 516836 275596
rect 526812 275544 526864 275596
rect 532332 275544 532384 275596
rect 629668 275544 629720 275596
rect 277492 275476 277544 275528
rect 285128 275476 285180 275528
rect 100116 275408 100168 275460
rect 71780 275272 71832 275324
rect 141056 275272 141108 275324
rect 156880 275408 156932 275460
rect 159456 275272 159508 275324
rect 163964 275408 164016 275460
rect 206376 275408 206428 275460
rect 221924 275408 221976 275460
rect 243544 275408 243596 275460
rect 256148 275408 256200 275460
rect 269396 275408 269448 275460
rect 285680 275408 285732 275460
rect 291200 275408 291252 275460
rect 358636 275408 358688 275460
rect 381452 275408 381504 275460
rect 385960 275408 386012 275460
rect 420460 275408 420512 275460
rect 435640 275408 435692 275460
rect 485044 275408 485096 275460
rect 485780 275408 485832 275460
rect 530400 275408 530452 275460
rect 537668 275408 537720 275460
rect 636752 275408 636804 275460
rect 299940 275340 299992 275392
rect 301136 275340 301188 275392
rect 200764 275272 200816 275324
rect 214840 275272 214892 275324
rect 239404 275272 239456 275324
rect 243176 275272 243228 275324
rect 256700 275272 256752 275324
rect 263232 275272 263284 275324
rect 273260 275272 273312 275324
rect 276296 275272 276348 275324
rect 283104 275272 283156 275324
rect 291660 275272 291712 275324
rect 295340 275272 295392 275324
rect 326436 275272 326488 275324
rect 335360 275272 335412 275324
rect 371056 275272 371108 275324
rect 399208 275272 399260 275324
rect 418804 275272 418856 275324
rect 466552 275272 466604 275324
rect 467564 275272 467616 275324
rect 537484 275272 537536 275324
rect 542084 275272 542136 275324
rect 643836 275272 643888 275324
rect 298744 275204 298796 275256
rect 300032 275204 300084 275256
rect 96620 275136 96672 275188
rect 149980 275136 150032 275188
rect 153384 275136 153436 275188
rect 169024 275136 169076 275188
rect 190000 275136 190052 275188
rect 222936 275136 222988 275188
rect 232504 275136 232556 275188
rect 240048 275136 240100 275188
rect 292856 275136 292908 275188
rect 295800 275136 295852 275188
rect 427084 275136 427136 275188
rect 477224 275136 477276 275188
rect 507492 275136 507544 275188
rect 594248 275136 594300 275188
rect 269212 275068 269264 275120
rect 274640 275068 274692 275120
rect 81256 275000 81308 275052
rect 145288 275000 145340 275052
rect 149796 275000 149848 275052
rect 189080 275000 189132 275052
rect 288072 275000 288124 275052
rect 292856 275000 292908 275052
rect 420552 275000 420604 275052
rect 470140 275000 470192 275052
rect 497924 275000 497976 275052
rect 579988 275000 580040 275052
rect 293960 274932 294012 274984
rect 297180 274932 297232 274984
rect 136824 274864 136876 274916
rect 137652 274864 137704 274916
rect 146208 274864 146260 274916
rect 185308 274864 185360 274916
rect 289268 274864 289320 274916
rect 292672 274864 292724 274916
rect 473084 274864 473136 274916
rect 544568 274864 544620 274916
rect 296352 274796 296404 274848
rect 298376 274796 298428 274848
rect 128544 274728 128596 274780
rect 167000 274728 167052 274780
rect 207756 274728 207808 274780
rect 210700 274728 210752 274780
rect 476764 274728 476816 274780
rect 523316 274728 523368 274780
rect 523684 274728 523736 274780
rect 533896 274728 533948 274780
rect 534724 274728 534776 274780
rect 540980 274728 541032 274780
rect 74172 274660 74224 274712
rect 76840 274660 76892 274712
rect 85948 274660 86000 274712
rect 90364 274660 90416 274712
rect 103704 274660 103756 274712
rect 104808 274660 104860 274712
rect 110788 274660 110840 274712
rect 111708 274660 111760 274712
rect 253848 274660 253900 274712
rect 256884 274660 256936 274712
rect 275100 274660 275152 274712
rect 278412 274660 278464 274712
rect 283380 274660 283432 274712
rect 289176 274660 289228 274712
rect 290464 274660 290516 274712
rect 294144 274660 294196 274712
rect 295156 274660 295208 274712
rect 296812 274660 296864 274712
rect 297548 274660 297600 274712
rect 299480 274660 299532 274712
rect 303436 274660 303488 274712
rect 303988 274660 304040 274712
rect 321192 274660 321244 274712
rect 328276 274660 328328 274712
rect 114376 274592 114428 274644
rect 171600 274592 171652 274644
rect 179328 274592 179380 274644
rect 214564 274592 214616 274644
rect 409788 274592 409840 274644
rect 453580 274592 453632 274644
rect 101312 274456 101364 274508
rect 160928 274456 160980 274508
rect 168748 274456 168800 274508
rect 208400 274456 208452 274508
rect 381544 274456 381596 274508
rect 392124 274456 392176 274508
rect 413836 274456 413888 274508
rect 460664 274592 460716 274644
rect 464436 274592 464488 274644
rect 480720 274592 480772 274644
rect 486792 274592 486844 274644
rect 563428 274592 563480 274644
rect 456064 274456 456116 274508
rect 465908 274456 465960 274508
rect 466092 274456 466144 274508
rect 485780 274456 485832 274508
rect 488356 274456 488408 274508
rect 567016 274456 567068 274508
rect 95424 274320 95476 274372
rect 157616 274320 157668 274372
rect 159272 274320 159324 274372
rect 202328 274320 202380 274372
rect 223120 274320 223172 274372
rect 247224 274320 247276 274372
rect 368940 274320 368992 274372
rect 387340 274320 387392 274372
rect 419080 274320 419132 274372
rect 467748 274320 467800 274372
rect 331956 274252 332008 274304
rect 337752 274252 337804 274304
rect 67088 274184 67140 274236
rect 130384 274184 130436 274236
rect 130844 274184 130896 274236
rect 182456 274184 182508 274236
rect 193496 274184 193548 274236
rect 226432 274184 226484 274236
rect 240048 274184 240100 274236
rect 253940 274184 253992 274236
rect 359464 274184 359516 274236
rect 380256 274184 380308 274236
rect 388996 274184 389048 274236
rect 425152 274184 425204 274236
rect 425704 274184 425756 274236
rect 474832 274320 474884 274372
rect 506204 274320 506256 274372
rect 591856 274320 591908 274372
rect 472256 274184 472308 274236
rect 77668 274048 77720 274100
rect 144920 274048 144972 274100
rect 154488 274048 154540 274100
rect 198096 274048 198148 274100
rect 210056 274048 210108 274100
rect 237840 274048 237892 274100
rect 249064 274048 249116 274100
rect 265256 274048 265308 274100
rect 266360 274048 266412 274100
rect 273536 274048 273588 274100
rect 278596 274048 278648 274100
rect 285864 274048 285916 274100
rect 337752 274048 337804 274100
rect 351920 274048 351972 274100
rect 353944 274048 353996 274100
rect 369584 274048 369636 274100
rect 373264 274048 373316 274100
rect 400312 274048 400364 274100
rect 401508 274048 401560 274100
rect 442908 274048 442960 274100
rect 451188 274048 451240 274100
rect 456064 274048 456116 274100
rect 456248 274048 456300 274100
rect 481364 274184 481416 274236
rect 485320 274184 485372 274236
rect 511632 274184 511684 274236
rect 598940 274184 598992 274236
rect 69388 273912 69440 273964
rect 139400 273912 139452 273964
rect 148600 273912 148652 273964
rect 194784 273912 194836 273964
rect 208860 273912 208912 273964
rect 237380 273912 237432 273964
rect 238484 273912 238536 273964
rect 88340 273776 88392 273828
rect 119344 273776 119396 273828
rect 120264 273776 120316 273828
rect 175280 273776 175332 273828
rect 192392 273776 192444 273828
rect 224960 273776 225012 273828
rect 271512 273912 271564 273964
rect 280344 273912 280396 273964
rect 322756 273912 322808 273964
rect 330576 273912 330628 273964
rect 335268 273912 335320 273964
rect 348332 273912 348384 273964
rect 350356 273912 350408 273964
rect 368480 273912 368532 273964
rect 377680 273912 377732 273964
rect 408592 273912 408644 273964
rect 422116 273912 422168 273964
rect 465724 273912 465776 273964
rect 465908 273912 465960 273964
rect 472256 273912 472308 273964
rect 513840 274048 513892 274100
rect 536748 274048 536800 274100
rect 634360 274048 634412 274100
rect 481916 273912 481968 273964
rect 258080 273776 258132 273828
rect 397000 273776 397052 273828
rect 435824 273776 435876 273828
rect 438124 273776 438176 273828
rect 473636 273776 473688 273828
rect 474648 273776 474700 273828
rect 545764 273912 545816 273964
rect 545948 273912 546000 273964
rect 639144 273912 639196 273964
rect 119068 273640 119120 273692
rect 173256 273640 173308 273692
rect 440884 273640 440936 273692
rect 132040 273504 132092 273556
rect 153844 273504 153896 273556
rect 259368 273504 259420 273556
rect 266360 273504 266412 273556
rect 447784 273504 447836 273556
rect 456248 273504 456300 273556
rect 457444 273504 457496 273556
rect 464436 273504 464488 273556
rect 465724 273640 465776 273692
rect 472440 273640 472492 273692
rect 484216 273640 484268 273692
rect 559932 273776 559984 273828
rect 485320 273640 485372 273692
rect 556344 273640 556396 273692
rect 556804 273640 556856 273692
rect 590660 273640 590712 273692
rect 471244 273504 471296 273556
rect 476028 273504 476080 273556
rect 549260 273504 549312 273556
rect 551284 273504 551336 273556
rect 583576 273504 583628 273556
rect 145288 273368 145340 273420
rect 147864 273368 147916 273420
rect 463240 273368 463292 273420
rect 466092 273368 466144 273420
rect 478696 273368 478748 273420
rect 552848 273368 552900 273420
rect 327724 273232 327776 273284
rect 329472 273232 329524 273284
rect 108396 273164 108448 273216
rect 165896 273164 165948 273216
rect 186412 273164 186464 273216
rect 218704 273164 218756 273216
rect 362776 273164 362828 273216
rect 386144 273164 386196 273216
rect 400036 273164 400088 273216
rect 439320 273164 439372 273216
rect 444012 273164 444064 273216
rect 102508 273028 102560 273080
rect 162860 273028 162912 273080
rect 172244 273028 172296 273080
rect 209780 273028 209832 273080
rect 219532 273028 219584 273080
rect 244556 273028 244608 273080
rect 280988 273028 281040 273080
rect 286324 273028 286376 273080
rect 361212 273028 361264 273080
rect 384948 273028 385000 273080
rect 385684 273028 385736 273080
rect 395620 273028 395672 273080
rect 404176 273028 404228 273080
rect 446496 273028 446548 273080
rect 446864 273028 446916 273080
rect 499488 273028 499540 273080
rect 499948 273164 500000 273216
rect 511448 273164 511500 273216
rect 503168 273028 503220 273080
rect 503352 273028 503404 273080
rect 507952 273028 508004 273080
rect 509700 273028 509752 273080
rect 515220 273164 515272 273216
rect 515404 273164 515456 273216
rect 519728 273164 519780 273216
rect 521476 273164 521528 273216
rect 614304 273164 614356 273216
rect 513564 273028 513616 273080
rect 518532 273028 518584 273080
rect 94228 272892 94280 272944
rect 155960 272892 156012 272944
rect 166356 272892 166408 272944
rect 207296 272892 207348 272944
rect 211252 272892 211304 272944
rect 220084 272892 220136 272944
rect 220728 272892 220780 272944
rect 245752 272892 245804 272944
rect 247868 272892 247920 272944
rect 264244 272892 264296 272944
rect 333796 272892 333848 272944
rect 345940 272892 345992 272944
rect 348424 272892 348476 272944
rect 362500 272892 362552 272944
rect 365444 272892 365496 272944
rect 390928 272892 390980 272944
rect 405556 272892 405608 272944
rect 448796 272892 448848 272944
rect 455328 272892 455380 272944
rect 461400 272892 461452 272944
rect 82452 272756 82504 272808
rect 148416 272756 148468 272808
rect 155684 272756 155736 272808
rect 200120 272756 200172 272808
rect 205364 272756 205416 272808
rect 234804 272756 234856 272808
rect 245384 272756 245436 272808
rect 72976 272620 73028 272672
rect 142160 272620 142212 272672
rect 142712 272620 142764 272672
rect 145564 272620 145616 272672
rect 147404 272620 147456 272672
rect 193220 272620 193272 272672
rect 195888 272620 195940 272672
rect 227904 272620 227956 272672
rect 228088 272620 228140 272672
rect 249064 272620 249116 272672
rect 262312 272756 262364 272808
rect 270960 272756 271012 272808
rect 273904 272756 273956 272808
rect 282920 272756 282972 272808
rect 325332 272756 325384 272808
rect 332968 272756 333020 272808
rect 344652 272756 344704 272808
rect 361396 272756 361448 272808
rect 362224 272756 362276 272808
rect 370780 272756 370832 272808
rect 262680 272620 262732 272672
rect 264428 272620 264480 272672
rect 269120 272620 269172 272672
rect 269396 272620 269448 272672
rect 270592 272620 270644 272672
rect 324044 272620 324096 272672
rect 331772 272620 331824 272672
rect 332324 272620 332376 272672
rect 343640 272620 343692 272672
rect 346216 272620 346268 272672
rect 363696 272620 363748 272672
rect 370504 272620 370556 272672
rect 396816 272756 396868 272808
rect 406844 272756 406896 272808
rect 449992 272756 450044 272808
rect 452292 272756 452344 272808
rect 515036 272892 515088 272944
rect 515220 272892 515272 272944
rect 562140 273028 562192 273080
rect 562324 273028 562376 273080
rect 601148 273028 601200 273080
rect 532516 272892 532568 272944
rect 376116 272620 376168 272672
rect 406292 272620 406344 272672
rect 412272 272620 412324 272672
rect 457076 272620 457128 272672
rect 457260 272620 457312 272672
rect 461032 272620 461084 272672
rect 461400 272620 461452 272672
rect 513564 272756 513616 272808
rect 513748 272756 513800 272808
rect 525616 272756 525668 272808
rect 529848 272756 529900 272808
rect 532884 272756 532936 272808
rect 533712 272756 533764 272808
rect 538680 272756 538732 272808
rect 539048 272892 539100 272944
rect 624976 273028 625028 273080
rect 618444 272892 618496 272944
rect 621388 272892 621440 272944
rect 628472 272756 628524 272808
rect 461860 272620 461912 272672
rect 319076 272552 319128 272604
rect 319628 272552 319680 272604
rect 466414 272620 466466 272672
rect 522120 272620 522172 272672
rect 526812 272620 526864 272672
rect 618444 272620 618496 272672
rect 620284 272620 620336 272672
rect 635556 272620 635608 272672
rect 65892 272484 65944 272536
rect 136824 272484 136876 272536
rect 137928 272484 137980 272536
rect 116676 272348 116728 272400
rect 172520 272348 172572 272400
rect 181720 272484 181772 272536
rect 187148 272484 187200 272536
rect 189080 272484 189132 272536
rect 196440 272484 196492 272536
rect 197084 272484 197136 272536
rect 229100 272484 229152 272536
rect 233700 272484 233752 272536
rect 254400 272484 254452 272536
rect 254952 272484 255004 272536
rect 269304 272484 269356 272536
rect 270316 272484 270368 272536
rect 280528 272484 280580 272536
rect 329748 272484 329800 272536
rect 338856 272484 338908 272536
rect 339224 272484 339276 272536
rect 354220 272484 354272 272536
rect 354496 272484 354548 272536
rect 375564 272484 375616 272536
rect 379428 272484 379480 272536
rect 410984 272484 411036 272536
rect 416596 272484 416648 272536
rect 463700 272484 463752 272536
rect 470554 272484 470606 272536
rect 470692 272484 470744 272536
rect 532700 272484 532752 272536
rect 532884 272484 532936 272536
rect 538496 272484 538548 272536
rect 538680 272484 538732 272536
rect 632060 272484 632112 272536
rect 634084 272484 634136 272536
rect 640340 272484 640392 272536
rect 318708 272416 318760 272468
rect 324688 272416 324740 272468
rect 187700 272348 187752 272400
rect 194968 272348 195020 272400
rect 227168 272348 227220 272400
rect 269120 272348 269172 272400
rect 276020 272348 276072 272400
rect 395988 272348 396040 272400
rect 434628 272348 434680 272400
rect 449716 272348 449768 272400
rect 499488 272348 499540 272400
rect 499672 272348 499724 272400
rect 513748 272348 513800 272400
rect 517428 272348 517480 272400
rect 600964 272348 601016 272400
rect 601148 272348 601200 272400
rect 620284 272348 620336 272400
rect 127348 272212 127400 272264
rect 179880 272212 179932 272264
rect 391848 272212 391900 272264
rect 428740 272212 428792 272264
rect 450544 272212 450596 272264
rect 510252 272212 510304 272264
rect 520096 272212 520148 272264
rect 610716 272212 610768 272264
rect 145104 272076 145156 272128
rect 192392 272076 192444 272128
rect 384948 272076 385000 272128
rect 418068 272076 418120 272128
rect 431684 272076 431736 272128
rect 480168 272076 480220 272128
rect 124956 271940 125008 271992
rect 151084 271940 151136 271992
rect 428464 271940 428516 271992
rect 470554 271940 470606 271992
rect 470692 271940 470744 271992
rect 489874 272076 489926 272128
rect 490012 272076 490064 272128
rect 552296 272076 552348 272128
rect 562324 272076 562376 272128
rect 600964 272076 601016 272128
rect 607220 272076 607272 272128
rect 483204 271940 483256 271992
rect 547512 271940 547564 271992
rect 547696 271940 547748 271992
rect 552848 271940 552900 271992
rect 558736 271940 558788 271992
rect 562140 271940 562192 271992
rect 569408 271940 569460 271992
rect 106004 271804 106056 271856
rect 164976 271804 165028 271856
rect 174268 271804 174320 271856
rect 189264 271804 189316 271856
rect 202972 271804 203024 271856
rect 233240 271804 233292 271856
rect 274640 271804 274692 271856
rect 279240 271804 279292 271856
rect 355324 271804 355376 271856
rect 356612 271804 356664 271856
rect 375288 271804 375340 271856
rect 403900 271804 403952 271856
rect 433156 271804 433208 271856
rect 97816 271668 97868 271720
rect 158812 271668 158864 271720
rect 169852 271668 169904 271720
rect 209964 271668 210016 271720
rect 225420 271668 225472 271720
rect 228364 271668 228416 271720
rect 351184 271668 351236 271720
rect 366088 271668 366140 271720
rect 382004 271668 382056 271720
rect 414572 271668 414624 271720
rect 87144 271532 87196 271584
rect 152004 271532 152056 271584
rect 165160 271532 165212 271584
rect 205640 271532 205692 271584
rect 215944 271532 215996 271584
rect 242072 271532 242124 271584
rect 337936 271532 337988 271584
rect 350724 271532 350776 271584
rect 360844 271532 360896 271584
rect 377864 271532 377916 271584
rect 387708 271532 387760 271584
rect 421656 271668 421708 271720
rect 430396 271668 430448 271720
rect 483020 271668 483072 271720
rect 485044 271804 485096 271856
rect 490012 271804 490064 271856
rect 496544 271804 496596 271856
rect 578884 271804 578936 271856
rect 486608 271668 486660 271720
rect 494704 271668 494756 271720
rect 501788 271668 501840 271720
rect 501972 271668 502024 271720
rect 585968 271668 586020 271720
rect 420184 271532 420236 271584
rect 431132 271532 431184 271584
rect 437204 271532 437256 271584
rect 493692 271532 493744 271584
rect 499304 271532 499356 271584
rect 582380 271532 582432 271584
rect 583024 271532 583076 271584
rect 611636 271532 611688 271584
rect 612004 271532 612056 271584
rect 618996 271532 619048 271584
rect 75368 271396 75420 271448
rect 142712 271396 142764 271448
rect 162676 271396 162728 271448
rect 204720 271396 204772 271448
rect 213644 271396 213696 271448
rect 240416 271396 240468 271448
rect 240784 271396 240836 271448
rect 259644 271396 259696 271448
rect 259828 271396 259880 271448
rect 272616 271396 272668 271448
rect 325516 271396 325568 271448
rect 334164 271396 334216 271448
rect 347688 271396 347740 271448
rect 364892 271396 364944 271448
rect 366364 271396 366416 271448
rect 383844 271396 383896 271448
rect 384764 271396 384816 271448
rect 419264 271396 419316 271448
rect 76840 271260 76892 271312
rect 143540 271260 143592 271312
rect 152188 271260 152240 271312
rect 197360 271260 197412 271312
rect 198280 271260 198332 271312
rect 229560 271260 229612 271312
rect 235264 271260 235316 271312
rect 255320 271260 255372 271312
rect 256700 271260 256752 271312
rect 261024 271260 261076 271312
rect 262036 271260 262088 271312
rect 274640 271260 274692 271312
rect 329564 271260 329616 271312
rect 340052 271260 340104 271312
rect 340604 271260 340656 271312
rect 355140 271260 355192 271312
rect 357164 271260 357216 271312
rect 379060 271260 379112 271312
rect 390284 271260 390336 271312
rect 426348 271396 426400 271448
rect 439964 271396 440016 271448
rect 497280 271396 497332 271448
rect 505008 271396 505060 271448
rect 589464 271396 589516 271448
rect 589924 271396 589976 271448
rect 633256 271396 633308 271448
rect 68192 271124 68244 271176
rect 138480 271124 138532 271176
rect 141516 271124 141568 271176
rect 189080 271124 189132 271176
rect 191196 271124 191248 271176
rect 225144 271124 225196 271176
rect 230204 271124 230256 271176
rect 252008 271124 252060 271176
rect 268016 271124 268068 271176
rect 278872 271124 278924 271176
rect 279792 271124 279844 271176
rect 287060 271124 287112 271176
rect 331128 271124 331180 271176
rect 342444 271124 342496 271176
rect 343548 271124 343600 271176
rect 360200 271124 360252 271176
rect 364156 271124 364208 271176
rect 389732 271124 389784 271176
rect 394332 271124 394384 271176
rect 432236 271260 432288 271312
rect 442908 271260 442960 271312
rect 500868 271260 500920 271312
rect 507676 271260 507728 271312
rect 593052 271260 593104 271312
rect 598204 271260 598256 271312
rect 645032 271260 645084 271312
rect 113456 270988 113508 271040
rect 169944 270988 169996 271040
rect 187424 270988 187476 271040
rect 216128 270988 216180 271040
rect 251456 270988 251508 271040
rect 266912 270988 266964 271040
rect 417424 270988 417476 271040
rect 437940 271124 437992 271176
rect 441344 271124 441396 271176
rect 445024 271124 445076 271176
rect 445668 271124 445720 271176
rect 504364 271124 504416 271176
rect 524052 271124 524104 271176
rect 617340 271124 617392 271176
rect 617524 271124 617576 271176
rect 626080 271124 626132 271176
rect 427452 270988 427504 271040
rect 479156 270988 479208 271040
rect 482284 270988 482336 271040
rect 494704 270988 494756 271040
rect 495256 270988 495308 271040
rect 575296 270988 575348 271040
rect 576124 270988 576176 271040
rect 604828 270988 604880 271040
rect 123760 270852 123812 270904
rect 177488 270852 177540 270904
rect 407764 270852 407816 270904
rect 440516 270852 440568 270904
rect 449164 270852 449216 270904
rect 490196 270852 490248 270904
rect 492496 270852 492548 270904
rect 571708 270852 571760 270904
rect 134432 270716 134484 270768
rect 185124 270716 185176 270768
rect 321376 270716 321428 270768
rect 327080 270716 327132 270768
rect 414480 270716 414532 270768
rect 450820 270716 450872 270768
rect 486976 270716 487028 270768
rect 564624 270716 564676 270768
rect 567844 270716 567896 270768
rect 597744 270716 597796 270768
rect 121460 270580 121512 270632
rect 168104 270580 168156 270632
rect 403624 270580 403676 270632
rect 433432 270580 433484 270632
rect 453304 270580 453356 270632
rect 487804 270580 487856 270632
rect 489644 270580 489696 270632
rect 568212 270580 568264 270632
rect 84108 270444 84160 270496
rect 137468 270444 137520 270496
rect 137652 270444 137704 270496
rect 186136 270444 186188 270496
rect 200764 270444 200816 270496
rect 201868 270444 201920 270496
rect 206836 270444 206888 270496
rect 235816 270444 235868 270496
rect 278412 270444 278464 270496
rect 283840 270444 283892 270496
rect 400864 270444 400916 270496
rect 441620 270444 441672 270496
rect 456432 270444 456484 270496
rect 520280 270444 520332 270496
rect 523132 270444 523184 270496
rect 532792 270444 532844 270496
rect 619640 270444 619692 270496
rect 78864 270308 78916 270360
rect 132500 270308 132552 270360
rect 133788 270308 133840 270360
rect 183652 270308 183704 270360
rect 185308 270308 185360 270360
rect 194416 270308 194468 270360
rect 199936 270308 199988 270360
rect 230848 270308 230900 270360
rect 233056 270308 233108 270360
rect 248236 270308 248288 270360
rect 283104 270308 283156 270360
rect 284668 270308 284720 270360
rect 355048 270308 355100 270360
rect 376944 270308 376996 270360
rect 380532 270308 380584 270360
rect 404360 270308 404412 270360
rect 409604 270308 409656 270360
rect 454040 270308 454092 270360
rect 458824 270308 458876 270360
rect 524420 270308 524472 270360
rect 525616 270308 525668 270360
rect 533528 270308 533580 270360
rect 626540 270308 626592 270360
rect 111984 270172 112036 270224
rect 168748 270172 168800 270224
rect 184848 270172 184900 270224
rect 219348 270172 219400 270224
rect 244372 270172 244424 270224
rect 262312 270172 262364 270224
rect 334348 270172 334400 270224
rect 346400 270172 346452 270224
rect 372252 270172 372304 270224
rect 397460 270172 397512 270224
rect 397920 270172 397972 270224
rect 412640 270172 412692 270224
rect 414664 270172 414716 270224
rect 461216 270172 461268 270224
rect 461400 270172 461452 270224
rect 527180 270172 527232 270224
rect 528376 270172 528428 270224
rect 533252 270172 533304 270224
rect 533528 270172 533580 270224
rect 623964 270172 624016 270224
rect 89628 270036 89680 270088
rect 153016 270036 153068 270088
rect 176568 270036 176620 270088
rect 211160 270036 211212 270088
rect 212448 270036 212500 270088
rect 239956 270036 240008 270088
rect 241888 270036 241940 270088
rect 260656 270036 260708 270088
rect 266176 270036 266228 270088
rect 277216 270036 277268 270088
rect 345296 270036 345348 270088
rect 358820 270036 358872 270088
rect 366640 270036 366692 270088
rect 393320 270036 393372 270088
rect 394700 270036 394752 270088
rect 408776 270036 408828 270088
rect 412456 270036 412508 270088
rect 458180 270036 458232 270088
rect 463516 270036 463568 270088
rect 530768 270036 530820 270088
rect 530952 270036 531004 270088
rect 532976 270036 533028 270088
rect 85488 269900 85540 269952
rect 149704 269900 149756 269952
rect 152832 269900 152884 269952
rect 157156 269900 157208 269952
rect 173808 269900 173860 269952
rect 212632 269900 212684 269952
rect 226616 269900 226668 269952
rect 249892 269900 249944 269952
rect 256884 269900 256936 269952
rect 268936 269900 268988 269952
rect 330208 269900 330260 269952
rect 340880 269900 340932 269952
rect 341800 269900 341852 269952
rect 357440 269900 357492 269952
rect 359188 269900 359240 269952
rect 382280 269900 382332 269952
rect 383016 269900 383068 269952
rect 411260 269900 411312 269952
rect 419632 269900 419684 269952
rect 467932 269900 467984 269952
rect 468484 269900 468536 269952
rect 538312 270036 538364 270088
rect 533988 269900 534040 269952
rect 630680 270036 630732 270088
rect 540520 269900 540572 269952
rect 640524 269900 640576 269952
rect 70584 269764 70636 269816
rect 79324 269764 79376 269816
rect 80060 269764 80112 269816
rect 146392 269764 146444 269816
rect 158628 269764 158680 269816
rect 201040 269764 201092 269816
rect 201684 269764 201736 269816
rect 232504 269764 232556 269816
rect 237196 269764 237248 269816
rect 257344 269764 257396 269816
rect 258540 269764 258592 269816
rect 272248 269764 272300 269816
rect 273076 269764 273128 269816
rect 282184 269764 282236 269816
rect 326896 269764 326948 269816
rect 335544 269764 335596 269816
rect 336004 269764 336056 269816
rect 349160 269764 349212 269816
rect 351736 269764 351788 269816
rect 371240 269764 371292 269816
rect 376576 269764 376628 269816
rect 407120 269764 407172 269816
rect 417148 269764 417200 269816
rect 465080 269764 465132 269816
rect 466000 269764 466052 269816
rect 532240 269764 532292 269816
rect 122748 269628 122800 269680
rect 176200 269628 176252 269680
rect 183468 269628 183520 269680
rect 205456 269628 205508 269680
rect 392032 269628 392084 269680
rect 401692 269628 401744 269680
rect 404360 269628 404412 269680
rect 423680 269628 423732 269680
rect 423864 269628 423916 269680
rect 451372 269628 451424 269680
rect 453580 269628 453632 269680
rect 509240 269628 509292 269680
rect 538864 269764 538916 269816
rect 539048 269764 539100 269816
rect 541624 269764 541676 269816
rect 541808 269764 541860 269816
rect 637580 269764 637632 269816
rect 129648 269492 129700 269544
rect 181168 269492 181220 269544
rect 204168 269492 204220 269544
rect 223488 269492 223540 269544
rect 401692 269492 401744 269544
rect 416780 269492 416832 269544
rect 424600 269492 424652 269544
rect 475016 269492 475068 269544
rect 492772 269492 492824 269544
rect 532792 269628 532844 269680
rect 615684 269628 615736 269680
rect 509884 269492 509936 269544
rect 596180 269492 596232 269544
rect 126888 269356 126940 269408
rect 178316 269356 178368 269408
rect 408316 269356 408368 269408
rect 426532 269356 426584 269408
rect 441620 269356 441672 269408
rect 458456 269356 458508 269408
rect 470968 269356 471020 269408
rect 538680 269356 538732 269408
rect 538864 269356 538916 269408
rect 572720 269356 572772 269408
rect 143908 269220 143960 269272
rect 191104 269220 191156 269272
rect 282736 269220 282788 269272
rect 288808 269220 288860 269272
rect 474280 269220 474332 269272
rect 546500 269220 546552 269272
rect 319444 269084 319496 269136
rect 325700 269084 325752 269136
rect 118608 269016 118660 269068
rect 174544 269016 174596 269068
rect 175096 269016 175148 269068
rect 177672 269016 177724 269068
rect 273260 269016 273312 269068
rect 275560 269016 275612 269068
rect 436560 269016 436612 269068
rect 491668 269016 491720 269068
rect 493324 269016 493376 269068
rect 574100 269016 574152 269068
rect 115848 268880 115900 268932
rect 110328 268744 110380 268796
rect 104992 268608 105044 268660
rect 163780 268608 163832 268660
rect 99288 268472 99340 268524
rect 160468 268472 160520 268524
rect 188896 268880 188948 268932
rect 190552 268880 190604 268932
rect 382372 268880 382424 268932
rect 415400 268880 415452 268932
rect 433708 268880 433760 268932
rect 488540 268880 488592 268932
rect 498292 268880 498344 268932
rect 581000 268880 581052 268932
rect 167000 268744 167052 268796
rect 181996 268744 182048 268796
rect 200580 268744 200632 268796
rect 231308 268744 231360 268796
rect 387340 268744 387392 268796
rect 422300 268744 422352 268796
rect 438676 268744 438728 268796
rect 495440 268744 495492 268796
rect 500776 268744 500828 268796
rect 583760 268744 583812 268796
rect 171232 268608 171284 268660
rect 176936 268608 176988 268660
rect 215116 268608 215168 268660
rect 224224 268608 224276 268660
rect 243268 268608 243320 268660
rect 352564 268608 352616 268660
rect 372620 268608 372672 268660
rect 393320 268608 393372 268660
rect 429200 268608 429252 268660
rect 441160 268608 441212 268660
rect 500132 268608 500184 268660
rect 503260 268608 503312 268660
rect 587900 268608 587952 268660
rect 167920 268472 167972 268524
rect 180616 268472 180668 268524
rect 217600 268472 217652 268524
rect 231676 268472 231728 268524
rect 253204 268472 253256 268524
rect 338488 268472 338540 268524
rect 352104 268472 352156 268524
rect 367468 268472 367520 268524
rect 393504 268472 393556 268524
rect 397276 268472 397328 268524
rect 436100 268472 436152 268524
rect 446128 268472 446180 268524
rect 506480 268472 506532 268524
rect 508228 268472 508280 268524
rect 594800 268472 594852 268524
rect 92388 268336 92440 268388
rect 155500 268336 155552 268388
rect 161572 268336 161624 268388
rect 203524 268336 203576 268388
rect 210700 268336 210752 268388
rect 236644 268336 236696 268388
rect 252652 268336 252704 268388
rect 268108 268336 268160 268388
rect 348792 268336 348844 268388
rect 367100 268336 367152 268388
rect 372436 268336 372488 268388
rect 400496 268336 400548 268388
rect 402244 268336 402296 268388
rect 443092 268336 443144 268388
rect 461860 268336 461912 268388
rect 528560 268336 528612 268388
rect 541348 268336 541400 268388
rect 641720 268336 641772 268388
rect 140688 268200 140740 268252
rect 188620 268200 188672 268252
rect 416228 268200 416280 268252
rect 447140 268200 447192 268252
rect 448428 268200 448480 268252
rect 494060 268200 494112 268252
rect 495808 268200 495860 268252
rect 576860 268200 576912 268252
rect 151728 268064 151780 268116
rect 196072 268064 196124 268116
rect 422300 268064 422352 268116
rect 444380 268064 444432 268116
rect 527180 268064 527232 268116
rect 607404 268064 607456 268116
rect 490840 267928 490892 267980
rect 569960 267928 570012 267980
rect 135628 267792 135680 267844
rect 130384 267656 130436 267708
rect 138112 267656 138164 267708
rect 276480 267724 276532 267776
rect 278044 267724 278096 267776
rect 186964 267656 187016 267708
rect 187148 267656 187200 267708
rect 195244 267656 195296 267708
rect 353392 267656 353444 267708
rect 374460 267656 374512 267708
rect 378232 267656 378284 267708
rect 394700 267656 394752 267708
rect 408040 267656 408092 267708
rect 423864 267656 423916 267708
rect 445300 267656 445352 267708
rect 498844 267656 498896 267708
rect 509884 267656 509936 267708
rect 567844 267656 567896 267708
rect 111708 267520 111760 267572
rect 169576 267520 169628 267572
rect 178684 267520 178736 267572
rect 209320 267520 209372 267572
rect 368296 267520 368348 267572
rect 385684 267520 385736 267572
rect 403072 267520 403124 267572
rect 422300 267520 422352 267572
rect 428740 267520 428792 267572
rect 447784 267520 447836 267572
rect 450268 267520 450320 267572
rect 505744 267520 505796 267572
rect 514852 267520 514904 267572
rect 576124 267520 576176 267572
rect 86224 267384 86276 267436
rect 144736 267384 144788 267436
rect 153844 267384 153896 267436
rect 184480 267384 184532 267436
rect 190552 267384 190604 267436
rect 104808 267248 104860 267300
rect 164608 267248 164660 267300
rect 79324 267112 79376 267164
rect 140596 267112 140648 267164
rect 145564 267112 145616 267164
rect 191932 267248 191984 267300
rect 195244 267384 195296 267436
rect 219256 267384 219308 267436
rect 223488 267384 223540 267436
rect 234160 267384 234212 267436
rect 243728 267384 243780 267436
rect 251548 267384 251600 267436
rect 315304 267384 315356 267436
rect 319076 267384 319128 267436
rect 340972 267384 341024 267436
rect 355324 267384 355376 267436
rect 371608 267384 371660 267436
rect 373264 267384 373316 267436
rect 380716 267384 380768 267436
rect 397920 267384 397972 267436
rect 404728 267384 404780 267436
rect 416228 267384 416280 267436
rect 421288 267384 421340 267436
rect 440884 267384 440936 267436
rect 447784 267384 447836 267436
rect 456064 267384 456116 267436
rect 460204 267384 460256 267436
rect 516784 267384 516836 267436
rect 519820 267384 519872 267436
rect 583024 267384 583076 267436
rect 224224 267248 224276 267300
rect 233884 267248 233936 267300
rect 244096 267248 244148 267300
rect 249064 267248 249116 267300
rect 250720 267248 250772 267300
rect 321928 267248 321980 267300
rect 327724 267248 327776 267300
rect 350908 267248 350960 267300
rect 362224 267248 362276 267300
rect 373264 267248 373316 267300
rect 392032 267248 392084 267300
rect 398104 267248 398156 267300
rect 417424 267248 417476 267300
rect 432880 267248 432932 267300
rect 453304 267248 453356 267300
rect 459376 267248 459428 267300
rect 460848 267248 460900 267300
rect 465172 267248 465224 267300
rect 523684 267248 523736 267300
rect 524788 267248 524840 267300
rect 612004 267248 612056 267300
rect 199384 267112 199436 267164
rect 204352 267112 204404 267164
rect 205456 267112 205508 267164
rect 218428 267112 218480 267164
rect 220084 267112 220136 267164
rect 239128 267112 239180 267164
rect 246948 267112 247000 267164
rect 263968 267112 264020 267164
rect 313648 267112 313700 267164
rect 317420 267112 317472 267164
rect 365812 267112 365864 267164
rect 381544 267112 381596 267164
rect 383200 267112 383252 267164
rect 401692 267112 401744 267164
rect 413008 267112 413060 267164
rect 441620 267112 441672 267164
rect 455144 267112 455196 267164
rect 515404 267112 515456 267164
rect 517244 267112 517296 267164
rect 527180 267112 527232 267164
rect 529664 267112 529716 267164
rect 617524 267112 617576 267164
rect 90364 266976 90416 267028
rect 151360 266976 151412 267028
rect 159456 266976 159508 267028
rect 162124 266976 162176 267028
rect 168104 266976 168156 267028
rect 177028 266976 177080 267028
rect 177672 266976 177724 267028
rect 214288 266976 214340 267028
rect 218704 266976 218756 267028
rect 220912 266976 220964 267028
rect 228364 266976 228416 267028
rect 249064 266976 249116 267028
rect 255964 266976 256016 267028
rect 259000 266976 259052 267028
rect 286324 266976 286376 267028
rect 287980 266976 288032 267028
rect 312820 266976 312872 267028
rect 316040 266976 316092 267028
rect 317788 266976 317840 267028
rect 322940 266976 322992 267028
rect 393136 266976 393188 267028
rect 420184 266976 420236 267028
rect 434352 266976 434404 267028
rect 457444 266976 457496 267028
rect 469312 266976 469364 267028
rect 470416 266976 470468 267028
rect 470600 266976 470652 267028
rect 534724 266976 534776 267028
rect 535552 266976 535604 267028
rect 536748 266976 536800 267028
rect 539692 266976 539744 267028
rect 634084 266976 634136 267028
rect 119344 266840 119396 266892
rect 153844 266840 153896 266892
rect 169024 266840 169076 266892
rect 199384 266840 199436 266892
rect 216128 266840 216180 266892
rect 222568 266840 222620 266892
rect 314476 266840 314528 266892
rect 319260 266840 319312 266892
rect 332692 266840 332744 266892
rect 343824 266840 343876 266892
rect 362500 266840 362552 266892
rect 368940 266840 368992 266892
rect 390652 266840 390704 266892
rect 408316 266840 408368 266892
rect 422944 266840 422996 266892
rect 438124 266840 438176 266892
rect 442724 266840 442776 266892
rect 137468 266704 137520 266756
rect 150532 266704 150584 266756
rect 151084 266704 151136 266756
rect 179512 266704 179564 266756
rect 347504 266704 347556 266756
rect 351184 266704 351236 266756
rect 360016 266704 360068 266756
rect 366364 266704 366416 266756
rect 388168 266704 388220 266756
rect 404360 266704 404412 266756
rect 407212 266704 407264 266756
rect 414480 266704 414532 266756
rect 434536 266704 434588 266756
rect 449164 266704 449216 266756
rect 457720 266704 457772 266756
rect 476764 266704 476816 266756
rect 308680 266636 308732 266688
rect 310612 266636 310664 266688
rect 316960 266636 317012 266688
rect 321560 266636 321612 266688
rect 427912 266636 427964 266688
rect 434352 266636 434404 266688
rect 132500 266568 132552 266620
rect 147220 266568 147272 266620
rect 149980 266568 150032 266620
rect 159640 266568 159692 266620
rect 345112 266568 345164 266620
rect 348424 266568 348476 266620
rect 399760 266568 399812 266620
rect 407764 266568 407816 266620
rect 437848 266568 437900 266620
rect 448428 266568 448480 266620
rect 499948 266840 500000 266892
rect 507860 266840 507912 266892
rect 534724 266840 534776 266892
rect 589924 266840 589976 266892
rect 490012 266704 490064 266756
rect 509700 266704 509752 266756
rect 510712 266704 510764 266756
rect 511632 266704 511684 266756
rect 512368 266704 512420 266756
rect 513196 266704 513248 266756
rect 516508 266704 516560 266756
rect 517428 266704 517480 266756
rect 518992 266704 519044 266756
rect 520096 266704 520148 266756
rect 527272 266704 527324 266756
rect 528192 266704 528244 266756
rect 528928 266704 528980 266756
rect 529848 266704 529900 266756
rect 531412 266704 531464 266756
rect 532608 266704 532660 266756
rect 533068 266704 533120 266756
rect 533988 266704 534040 266756
rect 543004 266704 543056 266756
rect 598204 266704 598256 266756
rect 482284 266568 482336 266620
rect 482560 266568 482612 266620
rect 485044 266568 485096 266620
rect 504824 266568 504876 266620
rect 556804 266568 556856 266620
rect 310336 266500 310388 266552
rect 311900 266500 311952 266552
rect 312360 266500 312412 266552
rect 314660 266500 314712 266552
rect 316132 266500 316184 266552
rect 320180 266500 320232 266552
rect 327724 266500 327776 266552
rect 331956 266500 332008 266552
rect 350080 266500 350132 266552
rect 353944 266500 353996 266552
rect 355876 266500 355928 266552
rect 360844 266500 360896 266552
rect 369952 266500 370004 266552
rect 372252 266500 372304 266552
rect 374920 266500 374972 266552
rect 380532 266500 380584 266552
rect 423772 266500 423824 266552
rect 425704 266500 425756 266552
rect 426256 266500 426308 266552
rect 428464 266500 428516 266552
rect 452752 266500 452804 266552
rect 462964 266500 463016 266552
rect 475108 266500 475160 266552
rect 479524 266500 479576 266552
rect 342628 266432 342680 266484
rect 345296 266432 345348 266484
rect 163504 266364 163556 266416
rect 167092 266364 167144 266416
rect 211160 266364 211212 266416
rect 213460 266364 213512 266416
rect 214564 266364 214616 266416
rect 215944 266364 215996 266416
rect 239404 266364 239456 266416
rect 241612 266364 241664 266416
rect 243544 266364 243596 266416
rect 246580 266364 246632 266416
rect 250444 266364 250496 266416
rect 256516 266364 256568 266416
rect 300952 266364 301004 266416
rect 302056 266364 302108 266416
rect 303712 266364 303764 266416
rect 304540 266364 304592 266416
rect 307852 266364 307904 266416
rect 309140 266364 309192 266416
rect 309508 266364 309560 266416
rect 310980 266364 311032 266416
rect 311164 266364 311216 266416
rect 313280 266364 313332 266416
rect 320272 266364 320324 266416
rect 321376 266364 321428 266416
rect 324412 266364 324464 266416
rect 325332 266364 325384 266416
rect 328552 266364 328604 266416
rect 329748 266364 329800 266416
rect 336832 266364 336884 266416
rect 337936 266364 337988 266416
rect 346768 266364 346820 266416
rect 347688 266364 347740 266416
rect 349252 266364 349304 266416
rect 350356 266364 350408 266416
rect 357532 266364 357584 266416
rect 359464 266364 359516 266416
rect 361672 266364 361724 266416
rect 362776 266364 362828 266416
rect 369124 266364 369176 266416
rect 370504 266364 370556 266416
rect 374092 266364 374144 266416
rect 375288 266364 375340 266416
rect 379888 266364 379940 266416
rect 383016 266364 383068 266416
rect 384028 266364 384080 266416
rect 384948 266364 385000 266416
rect 386512 266364 386564 266416
rect 387708 266364 387760 266416
rect 392308 266364 392360 266416
rect 393320 266364 393372 266416
rect 394792 266364 394844 266416
rect 398932 266364 398984 266416
rect 400036 266364 400088 266416
rect 403624 266432 403676 266484
rect 483388 266432 483440 266484
rect 484216 266432 484268 266484
rect 485872 266432 485924 266484
rect 486792 266432 486844 266484
rect 491668 266432 491720 266484
rect 492404 266432 492456 266484
rect 494152 266432 494204 266484
rect 495256 266432 495308 266484
rect 502432 266432 502484 266484
rect 503536 266432 503588 266484
rect 504088 266432 504140 266484
rect 505008 266432 505060 266484
rect 506572 266432 506624 266484
rect 507676 266432 507728 266484
rect 507860 266432 507912 266484
rect 551284 266432 551336 266484
rect 408868 266364 408920 266416
rect 409788 266364 409840 266416
rect 411352 266364 411404 266416
rect 412272 266364 412324 266416
rect 415492 266364 415544 266416
rect 416412 266364 416464 266416
rect 417976 266364 418028 266416
rect 418804 266364 418856 266416
rect 425428 266364 425480 266416
rect 427084 266364 427136 266416
rect 429568 266364 429620 266416
rect 430396 266364 430448 266416
rect 432052 266364 432104 266416
rect 433156 266364 433208 266416
rect 440332 266364 440384 266416
rect 441344 266364 441396 266416
rect 441988 266364 442040 266416
rect 442908 266364 442960 266416
rect 444472 266364 444524 266416
rect 445668 266364 445720 266416
rect 448612 266364 448664 266416
rect 450544 266364 450596 266416
rect 454408 266364 454460 266416
rect 455328 266364 455380 266416
rect 473452 266364 473504 266416
rect 474648 266364 474700 266416
rect 477592 266364 477644 266416
rect 478512 266364 478564 266416
rect 480076 266296 480128 266348
rect 554780 266296 554832 266348
rect 487528 266160 487580 266212
rect 565820 266160 565872 266212
rect 511540 266024 511592 266076
rect 599124 266024 599176 266076
rect 513196 265888 513248 265940
rect 601700 265888 601752 265940
rect 515680 265752 515732 265804
rect 605840 265752 605892 265804
rect 189080 265616 189132 265668
rect 189908 265616 189960 265668
rect 209780 265616 209832 265668
rect 210700 265616 210752 265668
rect 224960 265616 225012 265668
rect 225604 265616 225656 265668
rect 280344 265616 280396 265668
rect 280988 265616 281040 265668
rect 292672 265616 292724 265668
rect 293500 265616 293552 265668
rect 296812 265616 296864 265668
rect 297548 265616 297600 265668
rect 518164 265616 518216 265668
rect 608600 265616 608652 265668
rect 481732 265480 481784 265532
rect 557540 265480 557592 265532
rect 476764 265344 476816 265396
rect 549444 265344 549496 265396
rect 471796 265208 471848 265260
rect 542360 265208 542412 265260
rect 466828 265072 466880 265124
rect 535736 265072 535788 265124
rect 570604 261468 570656 261520
rect 645860 261468 645912 261520
rect 554412 260856 554464 260908
rect 568580 260856 568632 260908
rect 554320 259428 554372 259480
rect 560944 259428 560996 259480
rect 675852 259428 675904 259480
rect 676404 259428 676456 259480
rect 35808 256708 35860 256760
rect 40684 256708 40736 256760
rect 553952 256708 554004 256760
rect 563704 256708 563756 256760
rect 553492 255552 553544 255604
rect 555424 255552 555476 255604
rect 35808 255416 35860 255468
rect 39396 255416 39448 255468
rect 35808 254192 35860 254244
rect 39396 254192 39448 254244
rect 42064 253988 42116 254040
rect 43168 253988 43220 254040
rect 35532 253920 35584 253972
rect 41696 253920 41748 253972
rect 35808 252764 35860 252816
rect 41696 252696 41748 252748
rect 42064 252696 42116 252748
rect 42708 252696 42760 252748
rect 35808 252560 35860 252612
rect 41696 252560 41748 252612
rect 554412 252560 554464 252612
rect 562324 252560 562376 252612
rect 675852 252492 675904 252544
rect 679624 252492 679676 252544
rect 675484 251336 675536 251388
rect 554136 251200 554188 251252
rect 556804 251200 556856 251252
rect 675484 250724 675536 250776
rect 674840 250588 674892 250640
rect 675300 250588 675352 250640
rect 35808 249908 35860 249960
rect 39580 249908 39632 249960
rect 35808 248480 35860 248532
rect 40316 248480 40368 248532
rect 35808 247188 35860 247240
rect 40960 247188 41012 247240
rect 35808 247052 35860 247104
rect 39396 247052 39448 247104
rect 558184 246304 558236 246356
rect 647240 246304 647292 246356
rect 553860 245624 553912 245676
rect 596824 245624 596876 245676
rect 554504 244264 554556 244316
rect 573364 244264 573416 244316
rect 674472 243652 674524 243704
rect 675208 243652 675260 243704
rect 674380 242836 674432 242888
rect 675208 242836 675260 242888
rect 576124 242156 576176 242208
rect 648620 242156 648672 242208
rect 553676 241476 553728 241528
rect 629944 241476 629996 241528
rect 554504 240116 554556 240168
rect 577504 240116 577556 240168
rect 554320 238688 554372 238740
rect 576124 238688 576176 238740
rect 672080 236988 672132 237040
rect 671896 236852 671948 236904
rect 672954 236716 673006 236768
rect 673184 236444 673236 236496
rect 673092 236172 673144 236224
rect 554504 236036 554556 236088
rect 558184 236036 558236 236088
rect 671068 235900 671120 235952
rect 671252 235764 671304 235816
rect 669320 235560 669372 235612
rect 670884 235424 670936 235476
rect 669780 235084 669832 235136
rect 672080 234812 672132 234864
rect 554412 234540 554464 234592
rect 570604 234540 570656 234592
rect 668216 234540 668268 234592
rect 668032 234404 668084 234456
rect 670332 234132 670384 234184
rect 42248 233928 42300 233980
rect 43260 233928 43312 233980
rect 675852 233928 675904 233980
rect 683304 233996 683356 234048
rect 652392 233860 652444 233912
rect 675484 233860 675536 233912
rect 675852 233724 675904 233776
rect 678244 233724 678296 233776
rect 669596 233180 669648 233232
rect 672080 233180 672132 233232
rect 663064 232636 663116 232688
rect 675484 232704 675536 232756
rect 675852 232636 675904 232688
rect 683672 232636 683724 232688
rect 652208 232500 652260 232552
rect 675484 232364 675536 232416
rect 675852 232364 675904 232416
rect 679256 232364 679308 232416
rect 137928 231752 137980 231804
rect 152372 231752 152424 231804
rect 91744 231616 91796 231668
rect 168564 231616 168616 231668
rect 662328 231616 662380 231668
rect 668400 231616 668452 231668
rect 669136 231616 669188 231668
rect 675392 231616 675444 231668
rect 128268 231480 128320 231532
rect 195888 231480 195940 231532
rect 596824 231480 596876 231532
rect 633624 231480 633676 231532
rect 664996 231480 665048 231532
rect 57244 231344 57296 231396
rect 669136 231344 669188 231396
rect 64144 231208 64196 231260
rect 667204 231208 667256 231260
rect 58624 231072 58676 231124
rect 674932 231072 674984 231124
rect 668400 230936 668452 230988
rect 97908 230868 97960 230920
rect 173992 230868 174044 230920
rect 668400 230800 668452 230852
rect 668952 230800 669004 230852
rect 672080 230800 672132 230852
rect 110328 230732 110380 230784
rect 184296 230732 184348 230784
rect 118608 230596 118660 230648
rect 188160 230596 188212 230648
rect 195060 230596 195112 230648
rect 196900 230596 196952 230648
rect 665824 230596 665876 230648
rect 439320 230528 439372 230580
rect 152372 230460 152424 230512
rect 203616 230460 203668 230512
rect 130384 230392 130436 230444
rect 142620 230392 142672 230444
rect 142804 230392 142856 230444
rect 150808 230392 150860 230444
rect 206284 230392 206336 230444
rect 256424 230392 256476 230444
rect 276296 230392 276348 230444
rect 292488 230392 292540 230444
rect 308404 230392 308456 230444
rect 334992 230392 335044 230444
rect 440700 230392 440752 230444
rect 441896 230392 441948 230444
rect 443460 230392 443512 230444
rect 526904 230392 526956 230444
rect 536104 230392 536156 230444
rect 673460 230392 673512 230444
rect 42156 230324 42208 230376
rect 43076 230324 43128 230376
rect 387432 230324 387484 230376
rect 388444 230324 388496 230376
rect 398104 230324 398156 230376
rect 399392 230324 399444 230376
rect 438676 230324 438728 230376
rect 439320 230324 439372 230376
rect 443828 230324 443880 230376
rect 444840 230324 444892 230376
rect 449624 230324 449676 230376
rect 450544 230324 450596 230376
rect 452844 230324 452896 230376
rect 454316 230324 454368 230376
rect 455420 230324 455472 230376
rect 457168 230324 457220 230376
rect 463792 230324 463844 230376
rect 465724 230324 465776 230376
rect 470876 230324 470928 230376
rect 471888 230324 471940 230376
rect 472164 230324 472216 230376
rect 473176 230324 473228 230376
rect 487620 230324 487672 230376
rect 488448 230324 488500 230376
rect 493416 230324 493468 230376
rect 496360 230324 496412 230376
rect 497280 230324 497332 230376
rect 498108 230324 498160 230376
rect 510804 230324 510856 230376
rect 511908 230324 511960 230376
rect 133788 230256 133840 230308
rect 202328 230256 202380 230308
rect 210424 230256 210476 230308
rect 261576 230256 261628 230308
rect 275652 230256 275704 230308
rect 313096 230256 313148 230308
rect 436100 230256 436152 230308
rect 436836 230256 436888 230308
rect 528836 230256 528888 230308
rect 539600 230256 539652 230308
rect 388444 230188 388496 230240
rect 391664 230188 391716 230240
rect 444472 230188 444524 230240
rect 447600 230188 447652 230240
rect 451556 230188 451608 230240
rect 453304 230188 453356 230240
rect 453488 230188 453540 230240
rect 455788 230188 455840 230240
rect 468300 230188 468352 230240
rect 469128 230188 469180 230240
rect 490196 230188 490248 230240
rect 493784 230188 493836 230240
rect 511448 230188 511500 230240
rect 517520 230188 517572 230240
rect 674288 230188 674340 230240
rect 95240 230120 95292 230172
rect 157294 230120 157346 230172
rect 157432 230120 157484 230172
rect 161112 230120 161164 230172
rect 176752 230120 176804 230172
rect 235816 230120 235868 230172
rect 264244 230120 264296 230172
rect 302792 230120 302844 230172
rect 302976 230120 303028 230172
rect 329840 230120 329892 230172
rect 334256 230120 334308 230172
rect 355600 230120 355652 230172
rect 521108 230120 521160 230172
rect 529204 230120 529256 230172
rect 532700 230120 532752 230172
rect 547144 230120 547196 230172
rect 454132 230052 454184 230104
rect 455328 230052 455380 230104
rect 491484 230052 491536 230104
rect 492496 230052 492548 230104
rect 126888 229984 126940 230036
rect 195060 229984 195112 230036
rect 195428 229984 195480 230036
rect 214748 229984 214800 230036
rect 219992 229984 220044 230036
rect 230664 229984 230716 230036
rect 242532 229984 242584 230036
rect 287336 229984 287388 230036
rect 287520 229984 287572 230036
rect 307944 229984 307996 230036
rect 312636 229984 312688 230036
rect 340144 229984 340196 230036
rect 354956 229984 355008 230036
rect 371056 229984 371108 230036
rect 457352 229984 457404 230036
rect 463884 229984 463936 230036
rect 515312 229984 515364 230036
rect 524604 229984 524656 230036
rect 534632 229984 534684 230036
rect 549260 229984 549312 230036
rect 674104 229984 674156 230036
rect 86224 229848 86276 229900
rect 156696 229848 156748 229900
rect 68284 229712 68336 229764
rect 142804 229712 142856 229764
rect 142988 229712 143040 229764
rect 145656 229712 145708 229764
rect 145840 229712 145892 229764
rect 158536 229848 158588 229900
rect 158720 229848 158772 229900
rect 163688 229848 163740 229900
rect 163964 229848 164016 229900
rect 225512 229848 225564 229900
rect 230480 229848 230532 229900
rect 277032 229848 277084 229900
rect 282552 229848 282604 229900
rect 318248 229848 318300 229900
rect 324228 229848 324280 229900
rect 350448 229848 350500 229900
rect 366732 229848 366784 229900
rect 383936 229848 383988 229900
rect 467012 229848 467064 229900
rect 474004 229848 474056 229900
rect 476672 229848 476724 229900
rect 481640 229848 481692 229900
rect 481824 229848 481876 229900
rect 489920 229848 489972 229900
rect 495992 229848 496044 229900
rect 507124 229848 507176 229900
rect 509516 229848 509568 229900
rect 515404 229848 515456 229900
rect 517244 229848 517296 229900
rect 526444 229848 526496 229900
rect 536564 229848 536616 229900
rect 559564 229848 559616 229900
rect 433524 229780 433576 229832
rect 434168 229780 434220 229832
rect 157294 229712 157346 229764
rect 166264 229712 166316 229764
rect 171048 229712 171100 229764
rect 219992 229712 220044 229764
rect 82084 229576 82136 229628
rect 102140 229440 102192 229492
rect 139860 229440 139912 229492
rect 149060 229576 149112 229628
rect 153384 229576 153436 229628
rect 153844 229576 153896 229628
rect 157708 229576 157760 229628
rect 157984 229576 158036 229628
rect 111064 229304 111116 229356
rect 140320 229304 140372 229356
rect 142988 229304 143040 229356
rect 144184 229304 144236 229356
rect 146944 229304 146996 229356
rect 149612 229440 149664 229492
rect 149980 229440 150032 229492
rect 210056 229440 210108 229492
rect 214748 229576 214800 229628
rect 246120 229712 246172 229764
rect 256516 229712 256568 229764
rect 297640 229712 297692 229764
rect 318064 229712 318116 229764
rect 220360 229440 220412 229492
rect 220728 229440 220780 229492
rect 266728 229576 266780 229628
rect 296996 229576 297048 229628
rect 323400 229576 323452 229628
rect 345020 229712 345072 229764
rect 360752 229712 360804 229764
rect 361212 229712 361264 229764
rect 378784 229712 378836 229764
rect 391204 229712 391256 229764
rect 398748 229712 398800 229764
rect 399852 229712 399904 229764
rect 409696 229712 409748 229764
rect 410892 229712 410944 229764
rect 417424 229712 417476 229764
rect 465448 229712 465500 229764
rect 467472 229712 467524 229764
rect 469588 229712 469640 229764
rect 476764 229712 476816 229764
rect 479248 229712 479300 229764
rect 488080 229712 488132 229764
rect 492128 229712 492180 229764
rect 505100 229712 505152 229764
rect 507584 229712 507636 229764
rect 516784 229712 516836 229764
rect 523040 229712 523092 229764
rect 534816 229712 534868 229764
rect 538496 229712 538548 229764
rect 566464 229712 566516 229764
rect 660948 229712 661000 229764
rect 672080 229712 672132 229764
rect 674452 229916 674504 229968
rect 674334 229780 674386 229832
rect 345296 229576 345348 229628
rect 530124 229576 530176 229628
rect 531136 229576 531188 229628
rect 384304 229508 384356 229560
rect 389088 229508 389140 229560
rect 448980 229508 449032 229560
rect 451924 229508 451976 229560
rect 231124 229440 231176 229492
rect 271880 229440 271932 229492
rect 476028 229440 476080 229492
rect 478604 229440 478656 229492
rect 530768 229440 530820 229492
rect 538312 229576 538364 229628
rect 446404 229372 446456 229424
rect 448796 229372 448848 229424
rect 450912 229372 450964 229424
rect 453028 229372 453080 229424
rect 505652 229372 505704 229424
rect 510988 229372 511040 229424
rect 674242 229508 674294 229560
rect 147864 229304 147916 229356
rect 151176 229304 151228 229356
rect 123484 229168 123536 229220
rect 149060 229168 149112 229220
rect 149612 229168 149664 229220
rect 155960 229168 156012 229220
rect 156328 229304 156380 229356
rect 215208 229304 215260 229356
rect 246488 229304 246540 229356
rect 282184 229304 282236 229356
rect 413836 229304 413888 229356
rect 420000 229304 420052 229356
rect 450268 229236 450320 229288
rect 451740 229236 451792 229288
rect 488264 229236 488316 229288
rect 490380 229236 490432 229288
rect 495348 229236 495400 229288
rect 500224 229236 500276 229288
rect 513380 229236 513432 229288
rect 519360 229236 519412 229288
rect 161756 229168 161808 229220
rect 164608 229168 164660 229220
rect 174268 229168 174320 229220
rect 184664 229168 184716 229220
rect 240968 229168 241020 229220
rect 423496 229100 423548 229152
rect 427728 229100 427780 229152
rect 441252 229100 441304 229152
rect 442080 229100 442132 229152
rect 503720 229100 503772 229152
rect 509884 229100 509936 229152
rect 519176 229100 519228 229152
rect 100668 229032 100720 229084
rect 106188 229032 106240 229084
rect 142988 229032 143040 229084
rect 143448 229032 143500 229084
rect 147128 229032 147180 229084
rect 147312 229032 147364 229084
rect 202880 229032 202932 229084
rect 204720 229032 204772 229084
rect 212356 229032 212408 229084
rect 214380 229032 214432 229084
rect 257068 229032 257120 229084
rect 257528 229032 257580 229084
rect 296352 229032 296404 229084
rect 302148 229032 302200 229084
rect 331128 229032 331180 229084
rect 524972 229100 525024 229152
rect 529940 229100 529992 229152
rect 673736 229100 673788 229152
rect 164608 228896 164660 228948
rect 167368 228896 167420 228948
rect 169484 228896 169536 228948
rect 179788 228896 179840 228948
rect 180156 228896 180208 228948
rect 93768 228760 93820 228812
rect 166816 228760 166868 228812
rect 166954 228760 167006 228812
rect 174820 228760 174872 228812
rect 219808 228760 219860 228812
rect 220360 228896 220412 228948
rect 246764 228896 246816 228948
rect 257712 228896 257764 228948
rect 299572 228896 299624 228948
rect 300676 228896 300728 228948
rect 330484 228896 330536 228948
rect 226156 228760 226208 228812
rect 238576 228760 238628 228812
rect 282828 228760 282880 228812
rect 296628 228760 296680 228812
rect 329196 228760 329248 228812
rect 336464 228760 336516 228812
rect 358820 228760 358872 228812
rect 359924 228760 359976 228812
rect 376852 228760 376904 228812
rect 478880 228760 478932 228812
rect 490196 228760 490248 228812
rect 499856 228760 499908 228812
rect 517704 228896 517756 228948
rect 543188 228896 543240 228948
rect 67548 228624 67600 228676
rect 61660 228488 61712 228540
rect 142436 228488 142488 228540
rect 57244 228352 57296 228404
rect 141148 228352 141200 228404
rect 142988 228624 143040 228676
rect 152464 228624 152516 228676
rect 153108 228624 153160 228676
rect 146116 228488 146168 228540
rect 210700 228488 210752 228540
rect 212356 228624 212408 228676
rect 220360 228624 220412 228676
rect 220544 228624 220596 228676
rect 264796 228624 264848 228676
rect 285496 228624 285548 228676
rect 318892 228624 318944 228676
rect 325516 228624 325568 228676
rect 349160 228624 349212 228676
rect 350172 228624 350224 228676
rect 369124 228624 369176 228676
rect 377772 228624 377824 228676
rect 390376 228624 390428 228676
rect 498568 228624 498620 228676
rect 515772 228760 515824 228812
rect 518532 228760 518584 228812
rect 541624 228760 541676 228812
rect 512092 228624 512144 228676
rect 215852 228488 215904 228540
rect 216220 228488 216272 228540
rect 219624 228488 219676 228540
rect 219992 228488 220044 228540
rect 260288 228488 260340 228540
rect 268936 228488 268988 228540
rect 306012 228488 306064 228540
rect 313924 228488 313976 228540
rect 320824 228488 320876 228540
rect 326896 228488 326948 228540
rect 351092 228488 351144 228540
rect 354588 228488 354640 228540
rect 372344 228488 372396 228540
rect 373448 228488 373500 228540
rect 387156 228488 387208 228540
rect 390468 228488 390520 228540
rect 400036 228488 400088 228540
rect 148876 228352 148928 228404
rect 152464 228352 152516 228404
rect 166816 228352 166868 228404
rect 166954 228352 167006 228404
rect 214564 228352 214616 228404
rect 217508 228352 217560 228404
rect 221464 228352 221516 228404
rect 224592 228352 224644 228404
rect 273812 228352 273864 228404
rect 274272 228352 274324 228404
rect 312452 228352 312504 228404
rect 320088 228352 320140 228404
rect 346860 228352 346912 228404
rect 347044 228352 347096 228404
rect 365904 228352 365956 228404
rect 371148 228352 371200 228404
rect 385224 228352 385276 228404
rect 386236 228352 386288 228404
rect 397460 228352 397512 228404
rect 112812 228216 112864 228268
rect 184940 228216 184992 228268
rect 189724 228216 189776 228268
rect 239036 228216 239088 228268
rect 254952 228216 255004 228268
rect 295708 228216 295760 228268
rect 407764 228488 407816 228540
rect 409788 228488 409840 228540
rect 415492 228488 415544 228540
rect 485688 228488 485740 228540
rect 498292 228488 498344 228540
rect 502432 228488 502484 228540
rect 402796 228352 402848 228404
rect 411628 228352 411680 228404
rect 474464 228352 474516 228404
rect 484584 228352 484636 228404
rect 485044 228352 485096 228404
rect 498568 228352 498620 228404
rect 507124 228352 507176 228404
rect 512736 228352 512788 228404
rect 517888 228624 517940 228676
rect 539416 228624 539468 228676
rect 539600 228624 539652 228676
rect 555976 228624 556028 228676
rect 527548 228488 527600 228540
rect 553308 228488 553360 228540
rect 555424 228488 555476 228540
rect 571340 228488 571392 228540
rect 533344 228352 533396 228404
rect 537208 228352 537260 228404
rect 565636 228352 565688 228404
rect 520924 228216 520976 228268
rect 539416 228216 539468 228268
rect 540796 228216 540848 228268
rect 119988 228080 120040 228132
rect 190092 228080 190144 228132
rect 193036 228080 193088 228132
rect 204720 228080 204772 228132
rect 214564 228080 214616 228132
rect 126704 227944 126756 227996
rect 195244 227944 195296 227996
rect 205456 227944 205508 227996
rect 214380 227944 214432 227996
rect 219808 228080 219860 228132
rect 231308 228080 231360 228132
rect 233884 228080 233936 228132
rect 272524 228080 272576 228132
rect 400128 228080 400180 228132
rect 415032 228012 415084 228064
rect 421932 228012 421984 228064
rect 221004 227944 221056 227996
rect 221464 227944 221516 227996
rect 251272 227944 251324 227996
rect 416688 227876 416740 227928
rect 420644 227876 420696 227928
rect 447048 227876 447100 227928
rect 450544 227876 450596 227928
rect 88248 227808 88300 227860
rect 95240 227808 95292 227860
rect 133512 227808 133564 227860
rect 200396 227808 200448 227860
rect 203524 227808 203576 227860
rect 64788 227672 64840 227724
rect 111064 227672 111116 227724
rect 117228 227672 117280 227724
rect 110144 227536 110196 227588
rect 182364 227536 182416 227588
rect 185400 227672 185452 227724
rect 192668 227672 192720 227724
rect 200028 227672 200080 227724
rect 204904 227672 204956 227724
rect 210976 227808 211028 227860
rect 219992 227808 220044 227860
rect 226156 227808 226208 227860
rect 233884 227808 233936 227860
rect 239312 227808 239364 227860
rect 243544 227808 243596 227860
rect 246304 227808 246356 227860
rect 248696 227808 248748 227860
rect 249064 227808 249116 227860
rect 253848 227808 253900 227860
rect 331036 227740 331088 227792
rect 334256 227740 334308 227792
rect 351092 227740 351144 227792
rect 353024 227740 353076 227792
rect 371792 227740 371844 227792
rect 373632 227740 373684 227792
rect 409052 227740 409104 227792
rect 410340 227740 410392 227792
rect 411904 227740 411956 227792
rect 413560 227740 413612 227792
rect 420644 227740 420696 227792
rect 423864 227740 423916 227792
rect 471520 227740 471572 227792
rect 479524 227740 479576 227792
rect 489920 227740 489972 227792
rect 494704 227740 494756 227792
rect 664904 227740 664956 227792
rect 665272 227740 665324 227792
rect 669136 227740 669188 227792
rect 673644 227740 673696 227792
rect 217784 227672 217836 227724
rect 219808 227672 219860 227724
rect 228732 227672 228784 227724
rect 228916 227672 228968 227724
rect 268016 227672 268068 227724
rect 293776 227672 293828 227724
rect 325332 227672 325384 227724
rect 465908 227604 465960 227656
rect 469864 227604 469916 227656
rect 187516 227536 187568 227588
rect 60648 227400 60700 227452
rect 102140 227400 102192 227452
rect 103428 227400 103480 227452
rect 171232 227400 171284 227452
rect 172152 227400 172204 227452
rect 177212 227400 177264 227452
rect 181352 227400 181404 227452
rect 96436 227264 96488 227316
rect 89628 227128 89680 227180
rect 156696 227128 156748 227180
rect 169484 227264 169536 227316
rect 160192 227128 160244 227180
rect 185584 227264 185636 227316
rect 186136 227400 186188 227452
rect 214748 227536 214800 227588
rect 214932 227536 214984 227588
rect 262220 227536 262272 227588
rect 281356 227536 281408 227588
rect 317604 227536 317656 227588
rect 337752 227536 337804 227588
rect 345020 227536 345072 227588
rect 524604 227536 524656 227588
rect 537484 227536 537536 227588
rect 189908 227400 189960 227452
rect 204720 227400 204772 227452
rect 204904 227400 204956 227452
rect 251916 227400 251968 227452
rect 264796 227400 264848 227452
rect 304724 227400 304776 227452
rect 315488 227400 315540 227452
rect 341432 227400 341484 227452
rect 352564 227400 352616 227452
rect 363328 227400 363380 227452
rect 495072 227400 495124 227452
rect 511172 227400 511224 227452
rect 514024 227400 514076 227452
rect 535736 227400 535788 227452
rect 536104 227400 536156 227452
rect 552480 227400 552532 227452
rect 219532 227264 219584 227316
rect 219992 227264 220044 227316
rect 241612 227264 241664 227316
rect 249432 227264 249484 227316
rect 290556 227264 290608 227316
rect 291016 227264 291068 227316
rect 322112 227264 322164 227316
rect 322296 227264 322348 227316
rect 332416 227264 332468 227316
rect 333888 227264 333940 227316
rect 356244 227264 356296 227316
rect 357256 227264 357308 227316
rect 374276 227264 374328 227316
rect 382096 227264 382148 227316
rect 392952 227264 393004 227316
rect 171600 227128 171652 227180
rect 219808 227128 219860 227180
rect 56508 226992 56560 227044
rect 142160 226992 142212 227044
rect 143264 226992 143316 227044
rect 204076 226992 204128 227044
rect 122748 226856 122800 226908
rect 185400 226856 185452 226908
rect 185584 226856 185636 226908
rect 214104 226992 214156 227044
rect 233700 227128 233752 227180
rect 241152 227128 241204 227180
rect 286692 227128 286744 227180
rect 306196 227128 306248 227180
rect 336924 227128 336976 227180
rect 340696 227128 340748 227180
rect 361396 227128 361448 227180
rect 363512 227128 363564 227180
rect 368480 227128 368532 227180
rect 376668 227128 376720 227180
rect 389732 227128 389784 227180
rect 393136 227128 393188 227180
rect 402612 227264 402664 227316
rect 510988 227264 511040 227316
rect 524420 227264 524472 227316
rect 526260 227264 526312 227316
rect 551560 227264 551612 227316
rect 402244 227128 402296 227180
rect 408408 227128 408460 227180
rect 478604 227128 478656 227180
rect 486792 227128 486844 227180
rect 490380 227128 490432 227180
rect 503168 227128 503220 227180
rect 504916 227128 504968 227180
rect 523040 227128 523092 227180
rect 523684 227128 523736 227180
rect 548524 227128 548576 227180
rect 556804 227128 556856 227180
rect 570604 227128 570656 227180
rect 221832 226992 221884 227044
rect 271236 226992 271288 227044
rect 271788 226992 271840 227044
rect 308588 226992 308640 227044
rect 310336 226992 310388 227044
rect 338212 226992 338264 227044
rect 338672 226992 338724 227044
rect 360108 226992 360160 227044
rect 362776 226992 362828 227044
rect 379060 226992 379112 227044
rect 391756 226992 391808 227044
rect 403532 226992 403584 227044
rect 412548 226992 412600 227044
rect 419356 226992 419408 227044
rect 486976 226992 487028 227044
rect 500960 226992 501012 227044
rect 506296 226992 506348 227044
rect 526628 226992 526680 227044
rect 533712 226992 533764 227044
rect 560760 226992 560812 227044
rect 652024 226992 652076 227044
rect 129556 226720 129608 226772
rect 197452 226720 197504 226772
rect 204720 226720 204772 226772
rect 214748 226856 214800 226908
rect 219992 226856 220044 226908
rect 214104 226720 214156 226772
rect 218428 226720 218480 226772
rect 219348 226720 219400 226772
rect 267372 226856 267424 226908
rect 378784 226788 378836 226840
rect 385868 226788 385920 226840
rect 668952 226992 669004 227044
rect 673460 226992 673512 227044
rect 673552 226788 673604 226840
rect 676036 226788 676088 226840
rect 678244 226788 678296 226840
rect 235816 226720 235868 226772
rect 280252 226720 280304 226772
rect 136548 226584 136600 226636
rect 203156 226584 203208 226636
rect 204076 226584 204128 226636
rect 208124 226584 208176 226636
rect 212172 226584 212224 226636
rect 214932 226584 214984 226636
rect 219532 226584 219584 226636
rect 223580 226584 223632 226636
rect 225604 226584 225656 226636
rect 238392 226584 238444 226636
rect 259368 226584 259420 226636
rect 298284 226584 298336 226636
rect 673736 226516 673788 226568
rect 106924 226448 106976 226500
rect 146300 226448 146352 226500
rect 150072 226448 150124 226500
rect 213276 226448 213328 226500
rect 216404 226448 216456 226500
rect 220544 226448 220596 226500
rect 220728 226448 220780 226500
rect 228916 226448 228968 226500
rect 369124 226448 369176 226500
rect 376208 226448 376260 226500
rect 403992 226448 404044 226500
rect 412272 226448 412324 226500
rect 474740 226448 474792 226500
rect 482744 226448 482796 226500
rect 386052 226380 386104 226432
rect 391204 226380 391256 226432
rect 672724 226380 672776 226432
rect 407764 226312 407816 226364
rect 408684 226312 408736 226364
rect 481640 226312 481692 226364
rect 487804 226312 487856 226364
rect 488080 226312 488132 226364
rect 490012 226312 490064 226364
rect 122564 226244 122616 226296
rect 193956 226244 194008 226296
rect 195244 226244 195296 226296
rect 201684 226244 201736 226296
rect 203156 226244 203208 226296
rect 209412 226244 209464 226296
rect 209596 226244 209648 226296
rect 255136 226244 255188 226296
rect 260656 226244 260708 226296
rect 298928 226244 298980 226296
rect 308864 226244 308916 226296
rect 336280 226244 336332 226296
rect 388628 226244 388680 226296
rect 394240 226244 394292 226296
rect 458640 226244 458692 226296
rect 462964 226244 463016 226296
rect 72424 226108 72476 226160
rect 141148 226108 141200 226160
rect 141516 226108 141568 226160
rect 145012 226108 145064 226160
rect 145196 226108 145248 226160
rect 147496 226108 147548 226160
rect 148968 226108 149020 226160
rect 214564 226108 214616 226160
rect 222016 226108 222068 226160
rect 269948 226108 270000 226160
rect 270224 226108 270276 226160
rect 287520 226108 287572 226160
rect 288072 226108 288124 226160
rect 322756 226108 322808 226160
rect 526444 226108 526496 226160
rect 539968 226244 540020 226296
rect 563704 226244 563756 226296
rect 568120 226244 568172 226296
rect 83464 225972 83516 226024
rect 163044 225972 163096 226024
rect 193772 225972 193824 226024
rect 199292 225972 199344 226024
rect 199476 225972 199528 226024
rect 236460 225972 236512 226024
rect 252468 225972 252520 226024
rect 293132 225972 293184 226024
rect 299388 225972 299440 226024
rect 328552 225972 328604 226024
rect 335176 225972 335228 226024
rect 356888 225972 356940 226024
rect 361212 225972 361264 226024
rect 377496 225972 377548 226024
rect 498108 225972 498160 226024
rect 514300 225972 514352 226024
rect 516600 225972 516652 226024
rect 538496 226108 538548 226160
rect 672604 226108 672656 226160
rect 671252 226040 671304 226092
rect 538312 225972 538364 226024
rect 556160 225972 556212 226024
rect 557448 225972 557500 226024
rect 76564 225836 76616 225888
rect 158260 225836 158312 225888
rect 169668 225836 169720 225888
rect 171600 225836 171652 225888
rect 171784 225836 171836 225888
rect 204536 225836 204588 225888
rect 204720 225836 204772 225888
rect 249248 225836 249300 225888
rect 261852 225836 261904 225888
rect 300860 225836 300912 225888
rect 312912 225836 312964 225888
rect 341708 225836 341760 225888
rect 341984 225836 342036 225888
rect 365260 225836 365312 225888
rect 375012 225836 375064 225888
rect 387800 225836 387852 225888
rect 394332 225836 394384 225888
rect 403256 225836 403308 225888
rect 501144 225836 501196 225888
rect 519176 225836 519228 225888
rect 521752 225836 521804 225888
rect 545764 225836 545816 225888
rect 672264 225836 672316 225888
rect 66168 225700 66220 225752
rect 149796 225700 149848 225752
rect 151268 225700 151320 225752
rect 58992 225564 59044 225616
rect 141516 225564 141568 225616
rect 141792 225564 141844 225616
rect 203156 225564 203208 225616
rect 204904 225700 204956 225752
rect 244188 225700 244240 225752
rect 251088 225700 251140 225752
rect 294420 225700 294472 225752
rect 296444 225700 296496 225752
rect 327908 225700 327960 225752
rect 329748 225700 329800 225752
rect 353668 225700 353720 225752
rect 365352 225700 365404 225752
rect 383292 225700 383344 225752
rect 387708 225700 387760 225752
rect 397828 225700 397880 225752
rect 481180 225700 481232 225752
rect 492680 225700 492732 225752
rect 493784 225700 493836 225752
rect 505284 225700 505336 225752
rect 508872 225700 508924 225752
rect 529204 225700 529256 225752
rect 535920 225700 535972 225752
rect 563060 225700 563112 225752
rect 217140 225564 217192 225616
rect 219992 225564 220044 225616
rect 266084 225564 266136 225616
rect 267004 225564 267056 225616
rect 274456 225564 274508 225616
rect 278412 225564 278464 225616
rect 313280 225564 313332 225616
rect 327724 225564 327776 225616
rect 352380 225564 352432 225616
rect 352932 225564 352984 225616
rect 371608 225564 371660 225616
rect 382924 225564 382976 225616
rect 396172 225564 396224 225616
rect 410984 225564 411036 225616
rect 416136 225564 416188 225616
rect 467656 225564 467708 225616
rect 476580 225564 476632 225616
rect 477316 225564 477368 225616
rect 488724 225564 488776 225616
rect 489368 225564 489420 225616
rect 502984 225564 503036 225616
rect 510160 225564 510212 225616
rect 530952 225564 531004 225616
rect 531412 225564 531464 225616
rect 558184 225564 558236 225616
rect 672264 225496 672316 225548
rect 125232 225428 125284 225480
rect 196164 225428 196216 225480
rect 198004 225428 198056 225480
rect 204720 225428 204772 225480
rect 205088 225428 205140 225480
rect 209320 225428 209372 225480
rect 209504 225428 209556 225480
rect 259644 225428 259696 225480
rect 297364 225428 297416 225480
rect 310520 225428 310572 225480
rect 463148 225360 463200 225412
rect 467288 225360 467340 225412
rect 129372 225292 129424 225344
rect 199108 225292 199160 225344
rect 199292 225292 199344 225344
rect 204904 225292 204956 225344
rect 62028 225156 62080 225208
rect 130384 225156 130436 225208
rect 132408 225156 132460 225208
rect 195244 225156 195296 225208
rect 196624 225156 196676 225208
rect 199476 225156 199528 225208
rect 202788 225156 202840 225208
rect 135168 225020 135220 225072
rect 204260 225020 204312 225072
rect 204628 225156 204680 225208
rect 222936 225292 222988 225344
rect 242900 225292 242952 225344
rect 285036 225292 285088 225344
rect 672156 225292 672208 225344
rect 672034 225224 672086 225276
rect 254492 225156 254544 225208
rect 215208 225020 215260 225072
rect 219992 225020 220044 225072
rect 666468 225020 666520 225072
rect 355232 224952 355284 225004
rect 358176 224952 358228 225004
rect 404176 224952 404228 225004
rect 410616 224952 410668 225004
rect 416504 224952 416556 225004
rect 422208 224952 422260 225004
rect 96252 224884 96304 224936
rect 172980 224884 173032 224936
rect 176844 224884 176896 224936
rect 89444 224748 89496 224800
rect 168196 224748 168248 224800
rect 170864 224748 170916 224800
rect 178500 224748 178552 224800
rect 179328 224884 179380 224936
rect 185584 224884 185636 224936
rect 185768 224884 185820 224936
rect 199752 224884 199804 224936
rect 199936 224884 199988 224936
rect 248052 224884 248104 224936
rect 272524 224884 272576 224936
rect 309876 224884 309928 224936
rect 319812 224884 319864 224936
rect 345940 224884 345992 224936
rect 460572 224884 460624 224936
rect 463148 224884 463200 224936
rect 519360 224884 519412 224936
rect 535000 224884 535052 224936
rect 621020 224884 621072 224936
rect 350356 224816 350408 224868
rect 354956 224816 355008 224868
rect 670700 224816 670752 224868
rect 232596 224748 232648 224800
rect 245476 224748 245528 224800
rect 287704 224748 287756 224800
rect 311532 224748 311584 224800
rect 338856 224748 338908 224800
rect 462504 224748 462556 224800
rect 469312 224748 469364 224800
rect 506940 224748 506992 224800
rect 526352 224748 526404 224800
rect 529940 224748 529992 224800
rect 543004 224748 543056 224800
rect 543188 224748 543240 224800
rect 548616 224748 548668 224800
rect 548984 224748 549036 224800
rect 549996 224748 550048 224800
rect 85488 224612 85540 224664
rect 165620 224612 165672 224664
rect 79968 224476 80020 224528
rect 160468 224476 160520 224528
rect 165528 224476 165580 224528
rect 171784 224612 171836 224664
rect 171968 224612 172020 224664
rect 185400 224612 185452 224664
rect 185584 224612 185636 224664
rect 237748 224612 237800 224664
rect 248328 224612 248380 224664
rect 291844 224612 291896 224664
rect 294880 224612 294932 224664
rect 325976 224612 326028 224664
rect 346308 224612 346360 224664
rect 366548 224612 366600 224664
rect 494060 224612 494112 224664
rect 510160 224612 510212 224664
rect 520464 224612 520516 224664
rect 544568 224612 544620 224664
rect 548064 224612 548116 224664
rect 550640 224612 550692 224664
rect 554964 224748 555016 224800
rect 555976 224748 556028 224800
rect 557264 224748 557316 224800
rect 557448 224748 557500 224800
rect 558552 224748 558604 224800
rect 561404 224748 561456 224800
rect 562692 224748 562744 224800
rect 571708 224748 571760 224800
rect 73712 224340 73764 224392
rect 155316 224340 155368 224392
rect 157248 224340 157300 224392
rect 157984 224340 158036 224392
rect 162768 224340 162820 224392
rect 224868 224476 224920 224528
rect 228732 224476 228784 224528
rect 274916 224476 274968 224528
rect 275100 224476 275152 224528
rect 311164 224476 311216 224528
rect 322848 224476 322900 224528
rect 349804 224476 349856 224528
rect 359464 224476 359516 224528
rect 378140 224476 378192 224528
rect 379244 224476 379296 224528
rect 393596 224476 393648 224528
rect 456064 224476 456116 224528
rect 459744 224476 459796 224528
rect 491300 224476 491352 224528
rect 506020 224476 506072 224528
rect 515956 224476 516008 224528
rect 539508 224476 539560 224528
rect 543004 224476 543056 224528
rect 548984 224476 549036 224528
rect 549260 224476 549312 224528
rect 555792 224476 555844 224528
rect 626540 224612 626592 224664
rect 166172 224340 166224 224392
rect 68928 224204 68980 224256
rect 152740 224204 152792 224256
rect 155868 224204 155920 224256
rect 160192 224204 160244 224256
rect 168012 224340 168064 224392
rect 171554 224340 171606 224392
rect 172152 224340 172204 224392
rect 227444 224340 227496 224392
rect 233148 224340 233200 224392
rect 277676 224340 277728 224392
rect 286324 224340 286376 224392
rect 289912 224340 289964 224392
rect 290832 224340 290884 224392
rect 324044 224340 324096 224392
rect 342168 224340 342220 224392
rect 362040 224340 362092 224392
rect 366732 224340 366784 224392
rect 381636 224340 381688 224392
rect 394516 224340 394568 224392
rect 404544 224340 404596 224392
rect 480536 224340 480588 224392
rect 492864 224340 492916 224392
rect 499212 224340 499264 224392
rect 516600 224340 516652 224392
rect 525616 224340 525668 224392
rect 548064 224340 548116 224392
rect 548616 224340 548668 224392
rect 556160 224340 556212 224392
rect 557356 224340 557408 224392
rect 562600 224476 562652 224528
rect 563152 224476 563204 224528
rect 625252 224476 625304 224528
rect 562784 224340 562836 224392
rect 565176 224272 565228 224324
rect 625988 224340 626040 224392
rect 667020 224340 667072 224392
rect 671482 224612 671534 224664
rect 171968 224204 172020 224256
rect 172152 224204 172204 224256
rect 176292 224204 176344 224256
rect 102048 224068 102100 224120
rect 170864 224068 170916 224120
rect 171784 224068 171836 224120
rect 230020 224204 230072 224256
rect 231676 224204 231728 224256
rect 278964 224204 279016 224256
rect 289636 224204 289688 224256
rect 296996 224204 297048 224256
rect 299112 224204 299164 224256
rect 331772 224204 331824 224256
rect 339408 224204 339460 224256
rect 362316 224204 362368 224256
rect 372528 224204 372580 224256
rect 387432 224204 387484 224256
rect 390192 224204 390244 224256
rect 401968 224204 402020 224256
rect 405556 224204 405608 224256
rect 414204 224204 414256 224256
rect 470232 224204 470284 224256
rect 480352 224204 480404 224256
rect 483756 224204 483808 224256
rect 496912 224204 496964 224256
rect 177488 224068 177540 224120
rect 106004 223932 106056 223984
rect 181076 223932 181128 223984
rect 185400 224068 185452 224120
rect 194600 224068 194652 224120
rect 195888 224068 195940 224120
rect 250628 224068 250680 224120
rect 266268 224068 266320 224120
rect 303436 224068 303488 224120
rect 304264 224068 304316 224120
rect 315304 224068 315356 224120
rect 504364 224068 504416 224120
rect 523500 224204 523552 224256
rect 535276 224204 535328 224256
rect 562692 224204 562744 224256
rect 562876 224136 562928 224188
rect 610440 224136 610492 224188
rect 610624 224136 610676 224188
rect 617064 224136 617116 224188
rect 670792 224136 670844 224188
rect 524420 224000 524472 224052
rect 525064 224000 525116 224052
rect 619640 224000 619692 224052
rect 666836 224000 666888 224052
rect 185768 223932 185820 223984
rect 191564 223932 191616 223984
rect 199844 223932 199896 223984
rect 201408 223932 201460 223984
rect 255780 223932 255832 223984
rect 331864 223932 331916 223984
rect 337568 223932 337620 223984
rect 279424 223864 279476 223916
rect 284760 223864 284812 223916
rect 517704 223864 517756 223916
rect 610624 223864 610676 223916
rect 610808 223864 610860 223916
rect 622492 223864 622544 223916
rect 108672 223796 108724 223848
rect 183836 223796 183888 223848
rect 184388 223796 184440 223848
rect 207480 223796 207532 223848
rect 227536 223796 227588 223848
rect 273168 223796 273220 223848
rect 505100 223728 505152 223780
rect 507676 223728 507728 223780
rect 539968 223728 540020 223780
rect 622676 223728 622728 223780
rect 667020 223728 667072 223780
rect 115296 223660 115348 223712
rect 188804 223660 188856 223712
rect 207664 223660 207716 223712
rect 228088 223660 228140 223712
rect 505284 223592 505336 223644
rect 614948 223592 615000 223644
rect 670792 223592 670844 223644
rect 87972 223524 88024 223576
rect 164976 223524 165028 223576
rect 171784 223524 171836 223576
rect 181720 223524 181772 223576
rect 183192 223524 183244 223576
rect 184664 223524 184716 223576
rect 184848 223524 184900 223576
rect 239680 223524 239732 223576
rect 249432 223524 249484 223576
rect 276296 223524 276348 223576
rect 278596 223524 278648 223576
rect 315028 223524 315080 223576
rect 406752 223524 406804 223576
rect 414848 223524 414900 223576
rect 454868 223524 454920 223576
rect 460480 223524 460532 223576
rect 473452 223524 473504 223576
rect 475568 223524 475620 223576
rect 99288 223388 99340 223440
rect 176016 223388 176068 223440
rect 187332 223388 187384 223440
rect 242256 223388 242308 223440
rect 244096 223388 244148 223440
rect 286048 223388 286100 223440
rect 81348 223252 81400 223304
rect 151912 223252 151964 223304
rect 68744 223116 68796 223168
rect 146484 223116 146536 223168
rect 146668 223116 146720 223168
rect 156420 223252 156472 223304
rect 156604 223252 156656 223304
rect 161940 223252 161992 223304
rect 162124 223252 162176 223304
rect 186872 223252 186924 223304
rect 188896 223252 188948 223304
rect 245108 223252 245160 223304
rect 250904 223252 250956 223304
rect 291200 223388 291252 223440
rect 316684 223388 316736 223440
rect 327264 223388 327316 223440
rect 517520 223388 517572 223440
rect 532516 223388 532568 223440
rect 534816 223388 534868 223440
rect 547420 223388 547472 223440
rect 297548 223320 297600 223372
rect 305368 223320 305420 223372
rect 288992 223252 289044 223304
rect 295064 223252 295116 223304
rect 307668 223252 307720 223304
rect 335636 223252 335688 223304
rect 337936 223252 337988 223304
rect 359188 223252 359240 223304
rect 493048 223252 493100 223304
rect 508504 223252 508556 223304
rect 514668 223252 514720 223304
rect 535460 223252 535512 223304
rect 75828 222980 75880 223032
rect 154948 223116 155000 223168
rect 156420 223116 156472 223168
rect 176108 223116 176160 223168
rect 181996 223116 182048 223168
rect 240324 223116 240376 223168
rect 241336 223116 241388 223168
rect 283472 223116 283524 223168
rect 288256 223116 288308 223168
rect 321468 223116 321520 223168
rect 323952 223116 324004 223168
rect 348516 223116 348568 223168
rect 358544 223116 358596 223168
rect 374644 223116 374696 223168
rect 483112 223116 483164 223168
rect 496084 223116 496136 223168
rect 503352 223116 503404 223168
rect 521752 223116 521804 223168
rect 529480 223116 529532 223168
rect 555700 223116 555752 223168
rect 152372 222980 152424 223032
rect 71412 222844 71464 222896
rect 151636 222844 151688 222896
rect 151774 222844 151826 222896
rect 156420 222844 156472 222896
rect 158076 222980 158128 223032
rect 219072 222980 219124 223032
rect 245292 222980 245344 223032
rect 289268 222980 289320 223032
rect 291660 222980 291712 223032
rect 300216 222980 300268 223032
rect 315672 222980 315724 223032
rect 344652 222980 344704 223032
rect 171784 222844 171836 222896
rect 172888 222844 172940 222896
rect 212632 222844 212684 222896
rect 213184 222844 213236 222896
rect 233332 222844 233384 222896
rect 234528 222844 234580 222896
rect 281540 222844 281592 222896
rect 282736 222844 282788 222896
rect 316316 222844 316368 222896
rect 321468 222844 321520 222896
rect 346584 222980 346636 223032
rect 349068 222980 349120 223032
rect 367192 222980 367244 223032
rect 368388 222980 368440 223032
rect 382648 222980 382700 223032
rect 383568 222980 383620 223032
rect 394884 222980 394936 223032
rect 486608 222980 486660 223032
rect 500040 222980 500092 223032
rect 508228 222980 508280 223032
rect 527732 222980 527784 223032
rect 532056 222980 532108 223032
rect 559012 222980 559064 223032
rect 670792 223116 670844 223168
rect 345296 222844 345348 222896
rect 347872 222844 347924 222896
rect 78588 222708 78640 222760
rect 127624 222708 127676 222760
rect 127808 222708 127860 222760
rect 191380 222708 191432 222760
rect 197176 222708 197228 222760
rect 249984 222708 250036 222760
rect 284208 222708 284260 222760
rect 316960 222708 317012 222760
rect 347228 222708 347280 222760
rect 367836 222844 367888 222896
rect 375196 222844 375248 222896
rect 391020 222844 391072 222896
rect 395804 222844 395856 222896
rect 406476 222844 406528 222896
rect 420828 222844 420880 222896
rect 425152 222844 425204 222896
rect 459928 222844 459980 222896
rect 467104 222844 467156 222896
rect 467472 222844 467524 222896
rect 473728 222844 473780 222896
rect 479892 222844 479944 222896
rect 492036 222844 492088 222896
rect 500776 222844 500828 222896
rect 517520 222844 517572 222896
rect 519820 222844 519872 222896
rect 543372 222844 543424 222896
rect 554044 222844 554096 222896
rect 632704 222844 632756 222896
rect 651288 222844 651340 222896
rect 666468 222844 666520 222896
rect 532516 222708 532568 222760
rect 543004 222708 543056 222760
rect 558184 222708 558236 222760
rect 426440 222640 426492 222692
rect 426992 222640 427044 222692
rect 85304 222572 85356 222624
rect 156604 222572 156656 222624
rect 166356 222572 166408 222624
rect 192024 222572 192076 222624
rect 194508 222572 194560 222624
rect 247408 222572 247460 222624
rect 482744 222572 482796 222624
rect 593972 222572 594024 222624
rect 630680 222572 630732 222624
rect 118424 222436 118476 222488
rect 127624 222436 127676 222488
rect 146668 222436 146720 222488
rect 127808 222300 127860 222352
rect 139124 222300 139176 222352
rect 206836 222436 206888 222488
rect 207848 222436 207900 222488
rect 258356 222436 258408 222488
rect 500224 222436 500276 222488
rect 542820 222436 542872 222488
rect 543004 222436 543056 222488
rect 621204 222436 621256 222488
rect 490012 222368 490064 222420
rect 147128 222300 147180 222352
rect 211988 222300 212040 222352
rect 237012 222300 237064 222352
rect 280896 222300 280948 222352
rect 484584 222300 484636 222352
rect 629852 222300 629904 222352
rect 500224 222164 500276 222216
rect 542820 222164 542872 222216
rect 558184 222164 558236 222216
rect 558552 222164 558604 222216
rect 559932 222164 559984 222216
rect 627092 222164 627144 222216
rect 111984 222096 112036 222148
rect 185952 222096 186004 222148
rect 200396 222096 200448 222148
rect 252928 222096 252980 222148
rect 258080 222096 258132 222148
rect 263876 222096 263928 222148
rect 270040 222096 270092 222148
rect 306380 222096 306432 222148
rect 310704 222096 310756 222148
rect 312636 222096 312688 222148
rect 331404 222096 331456 222148
rect 353944 222096 353996 222148
rect 424968 222096 425020 222148
rect 429292 222096 429344 222148
rect 452568 222096 452620 222148
rect 455604 222096 455656 222148
rect 462136 222096 462188 222148
rect 468760 222096 468812 222148
rect 471888 222096 471940 222148
rect 477868 222096 477920 222148
rect 533160 222096 533212 222148
rect 538680 222096 538732 222148
rect 539508 222096 539560 222148
rect 542268 222096 542320 222148
rect 670792 222096 670844 222148
rect 543832 222028 543884 222080
rect 605012 222028 605064 222080
rect 91284 221960 91336 222012
rect 167184 221960 167236 222012
rect 167460 221960 167512 222012
rect 172704 221960 172756 222012
rect 94596 221824 94648 221876
rect 161434 221824 161486 221876
rect 161572 221824 161624 221876
rect 164332 221824 164384 221876
rect 164516 221824 164568 221876
rect 169852 221824 169904 221876
rect 97724 221688 97776 221740
rect 167460 221688 167512 221740
rect 167644 221688 167696 221740
rect 73896 221552 73948 221604
rect 82084 221552 82136 221604
rect 86316 221552 86368 221604
rect 161480 221552 161532 221604
rect 161664 221552 161716 221604
rect 167828 221552 167880 221604
rect 168196 221688 168248 221740
rect 226524 221960 226576 222012
rect 232136 221960 232188 222012
rect 234712 221960 234764 222012
rect 261024 221960 261076 222012
rect 301688 221960 301740 222012
rect 313188 221960 313240 222012
rect 340420 221960 340472 222012
rect 516784 221960 516836 222012
rect 527548 221960 527600 222012
rect 527732 221960 527784 222012
rect 528192 221960 528244 222012
rect 533528 221960 533580 222012
rect 533988 221960 534040 222012
rect 543004 221960 543056 222012
rect 543372 221960 543424 222012
rect 543694 221960 543746 222012
rect 174084 221824 174136 221876
rect 231952 221824 232004 221876
rect 233700 221824 233752 221876
rect 277952 221824 278004 221876
rect 280068 221824 280120 221876
rect 313740 221824 313792 221876
rect 318248 221824 318300 221876
rect 343640 221824 343692 221876
rect 353300 221824 353352 221876
rect 372712 221824 372764 221876
rect 174912 221688 174964 221740
rect 185768 221688 185820 221740
rect 243084 221688 243136 221740
rect 182640 221552 182692 221604
rect 232136 221552 232188 221604
rect 263140 221688 263192 221740
rect 263508 221688 263560 221740
rect 301044 221688 301096 221740
rect 303252 221688 303304 221740
rect 332784 221688 332836 221740
rect 344652 221688 344704 221740
rect 364524 221688 364576 221740
rect 370964 221688 371016 221740
rect 380348 221824 380400 221876
rect 492496 221824 492548 221876
rect 506848 221824 506900 221876
rect 515772 221824 515824 221876
rect 600320 221824 600372 221876
rect 380072 221688 380124 221740
rect 386512 221688 386564 221740
rect 484768 221688 484820 221740
rect 497740 221688 497792 221740
rect 501328 221688 501380 221740
rect 519636 221688 519688 221740
rect 522672 221688 522724 221740
rect 542360 221688 542412 221740
rect 543004 221688 543056 221740
rect 543694 221688 543746 221740
rect 543832 221688 543884 221740
rect 601148 221688 601200 221740
rect 59360 221416 59412 221468
rect 141332 221416 141384 221468
rect 147588 221416 147640 221468
rect 204904 221416 204956 221468
rect 205088 221416 205140 221468
rect 220176 221416 220228 221468
rect 221004 221416 221056 221468
rect 243728 221552 243780 221604
rect 283748 221552 283800 221604
rect 302424 221552 302476 221604
rect 334072 221552 334124 221604
rect 348792 221552 348844 221604
rect 370044 221552 370096 221604
rect 373724 221552 373776 221604
rect 384304 221552 384356 221604
rect 391020 221552 391072 221604
rect 400312 221552 400364 221604
rect 401232 221552 401284 221604
rect 405832 221552 405884 221604
rect 475844 221552 475896 221604
rect 486148 221552 486200 221604
rect 496268 221552 496320 221604
rect 513564 221552 513616 221604
rect 524236 221552 524288 221604
rect 234068 221416 234120 221468
rect 276112 221416 276164 221468
rect 284024 221416 284076 221468
rect 320364 221416 320416 221468
rect 333612 221416 333664 221468
rect 357532 221416 357584 221468
rect 369492 221416 369544 221468
rect 384120 221416 384172 221468
rect 384396 221416 384448 221468
rect 395160 221416 395212 221468
rect 396816 221416 396868 221468
rect 407304 221416 407356 221468
rect 408408 221416 408460 221468
rect 416872 221416 416924 221468
rect 468944 221416 468996 221468
rect 476212 221416 476264 221468
rect 483756 221416 483808 221468
rect 533160 221416 533212 221468
rect 533528 221552 533580 221604
rect 600688 221552 600740 221604
rect 543740 221416 543792 221468
rect 544752 221416 544804 221468
rect 606116 221552 606168 221604
rect 601148 221416 601200 221468
rect 605932 221416 605984 221468
rect 104532 221280 104584 221332
rect 176476 221280 176528 221332
rect 111156 221144 111208 221196
rect 167644 221144 167696 221196
rect 167828 221144 167880 221196
rect 185860 221280 185912 221332
rect 234252 221280 234304 221332
rect 237840 221280 237892 221332
rect 243728 221280 243780 221332
rect 266820 221280 266872 221332
rect 303804 221280 303856 221332
rect 600688 221280 600740 221332
rect 603172 221280 603224 221332
rect 177304 221144 177356 221196
rect 185308 221144 185360 221196
rect 520924 221212 520976 221264
rect 600504 221212 600556 221264
rect 124404 221008 124456 221060
rect 193312 221008 193364 221060
rect 204904 221144 204956 221196
rect 211160 221144 211212 221196
rect 211528 221144 211580 221196
rect 260840 221144 260892 221196
rect 517520 221076 517572 221128
rect 518440 221076 518492 221128
rect 600688 221076 600740 221128
rect 205088 221008 205140 221060
rect 218060 221008 218112 221060
rect 221004 221008 221056 221060
rect 227904 221008 227956 221060
rect 234068 221008 234120 221060
rect 83004 220940 83056 220992
rect 151084 220872 151136 220924
rect 155040 220872 155092 220924
rect 158260 220872 158312 220924
rect 158444 220872 158496 220924
rect 222292 220872 222344 220924
rect 223488 220872 223540 220924
rect 268200 221008 268252 221060
rect 523500 220940 523552 220992
rect 601700 220940 601752 220992
rect 253388 220872 253440 220924
rect 258632 220872 258684 220924
rect 80520 220804 80572 220856
rect 86132 220804 86184 220856
rect 418344 220804 418396 220856
rect 424048 220804 424100 220856
rect 456708 220804 456760 220856
rect 462136 220804 462188 220856
rect 466092 220804 466144 220856
rect 471336 220804 471388 220856
rect 538496 220804 538548 220856
rect 539508 220804 539560 220856
rect 542360 220804 542412 220856
rect 107844 220736 107896 220788
rect 176476 220736 176528 220788
rect 176614 220736 176666 220788
rect 180524 220736 180576 220788
rect 180708 220736 180760 220788
rect 236736 220736 236788 220788
rect 246948 220736 247000 220788
rect 288624 220736 288676 220788
rect 340052 220736 340104 220788
rect 342352 220736 342404 220788
rect 414204 220736 414256 220788
rect 418160 220736 418212 220788
rect 474004 220736 474056 220788
rect 475384 220736 475436 220788
rect 476764 220736 476816 220788
rect 478696 220736 478748 220788
rect 500408 220736 500460 220788
rect 511816 220736 511868 220788
rect 544384 220804 544436 220856
rect 553400 220804 553452 220856
rect 559564 220804 559616 220856
rect 563060 220804 563112 220856
rect 563244 220804 563296 220856
rect 609428 220804 609480 220856
rect 455328 220668 455380 220720
rect 458824 220668 458876 220720
rect 465724 220668 465776 220720
rect 469588 220668 469640 220720
rect 546592 220668 546644 220720
rect 79692 220600 79744 220652
rect 154028 220600 154080 220652
rect 154212 220600 154264 220652
rect 156788 220600 156840 220652
rect 156972 220600 157024 220652
rect 158904 220600 158956 220652
rect 160836 220600 160888 220652
rect 221280 220600 221332 220652
rect 76380 220464 76432 220516
rect 156144 220464 156196 220516
rect 156604 220464 156656 220516
rect 166954 220464 167006 220516
rect 167092 220464 167144 220516
rect 223764 220600 223816 220652
rect 236184 220600 236236 220652
rect 246488 220600 246540 220652
rect 254400 220600 254452 220652
rect 296812 220600 296864 220652
rect 304908 220600 304960 220652
rect 333428 220600 333480 220652
rect 509884 220600 509936 220652
rect 522580 220600 522632 220652
rect 529020 220600 529072 220652
rect 223764 220464 223816 220516
rect 270592 220464 270644 220516
rect 292488 220464 292540 220516
rect 326160 220464 326212 220516
rect 328092 220464 328144 220516
rect 351276 220464 351328 220516
rect 364524 220464 364576 220516
rect 379704 220464 379756 220516
rect 469128 220464 469180 220516
rect 474556 220464 474608 220516
rect 488448 220464 488500 220516
rect 501880 220464 501932 220516
rect 511632 220464 511684 220516
rect 531688 220464 531740 220516
rect 540796 220464 540848 220516
rect 543556 220464 543608 220516
rect 558000 220600 558052 220652
rect 566464 220600 566516 220652
rect 566648 220600 566700 220652
rect 567292 220600 567344 220652
rect 568580 220600 568632 220652
rect 569776 220600 569828 220652
rect 569960 220600 570012 220652
rect 610532 220600 610584 220652
rect 544936 220464 544988 220516
rect 64604 220328 64656 220380
rect 141976 220328 142028 220380
rect 73068 220192 73120 220244
rect 151636 220328 151688 220380
rect 151774 220328 151826 220380
rect 208584 220328 208636 220380
rect 213828 220328 213880 220380
rect 262404 220328 262456 220380
rect 262680 220328 262732 220380
rect 264244 220328 264296 220380
rect 264612 220328 264664 220380
rect 269304 220328 269356 220380
rect 273444 220328 273496 220380
rect 309232 220328 309284 220380
rect 316500 220328 316552 220380
rect 342904 220328 342956 220380
rect 351276 220328 351328 220380
rect 369308 220328 369360 220380
rect 376944 220328 376996 220380
rect 388444 220328 388496 220380
rect 436284 220328 436336 220380
rect 437020 220328 437072 220380
rect 473176 220328 473228 220380
rect 481180 220328 481232 220380
rect 496452 220328 496504 220380
rect 509332 220328 509384 220380
rect 515404 220328 515456 220380
rect 530032 220328 530084 220380
rect 531136 220328 531188 220380
rect 553032 220464 553084 220516
rect 553860 220464 553912 220516
rect 608600 220464 608652 220516
rect 647240 220464 647292 220516
rect 651472 220464 651524 220516
rect 144276 220192 144328 220244
rect 146760 220192 146812 220244
rect 146944 220192 146996 220244
rect 156604 220192 156656 220244
rect 156788 220192 156840 220244
rect 215944 220192 215996 220244
rect 217140 220192 217192 220244
rect 265164 220192 265216 220244
rect 267648 220192 267700 220244
rect 306840 220192 306892 220244
rect 309048 220192 309100 220244
rect 339684 220192 339736 220244
rect 342996 220192 343048 220244
rect 363328 220192 363380 220244
rect 363696 220192 363748 220244
rect 381084 220192 381136 220244
rect 388444 220192 388496 220244
rect 400956 220192 401008 220244
rect 430120 220192 430172 220244
rect 432052 220192 432104 220244
rect 459468 220192 459520 220244
rect 465448 220192 465500 220244
rect 472992 220192 473044 220244
rect 482008 220192 482060 220244
rect 482928 220192 482980 220244
rect 495348 220192 495400 220244
rect 497464 220192 497516 220244
rect 515220 220192 515272 220244
rect 528376 220192 528428 220244
rect 554044 220328 554096 220380
rect 563060 220328 563112 220380
rect 610072 220328 610124 220380
rect 560760 220260 560812 220312
rect 562876 220260 562928 220312
rect 548708 220192 548760 220244
rect 101220 220056 101272 220108
rect 166954 220056 167006 220108
rect 167092 220056 167144 220108
rect 114468 219920 114520 219972
rect 180892 219920 180944 219972
rect 181536 220056 181588 220108
rect 229284 220056 229336 220108
rect 230204 220056 230256 220108
rect 275284 220056 275336 220108
rect 276756 220056 276808 220108
rect 311348 220056 311400 220108
rect 328920 220056 328972 220108
rect 354772 220056 354824 220108
rect 355416 220056 355468 220108
rect 375564 220056 375616 220108
rect 379428 220056 379480 220108
rect 392124 220056 392176 220108
rect 395988 220056 396040 220108
rect 404728 220056 404780 220108
rect 421656 220056 421708 220108
rect 426716 220056 426768 220108
rect 431960 220056 432012 220108
rect 434812 220056 434864 220108
rect 478328 220056 478380 220108
rect 489460 220056 489512 220108
rect 489644 220056 489696 220108
rect 504364 220056 504416 220108
rect 513104 220056 513156 220108
rect 534172 220056 534224 220108
rect 538128 220056 538180 220108
rect 558000 220056 558052 220108
rect 576768 220192 576820 220244
rect 611636 220192 611688 220244
rect 668952 220192 669004 220244
rect 558368 220124 558420 220176
rect 576584 220124 576636 220176
rect 582472 220056 582524 220108
rect 633440 220056 633492 220108
rect 576768 219988 576820 220040
rect 576952 219988 577004 220040
rect 581644 219988 581696 220040
rect 581828 219988 581880 220040
rect 582334 219988 582386 220040
rect 669136 219988 669188 220040
rect 190460 219920 190512 219972
rect 190644 219920 190696 219972
rect 244464 219920 244516 219972
rect 253572 219920 253624 219972
rect 293316 219920 293368 219972
rect 530032 219852 530084 219904
rect 558368 219852 558420 219904
rect 558736 219852 558788 219904
rect 600964 219852 601016 219904
rect 601148 219852 601200 219904
rect 619824 219852 619876 219904
rect 121092 219784 121144 219836
rect 134340 219784 134392 219836
rect 140780 219784 140832 219836
rect 140964 219784 141016 219836
rect 141976 219784 142028 219836
rect 142160 219784 142212 219836
rect 200212 219784 200264 219836
rect 200580 219784 200632 219836
rect 252744 219784 252796 219836
rect 286692 219784 286744 219836
rect 319076 219784 319128 219836
rect 527548 219716 527600 219768
rect 548708 219716 548760 219768
rect 548892 219716 548944 219768
rect 146944 219648 146996 219700
rect 69756 219512 69808 219564
rect 142160 219512 142212 219564
rect 142344 219512 142396 219564
rect 205824 219648 205876 219700
rect 207204 219648 207256 219700
rect 257252 219648 257304 219700
rect 464988 219580 465040 219632
rect 472072 219580 472124 219632
rect 506020 219580 506072 219632
rect 576768 219580 576820 219632
rect 581644 219580 581696 219632
rect 582380 219580 582432 219632
rect 582656 219580 582708 219632
rect 601148 219580 601200 219632
rect 601516 219716 601568 219768
rect 620008 219716 620060 219768
rect 607496 219580 607548 219632
rect 147772 219512 147824 219564
rect 150716 219512 150768 219564
rect 150900 219512 150952 219564
rect 214012 219512 214064 219564
rect 270776 219512 270828 219564
rect 279148 219512 279200 219564
rect 289820 219512 289872 219564
rect 63960 219376 64012 219428
rect 64880 219376 64932 219428
rect 105820 219394 105872 219446
rect 147128 219376 147180 219428
rect 159824 219376 159876 219428
rect 204536 219376 204588 219428
rect 209688 219376 209740 219428
rect 210424 219376 210476 219428
rect 213000 219376 213052 219428
rect 258080 219376 258132 219428
rect 272892 219376 272944 219428
rect 366732 219512 366784 219564
rect 405924 219444 405976 219496
rect 412732 219444 412784 219496
rect 63132 219104 63184 219156
rect 106924 219240 106976 219292
rect 113640 219240 113692 219292
rect 156236 219240 156288 219292
rect 162492 219240 162544 219292
rect 166540 219240 166592 219292
rect 167460 219240 167512 219292
rect 168196 219240 168248 219292
rect 169116 219240 169168 219292
rect 169668 219240 169720 219292
rect 169944 219240 169996 219292
rect 171048 219240 171100 219292
rect 171600 219240 171652 219292
rect 172152 219240 172204 219292
rect 172428 219240 172480 219292
rect 173164 219240 173216 219292
rect 182364 219240 182416 219292
rect 189724 219240 189776 219292
rect 192852 219240 192904 219292
rect 198188 219240 198240 219292
rect 198924 219240 198976 219292
rect 200028 219240 200080 219292
rect 202604 219240 202656 219292
rect 207664 219240 207716 219292
rect 211344 219240 211396 219292
rect 218060 219240 218112 219292
rect 239496 219240 239548 219292
rect 272708 219240 272760 219292
rect 70584 219104 70636 219156
rect 117964 219104 118016 219156
rect 132592 219104 132644 219156
rect 177488 219104 177540 219156
rect 179052 219104 179104 219156
rect 196624 219104 196676 219156
rect 199752 219104 199804 219156
rect 243544 219104 243596 219156
rect 272340 219104 272392 219156
rect 289820 219240 289872 219292
rect 297548 219376 297600 219428
rect 304080 219376 304132 219428
rect 308404 219376 308456 219428
rect 320640 219376 320692 219428
rect 279056 219104 279108 219156
rect 286324 219104 286376 219156
rect 292028 219240 292080 219292
rect 313924 219240 313976 219292
rect 341340 219376 341392 219428
rect 342260 219376 342312 219428
rect 343824 219376 343876 219428
rect 347044 219376 347096 219428
rect 366180 219376 366232 219428
rect 399300 219376 399352 219428
rect 400220 219376 400272 219428
rect 415860 219376 415912 219428
rect 416780 219376 416832 219428
rect 417516 219376 417568 219428
rect 421012 219444 421064 219496
rect 501052 219444 501104 219496
rect 577136 219394 577188 219446
rect 582656 219308 582708 219360
rect 591948 219444 592000 219496
rect 600136 219444 600188 219496
rect 600964 219444 601016 219496
rect 607312 219444 607364 219496
rect 596824 219308 596876 219360
rect 345296 219240 345348 219292
rect 419172 219240 419224 219292
rect 422668 219240 422720 219292
rect 552480 219240 552532 219292
rect 574744 219240 574796 219292
rect 582472 219172 582524 219224
rect 597928 219172 597980 219224
rect 62304 218968 62356 219020
rect 72424 218968 72476 219020
rect 77208 218968 77260 219020
rect 140044 218968 140096 219020
rect 142436 218968 142488 219020
rect 143724 218968 143776 219020
rect 146760 218968 146812 219020
rect 150440 218968 150492 219020
rect 153384 218968 153436 219020
rect 203524 218968 203576 219020
rect 206376 218968 206428 219020
rect 253388 218968 253440 219020
rect 259184 218968 259236 219020
rect 291660 218968 291712 219020
rect 295800 219104 295852 219156
rect 296720 219104 296772 219156
rect 300492 219104 300544 219156
rect 322112 219104 322164 219156
rect 325332 219104 325384 219156
rect 327724 219104 327776 219156
rect 340512 219104 340564 219156
rect 352564 219104 352616 219156
rect 362040 219104 362092 219156
rect 370964 219104 371016 219156
rect 543740 219104 543792 219156
rect 549076 219104 549128 219156
rect 553032 219104 553084 219156
rect 556620 219104 556672 219156
rect 561680 219104 561732 219156
rect 562416 219104 562468 219156
rect 571340 219104 571392 219156
rect 571524 219104 571576 219156
rect 297364 218968 297416 219020
rect 307392 218968 307444 219020
rect 331864 218968 331916 219020
rect 333428 218968 333480 219020
rect 355232 218968 355284 219020
rect 357072 218968 357124 219020
rect 369124 218968 369176 219020
rect 370320 218968 370372 219020
rect 380072 218968 380124 219020
rect 380256 218968 380308 219020
rect 388628 218968 388680 219020
rect 50712 218832 50764 218884
rect 62672 218832 62724 218884
rect 83832 218832 83884 218884
rect 153844 218832 153896 218884
rect 156236 218832 156288 218884
rect 162124 218832 162176 218884
rect 165804 218832 165856 218884
rect 59820 218696 59872 218748
rect 142436 218696 142488 218748
rect 142620 218696 142672 218748
rect 143264 218696 143316 218748
rect 145104 218696 145156 218748
rect 145932 218696 145984 218748
rect 148416 218696 148468 218748
rect 148968 218696 149020 218748
rect 149244 218696 149296 218748
rect 150072 218696 150124 218748
rect 150440 218696 150492 218748
rect 166540 218832 166592 218884
rect 171140 218832 171192 218884
rect 180064 218832 180116 218884
rect 100392 218560 100444 218612
rect 105820 218560 105872 218612
rect 107016 218560 107068 218612
rect 152372 218560 152424 218612
rect 152556 218560 152608 218612
rect 153108 218560 153160 218612
rect 156696 218560 156748 218612
rect 157248 218560 157300 218612
rect 157524 218560 157576 218612
rect 158260 218560 158312 218612
rect 159180 218560 159232 218612
rect 160008 218560 160060 218612
rect 161480 218560 161532 218612
rect 166080 218560 166132 218612
rect 120264 218424 120316 218476
rect 166080 218424 166132 218476
rect 175740 218696 175792 218748
rect 181168 218696 181220 218748
rect 184388 218696 184440 218748
rect 186504 218832 186556 218884
rect 239312 218832 239364 218884
rect 246120 218832 246172 218884
rect 279056 218832 279108 218884
rect 279240 218832 279292 218884
rect 189908 218696 189960 218748
rect 191932 218696 191984 218748
rect 195244 218696 195296 218748
rect 195612 218696 195664 218748
rect 198004 218696 198056 218748
rect 198188 218696 198240 218748
rect 246304 218696 246356 218748
rect 252744 218696 252796 218748
rect 166632 218560 166684 218612
rect 202604 218560 202656 218612
rect 203064 218560 203116 218612
rect 206192 218560 206244 218612
rect 208032 218560 208084 218612
rect 170956 218424 171008 218476
rect 171140 218424 171192 218476
rect 181352 218424 181404 218476
rect 189816 218424 189868 218476
rect 191932 218424 191984 218476
rect 117964 218288 118016 218340
rect 123484 218288 123536 218340
rect 131856 218288 131908 218340
rect 132408 218288 132460 218340
rect 136824 218288 136876 218340
rect 139492 218288 139544 218340
rect 140136 218288 140188 218340
rect 181168 218288 181220 218340
rect 181536 218288 181588 218340
rect 181996 218288 182048 218340
rect 184020 218288 184072 218340
rect 184940 218288 184992 218340
rect 185676 218288 185728 218340
rect 186136 218288 186188 218340
rect 188160 218288 188212 218340
rect 188896 218288 188948 218340
rect 189080 218288 189132 218340
rect 193772 218424 193824 218476
rect 198096 218424 198148 218476
rect 200396 218424 200448 218476
rect 202236 218424 202288 218476
rect 202788 218424 202840 218476
rect 204720 218424 204772 218476
rect 207848 218424 207900 218476
rect 208860 218424 208912 218476
rect 209504 218424 209556 218476
rect 210148 218560 210200 218612
rect 217324 218560 217376 218612
rect 219624 218560 219676 218612
rect 264612 218560 264664 218612
rect 265992 218560 266044 218612
rect 272340 218560 272392 218612
rect 272708 218560 272760 218612
rect 279424 218560 279476 218612
rect 211528 218424 211580 218476
rect 217968 218424 218020 218476
rect 223488 218424 223540 218476
rect 225972 218424 226024 218476
rect 267004 218424 267056 218476
rect 285864 218832 285916 218884
rect 292028 218832 292080 218884
rect 314016 218832 314068 218884
rect 340052 218832 340104 218884
rect 347044 218832 347096 218884
rect 363512 218832 363564 218884
rect 368664 218832 368716 218884
rect 378784 218832 378836 218884
rect 382740 218832 382792 218884
rect 383568 218832 383620 218884
rect 386880 218832 386932 218884
rect 398104 218832 398156 218884
rect 402612 218832 402664 218884
rect 409052 218832 409104 218884
rect 411720 218832 411772 218884
rect 412548 218832 412600 218884
rect 291660 218696 291712 218748
rect 324596 218696 324648 218748
rect 327264 218696 327316 218748
rect 351092 218696 351144 218748
rect 353760 218696 353812 218748
rect 371792 218696 371844 218748
rect 383568 218696 383620 218748
rect 396264 218696 396316 218748
rect 412548 218696 412600 218748
rect 417148 218696 417200 218748
rect 429936 218696 429988 218748
rect 432696 218696 432748 218748
rect 471336 218696 471388 218748
rect 472900 218696 472952 218748
rect 482744 218696 482796 218748
rect 485320 218696 485372 218748
rect 542820 218696 542872 218748
rect 304264 218560 304316 218612
rect 398472 218560 398524 218612
rect 407764 218560 407816 218612
rect 469864 218560 469916 218612
rect 471244 218560 471296 218612
rect 475568 218560 475620 218612
rect 482836 218560 482888 218612
rect 537484 218560 537536 218612
rect 543004 218560 543056 218612
rect 572076 218968 572128 219020
rect 544936 218832 544988 218884
rect 555976 218832 556028 218884
rect 547420 218696 547472 218748
rect 567660 218832 567712 218884
rect 568212 218832 568264 218884
rect 575480 218968 575532 219020
rect 626356 218832 626408 218884
rect 556436 218696 556488 218748
rect 567844 218696 567896 218748
rect 568028 218696 568080 218748
rect 570972 218696 571024 218748
rect 572536 218696 572588 218748
rect 601884 218696 601936 218748
rect 644940 218696 644992 218748
rect 656164 218696 656216 218748
rect 555976 218560 556028 218612
rect 598848 218560 598900 218612
rect 288992 218424 289044 218476
rect 294144 218424 294196 218476
rect 316684 218424 316736 218476
rect 500040 218424 500092 218476
rect 609888 218424 609940 218476
rect 458180 218356 458232 218408
rect 192300 218288 192352 218340
rect 193036 218288 193088 218340
rect 193956 218288 194008 218340
rect 194508 218288 194560 218340
rect 194784 218288 194836 218340
rect 195888 218288 195940 218340
rect 196440 218288 196492 218340
rect 210148 218288 210200 218340
rect 210332 218288 210384 218340
rect 213184 218288 213236 218340
rect 222936 218288 222988 218340
rect 231032 218288 231084 218340
rect 232872 218288 232924 218340
rect 270776 218288 270828 218340
rect 426624 218288 426676 218340
rect 429568 218288 429620 218340
rect 450728 218288 450780 218340
rect 453856 218288 453908 218340
rect 461308 218288 461360 218340
rect 503168 218288 503220 218340
rect 55680 218152 55732 218204
rect 56508 218152 56560 218204
rect 57428 218152 57480 218204
rect 61660 218152 61712 218204
rect 67272 218152 67324 218204
rect 68284 218152 68336 218204
rect 75552 218152 75604 218204
rect 76564 218152 76616 218204
rect 123576 218152 123628 218204
rect 161480 218152 161532 218204
rect 161664 218152 161716 218204
rect 162768 218152 162820 218204
rect 163320 218152 163372 218204
rect 163964 218152 164016 218204
rect 164976 218152 165028 218204
rect 165528 218152 165580 218204
rect 56508 218016 56560 218068
rect 57244 218016 57296 218068
rect 58164 218016 58216 218068
rect 59360 218016 59412 218068
rect 61476 218016 61528 218068
rect 62028 218016 62080 218068
rect 65616 218016 65668 218068
rect 66168 218016 66220 218068
rect 66444 218016 66496 218068
rect 67548 218016 67600 218068
rect 68100 218016 68152 218068
rect 68744 218016 68796 218068
rect 72240 218016 72292 218068
rect 73712 218016 73764 218068
rect 74724 218016 74776 218068
rect 75828 218016 75880 218068
rect 78036 218016 78088 218068
rect 78588 218016 78640 218068
rect 78864 218016 78916 218068
rect 79968 218016 80020 218068
rect 82176 218016 82228 218068
rect 83464 218016 83516 218068
rect 84660 218016 84712 218068
rect 85304 218016 85356 218068
rect 87144 218016 87196 218068
rect 88248 218016 88300 218068
rect 88800 218016 88852 218068
rect 89444 218016 89496 218068
rect 90456 218016 90508 218068
rect 91744 218016 91796 218068
rect 92940 218016 92992 218068
rect 93768 218016 93820 218068
rect 95424 218016 95476 218068
rect 96252 218016 96304 218068
rect 97080 218016 97132 218068
rect 98000 218016 98052 218068
rect 98736 218016 98788 218068
rect 99288 218016 99340 218068
rect 99564 218016 99616 218068
rect 100668 218016 100720 218068
rect 102876 218016 102928 218068
rect 103428 218016 103480 218068
rect 105360 218016 105412 218068
rect 106004 218016 106056 218068
rect 109500 218016 109552 218068
rect 110144 218016 110196 218068
rect 116124 218016 116176 218068
rect 117228 218016 117280 218068
rect 117780 218016 117832 218068
rect 118700 218016 118752 218068
rect 119436 218016 119488 218068
rect 119988 218016 120040 218068
rect 121920 218016 121972 218068
rect 122564 218016 122616 218068
rect 126060 218016 126112 218068
rect 126704 218016 126756 218068
rect 127716 218016 127768 218068
rect 128268 218016 128320 218068
rect 128544 218016 128596 218068
rect 129372 218016 129424 218068
rect 130200 218016 130252 218068
rect 132500 218016 132552 218068
rect 132684 218016 132736 218068
rect 133512 218016 133564 218068
rect 135996 218016 136048 218068
rect 136548 218016 136600 218068
rect 138480 218016 138532 218068
rect 139124 218016 139176 218068
rect 139492 218016 139544 218068
rect 171416 218152 171468 218204
rect 173256 218152 173308 218204
rect 170772 218016 170824 218068
rect 176476 218016 176528 218068
rect 178224 218016 178276 218068
rect 179328 218016 179380 218068
rect 179880 218152 179932 218204
rect 225604 218152 225656 218204
rect 241980 218152 242032 218204
rect 242900 218152 242952 218204
rect 243544 218152 243596 218204
rect 249064 218152 249116 218204
rect 297456 218152 297508 218204
rect 302884 218152 302936 218204
rect 333060 218152 333112 218204
rect 333888 218152 333940 218204
rect 335544 218152 335596 218204
rect 338672 218152 338724 218204
rect 358728 218152 358780 218204
rect 359464 218152 359516 218204
rect 381912 218152 381964 218204
rect 382924 218152 382976 218204
rect 400956 218152 401008 218204
rect 402244 218152 402296 218204
rect 407580 218152 407632 218204
rect 411904 218152 411956 218204
rect 422484 218152 422536 218204
rect 425428 218152 425480 218204
rect 425796 218152 425848 218204
rect 427912 218152 427964 218204
rect 428464 218152 428516 218204
rect 430120 218152 430172 218204
rect 433248 218152 433300 218204
rect 435272 218152 435324 218204
rect 435732 218152 435784 218204
rect 436652 218152 436704 218204
rect 461952 218152 462004 218204
rect 466276 218152 466328 218204
rect 507676 218152 507728 218204
rect 542820 218152 542872 218204
rect 543004 218152 543056 218204
rect 556436 218152 556488 218204
rect 562232 218288 562284 218340
rect 562876 218288 562928 218340
rect 614488 218288 614540 218340
rect 572674 218152 572726 218204
rect 615684 218152 615736 218204
rect 210332 218016 210384 218068
rect 210516 218016 210568 218068
rect 210976 218016 211028 218068
rect 214656 218016 214708 218068
rect 215208 218016 215260 218068
rect 215484 218016 215536 218068
rect 216128 218016 216180 218068
rect 218796 218016 218848 218068
rect 219348 218016 219400 218068
rect 221280 218016 221332 218068
rect 221832 218016 221884 218068
rect 225420 218016 225472 218068
rect 226156 218016 226208 218068
rect 227076 218016 227128 218068
rect 227536 218016 227588 218068
rect 229560 218016 229612 218068
rect 230480 218016 230532 218068
rect 231216 218016 231268 218068
rect 231676 218016 231728 218068
rect 232044 218016 232096 218068
rect 233148 218016 233200 218068
rect 235356 218016 235408 218068
rect 235816 218016 235868 218068
rect 240324 218016 240376 218068
rect 241336 218016 241388 218068
rect 243636 218016 243688 218068
rect 244096 218016 244148 218068
rect 244464 218016 244516 218068
rect 245292 218016 245344 218068
rect 247776 218016 247828 218068
rect 248328 218016 248380 218068
rect 248604 218016 248656 218068
rect 249248 218016 249300 218068
rect 250260 218016 250312 218068
rect 250904 218016 250956 218068
rect 251916 218016 251968 218068
rect 252468 218016 252520 218068
rect 256056 218016 256108 218068
rect 256516 218016 256568 218068
rect 256884 218016 256936 218068
rect 257528 218016 257580 218068
rect 258540 218016 258592 218068
rect 259368 218016 259420 218068
rect 260196 218016 260248 218068
rect 260748 218016 260800 218068
rect 264336 218016 264388 218068
rect 264796 218016 264848 218068
rect 265164 218016 265216 218068
rect 266268 218016 266320 218068
rect 268476 218016 268528 218068
rect 268936 218016 268988 218068
rect 269304 218016 269356 218068
rect 270224 218016 270276 218068
rect 270960 218016 271012 218068
rect 272524 218016 272576 218068
rect 277584 218016 277636 218068
rect 278596 218016 278648 218068
rect 280896 218016 280948 218068
rect 281448 218016 281500 218068
rect 281724 218016 281776 218068
rect 282736 218016 282788 218068
rect 283380 218016 283432 218068
rect 284300 218016 284352 218068
rect 285036 218016 285088 218068
rect 285496 218016 285548 218068
rect 287520 218016 287572 218068
rect 288072 218016 288124 218068
rect 289176 218016 289228 218068
rect 289636 218016 289688 218068
rect 290004 218016 290056 218068
rect 291108 218016 291160 218068
rect 293316 218016 293368 218068
rect 293776 218016 293828 218068
rect 298284 218016 298336 218068
rect 299388 218016 299440 218068
rect 299940 218016 299992 218068
rect 300676 218016 300728 218068
rect 301596 218016 301648 218068
rect 302148 218016 302200 218068
rect 305736 218016 305788 218068
rect 306196 218016 306248 218068
rect 306564 218016 306616 218068
rect 307668 218016 307720 218068
rect 308220 218016 308272 218068
rect 308864 218016 308916 218068
rect 309876 218016 309928 218068
rect 310336 218016 310388 218068
rect 312360 218016 312412 218068
rect 312912 218016 312964 218068
rect 314844 218016 314896 218068
rect 315488 218016 315540 218068
rect 317328 218016 317380 218068
rect 317972 218016 318024 218068
rect 318984 218016 319036 218068
rect 320088 218016 320140 218068
rect 322296 218016 322348 218068
rect 322848 218016 322900 218068
rect 323124 218016 323176 218068
rect 323952 218016 324004 218068
rect 324780 218016 324832 218068
rect 325516 218016 325568 218068
rect 326436 218016 326488 218068
rect 326896 218016 326948 218068
rect 330576 218016 330628 218068
rect 331036 218016 331088 218068
rect 332232 218016 332284 218068
rect 333612 218016 333664 218068
rect 334716 218016 334768 218068
rect 335176 218016 335228 218068
rect 337200 218016 337252 218068
rect 337752 218016 337804 218068
rect 338856 218016 338908 218068
rect 339408 218016 339460 218068
rect 339684 218016 339736 218068
rect 340696 218016 340748 218068
rect 345480 218016 345532 218068
rect 347228 218016 347280 218068
rect 347964 218016 348016 218068
rect 349068 218016 349120 218068
rect 349620 218016 349672 218068
rect 350172 218016 350224 218068
rect 352104 218016 352156 218068
rect 353300 218016 353352 218068
rect 356244 218016 356296 218068
rect 357256 218016 357308 218068
rect 357900 218016 357952 218068
rect 358544 218016 358596 218068
rect 359556 218016 359608 218068
rect 360108 218016 360160 218068
rect 360384 218016 360436 218068
rect 361028 218016 361080 218068
rect 367836 218016 367888 218068
rect 368388 218016 368440 218068
rect 371976 218016 372028 218068
rect 372528 218016 372580 218068
rect 372804 218016 372856 218068
rect 373540 218016 373592 218068
rect 374460 218016 374512 218068
rect 375012 218016 375064 218068
rect 376116 218016 376168 218068
rect 376668 218016 376720 218068
rect 378600 218016 378652 218068
rect 379244 218016 379296 218068
rect 381084 218016 381136 218068
rect 382096 218016 382148 218068
rect 385224 218016 385276 218068
rect 386052 218016 386104 218068
rect 389364 218016 389416 218068
rect 390468 218016 390520 218068
rect 392676 218016 392728 218068
rect 393136 218016 393188 218068
rect 393504 218016 393556 218068
rect 394516 218016 394568 218068
rect 395160 218016 395212 218068
rect 395804 218016 395856 218068
rect 397644 218016 397696 218068
rect 401232 218016 401284 218068
rect 401784 218016 401836 218068
rect 402796 218016 402848 218068
rect 403440 218016 403492 218068
rect 403992 218016 404044 218068
rect 405096 218016 405148 218068
rect 405556 218016 405608 218068
rect 409236 218016 409288 218068
rect 409788 218016 409840 218068
rect 410064 218016 410116 218068
rect 410708 218016 410760 218068
rect 413376 218016 413428 218068
rect 413836 218016 413888 218068
rect 420000 218016 420052 218068
rect 420920 218016 420972 218068
rect 424140 218016 424192 218068
rect 426992 218016 427044 218068
rect 427452 218016 427504 218068
rect 428280 218016 428332 218068
rect 429108 218016 429160 218068
rect 430580 218016 430632 218068
rect 432420 218016 432472 218068
rect 433800 218016 433852 218068
rect 434904 218016 434956 218068
rect 436284 218016 436336 218068
rect 436560 218016 436612 218068
rect 437480 218016 437532 218068
rect 438216 218016 438268 218068
rect 438860 218016 438912 218068
rect 439872 218016 439924 218068
rect 440332 218016 440384 218068
rect 453304 218016 453356 218068
rect 455420 218016 455472 218068
rect 455604 218016 455656 218068
rect 457168 218016 457220 218068
rect 463148 218016 463200 218068
rect 464620 218016 464672 218068
rect 467288 218016 467340 218068
rect 467932 218016 467984 218068
rect 492036 218016 492088 218068
rect 505652 218016 505704 218068
rect 512736 218016 512788 218068
rect 572444 218084 572496 218136
rect 572628 218016 572680 218068
rect 604644 218016 604696 218068
rect 563612 217948 563664 218000
rect 572444 217948 572496 218000
rect 675852 217948 675904 218000
rect 676680 217948 676732 218000
rect 131028 217812 131080 217864
rect 197728 217812 197780 217864
rect 523040 217812 523092 217864
rect 524236 217812 524288 217864
rect 535460 217812 535512 217864
rect 536656 217812 536708 217864
rect 116952 217676 117004 217728
rect 189264 217676 189316 217728
rect 525984 217676 526036 217728
rect 526536 217676 526588 217728
rect 533436 217676 533488 217728
rect 598296 217812 598348 217864
rect 602988 217812 603040 217864
rect 603356 217812 603408 217864
rect 613384 217812 613436 217864
rect 103704 217540 103756 217592
rect 178408 217540 178460 217592
rect 530952 217540 531004 217592
rect 598664 217676 598716 217728
rect 604276 217676 604328 217728
rect 604644 217676 604696 217728
rect 616880 217676 616932 217728
rect 538220 217540 538272 217592
rect 539140 217540 539192 217592
rect 545764 217540 545816 217592
rect 606760 217540 606812 217592
rect 92112 217404 92164 217456
rect 170312 217404 170364 217456
rect 526536 217404 526588 217456
rect 93768 217268 93820 217320
rect 171232 217268 171284 217320
rect 535828 217268 535880 217320
rect 598664 217268 598716 217320
rect 598848 217268 598900 217320
rect 601148 217268 601200 217320
rect 601884 217404 601936 217456
rect 628288 217404 628340 217456
rect 602344 217268 602396 217320
rect 602988 217268 603040 217320
rect 603448 217268 603500 217320
rect 436100 217200 436152 217252
rect 437342 217200 437394 217252
rect 447140 217200 447192 217252
rect 448106 217200 448158 217252
rect 448612 217200 448664 217252
rect 449762 217200 449814 217252
rect 469312 217200 469364 217252
rect 470462 217200 470514 217252
rect 489920 217200 489972 217252
rect 491162 217200 491214 217252
rect 498292 217200 498344 217252
rect 499442 217200 499494 217252
rect 502984 217200 503036 217252
rect 503582 217200 503634 217252
rect 511034 217132 511086 217184
rect 562232 217132 562284 217184
rect 562508 217132 562560 217184
rect 562692 217132 562744 217184
rect 563060 217132 563112 217184
rect 599032 217132 599084 217184
rect 600136 217132 600188 217184
rect 604000 217132 604052 217184
rect 503582 217064 503634 217116
rect 608968 216996 609020 217048
rect 609888 216996 609940 217048
rect 614120 216996 614172 217048
rect 574100 216860 574152 216912
rect 597560 216860 597612 216912
rect 598296 216860 598348 216912
rect 600136 216860 600188 216912
rect 594800 216724 594852 216776
rect 612280 216860 612332 216912
rect 601148 216724 601200 216776
rect 623872 216724 623924 216776
rect 675852 216452 675904 216504
rect 676956 216452 677008 216504
rect 649908 215908 649960 215960
rect 663064 215908 663116 215960
rect 676036 215296 676088 215348
rect 676588 215296 676640 215348
rect 575480 214820 575532 214872
rect 622308 214820 622360 214872
rect 574928 214684 574980 214736
rect 616696 214684 616748 214736
rect 617064 214684 617116 214736
rect 617800 214684 617852 214736
rect 619824 214684 619876 214736
rect 620560 214684 620612 214736
rect 621020 214684 621072 214736
rect 621664 214684 621716 214736
rect 622492 214684 622544 214736
rect 623320 214684 623372 214736
rect 630036 214684 630088 214736
rect 632888 214684 632940 214736
rect 574744 214548 574796 214600
rect 625528 214548 625580 214600
rect 600504 214412 600556 214464
rect 601240 214412 601292 214464
rect 605932 214412 605984 214464
rect 606300 214412 606352 214464
rect 607312 214412 607364 214464
rect 607864 214412 607916 214464
rect 611452 214412 611504 214464
rect 611820 214412 611872 214464
rect 616696 214412 616748 214464
rect 624424 214412 624476 214464
rect 653220 214412 653272 214464
rect 660212 214412 660264 214464
rect 663432 214412 663484 214464
rect 665824 214412 665876 214464
rect 626356 214276 626408 214328
rect 628840 214276 628892 214328
rect 35808 214208 35860 214260
rect 39672 214208 39724 214260
rect 646320 214208 646372 214260
rect 653404 214208 653456 214260
rect 627460 213936 627512 213988
rect 629392 213936 629444 213988
rect 663156 213868 663208 213920
rect 663616 213868 663668 213920
rect 646044 213528 646096 213580
rect 646504 213528 646556 213580
rect 652116 213528 652168 213580
rect 654324 213528 654376 213580
rect 574100 213460 574152 213512
rect 594800 213460 594852 213512
rect 574376 213324 574428 213376
rect 612832 213324 612884 213376
rect 574560 213188 574612 213240
rect 616144 213188 616196 213240
rect 643836 213188 643888 213240
rect 666008 213324 666060 213376
rect 654600 213120 654652 213172
rect 657544 213120 657596 213172
rect 654140 212984 654192 213036
rect 654784 212984 654836 213036
rect 662052 212984 662104 213036
rect 664720 212984 664772 213036
rect 645492 212848 645544 212900
rect 651932 212848 651984 212900
rect 650460 212712 650512 212764
rect 651288 212712 651340 212764
rect 658740 212712 658792 212764
rect 659568 212712 659620 212764
rect 664260 212712 664312 212764
rect 665088 212712 665140 212764
rect 632704 212508 632756 212560
rect 634360 212508 634412 212560
rect 630680 212372 630732 212424
rect 631600 212372 631652 212424
rect 35808 211556 35860 211608
rect 41512 211420 41564 211472
rect 35624 211284 35676 211336
rect 41696 211284 41748 211336
rect 35808 211148 35860 211200
rect 40132 211148 40184 211200
rect 578332 211148 578384 211200
rect 580908 211148 580960 211200
rect 633440 211012 633492 211064
rect 633808 211012 633860 211064
rect 35808 209924 35860 209976
rect 40132 209924 40184 209976
rect 35532 209788 35584 209840
rect 40776 209788 40828 209840
rect 579528 209788 579580 209840
rect 582288 209788 582340 209840
rect 35808 208564 35860 208616
rect 40960 208564 41012 208616
rect 581644 208564 581696 208616
rect 632152 209516 632204 209568
rect 578884 208292 578936 208344
rect 589464 208292 589516 208344
rect 35808 207204 35860 207256
rect 40776 207204 40828 207256
rect 580908 206864 580960 206916
rect 589464 206864 589516 206916
rect 579528 205776 579580 205828
rect 581000 205776 581052 205828
rect 582288 205504 582340 205556
rect 589464 205504 589516 205556
rect 35808 204416 35860 204468
rect 41696 204416 41748 204468
rect 35624 204280 35676 204332
rect 41696 204280 41748 204332
rect 579712 204212 579764 204264
rect 589464 204212 589516 204264
rect 578332 202852 578384 202904
rect 580264 202852 580316 202904
rect 581000 202784 581052 202836
rect 589464 202784 589516 202836
rect 578792 200132 578844 200184
rect 590384 200132 590436 200184
rect 580264 199996 580316 200048
rect 589464 199996 589516 200048
rect 579528 198704 579580 198756
rect 589464 198704 589516 198756
rect 578516 195984 578568 196036
rect 589280 195984 589332 196036
rect 579528 194556 579580 194608
rect 589464 194556 589516 194608
rect 579528 191836 579580 191888
rect 589464 191836 589516 191888
rect 579528 190476 579580 190528
rect 590568 190476 590620 190528
rect 579528 187688 579580 187740
rect 589464 187688 589516 187740
rect 579528 186260 579580 186312
rect 589648 186260 589700 186312
rect 579528 184832 579580 184884
rect 589464 184832 589516 184884
rect 42156 183472 42208 183524
rect 42984 183472 43036 183524
rect 42432 182112 42484 182164
rect 43168 182112 43220 182164
rect 579528 182112 579580 182164
rect 589464 182112 589516 182164
rect 578792 180752 578844 180804
rect 590568 180752 590620 180804
rect 578792 178032 578844 178084
rect 589464 178032 589516 178084
rect 579528 177896 579580 177948
rect 589648 177896 589700 177948
rect 579988 175244 580040 175296
rect 589464 175312 589516 175364
rect 668032 174700 668084 174752
rect 670332 174700 670384 174752
rect 578424 174496 578476 174548
rect 589648 174496 589700 174548
rect 667940 173068 667992 173120
rect 669596 173068 669648 173120
rect 578240 172864 578292 172916
rect 579988 172864 580040 172916
rect 580908 172524 580960 172576
rect 589464 172524 589516 172576
rect 580264 171096 580316 171148
rect 589464 171096 589516 171148
rect 578700 169736 578752 169788
rect 580908 169736 580960 169788
rect 582380 168376 582432 168428
rect 589464 168376 589516 168428
rect 668216 168172 668268 168224
rect 670792 168172 670844 168224
rect 578240 167288 578292 167340
rect 580264 167288 580316 167340
rect 579988 167016 580040 167068
rect 589464 167016 589516 167068
rect 579528 166268 579580 166320
rect 589648 166268 589700 166320
rect 579344 165180 579396 165232
rect 582380 165180 582432 165232
rect 667940 164908 667992 164960
rect 669780 164908 669832 164960
rect 582472 164228 582524 164280
rect 589464 164228 589516 164280
rect 578240 163616 578292 163668
rect 579988 163616 580040 163668
rect 580908 162868 580960 162920
rect 589464 162868 589516 162920
rect 578424 162664 578476 162716
rect 582472 162664 582524 162716
rect 675944 161712 675996 161764
rect 679624 161712 679676 161764
rect 580540 161440 580592 161492
rect 589464 161440 589516 161492
rect 580724 160080 580776 160132
rect 589464 160080 589516 160132
rect 578884 158720 578936 158772
rect 580908 158720 580960 158772
rect 585784 158720 585836 158772
rect 589464 158720 589516 158772
rect 587164 157360 587216 157412
rect 589280 157360 589332 157412
rect 578332 154776 578384 154828
rect 580540 154776 580592 154828
rect 584404 154572 584456 154624
rect 589464 154572 589516 154624
rect 583024 153212 583076 153264
rect 589464 153212 589516 153264
rect 578240 152736 578292 152788
rect 580724 152736 580776 152788
rect 580264 151784 580316 151836
rect 589464 151784 589516 151836
rect 578884 150560 578936 150612
rect 585784 150560 585836 150612
rect 585140 149064 585192 149116
rect 589464 149064 589516 149116
rect 668400 149064 668452 149116
rect 670792 149064 670844 149116
rect 579528 148316 579580 148368
rect 587164 148316 587216 148368
rect 578884 146276 578936 146328
rect 585140 146276 585192 146328
rect 584772 144916 584824 144968
rect 589464 144916 589516 144968
rect 579252 144644 579304 144696
rect 584404 144644 584456 144696
rect 585784 143556 585836 143608
rect 589464 143556 589516 143608
rect 579528 143420 579580 143472
rect 583024 143420 583076 143472
rect 587164 142400 587216 142452
rect 589832 142400 589884 142452
rect 580448 140768 580500 140820
rect 589464 140768 589516 140820
rect 578608 140700 578660 140752
rect 580264 140700 580316 140752
rect 668216 140632 668268 140684
rect 670792 140632 670844 140684
rect 583024 139408 583076 139460
rect 589464 139408 589516 139460
rect 578608 139272 578660 139324
rect 589924 139272 589976 139324
rect 579528 138660 579580 138712
rect 588544 138660 588596 138712
rect 668584 137980 668636 138032
rect 670148 137980 670200 138032
rect 579068 137300 579120 137352
rect 584772 137300 584824 137352
rect 584588 136620 584640 136672
rect 589464 136620 589516 136672
rect 580264 134512 580316 134564
rect 589464 134512 589516 134564
rect 585968 132472 586020 132524
rect 589464 132472 589516 132524
rect 581828 131248 581880 131300
rect 589464 131248 589516 131300
rect 578884 131112 578936 131164
rect 585784 131112 585836 131164
rect 667940 130636 667992 130688
rect 669964 130636 670016 130688
rect 583392 129140 583444 129192
rect 590384 129140 590436 129192
rect 579528 129004 579580 129056
rect 587164 129004 587216 129056
rect 668768 128596 668820 128648
rect 670792 128596 670844 128648
rect 587808 126964 587860 127016
rect 589464 126964 589516 127016
rect 578332 125604 578384 125656
rect 580448 125604 580500 125656
rect 676036 125400 676088 125452
rect 676404 125400 676456 125452
rect 579068 124856 579120 124908
rect 587808 124856 587860 124908
rect 578700 124108 578752 124160
rect 583024 124108 583076 124160
rect 584404 122816 584456 122868
rect 589464 122816 589516 122868
rect 578884 122136 578936 122188
rect 584588 122136 584640 122188
rect 580632 122000 580684 122052
rect 590108 122000 590160 122052
rect 587348 121456 587400 121508
rect 589280 121456 589332 121508
rect 583208 120708 583260 120760
rect 590568 120708 590620 120760
rect 578516 118532 578568 118584
rect 580264 118532 580316 118584
rect 579528 116900 579580 116952
rect 583392 116900 583444 116952
rect 675852 116628 675904 116680
rect 678244 116628 678296 116680
rect 585784 115948 585836 116000
rect 589464 115948 589516 116000
rect 584588 115200 584640 115252
rect 589648 115200 589700 115252
rect 579252 114452 579304 114504
rect 581644 114452 581696 114504
rect 583024 113160 583076 113212
rect 589464 113160 589516 113212
rect 579528 112820 579580 112872
rect 585968 112820 586020 112872
rect 586152 112412 586204 112464
rect 590108 112412 590160 112464
rect 581644 110440 581696 110492
rect 589464 110440 589516 110492
rect 579344 110236 579396 110288
rect 581828 110236 581880 110288
rect 580448 109080 580500 109132
rect 589464 109080 589516 109132
rect 578332 108944 578384 108996
rect 580632 108944 580684 108996
rect 667940 107992 667992 108044
rect 670148 107992 670200 108044
rect 582288 107652 582340 107704
rect 589464 107652 589516 107704
rect 580264 106292 580316 106344
rect 589464 106292 589516 106344
rect 668400 106156 668452 106208
rect 670792 106156 670844 106208
rect 579344 105612 579396 105664
rect 582288 105612 582340 105664
rect 587164 104864 587216 104916
rect 589832 104864 589884 104916
rect 668308 104796 668360 104848
rect 670792 104796 670844 104848
rect 578516 103368 578568 103420
rect 588728 103368 588780 103420
rect 579160 102076 579212 102128
rect 584404 102076 584456 102128
rect 584404 100104 584456 100156
rect 589464 100104 589516 100156
rect 578608 99968 578660 100020
rect 587348 99968 587400 100020
rect 592684 99968 592736 100020
rect 667940 99968 667992 100020
rect 622308 99288 622360 99340
rect 630772 99288 630824 99340
rect 579528 99220 579580 99272
rect 583208 99220 583260 99272
rect 623688 99152 623740 99204
rect 633440 99152 633492 99204
rect 577504 99084 577556 99136
rect 595260 99084 595312 99136
rect 624608 99016 624660 99068
rect 635004 99016 635056 99068
rect 625068 98880 625120 98932
rect 636292 98880 636344 98932
rect 629024 98744 629076 98796
rect 643652 98744 643704 98796
rect 647148 98744 647200 98796
rect 661960 98744 662012 98796
rect 630496 98608 630548 98660
rect 646596 98608 646648 98660
rect 631416 98268 631468 98320
rect 642180 98268 642232 98320
rect 633624 98132 633676 98184
rect 640708 98132 640760 98184
rect 618720 97928 618772 97980
rect 625804 97928 625856 97980
rect 629760 97928 629812 97980
rect 645308 97996 645360 98048
rect 659200 97928 659252 97980
rect 664168 97928 664220 97980
rect 628288 97792 628340 97844
rect 631416 97792 631468 97844
rect 632704 97792 632756 97844
rect 647516 97792 647568 97844
rect 655244 97792 655296 97844
rect 659752 97792 659804 97844
rect 659936 97792 659988 97844
rect 665364 97792 665416 97844
rect 631232 97656 631284 97708
rect 647332 97656 647384 97708
rect 651840 97656 651892 97708
rect 659568 97656 659620 97708
rect 627552 97520 627604 97572
rect 633624 97520 633676 97572
rect 633808 97520 633860 97572
rect 637764 97520 637816 97572
rect 643008 97520 643060 97572
rect 655244 97520 655296 97572
rect 655428 97520 655480 97572
rect 662512 97520 662564 97572
rect 605472 97384 605524 97436
rect 611912 97384 611964 97436
rect 612648 97384 612700 97436
rect 620284 97384 620336 97436
rect 621664 97384 621716 97436
rect 629300 97384 629352 97436
rect 631968 97384 632020 97436
rect 648620 97384 648672 97436
rect 653956 97384 654008 97436
rect 655244 97384 655296 97436
rect 658188 97384 658240 97436
rect 663064 97384 663116 97436
rect 623136 97248 623188 97300
rect 632060 97248 632112 97300
rect 633256 97248 633308 97300
rect 620100 97112 620152 97164
rect 626448 97112 626500 97164
rect 634176 97112 634228 97164
rect 649080 97112 649132 97164
rect 650368 97248 650420 97300
rect 658280 97248 658332 97300
rect 650552 97112 650604 97164
rect 656808 97112 656860 97164
rect 661408 97112 661460 97164
rect 626080 96976 626132 97028
rect 633808 96976 633860 97028
rect 634728 96976 634780 97028
rect 647056 96976 647108 97028
rect 597652 96908 597704 96960
rect 598204 96908 598256 96960
rect 600320 96908 600372 96960
rect 601148 96908 601200 96960
rect 606208 96908 606260 96960
rect 607128 96908 607180 96960
rect 615776 96908 615828 96960
rect 616788 96908 616840 96960
rect 656716 96908 656768 96960
rect 660120 96908 660172 96960
rect 612096 96840 612148 96892
rect 612648 96840 612700 96892
rect 617248 96840 617300 96892
rect 618168 96840 618220 96892
rect 626816 96840 626868 96892
rect 639236 96840 639288 96892
rect 644296 96840 644348 96892
rect 658832 96772 658884 96824
rect 609152 96704 609204 96756
rect 609704 96704 609756 96756
rect 654784 96704 654836 96756
rect 655428 96704 655480 96756
rect 640064 96568 640116 96620
rect 645124 96568 645176 96620
rect 646412 96568 646464 96620
rect 652208 96568 652260 96620
rect 652576 96568 652628 96620
rect 664352 96568 664404 96620
rect 638592 96432 638644 96484
rect 641352 96432 641404 96484
rect 641536 96432 641588 96484
rect 648068 96432 648120 96484
rect 648896 96432 648948 96484
rect 664536 96432 664588 96484
rect 637580 96296 637632 96348
rect 660672 96296 660724 96348
rect 645492 96160 645544 96212
rect 647884 96160 647936 96212
rect 649264 96160 649316 96212
rect 663800 96160 663852 96212
rect 640524 96092 640576 96144
rect 644940 96092 644992 96144
rect 591304 96024 591356 96076
rect 602620 96024 602672 96076
rect 610624 96024 610676 96076
rect 621664 96024 621716 96076
rect 645768 96024 645820 96076
rect 648068 96024 648120 96076
rect 648620 96024 648672 96076
rect 663984 96024 664036 96076
rect 594064 95888 594116 95940
rect 668124 95888 668176 95940
rect 598940 95752 598992 95804
rect 599676 95752 599728 95804
rect 639052 95752 639104 95804
rect 648620 95752 648672 95804
rect 653312 95752 653364 95804
rect 665180 95752 665232 95804
rect 645124 95616 645176 95668
rect 652024 95616 652076 95668
rect 641352 95412 641404 95464
rect 643468 95412 643520 95464
rect 647884 95412 647936 95464
rect 648068 95344 648120 95396
rect 656164 95480 656216 95532
rect 647700 95276 647752 95328
rect 578332 95140 578384 95192
rect 584588 95140 584640 95192
rect 620928 95140 620980 95192
rect 625436 95140 625488 95192
rect 647056 95140 647108 95192
rect 650276 95140 650328 95192
rect 616512 94936 616564 94988
rect 624976 94936 625028 94988
rect 607680 94460 607732 94512
rect 620652 94460 620704 94512
rect 619548 93780 619600 93832
rect 626264 93780 626316 93832
rect 647516 93712 647568 93764
rect 648252 93712 648304 93764
rect 651288 93576 651340 93628
rect 654692 93576 654744 93628
rect 579252 93372 579304 93424
rect 586152 93372 586204 93424
rect 609704 93100 609756 93152
rect 618628 93100 618680 93152
rect 617984 92420 618036 92472
rect 626448 92420 626500 92472
rect 647700 92420 647752 92472
rect 655428 92420 655480 92472
rect 606944 91740 606996 91792
rect 622400 91740 622452 91792
rect 578608 91128 578660 91180
rect 585784 91128 585836 91180
rect 618168 91128 618220 91180
rect 611268 90992 611320 91044
rect 618168 90992 618220 91044
rect 626448 90992 626500 91044
rect 648620 90788 648672 90840
rect 655428 90788 655480 90840
rect 620652 89632 620704 89684
rect 625436 89632 625488 89684
rect 649724 88748 649776 88800
rect 658556 88748 658608 88800
rect 662328 88748 662380 88800
rect 664168 88748 664220 88800
rect 656164 88612 656216 88664
rect 657452 88612 657504 88664
rect 579252 88272 579304 88324
rect 589924 88272 589976 88324
rect 622400 88272 622452 88324
rect 626448 88272 626500 88324
rect 655244 88272 655296 88324
rect 658464 88272 658516 88324
rect 618168 88136 618220 88188
rect 626264 88136 626316 88188
rect 648436 86980 648488 87032
rect 662512 86980 662564 87032
rect 578332 86912 578384 86964
rect 580448 86912 580500 86964
rect 656716 86844 656768 86896
rect 659568 86844 659620 86896
rect 652024 86708 652076 86760
rect 660120 86708 660172 86760
rect 647884 86572 647936 86624
rect 661408 86572 661460 86624
rect 652208 86436 652260 86488
rect 657176 86436 657228 86488
rect 621664 86300 621716 86352
rect 626448 86300 626500 86352
rect 656348 86300 656400 86352
rect 660672 86300 660724 86352
rect 609888 85484 609940 85536
rect 626448 85484 626500 85536
rect 618628 85348 618680 85400
rect 625252 85348 625304 85400
rect 608508 84124 608560 84176
rect 626448 84124 626500 84176
rect 579252 83988 579304 84040
rect 581644 83988 581696 84040
rect 578884 82764 578936 82816
rect 583024 82764 583076 82816
rect 579252 82084 579304 82136
rect 587164 82084 587216 82136
rect 628748 81064 628800 81116
rect 642456 81064 642508 81116
rect 615408 80928 615460 80980
rect 646320 80928 646372 80980
rect 613844 80792 613896 80844
rect 647332 80792 647384 80844
rect 595444 80656 595496 80708
rect 636752 80656 636804 80708
rect 629208 79976 629260 80028
rect 633440 79976 633492 80028
rect 614028 79432 614080 79484
rect 646044 79432 646096 79484
rect 583024 79296 583076 79348
rect 600320 79296 600372 79348
rect 612648 79296 612700 79348
rect 648620 79296 648672 79348
rect 578240 78072 578292 78124
rect 580264 78072 580316 78124
rect 633440 78072 633492 78124
rect 645308 78072 645360 78124
rect 631048 77936 631100 77988
rect 643100 77936 643152 77988
rect 628472 77596 628524 77648
rect 632796 77596 632848 77648
rect 624424 77256 624476 77308
rect 628472 77392 628524 77444
rect 625804 77256 625856 77308
rect 631048 77256 631100 77308
rect 620284 76780 620336 76832
rect 648988 76780 649040 76832
rect 612004 76644 612056 76696
rect 662420 76644 662472 76696
rect 587164 76508 587216 76560
rect 668216 76508 668268 76560
rect 616788 75420 616840 75472
rect 646688 75420 646740 75472
rect 607128 75284 607180 75336
rect 646504 75284 646556 75336
rect 578884 75148 578936 75200
rect 666560 75148 666612 75200
rect 579528 73108 579580 73160
rect 588544 73108 588596 73160
rect 578516 71544 578568 71596
rect 584404 71544 584456 71596
rect 579528 66852 579580 66904
rect 625988 66852 626040 66904
rect 579528 64812 579580 64864
rect 592684 64812 592736 64864
rect 579528 62024 579580 62076
rect 587164 62024 587216 62076
rect 578332 59984 578384 60036
rect 624424 59984 624476 60036
rect 576124 58760 576176 58812
rect 603080 58760 603132 58812
rect 577504 58624 577556 58676
rect 604460 58624 604512 58676
rect 579528 57876 579580 57928
rect 594064 57876 594116 57928
rect 574928 57196 574980 57248
rect 600504 57196 600556 57248
rect 574744 55972 574796 56024
rect 598940 55972 598992 56024
rect 574468 55836 574520 55888
rect 601884 55836 601936 55888
rect 596456 55156 596508 55208
rect 597836 55020 597888 55072
rect 597652 54884 597704 54936
rect 599124 54748 599176 54800
rect 623044 54612 623096 54664
rect 463884 53592 463936 53644
rect 464528 53592 464580 53644
rect 463608 53456 463660 53508
rect 464804 53592 464856 53644
rect 625804 54476 625856 54528
rect 596180 54340 596232 54392
rect 474280 53592 474332 53644
rect 474464 53592 474516 53644
rect 464988 53456 465040 53508
rect 583024 54204 583076 54256
rect 580448 54068 580500 54120
rect 574744 53932 574796 53984
rect 475200 53592 475252 53644
rect 475384 53592 475436 53644
rect 480076 53592 480128 53644
rect 462228 53320 462280 53372
rect 574928 53796 574980 53848
rect 48964 53184 49016 53236
rect 129004 53184 129056 53236
rect 463148 53184 463200 53236
rect 468300 53184 468352 53236
rect 312360 53116 312412 53168
rect 313740 53116 313792 53168
rect 316316 53116 316368 53168
rect 317696 53116 317748 53168
rect 46204 53048 46256 53100
rect 130384 53048 130436 53100
rect 461308 53048 461360 53100
rect 480076 53048 480128 53100
rect 460388 52912 460440 52964
rect 474464 52912 474516 52964
rect 459146 52776 459198 52828
rect 464804 52776 464856 52828
rect 465126 52776 465178 52828
rect 475384 52776 475436 52828
rect 465908 52640 465960 52692
rect 474280 52640 474332 52692
rect 51724 51960 51776 52012
rect 129372 51960 129424 52012
rect 50528 51824 50580 51876
rect 130568 51824 130620 51876
rect 47584 51688 47636 51740
rect 129188 51688 129240 51740
rect 145380 51688 145432 51740
rect 306012 51688 306064 51740
rect 318340 50464 318392 50516
rect 458364 50464 458416 50516
rect 45468 50328 45520 50380
rect 129648 50328 129700 50380
rect 314016 50328 314068 50380
rect 458180 50328 458232 50380
rect 522948 50328 523000 50380
rect 544016 50328 544068 50380
rect 49148 48968 49200 49020
rect 131028 48968 131080 49020
rect 129188 47812 129240 47864
rect 131580 47812 131632 47864
rect 625988 46452 626040 46504
rect 661776 46452 661828 46504
rect 129648 46044 129700 46096
rect 132040 46044 132092 46096
rect 130384 45500 130436 45552
rect 132224 45500 132276 45552
rect 131304 45364 131356 45416
rect 132960 45364 133012 45416
rect 129372 45296 129424 45348
rect 130936 45296 130988 45348
rect 43812 45160 43864 45212
rect 130936 45064 130988 45116
rect 129372 44956 129424 45008
rect 128360 44820 128412 44872
rect 131396 44684 131448 44736
rect 129004 44616 129056 44668
rect 50344 44412 50396 44464
rect 128360 44412 128412 44464
rect 43628 44276 43680 44328
rect 131580 44276 131632 44328
rect 132040 44208 132092 44260
rect 132224 44208 132276 44260
rect 132592 44364 132644 44416
rect 132960 44252 133012 44304
rect 43444 44140 43496 44192
rect 131396 44140 131448 44192
rect 129372 44004 129424 44056
rect 440240 43800 440292 43852
rect 441068 43800 441120 43852
rect 410892 42848 410944 42900
rect 415584 42848 415636 42900
rect 187332 42780 187384 42832
rect 255872 42780 255924 42832
rect 310428 42712 310480 42764
rect 364524 42712 364576 42764
rect 361764 42440 361816 42492
rect 431224 42712 431276 42764
rect 441068 42712 441120 42764
rect 449164 42712 449216 42764
rect 453580 42712 453632 42764
rect 464344 42712 464396 42764
rect 364892 42576 364944 42628
rect 427084 42576 427136 42628
rect 441252 42576 441304 42628
rect 446404 42576 446456 42628
rect 454684 42576 454736 42628
rect 462964 42576 463016 42628
rect 364524 42304 364576 42356
rect 410892 42440 410944 42492
rect 415584 42304 415636 42356
rect 429108 42440 429160 42492
rect 454500 42440 454552 42492
rect 463700 42440 463752 42492
rect 661408 42129 661460 42181
rect 427084 41964 427136 42016
rect 431224 41964 431276 42016
rect 441068 41964 441120 42016
rect 446404 41964 446456 42016
rect 454500 41964 454552 42016
rect 441252 41828 441304 41880
rect 429108 41692 429160 41744
rect 454684 41828 454736 41880
rect 449164 41692 449216 41744
rect 453580 41692 453632 41744
<< metal2 >>
rect 703694 897668 703722 897804
rect 704154 897668 704182 897804
rect 704614 897668 704642 897804
rect 705074 897668 705102 897804
rect 705534 897668 705562 897804
rect 705994 897668 706022 897804
rect 706454 897668 706482 897804
rect 706914 897668 706942 897804
rect 707374 897668 707402 897804
rect 707834 897668 707862 897804
rect 708294 897668 708322 897804
rect 708754 897668 708782 897804
rect 709214 897668 709242 897804
rect 676034 897152 676090 897161
rect 676034 897087 676036 897096
rect 676088 897087 676090 897096
rect 676036 897058 676088 897064
rect 652024 897048 652076 897054
rect 652024 896990 652076 896996
rect 651472 868896 651524 868902
rect 651472 868838 651524 868844
rect 651484 868601 651512 868838
rect 651470 868592 651526 868601
rect 651470 868527 651526 868536
rect 652036 867649 652064 896990
rect 675850 896744 675906 896753
rect 675850 896679 675906 896688
rect 675864 895830 675892 896679
rect 676034 896336 676090 896345
rect 676034 896271 676090 896280
rect 654784 895824 654836 895830
rect 654784 895766 654836 895772
rect 675852 895824 675904 895830
rect 675852 895766 675904 895772
rect 653404 880524 653456 880530
rect 653404 880466 653456 880472
rect 652022 867640 652078 867649
rect 652022 867575 652078 867584
rect 651472 866652 651524 866658
rect 651472 866594 651524 866600
rect 651484 866289 651512 866594
rect 651470 866280 651526 866289
rect 651470 866215 651526 866224
rect 653416 865230 653444 880466
rect 654796 868902 654824 895766
rect 676048 895694 676076 896271
rect 672724 895688 672776 895694
rect 672724 895630 672776 895636
rect 676036 895688 676088 895694
rect 676036 895630 676088 895636
rect 672172 894464 672224 894470
rect 672172 894406 672224 894412
rect 671988 893036 672040 893042
rect 671988 892978 672040 892984
rect 670976 892900 671028 892906
rect 670976 892842 671028 892848
rect 657544 869440 657596 869446
rect 657544 869382 657596 869388
rect 654784 868896 654836 868902
rect 654784 868838 654836 868844
rect 654140 868080 654192 868086
rect 654140 868022 654192 868028
rect 651380 865224 651432 865230
rect 651378 865192 651380 865201
rect 653404 865224 653456 865230
rect 651432 865192 651434 865201
rect 653404 865166 653456 865172
rect 651378 865127 651434 865136
rect 651472 863864 651524 863870
rect 651470 863832 651472 863841
rect 651524 863832 651526 863841
rect 651470 863767 651526 863776
rect 654152 862510 654180 868022
rect 657556 863870 657584 869382
rect 657544 863864 657596 863870
rect 657544 863806 657596 863812
rect 651472 862504 651524 862510
rect 651472 862446 651524 862452
rect 654140 862504 654192 862510
rect 654140 862446 654192 862452
rect 651484 862345 651512 862446
rect 651470 862336 651526 862345
rect 651470 862271 651526 862280
rect 8588 818380 8616 818516
rect 9048 818380 9076 818516
rect 9508 818380 9536 818516
rect 9968 818380 9996 818516
rect 10428 818380 10456 818516
rect 10888 818380 10916 818516
rect 11348 818380 11376 818516
rect 11808 818380 11836 818516
rect 12268 818380 12296 818516
rect 12728 818380 12756 818516
rect 13188 818380 13216 818516
rect 13648 818380 13676 818516
rect 14108 818380 14136 818516
rect 35622 818000 35678 818009
rect 35622 817935 35678 817944
rect 35636 817154 35664 817935
rect 35806 817320 35862 817329
rect 35806 817255 35862 817264
rect 35820 817154 35848 817255
rect 35624 817148 35676 817154
rect 35624 817090 35676 817096
rect 35808 817148 35860 817154
rect 35808 817090 35860 817096
rect 44824 817148 44876 817154
rect 44824 817090 44876 817096
rect 35622 816912 35678 816921
rect 35622 816847 35678 816856
rect 35636 815794 35664 816847
rect 35806 816096 35862 816105
rect 35806 816031 35862 816040
rect 35624 815788 35676 815794
rect 35624 815730 35676 815736
rect 35820 815658 35848 816031
rect 43444 815788 43496 815794
rect 43444 815730 43496 815736
rect 35808 815652 35860 815658
rect 35808 815594 35860 815600
rect 35622 815280 35678 815289
rect 35622 815215 35678 815224
rect 35636 814298 35664 815215
rect 35806 814464 35862 814473
rect 35806 814399 35808 814408
rect 35860 814399 35862 814408
rect 35808 814370 35860 814376
rect 35624 814292 35676 814298
rect 35624 814234 35676 814240
rect 41326 813648 41382 813657
rect 41326 813583 41382 813592
rect 41340 812870 41368 813583
rect 41328 812864 41380 812870
rect 31666 812832 31722 812841
rect 41328 812806 41380 812812
rect 43260 812864 43312 812870
rect 43260 812806 43312 812812
rect 31666 812767 31722 812776
rect 31022 809976 31078 809985
rect 31022 809911 31078 809920
rect 30286 809160 30342 809169
rect 30286 809095 30342 809104
rect 30300 805254 30328 809095
rect 30288 805248 30340 805254
rect 30288 805190 30340 805196
rect 31036 801106 31064 809911
rect 31680 809402 31708 812767
rect 41326 812424 41382 812433
rect 41326 812359 41382 812368
rect 35162 812016 35218 812025
rect 35162 811951 35218 811960
rect 32218 811200 32274 811209
rect 32218 811135 32274 811144
rect 31668 809396 31720 809402
rect 31668 809338 31720 809344
rect 32232 802466 32260 811135
rect 33782 809398 33838 809407
rect 33782 809333 33838 809342
rect 32220 802460 32272 802466
rect 32220 802402 32272 802408
rect 33796 801242 33824 809333
rect 35176 802505 35204 811951
rect 39302 811608 39358 811617
rect 39302 811543 39358 811552
rect 35162 802496 35218 802505
rect 35162 802431 35218 802440
rect 33784 801236 33836 801242
rect 33784 801178 33836 801184
rect 31024 801100 31076 801106
rect 31024 801042 31076 801048
rect 39316 800601 39344 811543
rect 41340 811510 41368 812359
rect 41328 811504 41380 811510
rect 41328 811446 41380 811452
rect 41788 811504 41840 811510
rect 41788 811446 41840 811452
rect 41800 811345 41828 811446
rect 41786 811336 41842 811345
rect 41786 811271 41842 811280
rect 41786 810792 41842 810801
rect 41786 810727 41842 810736
rect 41326 808752 41382 808761
rect 41326 808687 41328 808696
rect 41380 808687 41382 808696
rect 41328 808658 41380 808664
rect 41142 808344 41198 808353
rect 41142 808279 41198 808288
rect 41156 807362 41184 808279
rect 41326 807528 41382 807537
rect 41326 807463 41328 807472
rect 41380 807463 41382 807472
rect 41328 807434 41380 807440
rect 41144 807356 41196 807362
rect 41144 807298 41196 807304
rect 41142 806712 41198 806721
rect 41142 806647 41198 806656
rect 41156 806002 41184 806647
rect 41326 806304 41382 806313
rect 41326 806239 41382 806248
rect 41340 806138 41368 806239
rect 41328 806132 41380 806138
rect 41328 806074 41380 806080
rect 41144 805996 41196 806002
rect 41144 805938 41196 805944
rect 41800 805633 41828 810727
rect 42154 810384 42210 810393
rect 42154 810319 42210 810328
rect 41970 807936 42026 807945
rect 41970 807871 42026 807880
rect 41786 805624 41842 805633
rect 41786 805559 41842 805568
rect 41984 804817 42012 807871
rect 41970 804808 42026 804817
rect 41970 804743 42026 804752
rect 42168 804658 42196 810319
rect 42432 809396 42484 809402
rect 42432 809338 42484 809344
rect 42444 808694 42472 809338
rect 41984 804630 42196 804658
rect 42260 808666 42472 808694
rect 43076 808716 43128 808722
rect 41984 804545 42012 804630
rect 42260 804554 42288 808666
rect 43076 808658 43128 808664
rect 42892 807492 42944 807498
rect 42892 807434 42944 807440
rect 42708 805248 42760 805254
rect 42708 805190 42760 805196
rect 42720 804554 42748 805190
rect 41970 804536 42026 804545
rect 41970 804471 42026 804480
rect 42168 804526 42288 804554
rect 42444 804526 42748 804554
rect 41788 802460 41840 802466
rect 41788 802402 41840 802408
rect 40500 801100 40552 801106
rect 40500 801042 40552 801048
rect 40512 800737 40540 801042
rect 40498 800728 40554 800737
rect 40498 800663 40554 800672
rect 39302 800592 39358 800601
rect 39302 800527 39358 800536
rect 41800 800329 41828 802402
rect 42168 801794 42196 804526
rect 42168 801766 42380 801794
rect 41786 800320 41842 800329
rect 41786 800255 41842 800264
rect 41786 799912 41842 799921
rect 41786 799847 41842 799856
rect 41800 799445 41828 799847
rect 42352 797619 42380 801766
rect 42182 797591 42380 797619
rect 42154 797328 42210 797337
rect 42154 797263 42210 797272
rect 42168 796960 42196 797263
rect 42248 796884 42300 796890
rect 42248 796826 42300 796832
rect 42260 795779 42288 796826
rect 42444 795954 42472 804526
rect 42616 801236 42668 801242
rect 42616 801178 42668 801184
rect 42628 796890 42656 801178
rect 42616 796884 42668 796890
rect 42616 796826 42668 796832
rect 42182 795751 42288 795779
rect 42352 795926 42472 795954
rect 42154 795424 42210 795433
rect 42154 795359 42210 795368
rect 42168 795124 42196 795359
rect 41786 794880 41842 794889
rect 41786 794815 41842 794824
rect 41800 794580 41828 794815
rect 42352 794458 42380 795926
rect 42708 794776 42760 794782
rect 42708 794718 42760 794724
rect 42168 794430 42380 794458
rect 42168 793900 42196 794430
rect 42720 793529 42748 794718
rect 42062 793520 42118 793529
rect 42062 793455 42118 793464
rect 42706 793520 42762 793529
rect 42706 793455 42762 793464
rect 42076 793288 42104 793455
rect 41786 793112 41842 793121
rect 41786 793047 41842 793056
rect 41800 792744 41828 793047
rect 42430 792704 42486 792713
rect 42430 792639 42486 792648
rect 42246 791344 42302 791353
rect 42246 791279 42302 791288
rect 42062 790664 42118 790673
rect 42062 790599 42118 790608
rect 42076 790228 42104 790599
rect 42260 789750 42288 791279
rect 42248 789744 42300 789750
rect 42248 789686 42300 789692
rect 42444 789630 42472 792639
rect 42614 791616 42670 791625
rect 42614 791551 42670 791560
rect 42182 789602 42472 789630
rect 42248 789540 42300 789546
rect 42248 789482 42300 789488
rect 42260 789290 42288 789482
rect 42628 789426 42656 791551
rect 42168 789262 42288 789290
rect 42352 789398 42656 789426
rect 42168 788936 42196 789262
rect 42352 788406 42380 789398
rect 42182 788378 42380 788406
rect 42246 788216 42302 788225
rect 42246 788151 42302 788160
rect 41786 786856 41842 786865
rect 41786 786791 41842 786800
rect 41800 786556 41828 786791
rect 41786 786176 41842 786185
rect 41786 786111 41842 786120
rect 41800 785944 41828 786111
rect 42260 785278 42288 788151
rect 42616 786684 42668 786690
rect 42616 786626 42668 786632
rect 42182 785250 42288 785278
rect 42628 784734 42656 786626
rect 42182 784706 42656 784734
rect 8588 775132 8616 775268
rect 9048 775132 9076 775268
rect 9508 775132 9536 775268
rect 9968 775132 9996 775268
rect 10428 775132 10456 775268
rect 10888 775132 10916 775268
rect 11348 775132 11376 775268
rect 11808 775132 11836 775268
rect 12268 775132 12296 775268
rect 12728 775132 12756 775268
rect 13188 775132 13216 775268
rect 13648 775132 13676 775268
rect 14108 775132 14136 775268
rect 35806 774752 35862 774761
rect 35806 774687 35862 774696
rect 35820 774246 35848 774687
rect 35808 774240 35860 774246
rect 35808 774182 35860 774188
rect 41696 774240 41748 774246
rect 42064 774240 42116 774246
rect 41748 774188 42064 774194
rect 41696 774182 42116 774188
rect 41708 774166 42104 774182
rect 35254 773936 35310 773945
rect 35254 773871 35310 773880
rect 35268 772886 35296 773871
rect 35622 773528 35678 773537
rect 35622 773463 35678 773472
rect 35440 773424 35492 773430
rect 35440 773366 35492 773372
rect 35452 773129 35480 773366
rect 35438 773120 35494 773129
rect 35438 773055 35494 773064
rect 35636 773022 35664 773463
rect 41512 773424 41564 773430
rect 41512 773366 41564 773372
rect 35808 773152 35860 773158
rect 35806 773120 35808 773129
rect 41524 773129 41552 773366
rect 41708 773226 42104 773242
rect 41696 773220 42116 773226
rect 41748 773214 42064 773220
rect 41696 773162 41748 773168
rect 42064 773162 42116 773168
rect 35860 773120 35862 773129
rect 35806 773055 35862 773064
rect 41510 773120 41566 773129
rect 41708 773090 42104 773106
rect 41510 773055 41566 773064
rect 41696 773084 42116 773090
rect 41748 773078 42064 773084
rect 41696 773026 41748 773032
rect 42064 773026 42116 773032
rect 35624 773016 35676 773022
rect 35624 772958 35676 772964
rect 35256 772880 35308 772886
rect 35256 772822 35308 772828
rect 41696 772880 41748 772886
rect 42064 772880 42116 772886
rect 41748 772828 42064 772834
rect 41696 772822 42116 772828
rect 41708 772806 42104 772822
rect 35622 772304 35678 772313
rect 35622 772239 35678 772248
rect 35636 771594 35664 772239
rect 35806 771896 35862 771905
rect 35806 771831 35808 771840
rect 35860 771831 35862 771840
rect 39488 771860 39540 771866
rect 35808 771802 35860 771808
rect 39488 771802 39540 771808
rect 35624 771588 35676 771594
rect 35624 771530 35676 771536
rect 35806 771488 35862 771497
rect 35806 771423 35808 771432
rect 35860 771423 35862 771432
rect 35808 771394 35860 771400
rect 35622 771080 35678 771089
rect 35622 771015 35678 771024
rect 35636 770098 35664 771015
rect 35806 770672 35862 770681
rect 35806 770607 35862 770616
rect 39118 770672 39174 770681
rect 39118 770607 39174 770616
rect 35820 770506 35848 770607
rect 39132 770506 39160 770607
rect 35808 770500 35860 770506
rect 35808 770442 35860 770448
rect 39120 770500 39172 770506
rect 39120 770442 39172 770448
rect 39500 770273 39528 771802
rect 42064 771656 42116 771662
rect 41708 771604 42064 771610
rect 41708 771598 42116 771604
rect 41708 771594 42104 771598
rect 41696 771588 42104 771594
rect 41748 771582 42104 771588
rect 41696 771530 41748 771536
rect 41708 771458 42104 771474
rect 41696 771452 42116 771458
rect 41748 771446 42064 771452
rect 41696 771394 41748 771400
rect 42904 771434 42932 807434
rect 43088 790673 43116 808658
rect 43074 790664 43130 790673
rect 43074 790599 43130 790608
rect 42064 771394 42116 771400
rect 42720 771406 42932 771434
rect 35806 770264 35862 770273
rect 35806 770199 35808 770208
rect 35860 770199 35862 770208
rect 39486 770264 39542 770273
rect 39486 770199 39542 770208
rect 39856 770228 39908 770234
rect 35808 770170 35860 770176
rect 39856 770170 39908 770176
rect 35624 770092 35676 770098
rect 35624 770034 35676 770040
rect 39868 769457 39896 770170
rect 41708 770098 42104 770114
rect 41696 770092 42116 770098
rect 41748 770086 42064 770092
rect 41696 770034 41748 770040
rect 42064 770034 42116 770040
rect 35806 769448 35862 769457
rect 35806 769383 35862 769392
rect 39854 769448 39910 769457
rect 39854 769383 39910 769392
rect 35622 769040 35678 769049
rect 35820 769010 35848 769383
rect 35622 768975 35678 768984
rect 35808 769004 35860 769010
rect 35636 768738 35664 768975
rect 35808 768946 35860 768952
rect 41696 769004 41748 769010
rect 41696 768946 41748 768952
rect 35808 768868 35860 768874
rect 35808 768810 35860 768816
rect 39764 768868 39816 768874
rect 39764 768810 39816 768816
rect 35624 768732 35676 768738
rect 35624 768674 35676 768680
rect 35820 768641 35848 768810
rect 35806 768632 35862 768641
rect 35806 768567 35862 768576
rect 35162 768224 35218 768233
rect 35162 768159 35218 768168
rect 32402 767816 32458 767825
rect 32402 767751 32458 767760
rect 32416 759694 32444 767751
rect 33782 767000 33838 767009
rect 33782 766935 33838 766944
rect 32404 759688 32456 759694
rect 32404 759630 32456 759636
rect 33796 758334 33824 766935
rect 35176 759830 35204 768159
rect 35806 767408 35862 767417
rect 35806 767343 35808 767352
rect 35860 767343 35862 767352
rect 36544 767372 36596 767378
rect 35808 767314 35860 767320
rect 36544 767314 36596 767320
rect 35806 766184 35862 766193
rect 35806 766119 35808 766128
rect 35860 766119 35862 766128
rect 35808 766090 35860 766096
rect 35806 765776 35862 765785
rect 35806 765711 35862 765720
rect 35820 764862 35848 765711
rect 35808 764856 35860 764862
rect 35808 764798 35860 764804
rect 35808 764584 35860 764590
rect 35806 764552 35808 764561
rect 35860 764552 35862 764561
rect 35806 764487 35862 764496
rect 35622 764144 35678 764153
rect 35622 764079 35678 764088
rect 35636 763434 35664 764079
rect 35806 763736 35862 763745
rect 35806 763671 35862 763680
rect 35624 763428 35676 763434
rect 35624 763370 35676 763376
rect 35820 763230 35848 763671
rect 35808 763224 35860 763230
rect 35808 763166 35860 763172
rect 35806 762920 35862 762929
rect 35806 762855 35862 762864
rect 35820 761938 35848 762855
rect 35808 761932 35860 761938
rect 35808 761874 35860 761880
rect 35164 759824 35216 759830
rect 35164 759766 35216 759772
rect 33784 758328 33836 758334
rect 33784 758270 33836 758276
rect 36556 757761 36584 767314
rect 39580 766148 39632 766154
rect 39580 766090 39632 766096
rect 39592 764561 39620 766090
rect 39578 764552 39634 764561
rect 39578 764487 39634 764496
rect 39776 764153 39804 768810
rect 40040 768732 40092 768738
rect 40040 768674 40092 768680
rect 40052 767009 40080 768674
rect 40038 767000 40094 767009
rect 40038 766935 40094 766944
rect 41708 765914 41736 768946
rect 41708 765886 42288 765914
rect 40132 764856 40184 764862
rect 40132 764798 40184 764804
rect 39762 764144 39818 764153
rect 39762 764079 39818 764088
rect 39948 761932 40000 761938
rect 39948 761874 40000 761880
rect 39960 758577 39988 761874
rect 40144 761841 40172 764798
rect 41696 764584 41748 764590
rect 42064 764584 42116 764590
rect 41748 764532 42064 764538
rect 41696 764526 42116 764532
rect 41708 764510 42104 764526
rect 40500 763360 40552 763366
rect 40498 763328 40500 763337
rect 42064 763360 42116 763366
rect 40552 763328 40554 763337
rect 40498 763263 40554 763272
rect 41708 763308 42064 763314
rect 41708 763302 42116 763308
rect 41708 763286 42104 763302
rect 41708 763230 41736 763286
rect 41696 763224 41748 763230
rect 41696 763166 41748 763172
rect 40130 761832 40186 761841
rect 40130 761767 40186 761776
rect 41696 759824 41748 759830
rect 41748 759772 42012 759778
rect 41696 759766 42012 759772
rect 41708 759750 42012 759766
rect 41604 759688 41656 759694
rect 41656 759636 41828 759642
rect 41604 759630 41828 759636
rect 41616 759614 41828 759630
rect 39946 758568 40002 758577
rect 39946 758503 40002 758512
rect 39856 758328 39908 758334
rect 39856 758270 39908 758276
rect 36542 757752 36598 757761
rect 36542 757687 36598 757696
rect 39868 757353 39896 758270
rect 39854 757344 39910 757353
rect 39854 757279 39910 757288
rect 41800 757081 41828 759614
rect 41984 757217 42012 759750
rect 41970 757208 42026 757217
rect 41970 757143 42026 757152
rect 41786 757072 41842 757081
rect 41786 757007 41842 757016
rect 41878 756664 41934 756673
rect 41878 756599 41934 756608
rect 41892 756226 41920 756599
rect 42260 754882 42288 765886
rect 42430 764144 42486 764153
rect 42430 764079 42486 764088
rect 42168 754854 42288 754882
rect 42168 754392 42196 754854
rect 42248 754316 42300 754322
rect 42248 754258 42300 754264
rect 42260 754202 42288 754258
rect 42076 754174 42288 754202
rect 42444 754186 42472 764079
rect 42720 761920 42748 771406
rect 43272 770681 43300 812806
rect 43456 807974 43484 815730
rect 44180 815652 44232 815658
rect 44180 815594 44232 815600
rect 43444 807968 43496 807974
rect 43444 807910 43496 807916
rect 43444 807356 43496 807362
rect 43444 807298 43496 807304
rect 43456 794782 43484 807298
rect 43812 806132 43864 806138
rect 43812 806074 43864 806080
rect 43628 799128 43680 799134
rect 43628 799070 43680 799076
rect 43640 797337 43668 799070
rect 43626 797328 43682 797337
rect 43626 797263 43682 797272
rect 43444 794776 43496 794782
rect 43444 794718 43496 794724
rect 43258 770672 43314 770681
rect 43258 770607 43314 770616
rect 43074 770264 43130 770273
rect 43074 770199 43130 770208
rect 42720 761892 42932 761920
rect 42614 761832 42670 761841
rect 42614 761767 42670 761776
rect 42432 754180 42484 754186
rect 42076 753780 42104 754174
rect 42432 754122 42484 754128
rect 42246 754080 42302 754089
rect 42246 754015 42302 754024
rect 42260 753494 42288 754015
rect 42628 753930 42656 761767
rect 42904 756922 42932 761892
rect 43088 756922 43116 770199
rect 43258 758568 43314 758577
rect 43258 758503 43314 758512
rect 42904 756894 43024 756922
rect 43088 756894 43208 756922
rect 42800 754180 42852 754186
rect 42800 754122 42852 754128
rect 42168 753466 42288 753494
rect 42352 753902 42656 753930
rect 42168 753409 42196 753466
rect 42154 753400 42210 753409
rect 42154 753335 42210 753344
rect 42062 752992 42118 753001
rect 42062 752927 42118 752936
rect 42076 752556 42104 752927
rect 42076 751641 42104 751944
rect 41878 751632 41934 751641
rect 41878 751567 41934 751576
rect 42062 751632 42118 751641
rect 42352 751618 42380 753902
rect 42614 753672 42670 753681
rect 42614 753607 42670 753616
rect 42628 753494 42656 753607
rect 42062 751567 42118 751576
rect 42260 751590 42380 751618
rect 42536 753466 42656 753494
rect 41892 751369 41920 751567
rect 42260 751534 42288 751590
rect 42248 751528 42300 751534
rect 42248 751470 42300 751476
rect 42248 751188 42300 751194
rect 42248 751130 42300 751136
rect 42260 750734 42288 751130
rect 42182 750706 42288 750734
rect 41970 750544 42026 750553
rect 41970 750479 42026 750488
rect 41984 750108 42012 750479
rect 41970 749728 42026 749737
rect 41970 749663 42026 749672
rect 41984 749529 42012 749663
rect 42246 749456 42302 749465
rect 42246 749391 42302 749400
rect 42260 747062 42288 749391
rect 42182 747034 42288 747062
rect 41786 746872 41842 746881
rect 41786 746807 41842 746816
rect 41800 746401 41828 746807
rect 42536 745770 42564 753466
rect 42182 745742 42564 745770
rect 42812 745657 42840 754122
rect 42996 752114 43024 756894
rect 42996 752086 43116 752114
rect 41970 745648 42026 745657
rect 41970 745583 42026 745592
rect 42798 745648 42854 745657
rect 42798 745583 42854 745592
rect 41984 745212 42012 745583
rect 42246 745376 42302 745385
rect 42246 745311 42302 745320
rect 41786 743744 41842 743753
rect 41786 743679 41842 743688
rect 41800 743376 41828 743679
rect 42260 743186 42288 745311
rect 42522 744424 42578 744433
rect 42168 743158 42288 743186
rect 42352 744382 42522 744410
rect 42168 742696 42196 743158
rect 42352 742098 42380 744382
rect 42522 744359 42578 744368
rect 42524 743912 42576 743918
rect 42524 743854 42576 743860
rect 42182 742070 42380 742098
rect 42536 741554 42564 743854
rect 43088 743834 43116 752086
rect 42182 741526 42564 741554
rect 42904 743806 43116 743834
rect 8588 731884 8616 732020
rect 9048 731884 9076 732020
rect 9508 731884 9536 732020
rect 9968 731884 9996 732020
rect 10428 731884 10456 732020
rect 10888 731884 10916 732020
rect 11348 731884 11376 732020
rect 11808 731884 11836 732020
rect 12268 731884 12296 732020
rect 12728 731884 12756 732020
rect 13188 731884 13216 732020
rect 13648 731884 13676 732020
rect 14108 731884 14136 732020
rect 41142 730960 41198 730969
rect 41142 730895 41198 730904
rect 41156 730250 41184 730895
rect 41696 730312 41748 730318
rect 42064 730312 42116 730318
rect 41748 730260 42064 730266
rect 41696 730254 42116 730260
rect 41144 730244 41196 730250
rect 41708 730238 42104 730254
rect 41144 730186 41196 730192
rect 41328 729088 41380 729094
rect 41328 729030 41380 729036
rect 41696 729088 41748 729094
rect 41696 729030 41748 729036
rect 41340 728691 41368 729030
rect 40774 728682 40830 728691
rect 40774 728617 40830 728626
rect 41326 728682 41382 728691
rect 41708 728668 41736 729030
rect 42064 728680 42116 728686
rect 41708 728640 42064 728668
rect 41326 728617 41382 728626
rect 42064 728622 42116 728628
rect 40788 727326 40816 728617
rect 41050 727458 41106 727467
rect 41050 727393 41106 727402
rect 41696 727456 41748 727462
rect 42064 727456 42116 727462
rect 41748 727416 42064 727444
rect 41696 727398 41748 727404
rect 42064 727398 42116 727404
rect 40776 727320 40828 727326
rect 40776 727262 40828 727268
rect 41696 727320 41748 727326
rect 42064 727320 42116 727326
rect 41748 727268 42064 727274
rect 41696 727262 42116 727268
rect 41708 727246 42104 727262
rect 41142 726880 41198 726889
rect 41142 726815 41198 726824
rect 40958 726234 41014 726243
rect 40958 726169 41014 726178
rect 35162 724840 35218 724849
rect 35162 724775 35218 724784
rect 33046 724432 33102 724441
rect 33046 724367 33102 724376
rect 33060 716825 33088 724367
rect 33782 723786 33838 723795
rect 33782 723721 33838 723730
rect 33046 716816 33102 716825
rect 33046 716751 33102 716760
rect 33796 715562 33824 723721
rect 35176 715698 35204 724775
rect 39302 723208 39358 723217
rect 39302 723143 39358 723152
rect 35164 715692 35216 715698
rect 35164 715634 35216 715640
rect 33784 715556 33836 715562
rect 33784 715498 33836 715504
rect 39316 714241 39344 723143
rect 40972 717641 41000 726169
rect 41156 725966 41184 726815
rect 41326 726234 41382 726243
rect 41326 726169 41382 726178
rect 41696 726232 41748 726238
rect 41748 726180 41828 726186
rect 41696 726174 41828 726180
rect 41708 726158 41828 726174
rect 41144 725960 41196 725966
rect 41144 725902 41196 725908
rect 41604 725960 41656 725966
rect 41800 725948 41828 726158
rect 42064 725960 42116 725966
rect 41800 725920 42064 725948
rect 41604 725902 41656 725908
rect 42064 725902 42116 725908
rect 42708 725960 42760 725966
rect 42708 725902 42760 725908
rect 41616 725778 41644 725902
rect 41786 725792 41842 725801
rect 41616 725750 41786 725778
rect 41786 725727 41842 725736
rect 41326 725656 41382 725665
rect 41326 725591 41382 725600
rect 41142 725248 41198 725257
rect 41142 725183 41198 725192
rect 40958 717632 41014 717641
rect 40958 717567 41014 717576
rect 40776 715556 40828 715562
rect 40776 715498 40828 715504
rect 40788 715329 40816 715498
rect 40774 715320 40830 715329
rect 40774 715255 40830 715264
rect 41156 714921 41184 725183
rect 41340 718865 41368 725591
rect 41786 722392 41842 722401
rect 41786 722327 41842 722336
rect 41326 718856 41382 718865
rect 41326 718791 41382 718800
rect 41800 718593 41828 722327
rect 42062 720352 42118 720361
rect 42062 720287 42118 720296
rect 42076 719030 42104 720287
rect 42064 719024 42116 719030
rect 42064 718966 42116 718972
rect 42062 718856 42118 718865
rect 42062 718791 42118 718800
rect 41786 718584 41842 718593
rect 41786 718519 41842 718528
rect 41512 715216 41564 715222
rect 41512 715158 41564 715164
rect 41142 714912 41198 714921
rect 41142 714847 41198 714856
rect 41524 714354 41552 715158
rect 42076 714649 42104 718791
rect 42720 717262 42748 725902
rect 42248 717256 42300 717262
rect 42248 717198 42300 717204
rect 42708 717256 42760 717262
rect 42708 717198 42760 717204
rect 42260 714728 42288 717198
rect 42430 715320 42486 715329
rect 42430 715255 42486 715264
rect 42444 715034 42472 715255
rect 42444 715006 42748 715034
rect 42522 714912 42578 714921
rect 42522 714854 42578 714856
rect 42522 714847 42656 714854
rect 42536 714826 42656 714847
rect 42260 714700 42564 714728
rect 42062 714640 42118 714649
rect 42062 714575 42118 714584
rect 41524 714326 42288 714354
rect 39302 714232 39358 714241
rect 39302 714167 39358 714176
rect 42260 713062 42288 714326
rect 42182 713034 42288 713062
rect 42536 711634 42564 714700
rect 42352 711606 42564 711634
rect 42352 711226 42380 711606
rect 42182 711198 42380 711226
rect 42154 710832 42210 710841
rect 42154 710767 42210 710776
rect 42168 710561 42196 710767
rect 41786 709880 41842 709889
rect 41786 709815 41842 709824
rect 41800 709376 41828 709815
rect 42076 708529 42104 708696
rect 41878 708520 41934 708529
rect 41878 708455 41934 708464
rect 42062 708520 42118 708529
rect 42062 708455 42118 708464
rect 41892 708152 41920 708455
rect 42062 707840 42118 707849
rect 42062 707775 42118 707784
rect 42076 707540 42104 707775
rect 41786 707432 41842 707441
rect 41786 707367 41842 707376
rect 41800 706860 41828 707367
rect 42628 706602 42656 714826
rect 42352 706574 42656 706602
rect 42352 706330 42380 706574
rect 42522 706480 42578 706489
rect 42522 706415 42578 706424
rect 42182 706302 42380 706330
rect 42248 705560 42300 705566
rect 42248 705502 42300 705508
rect 41786 704304 41842 704313
rect 41786 704239 41842 704248
rect 41800 703868 41828 704239
rect 42260 703746 42288 705502
rect 42536 705194 42564 706415
rect 42536 705166 42656 705194
rect 42076 703718 42288 703746
rect 42076 703188 42104 703718
rect 42246 703624 42302 703633
rect 42246 703559 42302 703568
rect 42062 703080 42118 703089
rect 42062 703015 42118 703024
rect 42076 702576 42104 703015
rect 41970 702264 42026 702273
rect 42260 702234 42288 703559
rect 42628 703202 42656 705166
rect 42536 703174 42656 703202
rect 42536 702273 42564 703174
rect 42720 703089 42748 715006
rect 42706 703080 42762 703089
rect 42706 703015 42762 703024
rect 42522 702264 42578 702273
rect 41970 702199 42026 702208
rect 42248 702228 42300 702234
rect 41984 702032 42012 702199
rect 42522 702199 42578 702208
rect 42248 702170 42300 702176
rect 42248 701956 42300 701962
rect 42248 701898 42300 701904
rect 42260 700179 42288 701898
rect 42522 701856 42578 701865
rect 42182 700151 42288 700179
rect 42352 701814 42522 701842
rect 42352 699530 42380 701814
rect 42522 701791 42578 701800
rect 42522 701584 42578 701593
rect 42522 701519 42578 701528
rect 42182 699502 42380 699530
rect 42536 699394 42564 701519
rect 42708 701140 42760 701146
rect 42708 701082 42760 701088
rect 42352 699366 42564 699394
rect 42352 698918 42380 699366
rect 42168 698850 42196 698904
rect 42260 698890 42380 698918
rect 42260 698850 42288 698890
rect 42168 698822 42288 698850
rect 42720 698339 42748 701082
rect 42182 698311 42748 698339
rect 8588 688772 8616 688908
rect 9048 688772 9076 688908
rect 9508 688772 9536 688908
rect 9968 688772 9996 688908
rect 10428 688772 10456 688908
rect 10888 688772 10916 688908
rect 11348 688772 11376 688908
rect 11808 688772 11836 688908
rect 12268 688772 12296 688908
rect 12728 688772 12756 688908
rect 13188 688772 13216 688908
rect 13648 688772 13676 688908
rect 14108 688772 14136 688908
rect 42706 688120 42762 688129
rect 42706 688055 42762 688064
rect 42720 687342 42748 688055
rect 42708 687336 42760 687342
rect 42708 687278 42760 687284
rect 40866 686896 40922 686905
rect 40866 686831 40922 686840
rect 40880 685914 40908 686831
rect 41142 686488 41198 686497
rect 41142 686423 41198 686432
rect 41156 686050 41184 686423
rect 41144 686044 41196 686050
rect 41144 685986 41196 685992
rect 41696 686044 41748 686050
rect 42064 686044 42116 686050
rect 41748 686004 42064 686032
rect 41696 685986 41748 685992
rect 42064 685986 42116 685992
rect 40868 685908 40920 685914
rect 40868 685850 40920 685856
rect 41050 685910 41106 685919
rect 41050 685845 41106 685854
rect 41696 685908 41748 685914
rect 42064 685908 42116 685914
rect 41748 685868 42064 685896
rect 41696 685850 41748 685856
rect 42064 685850 42116 685856
rect 41064 682990 41092 685845
rect 41326 683462 41382 683471
rect 41326 683397 41382 683406
rect 41696 683460 41748 683466
rect 41748 683420 41920 683448
rect 41696 683402 41748 683408
rect 41052 682984 41104 682990
rect 41052 682926 41104 682932
rect 41696 682984 41748 682990
rect 41696 682926 41748 682932
rect 35162 682000 35218 682009
rect 35162 681935 35218 681944
rect 31666 681592 31722 681601
rect 31666 681527 31722 681536
rect 31680 674150 31708 681527
rect 32402 681014 32458 681023
rect 32402 680949 32458 680958
rect 33782 681014 33838 681023
rect 33782 680949 33838 680958
rect 31668 674144 31720 674150
rect 31668 674086 31720 674092
rect 32416 672761 32444 680949
rect 32402 672752 32458 672761
rect 32402 672687 32458 672696
rect 33796 671362 33824 680949
rect 35176 672790 35204 681935
rect 41708 681057 41736 682926
rect 41694 681048 41750 681057
rect 41694 680983 41750 680992
rect 41892 678974 41920 683420
rect 42706 682408 42762 682417
rect 42706 682343 42762 682352
rect 41892 678946 42380 678974
rect 41142 677104 41198 677113
rect 41142 677039 41198 677048
rect 41156 676258 41184 677039
rect 41144 676252 41196 676258
rect 41144 676194 41196 676200
rect 41696 676252 41748 676258
rect 42064 676252 42116 676258
rect 41748 676212 42064 676240
rect 41696 676194 41748 676200
rect 42064 676194 42116 676200
rect 41512 674144 41564 674150
rect 41512 674086 41564 674092
rect 35164 672784 35216 672790
rect 35164 672726 35216 672732
rect 33784 671356 33836 671362
rect 33784 671298 33836 671304
rect 41524 671106 41552 674086
rect 41696 672784 41748 672790
rect 41748 672732 42104 672738
rect 41696 672726 42104 672732
rect 41708 672722 42104 672726
rect 41708 672716 42116 672722
rect 41708 672710 42064 672716
rect 42064 672658 42116 672664
rect 42352 671673 42380 678946
rect 42524 672716 42576 672722
rect 42524 672658 42576 672664
rect 42536 672602 42564 672658
rect 42536 672574 42656 672602
rect 42338 671664 42394 671673
rect 42338 671599 42394 671608
rect 41696 671356 41748 671362
rect 41748 671316 42564 671344
rect 41696 671298 41748 671304
rect 41524 671078 42288 671106
rect 42168 669746 42196 669868
rect 42260 669746 42288 671078
rect 42168 669718 42288 669746
rect 42340 669384 42392 669390
rect 42340 669326 42392 669332
rect 42062 668536 42118 668545
rect 42062 668471 42118 668480
rect 42076 668032 42104 668471
rect 42352 667366 42380 669326
rect 42182 667338 42380 667366
rect 42248 667276 42300 667282
rect 42248 667218 42300 667224
rect 42062 666632 42118 666641
rect 42062 666567 42118 666576
rect 42076 666165 42104 666567
rect 42260 665530 42288 667218
rect 42182 665502 42288 665530
rect 42340 665440 42392 665446
rect 42340 665382 42392 665388
rect 41786 665136 41842 665145
rect 41786 665071 41842 665080
rect 41800 664972 41828 665071
rect 42352 664339 42380 665382
rect 42182 664311 42380 664339
rect 41786 664048 41842 664057
rect 41786 663983 41842 663992
rect 41800 663680 41828 663983
rect 42536 663898 42564 671316
rect 42444 663882 42564 663898
rect 42432 663876 42564 663882
rect 42484 663870 42564 663876
rect 42432 663818 42484 663824
rect 42628 663218 42656 672574
rect 42352 663190 42656 663218
rect 42352 663150 42380 663190
rect 42182 663122 42380 663150
rect 42432 663060 42484 663066
rect 42432 663002 42484 663008
rect 42246 662824 42302 662833
rect 42246 662759 42302 662768
rect 42260 661042 42288 662759
rect 42168 661014 42288 661042
rect 42168 660620 42196 661014
rect 42156 660544 42208 660550
rect 42156 660486 42208 660492
rect 42168 660008 42196 660486
rect 42444 659371 42472 663002
rect 42182 659343 42472 659371
rect 42168 658838 42380 658866
rect 42168 658784 42196 658838
rect 42352 658798 42380 658838
rect 42720 658798 42748 682343
rect 42352 658770 42748 658798
rect 42522 658608 42578 658617
rect 42352 658566 42522 658594
rect 41800 658430 42288 658458
rect 41800 658345 41828 658430
rect 41786 658336 41842 658345
rect 41786 658271 41842 658280
rect 41786 657248 41842 657257
rect 41786 657183 41842 657192
rect 41800 656948 41828 657183
rect 42260 656350 42288 658430
rect 42182 656322 42288 656350
rect 42168 655710 42288 655738
rect 42168 655656 42196 655710
rect 42260 655670 42288 655710
rect 42352 655670 42380 658566
rect 42522 658543 42578 658552
rect 42524 657416 42576 657422
rect 42524 657358 42576 657364
rect 42260 655642 42380 655670
rect 42536 655126 42564 657358
rect 42182 655098 42564 655126
rect 8588 645524 8616 645660
rect 9048 645524 9076 645660
rect 9508 645524 9536 645660
rect 9968 645524 9996 645660
rect 10428 645524 10456 645660
rect 10888 645524 10916 645660
rect 11348 645524 11376 645660
rect 11808 645524 11836 645660
rect 12268 645524 12296 645660
rect 12728 645524 12756 645660
rect 13188 645524 13216 645660
rect 13648 645524 13676 645660
rect 14108 645524 14136 645660
rect 35806 644736 35862 644745
rect 35806 644671 35862 644680
rect 39486 644736 39542 644745
rect 39486 644671 39542 644680
rect 35820 644502 35848 644671
rect 35808 644496 35860 644502
rect 35808 644438 35860 644444
rect 38566 644328 38622 644337
rect 38566 644263 38622 644272
rect 35346 643920 35402 643929
rect 35346 643855 35402 643864
rect 35360 643142 35388 643855
rect 35808 643544 35860 643550
rect 35530 643512 35586 643521
rect 35530 643447 35586 643456
rect 35806 643512 35808 643521
rect 35860 643512 35862 643521
rect 35806 643447 35862 643456
rect 35544 643278 35572 643447
rect 35532 643272 35584 643278
rect 35532 643214 35584 643220
rect 35348 643136 35400 643142
rect 35348 643078 35400 643084
rect 35622 642696 35678 642705
rect 35622 642631 35678 642640
rect 35636 642054 35664 642631
rect 38580 642530 38608 644263
rect 38568 642524 38620 642530
rect 38568 642466 38620 642472
rect 35806 642288 35862 642297
rect 35806 642223 35862 642232
rect 35624 642048 35676 642054
rect 35624 641990 35676 641996
rect 35820 641782 35848 642223
rect 39500 642054 39528 644671
rect 41696 644496 41748 644502
rect 42064 644496 42116 644502
rect 41748 644446 42064 644474
rect 41696 644438 41748 644444
rect 42064 644438 42116 644444
rect 40500 643544 40552 643550
rect 40498 643512 40500 643521
rect 40552 643512 40554 643521
rect 40498 643447 40554 643456
rect 41708 643346 42104 643362
rect 41696 643340 42116 643346
rect 41748 643334 42064 643340
rect 41696 643282 41748 643288
rect 42064 643282 42116 643288
rect 41696 643136 41748 643142
rect 42064 643136 42116 643142
rect 41748 643084 42064 643090
rect 41696 643078 42116 643084
rect 41708 643062 42104 643078
rect 41696 642524 41748 642530
rect 41748 642484 42104 642512
rect 41696 642466 41748 642472
rect 42076 642394 42104 642484
rect 42064 642388 42116 642394
rect 42064 642330 42116 642336
rect 39488 642048 39540 642054
rect 39488 641990 39540 641996
rect 35808 641776 35860 641782
rect 35808 641718 35860 641724
rect 41696 641776 41748 641782
rect 42064 641776 42116 641782
rect 41748 641724 42064 641730
rect 41696 641718 42116 641724
rect 41708 641702 42104 641718
rect 35622 641472 35678 641481
rect 35622 641407 35678 641416
rect 35636 640354 35664 641407
rect 35806 641064 35862 641073
rect 35806 640999 35862 641008
rect 39578 641064 39634 641073
rect 39578 640999 39634 641008
rect 35820 640830 35848 640999
rect 35808 640824 35860 640830
rect 35808 640766 35860 640772
rect 39592 640762 39620 640999
rect 39580 640756 39632 640762
rect 39580 640698 39632 640704
rect 35806 640656 35862 640665
rect 35806 640591 35862 640600
rect 35820 640490 35848 640591
rect 35808 640484 35860 640490
rect 35808 640426 35860 640432
rect 39948 640484 40000 640490
rect 39948 640426 40000 640432
rect 35624 640348 35676 640354
rect 35624 640290 35676 640296
rect 39960 640257 39988 640426
rect 41696 640348 41748 640354
rect 42064 640348 42116 640354
rect 41748 640306 42064 640334
rect 41696 640290 41748 640296
rect 42064 640290 42116 640296
rect 39946 640248 40002 640257
rect 39946 640183 40002 640192
rect 35346 639840 35402 639849
rect 35346 639775 35402 639784
rect 35360 638246 35388 639775
rect 35530 639432 35586 639441
rect 35530 639367 35586 639376
rect 35806 639432 35862 639441
rect 35806 639367 35862 639376
rect 35544 638994 35572 639367
rect 35820 639130 35848 639367
rect 35808 639124 35860 639130
rect 35808 639066 35860 639072
rect 41696 639124 41748 639130
rect 41696 639066 41748 639072
rect 41708 639010 41736 639066
rect 35532 638988 35584 638994
rect 35532 638930 35584 638936
rect 37924 638988 37976 638994
rect 41708 638982 41920 639010
rect 37924 638930 37976 638936
rect 35622 638616 35678 638625
rect 35622 638551 35678 638560
rect 35348 638240 35400 638246
rect 35348 638182 35400 638188
rect 32402 637800 32458 637809
rect 32402 637735 32458 637744
rect 32416 629921 32444 637735
rect 35162 637392 35218 637401
rect 35162 637327 35218 637336
rect 32402 629912 32458 629921
rect 32402 629847 32458 629856
rect 35176 628726 35204 637327
rect 35636 637226 35664 638551
rect 35806 638208 35862 638217
rect 35806 638143 35862 638152
rect 35820 637634 35848 638143
rect 35808 637628 35860 637634
rect 35808 637570 35860 637576
rect 36544 637628 36596 637634
rect 36544 637570 36596 637576
rect 35624 637220 35676 637226
rect 35624 637162 35676 637168
rect 35622 636984 35678 636993
rect 35622 636919 35678 636928
rect 35636 636546 35664 636919
rect 35806 636576 35862 636585
rect 35624 636540 35676 636546
rect 35806 636511 35862 636520
rect 35624 636482 35676 636488
rect 35820 636274 35848 636511
rect 35808 636268 35860 636274
rect 35808 636210 35860 636216
rect 35806 635760 35862 635769
rect 35806 635695 35862 635704
rect 35820 634982 35848 635695
rect 35808 634976 35860 634982
rect 35808 634918 35860 634924
rect 35806 634536 35862 634545
rect 35806 634471 35862 634480
rect 35820 633894 35848 634471
rect 35808 633888 35860 633894
rect 35808 633830 35860 633836
rect 35622 633720 35678 633729
rect 35622 633655 35678 633664
rect 35636 633486 35664 633655
rect 35808 633616 35860 633622
rect 35808 633558 35860 633564
rect 35624 633480 35676 633486
rect 35624 633422 35676 633428
rect 35820 633321 35848 633558
rect 35806 633312 35862 633321
rect 35806 633247 35862 633256
rect 36556 630630 36584 637570
rect 36544 630624 36596 630630
rect 36544 630566 36596 630572
rect 37936 629241 37964 638930
rect 41696 638240 41748 638246
rect 41696 638182 41748 638188
rect 40408 636948 40460 636954
rect 40408 636890 40460 636896
rect 39856 636540 39908 636546
rect 39856 636482 39908 636488
rect 39028 636200 39080 636206
rect 39026 636168 39028 636177
rect 39080 636168 39082 636177
rect 39026 636103 39082 636112
rect 39868 635769 39896 636482
rect 39854 635760 39910 635769
rect 39854 635695 39910 635704
rect 39488 634976 39540 634982
rect 39488 634918 39540 634924
rect 39500 634545 39528 634918
rect 39486 634536 39542 634545
rect 39486 634471 39542 634480
rect 40132 633888 40184 633894
rect 40132 633830 40184 633836
rect 40144 633729 40172 633830
rect 40130 633720 40186 633729
rect 39764 633684 39816 633690
rect 40130 633655 40186 633664
rect 39764 633626 39816 633632
rect 39776 632913 39804 633626
rect 39762 632904 39818 632913
rect 39762 632839 39818 632848
rect 40420 632641 40448 636890
rect 41708 635066 41736 638182
rect 41708 635038 41828 635066
rect 41604 633480 41656 633486
rect 41604 633422 41656 633428
rect 41616 633321 41644 633422
rect 41602 633312 41658 633321
rect 41602 633247 41658 633256
rect 40406 632632 40462 632641
rect 40406 632567 40462 632576
rect 41800 630674 41828 635038
rect 41892 634930 41920 638982
rect 41892 634902 42380 634930
rect 42064 633480 42116 633486
rect 42064 633422 42116 633428
rect 42076 633321 42104 633422
rect 42062 633312 42118 633321
rect 42062 633247 42118 633256
rect 42352 630674 42380 634902
rect 42706 632632 42762 632641
rect 42706 632567 42762 632576
rect 41800 630646 42196 630674
rect 42352 630646 42564 630674
rect 41604 630624 41656 630630
rect 41656 630572 41828 630578
rect 41604 630566 41828 630572
rect 41616 630550 41828 630566
rect 37922 629232 37978 629241
rect 37922 629167 37978 629176
rect 35164 628720 35216 628726
rect 40500 628720 40552 628726
rect 35164 628662 35216 628668
rect 40498 628688 40500 628697
rect 40552 628688 40554 628697
rect 40498 628623 40554 628632
rect 41800 627473 41828 630550
rect 42168 628538 42196 630646
rect 42338 628688 42394 628697
rect 42338 628623 42394 628632
rect 42168 628510 42288 628538
rect 41786 627464 41842 627473
rect 41786 627399 41842 627408
rect 41786 627192 41842 627201
rect 41786 627127 41842 627136
rect 41800 626620 41828 627127
rect 42260 625274 42288 628510
rect 42352 627914 42380 628623
rect 42352 627886 42472 627914
rect 42076 625246 42288 625274
rect 42076 624784 42104 625246
rect 42062 624472 42118 624481
rect 42062 624407 42118 624416
rect 42076 624172 42104 624407
rect 41786 623384 41842 623393
rect 41786 623319 41842 623328
rect 41800 622948 41828 623319
rect 42168 622033 42196 622336
rect 41786 622024 41842 622033
rect 41786 621959 41842 621968
rect 42154 622024 42210 622033
rect 42154 621959 42210 621968
rect 41800 621792 41828 621959
rect 42248 621716 42300 621722
rect 42248 621658 42300 621664
rect 42260 621126 42288 621658
rect 42182 621098 42288 621126
rect 41786 620800 41842 620809
rect 41786 620735 41842 620744
rect 41800 620500 41828 620735
rect 42248 620424 42300 620430
rect 42248 620366 42300 620372
rect 42260 620242 42288 620366
rect 42076 620214 42288 620242
rect 42076 619956 42104 620214
rect 42248 619676 42300 619682
rect 42248 619618 42300 619624
rect 42260 619018 42288 619618
rect 42260 618990 42380 619018
rect 42352 617454 42380 618990
rect 42182 617426 42380 617454
rect 42248 617364 42300 617370
rect 42248 617306 42300 617312
rect 42260 617250 42288 617306
rect 42076 617222 42288 617250
rect 42076 616828 42104 617222
rect 42444 616298 42472 627886
rect 42536 620242 42564 630646
rect 42720 620430 42748 632567
rect 42708 620424 42760 620430
rect 42708 620366 42760 620372
rect 42536 620214 42748 620242
rect 42168 616270 42472 616298
rect 42168 616148 42196 616270
rect 41878 616040 41934 616049
rect 41934 615998 42288 616026
rect 41878 615975 41934 615984
rect 42062 615904 42118 615913
rect 42062 615839 42118 615848
rect 42076 615604 42104 615839
rect 42260 614122 42288 615998
rect 42720 615913 42748 620214
rect 42706 615904 42762 615913
rect 42706 615839 42762 615848
rect 42614 615496 42670 615505
rect 42614 615431 42670 615440
rect 42628 615346 42656 615431
rect 42168 614094 42288 614122
rect 42536 615318 42656 615346
rect 42168 613768 42196 614094
rect 41878 613456 41934 613465
rect 41878 613391 41934 613400
rect 41892 613121 41920 613391
rect 42536 612490 42564 615318
rect 42708 614168 42760 614174
rect 42708 614110 42760 614116
rect 42182 612462 42564 612490
rect 42720 612082 42748 614110
rect 42904 612814 42932 743806
rect 43180 736934 43208 756894
rect 43088 736906 43208 736934
rect 43088 729337 43116 736906
rect 43074 729328 43130 729337
rect 43074 729263 43130 729272
rect 43076 728680 43128 728686
rect 43076 728622 43128 728628
rect 43088 686089 43116 728622
rect 43074 686080 43130 686089
rect 43074 686015 43130 686024
rect 43074 680368 43130 680377
rect 43074 680303 43130 680312
rect 43088 660550 43116 680303
rect 43076 660544 43128 660550
rect 43076 660486 43128 660492
rect 43074 635760 43130 635769
rect 43074 635695 43130 635704
rect 43088 617370 43116 635695
rect 43076 617364 43128 617370
rect 43076 617306 43128 617312
rect 43076 616548 43128 616554
rect 43076 616490 43128 616496
rect 42892 612808 42944 612814
rect 42892 612750 42944 612756
rect 43088 612542 43116 616490
rect 43076 612536 43128 612542
rect 43076 612478 43128 612484
rect 43272 612241 43300 758503
rect 43442 731368 43498 731377
rect 43442 731303 43498 731312
rect 43456 730182 43484 731303
rect 43626 730552 43682 730561
rect 43626 730487 43682 730496
rect 43444 730176 43496 730182
rect 43444 730118 43496 730124
rect 43640 729366 43668 730487
rect 43628 729360 43680 729366
rect 43628 729302 43680 729308
rect 43442 723616 43498 723625
rect 43442 723551 43498 723560
rect 43456 705566 43484 723551
rect 43628 712156 43680 712162
rect 43628 712098 43680 712104
rect 43640 710841 43668 712098
rect 43626 710832 43682 710841
rect 43626 710767 43682 710776
rect 43628 709368 43680 709374
rect 43628 709310 43680 709316
rect 43640 707849 43668 709310
rect 43626 707840 43682 707849
rect 43626 707775 43682 707784
rect 43444 705560 43496 705566
rect 43444 705502 43496 705508
rect 43442 687304 43498 687313
rect 43442 687239 43498 687248
rect 43456 686526 43484 687239
rect 43444 686520 43496 686526
rect 43444 686462 43496 686468
rect 43626 679552 43682 679561
rect 43626 679487 43682 679496
rect 43442 676696 43498 676705
rect 43442 676631 43498 676640
rect 43456 630674 43484 676631
rect 43640 665446 43668 679487
rect 43628 665440 43680 665446
rect 43628 665382 43680 665388
rect 43626 633720 43682 633729
rect 43626 633655 43682 633664
rect 43456 630646 43576 630674
rect 43548 614718 43576 630646
rect 43640 616298 43668 633655
rect 43824 616554 43852 806074
rect 44192 773226 44220 815594
rect 44364 814428 44416 814434
rect 44364 814370 44416 814376
rect 44180 773220 44232 773226
rect 44180 773162 44232 773168
rect 44376 771458 44404 814370
rect 44548 814292 44600 814298
rect 44548 814234 44600 814240
rect 44560 771662 44588 814234
rect 44836 785194 44864 817090
rect 61384 817012 61436 817018
rect 61384 816954 61436 816960
rect 53104 799128 53156 799134
rect 53104 799070 53156 799076
rect 45008 797700 45060 797706
rect 45008 797642 45060 797648
rect 45020 795433 45048 797642
rect 45006 795424 45062 795433
rect 45006 795359 45062 795368
rect 53116 790770 53144 799070
rect 57244 797700 57296 797706
rect 57244 797642 57296 797648
rect 53104 790764 53156 790770
rect 53104 790706 53156 790712
rect 57256 789206 57284 797642
rect 57244 789200 57296 789206
rect 57244 789142 57296 789148
rect 61396 786185 61424 816954
rect 62764 807968 62816 807974
rect 62764 807910 62816 807916
rect 62212 790764 62264 790770
rect 62212 790706 62264 790712
rect 62224 790537 62252 790706
rect 62210 790528 62266 790537
rect 62210 790463 62266 790472
rect 62120 789200 62172 789206
rect 62118 789168 62120 789177
rect 62172 789168 62174 789177
rect 62118 789103 62174 789112
rect 62118 787400 62174 787409
rect 62118 787335 62174 787344
rect 62132 786690 62160 787335
rect 62776 787137 62804 807910
rect 64144 805996 64196 806002
rect 64144 805938 64196 805944
rect 62762 787128 62818 787137
rect 62762 787063 62818 787072
rect 62120 786684 62172 786690
rect 62120 786626 62172 786632
rect 61382 786176 61438 786185
rect 61382 786111 61438 786120
rect 44824 785188 44876 785194
rect 44824 785130 44876 785136
rect 62120 785188 62172 785194
rect 62120 785130 62172 785136
rect 62132 784961 62160 785130
rect 62118 784952 62174 784961
rect 62118 784887 62174 784896
rect 60004 774240 60056 774246
rect 60004 774182 60056 774188
rect 44914 773120 44970 773129
rect 44914 773055 44970 773064
rect 46204 773084 46256 773090
rect 44548 771656 44600 771662
rect 44548 771598 44600 771604
rect 44364 771452 44416 771458
rect 44364 771394 44416 771400
rect 44546 769448 44602 769457
rect 44546 769383 44602 769392
rect 44180 764584 44232 764590
rect 44180 764526 44232 764532
rect 44362 764552 44418 764561
rect 44192 751913 44220 764526
rect 44362 764487 44418 764496
rect 44376 753001 44404 764487
rect 44362 752992 44418 753001
rect 44362 752927 44418 752936
rect 44178 751904 44234 751913
rect 44178 751839 44234 751848
rect 44270 728104 44326 728113
rect 44270 728039 44326 728048
rect 44284 685273 44312 728039
rect 44560 727705 44588 769383
rect 44732 755540 44784 755546
rect 44732 755482 44784 755488
rect 44744 754322 44772 755482
rect 44732 754316 44784 754322
rect 44732 754258 44784 754264
rect 44928 730153 44956 773055
rect 46204 773026 46256 773032
rect 45376 770092 45428 770098
rect 45376 770034 45428 770040
rect 45098 751632 45154 751641
rect 45098 751567 45154 751576
rect 45112 746570 45140 751567
rect 45100 746564 45152 746570
rect 45100 746506 45152 746512
rect 44914 730144 44970 730153
rect 44914 730079 44970 730088
rect 45190 729736 45246 729745
rect 45190 729671 45246 729680
rect 44546 727696 44602 727705
rect 44546 727631 44602 727640
rect 45008 727456 45060 727462
rect 45008 727398 45060 727404
rect 44454 722800 44510 722809
rect 44454 722735 44510 722744
rect 44468 709374 44496 722735
rect 44638 721576 44694 721585
rect 44638 721511 44694 721520
rect 44456 709368 44508 709374
rect 44456 709310 44508 709316
rect 44652 708801 44680 721511
rect 44638 708792 44694 708801
rect 44638 708727 44694 708736
rect 44454 708520 44510 708529
rect 44454 708455 44510 708464
rect 44468 703798 44496 708455
rect 44456 703792 44508 703798
rect 44456 703734 44508 703740
rect 44822 687712 44878 687721
rect 44822 687647 44878 687656
rect 44270 685264 44326 685273
rect 44270 685199 44326 685208
rect 44638 684856 44694 684865
rect 44638 684791 44694 684800
rect 44454 684040 44510 684049
rect 44454 683975 44510 683984
rect 44270 681048 44326 681057
rect 44270 680983 44326 680992
rect 43994 677920 44050 677929
rect 43994 677855 44050 677864
rect 44008 649994 44036 677855
rect 44008 649966 44128 649994
rect 44100 618254 44128 649966
rect 44284 644745 44312 680983
rect 44270 644736 44326 644745
rect 44270 644671 44326 644680
rect 44468 641073 44496 683975
rect 44652 641782 44680 684791
rect 44836 655518 44864 687647
rect 45020 684457 45048 727398
rect 45204 685914 45232 729671
rect 45388 727326 45416 770034
rect 45558 763328 45614 763337
rect 45558 763263 45614 763272
rect 45376 727320 45428 727326
rect 45376 727262 45428 727268
rect 45376 686044 45428 686050
rect 45376 685986 45428 685992
rect 45192 685908 45244 685914
rect 45192 685850 45244 685856
rect 45006 684448 45062 684457
rect 45006 684383 45062 684392
rect 45006 679960 45062 679969
rect 45006 679895 45062 679904
rect 45020 666641 45048 679895
rect 45006 666632 45062 666641
rect 45006 666567 45062 666576
rect 44824 655512 44876 655518
rect 44824 655454 44876 655460
rect 45006 643512 45062 643521
rect 45006 643447 45062 643456
rect 44640 641776 44692 641782
rect 44640 641718 44692 641724
rect 44454 641064 44510 641073
rect 44454 640999 44510 641008
rect 44638 636168 44694 636177
rect 44638 636103 44694 636112
rect 44270 634536 44326 634545
rect 44270 634471 44326 634480
rect 44284 619682 44312 634471
rect 44456 625864 44508 625870
rect 44456 625806 44508 625812
rect 44468 624481 44496 625806
rect 44454 624472 44510 624481
rect 44454 624407 44510 624416
rect 44652 622146 44680 636103
rect 44822 632904 44878 632913
rect 44822 632839 44878 632848
rect 44836 627914 44864 632839
rect 44836 627886 44956 627914
rect 44560 622118 44680 622146
rect 44560 621722 44588 622118
rect 44730 622024 44786 622033
rect 44730 621959 44786 621968
rect 44548 621716 44600 621722
rect 44548 621658 44600 621664
rect 44272 619676 44324 619682
rect 44272 619618 44324 619624
rect 44100 618226 44220 618254
rect 43812 616548 43864 616554
rect 43812 616490 43864 616496
rect 43640 616270 43852 616298
rect 43536 614712 43588 614718
rect 43536 614654 43588 614660
rect 43824 613135 43852 616270
rect 43824 613107 43944 613135
rect 43916 612270 43944 613107
rect 43904 612264 43956 612270
rect 43258 612232 43314 612241
rect 43258 612167 43314 612176
rect 43764 612232 43820 612241
rect 43904 612206 43956 612212
rect 43764 612167 43766 612176
rect 43818 612167 43820 612176
rect 43766 612138 43818 612144
rect 42536 612054 42748 612082
rect 43873 612096 43929 612105
rect 42536 611946 42564 612054
rect 43873 612031 43929 612040
rect 42182 611918 42564 611946
rect 43887 611930 43915 612031
rect 43875 611924 43927 611930
rect 43875 611866 43927 611872
rect 44192 611266 44220 618226
rect 44744 616826 44772 621959
rect 44732 616820 44784 616826
rect 44732 616762 44784 616768
rect 44364 614712 44416 614718
rect 44364 614654 44416 614660
rect 44376 611658 44404 614654
rect 44548 612264 44600 612270
rect 44548 612206 44600 612212
rect 44364 611652 44416 611658
rect 44364 611594 44416 611600
rect 44192 611238 44358 611266
rect 44330 611182 44358 611238
rect 44318 611176 44370 611182
rect 44318 611118 44370 611124
rect 44560 611114 44588 612206
rect 44928 611354 44956 627886
rect 44836 611326 44956 611354
rect 44836 611250 44864 611326
rect 44824 611244 44876 611250
rect 44824 611186 44876 611192
rect 44548 611108 44600 611114
rect 44548 611050 44600 611056
rect 8588 602276 8616 602412
rect 9048 602276 9076 602412
rect 9508 602276 9536 602412
rect 9968 602276 9996 602412
rect 10428 602276 10456 602412
rect 10888 602276 10916 602412
rect 11348 602276 11376 602412
rect 11808 602276 11836 602412
rect 12268 602276 12296 602412
rect 12728 602276 12756 602412
rect 13188 602276 13216 602412
rect 13648 602276 13676 602412
rect 14108 602276 14136 602412
rect 33782 601760 33838 601769
rect 33782 601695 33838 601704
rect 32402 595232 32458 595241
rect 32402 595167 32458 595176
rect 31022 594416 31078 594425
rect 31022 594351 31078 594360
rect 31036 585818 31064 594351
rect 32416 585954 32444 595167
rect 33796 589393 33824 601695
rect 38566 601352 38622 601361
rect 38566 601287 38622 601296
rect 35438 595810 35494 595819
rect 35438 595745 35494 595754
rect 33782 589384 33838 589393
rect 33782 589319 33838 589328
rect 35452 587178 35480 595745
rect 38580 594182 38608 601287
rect 39946 600944 40002 600953
rect 39946 600879 40002 600888
rect 39960 595814 39988 600879
rect 45020 600545 45048 643447
rect 45388 643346 45416 685986
rect 45376 643340 45428 643346
rect 45376 643282 45428 643288
rect 45376 640348 45428 640354
rect 45376 640290 45428 640296
rect 45190 640248 45246 640257
rect 45190 640183 45246 640192
rect 45006 600536 45062 600545
rect 45006 600471 45062 600480
rect 44638 600128 44694 600137
rect 44638 600063 44694 600072
rect 42890 597680 42946 597689
rect 42890 597615 42946 597624
rect 42904 597446 42932 597615
rect 42892 597440 42944 597446
rect 42892 597382 42944 597388
rect 42892 597032 42944 597038
rect 42892 596974 42944 596980
rect 43074 597000 43130 597009
rect 42154 596864 42210 596873
rect 42154 596799 42210 596808
rect 39948 595808 40000 595814
rect 41696 595808 41748 595814
rect 39948 595750 40000 595756
rect 41694 595776 41696 595785
rect 41748 595776 41750 595785
rect 41694 595711 41750 595720
rect 39302 594824 39358 594833
rect 39302 594759 39358 594768
rect 38568 594176 38620 594182
rect 38568 594118 38620 594124
rect 36542 593600 36598 593609
rect 36542 593535 36598 593544
rect 35440 587172 35492 587178
rect 35440 587114 35492 587120
rect 36556 586158 36584 593535
rect 36544 586152 36596 586158
rect 36544 586094 36596 586100
rect 32404 585948 32456 585954
rect 32404 585890 32456 585896
rect 31024 585812 31076 585818
rect 31024 585754 31076 585760
rect 39316 585177 39344 594759
rect 41696 594176 41748 594182
rect 41694 594144 41696 594153
rect 41748 594144 41750 594153
rect 41694 594079 41750 594088
rect 41970 592784 42026 592793
rect 41970 592719 42026 592728
rect 41786 592376 41842 592385
rect 41524 592334 41786 592362
rect 41524 589121 41552 592334
rect 41786 592311 41842 592320
rect 41786 590336 41842 590345
rect 41786 590271 41842 590280
rect 41800 589274 41828 590271
rect 41984 589665 42012 592719
rect 41970 589656 42026 589665
rect 41970 589591 42026 589600
rect 41708 589246 41828 589274
rect 41708 589121 41736 589246
rect 41510 589112 41566 589121
rect 41510 589047 41566 589056
rect 41694 589112 41750 589121
rect 41694 589047 41750 589056
rect 41512 587172 41564 587178
rect 41512 587114 41564 587120
rect 41524 586945 41552 587114
rect 41510 586936 41566 586945
rect 41510 586871 41566 586880
rect 39672 586152 39724 586158
rect 39670 586120 39672 586129
rect 39724 586120 39726 586129
rect 39670 586055 39726 586064
rect 41696 585948 41748 585954
rect 42168 585936 42196 596799
rect 42706 596048 42762 596057
rect 42706 595983 42762 595992
rect 42720 592034 42748 595983
rect 42536 592006 42748 592034
rect 42904 592034 42932 596974
rect 43074 596935 43130 596944
rect 42904 592006 43024 592034
rect 42536 589274 42564 592006
rect 42536 589246 42656 589274
rect 42628 586072 42656 589246
rect 42798 586936 42854 586945
rect 42798 586871 42854 586880
rect 42536 586044 42656 586072
rect 42536 585936 42564 586044
rect 42168 585908 42380 585936
rect 41696 585890 41748 585896
rect 41708 585834 41736 585890
rect 39764 585812 39816 585818
rect 41708 585806 42288 585834
rect 39764 585754 39816 585760
rect 39302 585168 39358 585177
rect 39302 585103 39358 585112
rect 39776 584633 39804 585754
rect 39762 584624 39818 584633
rect 39762 584559 39818 584568
rect 42260 583454 42288 585806
rect 42182 583426 42288 583454
rect 42352 583250 42380 585908
rect 42444 585908 42564 585936
rect 42444 584474 42472 585908
rect 42614 584624 42670 584633
rect 42614 584559 42670 584568
rect 42444 584446 42564 584474
rect 42260 583222 42380 583250
rect 42260 581618 42288 583222
rect 42182 581590 42288 581618
rect 42338 581224 42394 581233
rect 42338 581159 42394 581168
rect 42076 580689 42104 580961
rect 42062 580680 42118 580689
rect 42062 580615 42118 580624
rect 41786 580272 41842 580281
rect 41786 580207 41842 580216
rect 41800 579768 41828 580207
rect 42182 579107 42288 579135
rect 42260 578921 42288 579107
rect 42352 579034 42380 581159
rect 42352 579006 42472 579034
rect 42246 578912 42302 578921
rect 42246 578847 42302 578856
rect 42168 578598 42288 578626
rect 42168 578544 42196 578598
rect 42260 578558 42288 578598
rect 42444 578558 42472 579006
rect 42260 578530 42472 578558
rect 42246 578096 42302 578105
rect 42246 578031 42302 578040
rect 42260 577946 42288 578031
rect 42182 577918 42288 577946
rect 41786 577824 41842 577833
rect 41786 577759 41842 577768
rect 41800 577281 41828 577759
rect 42536 577674 42564 584446
rect 42444 577658 42564 577674
rect 42432 577652 42564 577658
rect 42484 577646 42564 577652
rect 42432 577594 42484 577600
rect 42628 577590 42656 584559
rect 42616 577584 42668 577590
rect 42616 577526 42668 577532
rect 42616 577448 42668 577454
rect 42812 577425 42840 586871
rect 42616 577390 42668 577396
rect 42798 577416 42854 577425
rect 42340 577312 42392 577318
rect 42340 577254 42392 577260
rect 41970 577144 42026 577153
rect 41970 577079 42026 577088
rect 41984 576708 42012 577079
rect 41786 574696 41842 574705
rect 42352 574682 42380 577254
rect 41786 574631 41842 574640
rect 42260 574654 42380 574682
rect 41800 574260 41828 574631
rect 41786 573880 41842 573889
rect 41786 573815 41842 573824
rect 41800 573580 41828 573815
rect 42260 572982 42288 574654
rect 42182 572954 42288 572982
rect 42628 572438 42656 577390
rect 42798 577351 42854 577360
rect 42996 572714 43024 592006
rect 42168 572370 42196 572424
rect 42260 572410 42656 572438
rect 42812 572686 43024 572714
rect 42260 572370 42288 572410
rect 42168 572342 42288 572370
rect 42246 572248 42302 572257
rect 42246 572183 42302 572192
rect 41786 570888 41842 570897
rect 41786 570823 41842 570832
rect 41800 570588 41828 570823
rect 42260 569922 42288 572183
rect 42614 571976 42670 571985
rect 42614 571911 42670 571920
rect 42430 571432 42486 571441
rect 42430 571367 42486 571376
rect 42182 569894 42288 569922
rect 42444 569430 42472 571367
rect 42432 569424 42484 569430
rect 42432 569366 42484 569372
rect 42628 569310 42656 571911
rect 42168 569242 42196 569296
rect 42260 569282 42656 569310
rect 42260 569242 42288 569282
rect 42168 569214 42288 569242
rect 42432 569220 42484 569226
rect 42432 569162 42484 569168
rect 42444 568766 42472 569162
rect 42168 568698 42196 568752
rect 42260 568738 42472 568766
rect 42260 568698 42288 568738
rect 42168 568670 42288 568698
rect 8588 559164 8616 559300
rect 9048 559164 9076 559300
rect 9508 559164 9536 559300
rect 9968 559164 9996 559300
rect 10428 559164 10456 559300
rect 10888 559164 10916 559300
rect 11348 559164 11376 559300
rect 11808 559164 11836 559300
rect 12268 559164 12296 559300
rect 12728 559164 12756 559300
rect 13188 559164 13216 559300
rect 13648 559164 13676 559300
rect 14108 559164 14136 559300
rect 41142 558104 41198 558113
rect 41142 558039 41198 558048
rect 40038 553408 40094 553417
rect 40038 553343 40040 553352
rect 40092 553343 40094 553352
rect 40040 553318 40092 553324
rect 37922 552392 37978 552401
rect 37922 552327 37978 552336
rect 29642 551984 29698 551993
rect 29642 551919 29698 551928
rect 29656 544406 29684 551919
rect 29644 544400 29696 544406
rect 29644 544342 29696 544348
rect 37936 542337 37964 552327
rect 41156 550594 41184 558039
rect 42812 554849 42840 572686
rect 43088 556481 43116 596935
rect 44362 593192 44418 593201
rect 44362 593127 44418 593136
rect 44178 591968 44234 591977
rect 44178 591903 44234 591912
rect 43350 591560 43406 591569
rect 43350 591495 43406 591504
rect 43364 582374 43392 591495
rect 43626 589112 43682 589121
rect 43626 589047 43682 589056
rect 43364 582346 43484 582374
rect 43074 556472 43130 556481
rect 43074 556407 43130 556416
rect 42798 554840 42854 554849
rect 42798 554775 42854 554784
rect 41696 553376 41748 553382
rect 41748 553324 42380 553330
rect 41696 553318 42380 553324
rect 41708 553302 42380 553318
rect 41326 552800 41382 552809
rect 41326 552735 41382 552744
rect 41340 552158 41368 552735
rect 41328 552152 41380 552158
rect 41328 552094 41380 552100
rect 41696 552152 41748 552158
rect 41696 552094 41748 552100
rect 41708 551857 41736 552094
rect 41694 551848 41750 551857
rect 41694 551783 41750 551792
rect 41708 550594 42196 550610
rect 41144 550588 41196 550594
rect 41144 550530 41196 550536
rect 41696 550588 42196 550594
rect 41748 550582 42196 550588
rect 41696 550530 41748 550536
rect 41970 550352 42026 550361
rect 41970 550287 42026 550296
rect 41786 549944 41842 549953
rect 41786 549879 41842 549888
rect 41800 545465 41828 549879
rect 41984 545737 42012 550287
rect 42168 550225 42196 550582
rect 42154 550216 42210 550225
rect 42154 550151 42210 550160
rect 41970 545728 42026 545737
rect 41970 545663 42026 545672
rect 41786 545456 41842 545465
rect 41786 545391 41842 545400
rect 41696 544400 41748 544406
rect 41696 544342 41748 544348
rect 41708 543734 41736 544342
rect 41708 543706 42288 543734
rect 37922 542328 37978 542337
rect 37922 542263 37978 542272
rect 42260 540274 42288 543706
rect 42182 540246 42288 540274
rect 42352 539730 42380 553302
rect 42798 551168 42854 551177
rect 42798 551103 42854 551112
rect 42260 539702 42380 539730
rect 42168 538370 42196 538424
rect 42260 538370 42288 539702
rect 42430 539608 42486 539617
rect 42430 539543 42486 539552
rect 42168 538342 42288 538370
rect 42168 537798 42288 537826
rect 42168 537744 42196 537798
rect 42260 537758 42288 537798
rect 42444 537758 42472 539543
rect 42260 537730 42472 537758
rect 42522 537568 42578 537577
rect 42522 537503 42578 537512
rect 42338 537296 42394 537305
rect 42338 537231 42394 537240
rect 41786 537024 41842 537033
rect 41786 536959 41842 536968
rect 41800 536588 41828 536959
rect 42076 535809 42104 535908
rect 42062 535800 42118 535809
rect 42062 535735 42118 535744
rect 42154 535528 42210 535537
rect 42154 535463 42210 535472
rect 42168 535364 42196 535463
rect 42352 534766 42380 537231
rect 42168 534698 42196 534752
rect 42260 534738 42380 534766
rect 42260 534698 42288 534738
rect 42168 534670 42288 534698
rect 42536 534086 42564 537503
rect 42182 534058 42564 534086
rect 42430 533896 42486 533905
rect 42430 533831 42486 533840
rect 41786 533760 41842 533769
rect 41786 533695 41842 533704
rect 41800 533528 41828 533695
rect 42248 533452 42300 533458
rect 42248 533394 42300 533400
rect 42260 531434 42288 533394
rect 42076 531406 42288 531434
rect 42076 531045 42104 531406
rect 42444 530754 42472 533831
rect 42614 532944 42670 532953
rect 42614 532879 42670 532888
rect 42628 532522 42656 532879
rect 42168 530726 42472 530754
rect 42536 532494 42656 532522
rect 42168 530400 42196 530726
rect 42062 530224 42118 530233
rect 42062 530159 42118 530168
rect 42076 529757 42104 530159
rect 42536 530074 42564 532494
rect 42812 531434 42840 551103
rect 42982 549536 43038 549545
rect 42982 549471 43038 549480
rect 42996 533458 43024 549471
rect 42984 533452 43036 533458
rect 42984 533394 43036 533400
rect 42720 531406 42840 531434
rect 42720 530233 42748 531406
rect 42706 530224 42762 530233
rect 42706 530159 42762 530168
rect 42536 530046 42656 530074
rect 42338 529952 42394 529961
rect 42338 529887 42394 529896
rect 41878 529408 41934 529417
rect 41878 529343 41934 529352
rect 41892 529205 41920 529343
rect 42352 529122 42380 529887
rect 42260 529094 42380 529122
rect 42260 527762 42288 529094
rect 42430 529000 42486 529009
rect 42430 528935 42486 528944
rect 42168 527734 42288 527762
rect 42168 527340 42196 527734
rect 42444 526742 42472 528935
rect 42628 528554 42656 530046
rect 42182 526714 42472 526742
rect 42536 528526 42656 528554
rect 42536 526091 42564 528526
rect 42706 527232 42762 527241
rect 42706 527167 42762 527176
rect 42182 526063 42564 526091
rect 42720 525586 42748 527167
rect 42168 525558 42288 525586
rect 42168 525504 42196 525558
rect 42260 525518 42288 525558
rect 42536 525558 42748 525586
rect 42536 525518 42564 525558
rect 42260 525490 42564 525518
rect 8588 431596 8616 431664
rect 9048 431596 9076 431664
rect 9508 431596 9536 431664
rect 9968 431596 9996 431664
rect 10428 431596 10456 431664
rect 10888 431596 10916 431664
rect 11348 431596 11376 431664
rect 11808 431596 11836 431664
rect 12268 431596 12296 431664
rect 12728 431596 12756 431664
rect 13188 431596 13216 431664
rect 13648 431596 13676 431664
rect 14108 431596 14136 431664
rect 35806 430128 35862 430137
rect 35806 430063 35862 430072
rect 35820 429214 35848 430063
rect 35808 429208 35860 429214
rect 35808 429150 35860 429156
rect 41328 429208 41380 429214
rect 41328 429150 41380 429156
rect 41142 426048 41198 426057
rect 41142 425983 41198 425992
rect 35162 425402 35218 425411
rect 35162 425337 35218 425346
rect 39302 425402 39358 425411
rect 41156 425406 41184 425983
rect 39302 425337 39358 425346
rect 41144 425400 41196 425406
rect 41144 425342 41196 425348
rect 33046 424824 33102 424833
rect 33046 424759 33102 424768
rect 33060 415954 33088 424759
rect 33782 424008 33838 424017
rect 33782 423943 33838 423952
rect 33048 415948 33100 415954
rect 33048 415890 33100 415896
rect 33796 414633 33824 423943
rect 35176 414905 35204 425337
rect 39316 415313 39344 425337
rect 41340 425054 41368 429150
rect 41696 425400 41748 425406
rect 41748 425348 42012 425354
rect 41696 425342 42012 425348
rect 41708 425326 42012 425342
rect 41340 425026 41828 425054
rect 40958 424416 41014 424425
rect 40958 424351 41014 424360
rect 40972 420986 41000 424351
rect 41800 424017 41828 425026
rect 41786 424008 41842 424017
rect 41786 423943 41842 423952
rect 41786 421968 41842 421977
rect 41524 421926 41786 421954
rect 40960 420980 41012 420986
rect 40960 420922 41012 420928
rect 41524 418713 41552 421926
rect 41786 421903 41842 421912
rect 41696 420980 41748 420986
rect 41696 420922 41748 420928
rect 41510 418704 41566 418713
rect 41510 418639 41566 418648
rect 40590 415984 40646 415993
rect 40590 415919 40592 415928
rect 40644 415919 40646 415928
rect 40592 415890 40644 415896
rect 41708 415426 41736 420922
rect 41984 418154 42012 425326
rect 42154 424008 42210 424017
rect 42154 423943 42210 423952
rect 42168 422929 42196 423943
rect 42798 423600 42854 423609
rect 42798 423535 42854 423544
rect 42154 422920 42210 422929
rect 42154 422855 42210 422864
rect 41984 418126 42380 418154
rect 41708 415398 42288 415426
rect 39302 415304 39358 415313
rect 39302 415239 39358 415248
rect 35162 414896 35218 414905
rect 35162 414831 35218 414840
rect 33782 414624 33838 414633
rect 33782 414559 33838 414568
rect 42260 413114 42288 415398
rect 42168 413086 42288 413114
rect 42168 412624 42196 413086
rect 42352 411346 42380 418126
rect 42614 415984 42670 415993
rect 42614 415919 42670 415928
rect 42168 411318 42380 411346
rect 42168 410788 42196 411318
rect 42182 410162 42472 410190
rect 42246 409864 42302 409873
rect 42246 409799 42302 409808
rect 42260 408966 42288 409799
rect 42182 408938 42288 408966
rect 42168 408218 42196 408340
rect 42168 408190 42288 408218
rect 42062 408096 42118 408105
rect 42062 408031 42118 408040
rect 42076 407796 42104 408031
rect 41800 407017 41828 407116
rect 41786 407008 41842 407017
rect 41786 406943 41842 406952
rect 42062 406736 42118 406745
rect 42062 406671 42118 406680
rect 42076 406504 42104 406671
rect 42260 406094 42288 408190
rect 42444 407289 42472 410162
rect 42430 407280 42486 407289
rect 42430 407215 42486 407224
rect 42248 406088 42300 406094
rect 42248 406030 42300 406036
rect 42628 405943 42656 415919
rect 42182 405915 42656 405943
rect 42248 405680 42300 405686
rect 42248 405622 42300 405628
rect 42260 404569 42288 405622
rect 42246 404560 42302 404569
rect 42246 404495 42302 404504
rect 41786 403880 41842 403889
rect 41786 403815 41842 403824
rect 41800 403444 41828 403815
rect 42812 402974 42840 423535
rect 43258 420744 43314 420753
rect 43258 420679 43314 420688
rect 43074 419520 43130 419529
rect 43074 419455 43130 419464
rect 42536 402946 42840 402974
rect 42338 402928 42394 402937
rect 42168 402886 42338 402914
rect 42168 402801 42196 402886
rect 42338 402863 42394 402872
rect 42536 402166 42564 402946
rect 42182 402138 42564 402166
rect 41786 401976 41842 401985
rect 41786 401911 41842 401920
rect 41800 401608 41828 401911
rect 42430 399800 42486 399809
rect 42182 399758 42430 399786
rect 42430 399735 42486 399744
rect 41786 399392 41842 399401
rect 41786 399327 41842 399336
rect 41800 399121 41828 399327
rect 41786 398848 41842 398857
rect 41786 398783 41842 398792
rect 41800 398480 41828 398783
rect 42168 395729 42196 397936
rect 42154 395720 42210 395729
rect 42154 395655 42210 395664
rect 8588 388348 8616 388484
rect 9048 388348 9076 388484
rect 9508 388348 9536 388484
rect 9968 388348 9996 388484
rect 10428 388348 10456 388484
rect 10888 388348 10916 388484
rect 11348 388348 11376 388484
rect 11808 388348 11836 388484
rect 12268 388348 12296 388484
rect 12728 388348 12756 388484
rect 13188 388348 13216 388484
rect 13648 388348 13676 388484
rect 14108 388348 14136 388484
rect 41142 387152 41198 387161
rect 41142 387087 41198 387096
rect 40958 385928 41014 385937
rect 40958 385863 41014 385872
rect 40972 382265 41000 385863
rect 40222 382256 40278 382265
rect 40222 382191 40278 382200
rect 40958 382256 41014 382265
rect 40958 382191 41014 382200
rect 40038 381848 40094 381857
rect 40038 381783 40094 381792
rect 32402 381440 32458 381449
rect 32402 381375 32458 381384
rect 32416 373318 32444 381375
rect 37922 381032 37978 381041
rect 37922 380967 37978 380976
rect 35806 376544 35862 376553
rect 35806 376479 35862 376488
rect 35820 376145 35848 376479
rect 35806 376136 35862 376145
rect 35806 376071 35862 376080
rect 32404 373312 32456 373318
rect 32404 373254 32456 373260
rect 37936 372366 37964 380967
rect 40052 376961 40080 381783
rect 40236 379001 40264 382191
rect 41156 381857 41184 387087
rect 41326 386744 41382 386753
rect 41326 386679 41382 386688
rect 41340 385937 41368 386679
rect 41326 385928 41382 385937
rect 41326 385863 41382 385872
rect 41326 382664 41382 382673
rect 41326 382599 41382 382608
rect 41340 382430 41368 382599
rect 41328 382424 41380 382430
rect 41328 382366 41380 382372
rect 41696 382424 41748 382430
rect 41696 382366 41748 382372
rect 41142 381848 41198 381857
rect 41142 381783 41198 381792
rect 41708 379514 41736 382366
rect 42798 379944 42854 379953
rect 42798 379879 42854 379888
rect 41708 379486 42472 379514
rect 40222 378992 40278 379001
rect 40222 378927 40278 378936
rect 40038 376952 40094 376961
rect 40038 376887 40094 376896
rect 39026 376544 39082 376553
rect 39026 376479 39082 376488
rect 39040 376145 39068 376479
rect 39026 376136 39082 376145
rect 39026 376071 39082 376080
rect 41696 373312 41748 373318
rect 41748 373260 42104 373266
rect 41696 373254 42104 373260
rect 41708 373250 42104 373254
rect 41708 373244 42116 373250
rect 41708 373238 42064 373244
rect 42064 373186 42116 373192
rect 37924 372360 37976 372366
rect 37924 372302 37976 372308
rect 41696 372360 41748 372366
rect 41696 372302 41748 372308
rect 41708 372178 41736 372302
rect 41708 372150 42288 372178
rect 42260 369458 42288 372150
rect 42182 369430 42288 369458
rect 42444 367622 42472 379486
rect 42616 373244 42668 373250
rect 42616 373186 42668 373192
rect 42628 369854 42656 373186
rect 42628 369826 42748 369854
rect 42182 367594 42472 367622
rect 42182 366947 42472 366975
rect 41800 365673 41828 365772
rect 41786 365664 41842 365673
rect 41786 365599 41842 365608
rect 42182 365107 42288 365135
rect 41800 364313 41828 364548
rect 42260 364426 42288 365107
rect 42260 364398 42380 364426
rect 41786 364304 41842 364313
rect 41786 364239 41842 364248
rect 42154 364304 42210 364313
rect 42154 364239 42210 364248
rect 42168 363936 42196 364239
rect 41786 363760 41842 363769
rect 41786 363695 41842 363704
rect 41800 363256 41828 363695
rect 42352 363202 42380 364398
rect 42260 363174 42380 363202
rect 42260 362953 42288 363174
rect 42444 363089 42472 366947
rect 42430 363080 42486 363089
rect 42430 363015 42486 363024
rect 42246 362944 42302 362953
rect 42246 362879 42302 362888
rect 42168 362766 42288 362794
rect 42168 362712 42196 362766
rect 42260 362726 42288 362766
rect 42720 362726 42748 369826
rect 42260 362698 42748 362726
rect 42168 360210 42196 360264
rect 42260 360250 42472 360278
rect 42260 360210 42288 360250
rect 42168 360182 42288 360210
rect 42156 359984 42208 359990
rect 42156 359926 42208 359932
rect 42168 359584 42196 359926
rect 42062 359272 42118 359281
rect 42062 359207 42118 359216
rect 42076 358972 42104 359207
rect 42444 358737 42472 360250
rect 42812 359990 42840 379879
rect 42800 359984 42852 359990
rect 42800 359926 42852 359932
rect 41878 358728 41934 358737
rect 41878 358663 41934 358672
rect 42430 358728 42486 358737
rect 42430 358663 42486 358672
rect 41892 358428 41920 358663
rect 41786 356960 41842 356969
rect 41786 356895 41842 356904
rect 41800 356592 41828 356895
rect 42182 355898 42472 355926
rect 41878 355600 41934 355609
rect 41878 355535 41934 355544
rect 41892 355300 41920 355535
rect 42168 353297 42196 354725
rect 42154 353288 42210 353297
rect 42154 353223 42210 353232
rect 42444 353025 42472 355898
rect 43088 353977 43116 419455
rect 43074 353968 43130 353977
rect 43074 353903 43130 353912
rect 43272 353705 43300 420679
rect 43456 354674 43484 582346
rect 43640 379514 43668 589047
rect 44192 581233 44220 591903
rect 44178 581224 44234 581233
rect 44178 581159 44234 581168
rect 44376 578105 44404 593127
rect 44362 578096 44418 578105
rect 44362 578031 44418 578040
rect 44652 558793 44680 600063
rect 44914 598496 44970 598505
rect 44914 598431 44970 598440
rect 44638 558784 44694 558793
rect 44638 558719 44694 558728
rect 44546 556880 44602 556889
rect 44546 556815 44602 556824
rect 44362 551576 44418 551585
rect 44362 551511 44418 551520
rect 44178 549128 44234 549137
rect 44178 549063 44234 549072
rect 43810 548312 43866 548321
rect 43810 548247 43866 548256
rect 43824 379514 43852 548247
rect 43994 547088 44050 547097
rect 43994 547023 44050 547032
rect 43640 379486 43760 379514
rect 43824 379486 43944 379514
rect 43732 354674 43760 379486
rect 43916 354929 43944 379486
rect 44008 355042 44036 547023
rect 44192 537577 44220 549063
rect 44178 537568 44234 537577
rect 44178 537503 44234 537512
rect 44376 529009 44404 551511
rect 44362 529000 44418 529009
rect 44362 528935 44418 528944
rect 44560 429729 44588 556815
rect 44730 556064 44786 556073
rect 44730 555999 44786 556008
rect 44744 553394 44772 555999
rect 44928 555665 44956 598431
rect 45204 598097 45232 640183
rect 45388 598913 45416 640290
rect 45572 612105 45600 763263
rect 46216 743782 46244 773026
rect 58624 763224 58676 763230
rect 58624 763166 58676 763172
rect 46204 743776 46256 743782
rect 46204 743718 46256 743724
rect 46204 730312 46256 730318
rect 46204 730254 46256 730260
rect 46216 698222 46244 730254
rect 47214 721168 47270 721177
rect 47214 721103 47270 721112
rect 47030 719944 47086 719953
rect 47030 719879 47086 719888
rect 46204 698216 46256 698222
rect 46204 698158 46256 698164
rect 45558 612096 45614 612105
rect 47044 612066 47072 719879
rect 45558 612031 45614 612040
rect 47032 612060 47084 612066
rect 47032 612002 47084 612008
rect 47228 611930 47256 721103
rect 57244 719024 57296 719030
rect 57244 718966 57296 718972
rect 50344 712156 50396 712162
rect 50344 712098 50396 712104
rect 50356 705158 50384 712098
rect 50344 705152 50396 705158
rect 50344 705094 50396 705100
rect 55864 676252 55916 676258
rect 55864 676194 55916 676200
rect 53104 669384 53156 669390
rect 53104 669326 53156 669332
rect 53116 660958 53144 669326
rect 53104 660952 53156 660958
rect 53104 660894 53156 660900
rect 54484 644496 54536 644502
rect 54484 644438 54536 644444
rect 54496 612678 54524 644438
rect 54484 612672 54536 612678
rect 54484 612614 54536 612620
rect 47216 611924 47268 611930
rect 47216 611866 47268 611872
rect 45374 598904 45430 598913
rect 45374 598839 45430 598848
rect 45190 598088 45246 598097
rect 45190 598023 45246 598032
rect 45098 580680 45154 580689
rect 45098 580615 45154 580624
rect 45112 575482 45140 580615
rect 45558 578912 45614 578921
rect 45558 578847 45614 578856
rect 45100 575476 45152 575482
rect 45100 575418 45152 575424
rect 45572 574054 45600 578847
rect 45560 574048 45612 574054
rect 45560 573990 45612 573996
rect 54482 558512 54538 558521
rect 54482 558447 54538 558456
rect 44914 555656 44970 555665
rect 44914 555591 44970 555600
rect 45834 555248 45890 555257
rect 45834 555183 45890 555192
rect 45650 554432 45706 554441
rect 45650 554367 45706 554376
rect 44744 553366 44956 553394
rect 44730 535800 44786 535809
rect 44730 535735 44786 535744
rect 44744 531282 44772 535735
rect 44732 531276 44784 531282
rect 44732 531218 44784 531224
rect 44546 429720 44602 429729
rect 44546 429655 44602 429664
rect 44270 429312 44326 429321
rect 44270 429247 44326 429256
rect 44284 386481 44312 429247
rect 44928 428913 44956 553366
rect 45098 550760 45154 550769
rect 45098 550695 45154 550704
rect 45112 533905 45140 550695
rect 45282 548720 45338 548729
rect 45282 548655 45338 548664
rect 45296 535537 45324 548655
rect 45282 535528 45338 535537
rect 45282 535463 45338 535472
rect 45098 533896 45154 533905
rect 45098 533831 45154 533840
rect 45100 528624 45152 528630
rect 45100 528566 45152 528572
rect 45112 527241 45140 528566
rect 45098 527232 45154 527241
rect 45098 527167 45154 527176
rect 44914 428904 44970 428913
rect 44914 428839 44970 428848
rect 44638 428496 44694 428505
rect 44638 428431 44694 428440
rect 44454 421560 44510 421569
rect 44454 421495 44510 421504
rect 44468 406745 44496 421495
rect 44454 406736 44510 406745
rect 44454 406671 44510 406680
rect 44270 386472 44326 386481
rect 44270 386407 44326 386416
rect 44652 385665 44680 428431
rect 45664 427938 45692 554367
rect 45848 428097 45876 555183
rect 47582 547496 47638 547505
rect 47582 547431 47638 547440
rect 45834 428088 45890 428097
rect 45834 428023 45890 428032
rect 45664 427910 45784 427938
rect 45558 427680 45614 427689
rect 45558 427615 45614 427624
rect 44914 423192 44970 423201
rect 44914 423127 44970 423136
rect 44928 402937 44956 423127
rect 45098 422648 45154 422657
rect 45098 422583 45154 422592
rect 45112 409873 45140 422583
rect 45282 421152 45338 421161
rect 45282 421087 45338 421096
rect 45098 409864 45154 409873
rect 45098 409799 45154 409808
rect 45296 408105 45324 421087
rect 45282 408096 45338 408105
rect 45282 408031 45338 408040
rect 45098 407280 45154 407289
rect 45098 407215 45154 407224
rect 45112 404326 45140 407215
rect 45100 404320 45152 404326
rect 45100 404262 45152 404268
rect 44914 402928 44970 402937
rect 44914 402863 44970 402872
rect 44638 385656 44694 385665
rect 44638 385591 44694 385600
rect 45098 385248 45154 385257
rect 45098 385183 45154 385192
rect 44914 382256 44970 382265
rect 44914 382191 44970 382200
rect 44454 380352 44510 380361
rect 44454 380287 44510 380296
rect 44178 377496 44234 377505
rect 44178 377431 44234 377440
rect 44192 359122 44220 377431
rect 44468 359281 44496 380287
rect 44638 379400 44694 379409
rect 44638 379335 44694 379344
rect 44652 364313 44680 379335
rect 44638 364304 44694 364313
rect 44638 364239 44694 364248
rect 44928 360194 44956 382191
rect 45112 360194 45140 385183
rect 45572 384849 45600 427615
rect 45756 427281 45784 427910
rect 45742 427272 45798 427281
rect 45742 427207 45798 427216
rect 45926 426864 45982 426873
rect 45926 426799 45982 426808
rect 45742 426456 45798 426465
rect 45742 426391 45798 426400
rect 45756 399809 45784 426391
rect 45742 399800 45798 399809
rect 45742 399735 45798 399744
rect 45558 384840 45614 384849
rect 45558 384775 45614 384784
rect 45558 384432 45614 384441
rect 45558 384367 45614 384376
rect 45374 363080 45430 363089
rect 45374 363015 45430 363024
rect 45388 361554 45416 363015
rect 45376 361548 45428 361554
rect 45376 361490 45428 361496
rect 44836 360166 44956 360194
rect 45020 360166 45140 360194
rect 44454 359272 44510 359281
rect 44454 359207 44510 359216
rect 44192 359106 44680 359122
rect 44192 359100 44692 359106
rect 44192 359094 44640 359100
rect 44640 359042 44692 359048
rect 44008 355026 44680 355042
rect 44008 355020 44692 355026
rect 44008 355014 44640 355020
rect 44640 354962 44692 354968
rect 43902 354920 43958 354929
rect 43902 354855 43958 354864
rect 44640 354680 44692 354686
rect 43456 354646 43668 354674
rect 43732 354646 44640 354674
rect 43640 354498 43668 354646
rect 44836 354674 44864 360166
rect 45020 354674 45048 360166
rect 45376 359100 45428 359106
rect 45376 359042 45428 359048
rect 45190 354920 45246 354929
rect 45190 354855 45246 354864
rect 45204 354674 45232 354855
rect 45388 354674 45416 359042
rect 44836 354646 44956 354674
rect 45020 354646 45140 354674
rect 45204 354646 45324 354674
rect 45388 354646 45508 354674
rect 44640 354622 44692 354628
rect 43640 354482 44772 354498
rect 43640 354476 44784 354482
rect 43640 354470 44732 354476
rect 44732 354418 44784 354424
rect 43258 353696 43314 353705
rect 43258 353631 43314 353640
rect 42430 353016 42486 353025
rect 42430 352951 42486 352960
rect 8588 345100 8616 345236
rect 9048 345100 9076 345236
rect 9508 345100 9536 345236
rect 9968 345100 9996 345236
rect 10428 345100 10456 345236
rect 10888 345100 10916 345236
rect 11348 345100 11376 345236
rect 11808 345100 11836 345236
rect 12268 345100 12296 345236
rect 12728 345100 12756 345236
rect 13188 345100 13216 345236
rect 13648 345100 13676 345236
rect 14108 345100 14136 345236
rect 35808 344616 35860 344622
rect 35808 344558 35860 344564
rect 40040 344616 40092 344622
rect 40040 344558 40092 344564
rect 35820 344321 35848 344558
rect 35530 344312 35586 344321
rect 35530 344247 35586 344256
rect 35806 344312 35862 344321
rect 35806 344247 35862 344256
rect 39670 344312 39726 344321
rect 39670 344247 39726 344256
rect 35544 343806 35572 344247
rect 35532 343800 35584 343806
rect 35532 343742 35584 343748
rect 35806 343496 35862 343505
rect 35806 343431 35862 343440
rect 35820 342242 35848 343431
rect 35808 342236 35860 342242
rect 35808 342178 35860 342184
rect 39486 341864 39542 341873
rect 39486 341799 39542 341808
rect 35622 341456 35678 341465
rect 35622 341391 35678 341400
rect 35636 341086 35664 341391
rect 35808 341216 35860 341222
rect 35808 341158 35860 341164
rect 35624 341080 35676 341086
rect 35820 341057 35848 341158
rect 35624 341022 35676 341028
rect 35806 341048 35862 341057
rect 35806 340983 35862 340992
rect 39500 340241 39528 341799
rect 39684 341086 39712 344247
rect 39856 343800 39908 343806
rect 39856 343742 39908 343748
rect 39868 341465 39896 343742
rect 40052 341873 40080 344558
rect 44928 343369 44956 354646
rect 44914 343360 44970 343369
rect 44914 343295 44970 343304
rect 45112 342553 45140 354646
rect 45296 354414 45324 354646
rect 45284 354408 45336 354414
rect 45284 354350 45336 354356
rect 45282 353968 45338 353977
rect 45282 353903 45284 353912
rect 45336 353903 45338 353912
rect 45284 353874 45336 353880
rect 45303 353728 45355 353734
rect 45282 353696 45303 353705
rect 45338 353670 45355 353676
rect 45338 353654 45343 353670
rect 45282 353631 45338 353640
rect 45480 353274 45508 354646
rect 45434 353258 45508 353274
rect 45422 353252 45508 353258
rect 45474 353246 45508 353252
rect 45422 353194 45474 353200
rect 45572 344321 45600 384367
rect 45940 384033 45968 426799
rect 46110 404560 46166 404569
rect 46110 404495 46166 404504
rect 46124 402966 46152 404495
rect 46112 402960 46164 402966
rect 46112 402902 46164 402908
rect 47596 397458 47624 547431
rect 53102 539608 53158 539617
rect 53102 539543 53158 539552
rect 53116 531146 53144 539543
rect 53104 531140 53156 531146
rect 53104 531082 53156 531088
rect 54496 527134 54524 558447
rect 54484 527128 54536 527134
rect 54484 527070 54536 527076
rect 47950 430944 48006 430953
rect 47950 430879 48006 430888
rect 47766 419928 47822 419937
rect 47766 419863 47822 419872
rect 47584 397452 47636 397458
rect 47584 397394 47636 397400
rect 45926 384024 45982 384033
rect 45926 383959 45982 383968
rect 46202 383616 46258 383625
rect 46202 383551 46258 383560
rect 46018 380760 46074 380769
rect 46018 380695 46074 380704
rect 45834 376272 45890 376281
rect 45834 376207 45890 376216
rect 45848 353530 45876 376207
rect 45836 353524 45888 353530
rect 45836 353466 45888 353472
rect 46032 353138 46060 380695
rect 46216 369854 46244 383551
rect 46478 378720 46534 378729
rect 46478 378655 46534 378664
rect 45940 353110 46060 353138
rect 46124 369826 46244 369854
rect 45940 353025 45968 353110
rect 45926 353016 45982 353025
rect 45926 352951 45982 352960
rect 45558 344312 45614 344321
rect 45558 344247 45614 344256
rect 45098 342544 45154 342553
rect 45098 342479 45154 342488
rect 40222 342272 40278 342281
rect 40222 342207 40224 342216
rect 40276 342207 40278 342216
rect 45466 342272 45522 342281
rect 45466 342207 45468 342216
rect 40224 342178 40276 342184
rect 45520 342207 45522 342216
rect 45468 342178 45520 342184
rect 40038 341864 40094 341873
rect 40038 341799 40094 341808
rect 39854 341456 39910 341465
rect 39854 341391 39910 341400
rect 40224 341216 40276 341222
rect 40224 341158 40276 341164
rect 39672 341080 39724 341086
rect 40236 341057 40264 341158
rect 39672 341022 39724 341028
rect 40222 341048 40278 341057
rect 40222 340983 40278 340992
rect 46124 340785 46152 369826
rect 46492 358737 46520 378655
rect 47582 376680 47638 376689
rect 47582 376615 47638 376624
rect 46754 362672 46810 362681
rect 46754 362607 46810 362616
rect 46768 360194 46796 362607
rect 46756 360188 46808 360194
rect 46756 360130 46808 360136
rect 46478 358728 46534 358737
rect 46478 358663 46534 358672
rect 46110 340776 46166 340785
rect 46110 340711 46166 340720
rect 39486 340232 39542 340241
rect 39486 340167 39542 340176
rect 35530 339824 35586 339833
rect 35530 339759 35586 339768
rect 35806 339824 35862 339833
rect 35806 339759 35862 339768
rect 35544 339658 35572 339759
rect 35532 339652 35584 339658
rect 35532 339594 35584 339600
rect 35820 339522 35848 339759
rect 36544 339652 36596 339658
rect 36544 339594 36596 339600
rect 35808 339516 35860 339522
rect 35808 339458 35860 339464
rect 35162 338600 35218 338609
rect 35162 338535 35218 338544
rect 35176 330449 35204 338535
rect 35808 336252 35860 336258
rect 35808 336194 35860 336200
rect 35820 335753 35848 336194
rect 35530 335744 35586 335753
rect 35530 335679 35586 335688
rect 35806 335744 35862 335753
rect 35806 335679 35862 335688
rect 35544 335374 35572 335679
rect 35532 335368 35584 335374
rect 35532 335310 35584 335316
rect 35806 334520 35862 334529
rect 35806 334455 35862 334464
rect 35820 334150 35848 334455
rect 35808 334144 35860 334150
rect 35808 334086 35860 334092
rect 35806 332888 35862 332897
rect 35806 332823 35862 332832
rect 35820 331809 35848 332823
rect 35806 331800 35862 331809
rect 35806 331735 35862 331744
rect 36556 331265 36584 339594
rect 38568 339516 38620 339522
rect 38568 339458 38620 339464
rect 38580 335753 38608 339458
rect 45650 339280 45706 339289
rect 45650 339215 45706 339224
rect 45466 338056 45522 338065
rect 45466 337991 45522 338000
rect 40040 336252 40092 336258
rect 40040 336194 40092 336200
rect 38566 335744 38622 335753
rect 38566 335679 38622 335688
rect 40052 334529 40080 336194
rect 40224 335368 40276 335374
rect 40224 335310 40276 335316
rect 40038 334520 40094 334529
rect 40038 334455 40094 334464
rect 39764 334144 39816 334150
rect 39764 334086 39816 334092
rect 39776 332897 39804 334086
rect 39762 332888 39818 332897
rect 39762 332823 39818 332832
rect 40236 332489 40264 335310
rect 44178 334656 44234 334665
rect 44178 334591 44234 334600
rect 42798 334384 42854 334393
rect 42798 334319 42854 334328
rect 40222 332480 40278 332489
rect 40222 332415 40278 332424
rect 36542 331256 36598 331265
rect 36542 331191 36598 331200
rect 35162 330440 35218 330449
rect 35162 330375 35218 330384
rect 42430 327040 42486 327049
rect 42430 326975 42486 326984
rect 42444 326278 42472 326975
rect 42168 326210 42196 326264
rect 42260 326250 42472 326278
rect 42260 326210 42288 326250
rect 42168 326182 42288 326210
rect 41786 324864 41842 324873
rect 41786 324799 41842 324808
rect 41800 324428 41828 324799
rect 42182 323734 42472 323762
rect 41786 322824 41842 322833
rect 41786 322759 41842 322768
rect 41800 322592 41828 322759
rect 42182 321898 42288 321926
rect 42076 321201 42104 321368
rect 42062 321192 42118 321201
rect 42062 321127 42118 321136
rect 42168 320521 42196 320725
rect 42260 320634 42288 321898
rect 42444 320793 42472 323734
rect 42430 320784 42486 320793
rect 42430 320719 42486 320728
rect 42260 320606 42380 320634
rect 42154 320512 42210 320521
rect 42154 320447 42210 320456
rect 42352 320113 42380 320606
rect 42338 320104 42394 320113
rect 42168 319954 42196 320076
rect 42338 320039 42394 320048
rect 42168 319938 42288 319954
rect 42168 319932 42300 319938
rect 42168 319926 42248 319932
rect 42248 319874 42300 319880
rect 42430 319696 42486 319705
rect 42430 319631 42486 319640
rect 42444 319546 42472 319631
rect 42182 319518 42472 319546
rect 42812 317098 42840 334319
rect 42982 332888 43038 332897
rect 42982 332823 43038 332832
rect 42996 321201 43024 332823
rect 43166 332480 43222 332489
rect 43166 332415 43222 332424
rect 42982 321192 43038 321201
rect 42982 321127 43038 321136
rect 43180 320521 43208 332415
rect 43166 320512 43222 320521
rect 43166 320447 43222 320456
rect 44192 319954 44220 334591
rect 45282 327040 45338 327049
rect 45480 327026 45508 337991
rect 45664 331214 45692 339215
rect 46938 338464 46994 338473
rect 46938 338399 46994 338408
rect 45338 326998 45508 327026
rect 45572 331186 45692 331214
rect 45282 326975 45338 326984
rect 43364 319938 44220 319954
rect 43352 319932 44220 319938
rect 43404 319926 44220 319932
rect 43352 319874 43404 319880
rect 42536 317070 42840 317098
rect 42536 317059 42564 317070
rect 42182 317031 42564 317059
rect 41786 316840 41842 316849
rect 41786 316775 41842 316784
rect 41800 316404 41828 316775
rect 41786 316024 41842 316033
rect 41786 315959 41842 315968
rect 41800 315757 41828 315959
rect 41786 315616 41842 315625
rect 41786 315551 41842 315560
rect 41800 315180 41828 315551
rect 41786 313712 41842 313721
rect 41786 313647 41842 313656
rect 41800 313344 41828 313647
rect 42430 312760 42486 312769
rect 42182 312718 42430 312746
rect 42430 312695 42486 312704
rect 45572 312361 45600 331186
rect 46952 319705 46980 338399
rect 46938 319696 46994 319705
rect 46938 319631 46994 319640
rect 42154 312352 42210 312361
rect 42154 312287 42210 312296
rect 45558 312352 45614 312361
rect 45558 312287 45614 312296
rect 42168 312052 42196 312287
rect 42076 310457 42104 311508
rect 42062 310448 42118 310457
rect 42062 310383 42118 310392
rect 8588 301988 8616 302124
rect 9048 301988 9076 302124
rect 9508 301988 9536 302124
rect 9968 301988 9996 302124
rect 10428 301988 10456 302124
rect 10888 301988 10916 302124
rect 11348 301988 11376 302124
rect 11808 301988 11836 302124
rect 12268 301988 12296 302124
rect 12728 301988 12756 302124
rect 13188 301988 13216 302124
rect 13648 301988 13676 302124
rect 14108 301988 14136 302124
rect 47596 301782 47624 376615
rect 47584 301776 47636 301782
rect 47584 301718 47636 301724
rect 35622 300928 35678 300937
rect 35622 300863 35678 300872
rect 35636 298790 35664 300863
rect 46202 300520 46258 300529
rect 46202 300455 46258 300464
rect 44178 299704 44234 299713
rect 44178 299639 44234 299648
rect 35806 298888 35862 298897
rect 35806 298823 35862 298832
rect 35624 298784 35676 298790
rect 35624 298726 35676 298732
rect 35820 298314 35848 298823
rect 41604 298784 41656 298790
rect 41786 298752 41842 298761
rect 41656 298732 41786 298738
rect 41604 298726 41786 298732
rect 41616 298710 41786 298726
rect 41786 298687 41842 298696
rect 35808 298308 35860 298314
rect 35808 298250 35860 298256
rect 41604 298308 41656 298314
rect 41604 298250 41656 298256
rect 41616 297378 41644 298250
rect 41786 297392 41842 297401
rect 41616 297350 41786 297378
rect 41786 297327 41842 297336
rect 42798 297392 42854 297401
rect 42798 297327 42854 297336
rect 35806 297256 35862 297265
rect 35806 297191 35862 297200
rect 35820 296750 35848 297191
rect 35808 296744 35860 296750
rect 35808 296686 35860 296692
rect 41604 296744 41656 296750
rect 41604 296686 41656 296692
rect 41616 296562 41644 296686
rect 41786 296576 41842 296585
rect 41616 296534 41786 296562
rect 41786 296511 41842 296520
rect 35438 296440 35494 296449
rect 35438 296375 35494 296384
rect 31022 294808 31078 294817
rect 31022 294743 31078 294752
rect 31036 286346 31064 294743
rect 35452 294642 35480 296375
rect 35622 296032 35678 296041
rect 35622 295967 35678 295976
rect 35636 295526 35664 295967
rect 35806 295624 35862 295633
rect 35806 295559 35862 295568
rect 35624 295520 35676 295526
rect 35624 295462 35676 295468
rect 35820 295390 35848 295559
rect 39304 295520 39356 295526
rect 39304 295462 39356 295468
rect 35808 295384 35860 295390
rect 35808 295326 35860 295332
rect 35806 295216 35862 295225
rect 35806 295151 35862 295160
rect 35440 294636 35492 294642
rect 35440 294578 35492 294584
rect 35820 294030 35848 295151
rect 35808 294024 35860 294030
rect 35808 293966 35860 293972
rect 35806 293584 35862 293593
rect 35806 293519 35862 293528
rect 35820 292942 35848 293519
rect 35808 292936 35860 292942
rect 35808 292878 35860 292884
rect 35806 292768 35862 292777
rect 35806 292703 35862 292712
rect 35820 292602 35848 292703
rect 35808 292596 35860 292602
rect 35808 292538 35860 292544
rect 35806 290320 35862 290329
rect 35806 290255 35862 290264
rect 31024 286340 31076 286346
rect 31024 286282 31076 286288
rect 35820 284986 35848 290255
rect 35808 284980 35860 284986
rect 35808 284922 35860 284928
rect 39316 284345 39344 295462
rect 41328 295384 41380 295390
rect 41328 295326 41380 295332
rect 40040 294024 40092 294030
rect 40040 293966 40092 293972
rect 39856 292868 39908 292874
rect 39856 292810 39908 292816
rect 39868 291174 39896 292810
rect 40052 291378 40080 293966
rect 40774 292588 40830 292597
rect 40774 292523 40830 292532
rect 40788 292126 40816 292523
rect 41340 292482 41368 295326
rect 41696 294636 41748 294642
rect 41696 294578 41748 294584
rect 41708 294522 41736 294578
rect 41708 294494 41920 294522
rect 41892 292574 41920 294494
rect 41892 292546 42472 292574
rect 41786 292496 41842 292505
rect 41340 292454 41786 292482
rect 41786 292431 41842 292440
rect 41604 292392 41656 292398
rect 41604 292334 41656 292340
rect 41616 292210 41644 292334
rect 41786 292224 41842 292233
rect 41616 292182 41786 292210
rect 41786 292159 41842 292168
rect 40776 292120 40828 292126
rect 40776 292062 40828 292068
rect 41604 292120 41656 292126
rect 41604 292062 41656 292068
rect 41616 291938 41644 292062
rect 41786 291952 41842 291961
rect 41616 291910 41786 291938
rect 41786 291887 41842 291896
rect 40040 291372 40092 291378
rect 40040 291314 40092 291320
rect 41696 291372 41748 291378
rect 41696 291314 41748 291320
rect 42154 291374 42210 291383
rect 41708 291258 41736 291314
rect 42154 291309 42210 291318
rect 41708 291242 42104 291258
rect 41708 291236 42116 291242
rect 41708 291230 42064 291236
rect 42064 291178 42116 291184
rect 39856 291168 39908 291174
rect 39856 291110 39908 291116
rect 41604 291168 41656 291174
rect 41786 291136 41842 291145
rect 41656 291116 41786 291122
rect 41604 291110 41786 291116
rect 41616 291094 41786 291110
rect 41786 291071 41842 291080
rect 41512 286340 41564 286346
rect 41512 286282 41564 286288
rect 41524 284730 41552 286282
rect 41696 284980 41748 284986
rect 41696 284922 41748 284928
rect 41708 284866 41736 284922
rect 41708 284838 42380 284866
rect 41524 284702 42288 284730
rect 39302 284336 39358 284345
rect 39302 284271 39358 284280
rect 42260 283059 42288 284702
rect 42182 283031 42288 283059
rect 42352 281874 42380 284838
rect 42182 281846 42380 281874
rect 42168 281302 42288 281330
rect 42168 281180 42196 281302
rect 42260 281194 42288 281302
rect 42444 281194 42472 292546
rect 42616 291236 42668 291242
rect 42616 291178 42668 291184
rect 42260 281166 42472 281194
rect 42182 280554 42472 280582
rect 41786 279848 41842 279857
rect 41786 279783 41842 279792
rect 41800 279344 41828 279783
rect 42444 278769 42472 280554
rect 42430 278760 42486 278769
rect 42182 278718 42288 278746
rect 42062 278488 42118 278497
rect 42062 278423 42118 278432
rect 42076 278188 42104 278423
rect 42062 277944 42118 277953
rect 42062 277879 42118 277888
rect 42076 277508 42104 277879
rect 41786 277128 41842 277137
rect 41786 277063 41842 277072
rect 41800 276896 41828 277063
rect 42062 276720 42118 276729
rect 42062 276655 42118 276664
rect 42076 276352 42104 276655
rect 42260 275913 42288 278718
rect 42430 278695 42486 278704
rect 42628 276729 42656 291178
rect 42614 276720 42670 276729
rect 42614 276655 42670 276664
rect 42246 275904 42302 275913
rect 42246 275839 42302 275848
rect 41786 274272 41842 274281
rect 41786 274207 41842 274216
rect 41800 273836 41828 274207
rect 42168 273170 42196 273224
rect 42338 273184 42394 273193
rect 42168 273142 42338 273170
rect 42338 273119 42394 273128
rect 42430 272912 42486 272921
rect 42430 272847 42486 272856
rect 42444 272558 42472 272847
rect 42182 272530 42472 272558
rect 41786 272368 41842 272377
rect 41786 272303 41842 272312
rect 41800 272000 41828 272303
rect 41786 270464 41842 270473
rect 41786 270399 41842 270408
rect 42430 270464 42486 270473
rect 42430 270399 42486 270408
rect 41800 270164 41828 270399
rect 42444 269535 42472 270399
rect 42182 269507 42472 269535
rect 42062 269104 42118 269113
rect 42062 269039 42118 269048
rect 42076 268872 42104 269039
rect 40682 267064 40738 267073
rect 40682 266999 40738 267008
rect 8588 258740 8616 258876
rect 9048 258740 9076 258876
rect 9508 258740 9536 258876
rect 9968 258740 9996 258876
rect 10428 258740 10456 258876
rect 10888 258740 10916 258876
rect 11348 258740 11376 258876
rect 11808 258740 11836 258876
rect 12268 258740 12296 258876
rect 12728 258740 12756 258876
rect 13188 258740 13216 258876
rect 13648 258740 13676 258876
rect 14108 258740 14136 258876
rect 35806 257136 35862 257145
rect 35806 257071 35862 257080
rect 35820 256766 35848 257071
rect 40696 256766 40724 266999
rect 42168 266257 42196 268328
rect 42154 266248 42210 266257
rect 42154 266183 42210 266192
rect 35808 256760 35860 256766
rect 35808 256702 35860 256708
rect 40684 256760 40736 256766
rect 40684 256702 40736 256708
rect 42812 255921 42840 297327
rect 43166 296576 43222 296585
rect 43166 296511 43222 296520
rect 42982 292224 43038 292233
rect 42982 292159 43038 292168
rect 42996 277953 43024 292159
rect 42982 277944 43038 277953
rect 42982 277879 43038 277888
rect 35806 255912 35862 255921
rect 35806 255847 35862 255856
rect 39394 255912 39450 255921
rect 39394 255847 39450 255856
rect 42798 255912 42854 255921
rect 42798 255847 42854 255856
rect 35820 255474 35848 255847
rect 39408 255474 39436 255847
rect 35808 255468 35860 255474
rect 35808 255410 35860 255416
rect 39396 255468 39448 255474
rect 39396 255410 39448 255416
rect 35530 254280 35586 254289
rect 35530 254215 35586 254224
rect 35806 254280 35862 254289
rect 35806 254215 35808 254224
rect 35544 253978 35572 254215
rect 35860 254215 35862 254224
rect 39396 254244 39448 254250
rect 35808 254186 35860 254192
rect 39396 254186 39448 254192
rect 35532 253972 35584 253978
rect 35532 253914 35584 253920
rect 39408 253881 39436 254186
rect 43180 254046 43208 296511
rect 43352 291372 43404 291378
rect 43352 291314 43404 291320
rect 43364 282914 43392 291314
rect 43626 291136 43682 291145
rect 43626 291071 43682 291080
rect 43364 282886 43484 282914
rect 43456 263594 43484 282886
rect 43640 273193 43668 291071
rect 43626 273184 43682 273193
rect 43626 273119 43682 273128
rect 43456 263566 43576 263594
rect 42064 254040 42116 254046
rect 41708 253988 42064 253994
rect 41708 253982 42116 253988
rect 43168 254040 43220 254046
rect 43168 253982 43220 253988
rect 41708 253978 42104 253982
rect 41696 253972 42104 253978
rect 41748 253966 42104 253972
rect 41696 253914 41748 253920
rect 39394 253872 39450 253881
rect 39394 253807 39450 253816
rect 42890 253872 42946 253881
rect 42890 253807 42946 253816
rect 35806 253056 35862 253065
rect 35806 252991 35862 253000
rect 35820 252822 35848 252991
rect 35808 252816 35860 252822
rect 35808 252758 35860 252764
rect 41708 252754 42104 252770
rect 41696 252748 42116 252754
rect 41748 252742 42064 252748
rect 41696 252690 41748 252696
rect 42064 252690 42116 252696
rect 42708 252748 42760 252754
rect 42708 252690 42760 252696
rect 35806 252648 35862 252657
rect 35806 252583 35808 252592
rect 35860 252583 35862 252592
rect 41696 252612 41748 252618
rect 35808 252554 35860 252560
rect 41696 252554 41748 252560
rect 35806 250200 35862 250209
rect 35806 250135 35862 250144
rect 35820 249966 35848 250135
rect 35808 249960 35860 249966
rect 35808 249902 35860 249908
rect 39580 249960 39632 249966
rect 39580 249902 39632 249908
rect 35806 248568 35862 248577
rect 35806 248503 35808 248512
rect 35860 248503 35862 248512
rect 35808 248474 35860 248480
rect 35806 247752 35862 247761
rect 35806 247687 35862 247696
rect 35820 247246 35848 247687
rect 35808 247240 35860 247246
rect 35808 247182 35860 247188
rect 35808 247104 35860 247110
rect 35808 247046 35860 247052
rect 39396 247104 39448 247110
rect 39396 247046 39448 247052
rect 35820 246945 35848 247046
rect 35806 246936 35862 246945
rect 35806 246871 35862 246880
rect 39408 244769 39436 247046
rect 39394 244760 39450 244769
rect 39394 244695 39450 244704
rect 39592 244089 39620 249902
rect 40316 248532 40368 248538
rect 40316 248474 40368 248480
rect 40328 245721 40356 248474
rect 40958 247752 41014 247761
rect 40958 247687 41014 247696
rect 40972 247246 41000 247687
rect 40960 247240 41012 247246
rect 40960 247182 41012 247188
rect 40314 245712 40370 245721
rect 40314 245647 40370 245656
rect 41708 244274 41736 252554
rect 42522 244760 42578 244769
rect 42522 244695 42578 244704
rect 41708 244246 42288 244274
rect 39578 244080 39634 244089
rect 39578 244015 39634 244024
rect 42062 240136 42118 240145
rect 42062 240071 42118 240080
rect 42076 239836 42104 240071
rect 42260 238921 42288 244246
rect 42246 238912 42302 238921
rect 42246 238847 42302 238856
rect 42536 238663 42564 244695
rect 42720 244274 42748 252690
rect 42182 238635 42564 238663
rect 42628 244246 42748 244274
rect 42628 238082 42656 244246
rect 42904 240134 42932 253807
rect 43350 247752 43406 247761
rect 43350 247687 43406 247696
rect 43166 245712 43222 245721
rect 43166 245647 43222 245656
rect 43180 245562 43208 245647
rect 43180 245534 43300 245562
rect 43074 244080 43130 244089
rect 43074 244015 43130 244024
rect 42536 238054 42656 238082
rect 42812 240106 42932 240134
rect 42536 238014 42564 238054
rect 42182 237986 42564 238014
rect 41786 236600 41842 236609
rect 41786 236535 41842 236544
rect 41800 236164 41828 236535
rect 42430 235920 42486 235929
rect 42430 235855 42486 235864
rect 42444 234983 42472 235855
rect 42182 234955 42472 234983
rect 42182 234314 42472 234342
rect 42248 233980 42300 233986
rect 42248 233922 42300 233928
rect 42260 233695 42288 233922
rect 42182 233667 42288 233695
rect 42444 233345 42472 234314
rect 42430 233336 42486 233345
rect 42430 233271 42486 233280
rect 42168 233158 42288 233186
rect 42168 233104 42196 233158
rect 42260 233118 42288 233158
rect 42260 233090 42472 233118
rect 42444 231985 42472 233090
rect 42430 231976 42486 231985
rect 42430 231911 42486 231920
rect 42182 230642 42472 230670
rect 42156 230376 42208 230382
rect 42156 230318 42208 230324
rect 42168 229976 42196 230318
rect 41786 229664 41842 229673
rect 41786 229599 41842 229608
rect 41800 229364 41828 229599
rect 42444 228993 42472 230642
rect 42430 228984 42486 228993
rect 42430 228919 42486 228928
rect 42182 228806 42656 228834
rect 42430 227624 42486 227633
rect 42430 227559 42486 227568
rect 42444 226998 42472 227559
rect 42168 226930 42196 226984
rect 42260 226970 42472 226998
rect 42260 226930 42288 226970
rect 42168 226902 42288 226930
rect 42168 226358 42288 226386
rect 42168 226304 42196 226358
rect 42260 226318 42288 226358
rect 42260 226290 42472 226318
rect 41970 226128 42026 226137
rect 41970 226063 42026 226072
rect 41984 225692 42012 226063
rect 42168 223553 42196 225148
rect 42444 224913 42472 226290
rect 42628 226273 42656 228806
rect 42614 226264 42670 226273
rect 42614 226199 42670 226208
rect 42430 224904 42486 224913
rect 42430 224839 42486 224848
rect 42154 223544 42210 223553
rect 42154 223479 42210 223488
rect 35806 217968 35862 217977
rect 35806 217903 35862 217912
rect 8588 215492 8616 215628
rect 9048 215492 9076 215628
rect 9508 215492 9536 215628
rect 9968 215492 9996 215628
rect 10428 215492 10456 215628
rect 10888 215492 10916 215628
rect 11348 215492 11376 215628
rect 11808 215492 11836 215628
rect 12268 215492 12296 215628
rect 12728 215492 12756 215628
rect 13188 215492 13216 215628
rect 13648 215492 13676 215628
rect 14108 215492 14136 215628
rect 35820 214713 35848 217903
rect 35806 214704 35862 214713
rect 35806 214639 35862 214648
rect 35806 214296 35862 214305
rect 35806 214231 35808 214240
rect 35860 214231 35862 214240
rect 39670 214296 39726 214305
rect 39670 214231 39672 214240
rect 35808 214202 35860 214208
rect 39724 214231 39726 214240
rect 39672 214202 39724 214208
rect 35806 212256 35862 212265
rect 35806 212191 35862 212200
rect 35622 211848 35678 211857
rect 35622 211783 35678 211792
rect 35636 211342 35664 211783
rect 35820 211614 35848 212191
rect 42812 211857 42840 240106
rect 43088 230382 43116 244015
rect 43272 240134 43300 245534
rect 43180 240106 43300 240134
rect 43180 234002 43208 240106
rect 43364 235226 43392 247687
rect 43548 247058 43576 263566
rect 44192 256873 44220 299639
rect 44638 298072 44694 298081
rect 44638 298007 44694 298016
rect 44362 294400 44418 294409
rect 44362 294335 44418 294344
rect 44376 270473 44404 294335
rect 44362 270464 44418 270473
rect 44362 270399 44418 270408
rect 44178 256864 44234 256873
rect 44178 256799 44234 256808
rect 44362 256456 44418 256465
rect 44362 256391 44418 256400
rect 44178 254824 44234 254833
rect 44178 254759 44234 254768
rect 43456 247030 43576 247058
rect 43456 241514 43484 247030
rect 43456 241486 43668 241514
rect 43640 240134 43668 241486
rect 43640 240106 44036 240134
rect 43810 237960 43866 237969
rect 43810 237895 43866 237904
rect 43364 235198 43760 235226
rect 43180 233986 43300 234002
rect 43180 233980 43312 233986
rect 43180 233974 43260 233980
rect 43260 233922 43312 233928
rect 43442 230488 43498 230497
rect 43732 230474 43760 235198
rect 43442 230423 43498 230432
rect 43640 230446 43760 230474
rect 43076 230376 43128 230382
rect 43076 230318 43128 230324
rect 40130 211848 40186 211857
rect 40130 211783 40186 211792
rect 42798 211848 42854 211857
rect 42798 211783 42854 211792
rect 35808 211608 35860 211614
rect 35808 211550 35860 211556
rect 35806 211440 35862 211449
rect 35806 211375 35862 211384
rect 35624 211336 35676 211342
rect 35624 211278 35676 211284
rect 35820 211206 35848 211375
rect 40144 211206 40172 211783
rect 41512 211472 41564 211478
rect 41512 211414 41564 211420
rect 35808 211200 35860 211206
rect 35808 211142 35860 211148
rect 40132 211200 40184 211206
rect 40132 211142 40184 211148
rect 35530 210216 35586 210225
rect 35530 210151 35586 210160
rect 35806 210216 35862 210225
rect 35806 210151 35862 210160
rect 35544 209846 35572 210151
rect 35820 209982 35848 210151
rect 35808 209976 35860 209982
rect 35808 209918 35860 209924
rect 40132 209976 40184 209982
rect 40132 209918 40184 209924
rect 35532 209840 35584 209846
rect 35532 209782 35584 209788
rect 35806 209400 35862 209409
rect 35806 209335 35862 209344
rect 33046 208992 33102 209001
rect 33046 208927 33102 208936
rect 33060 202201 33088 208927
rect 35820 208622 35848 209335
rect 35808 208616 35860 208622
rect 35808 208558 35860 208564
rect 35806 207768 35862 207777
rect 35806 207703 35862 207712
rect 35820 207262 35848 207703
rect 40144 207369 40172 209918
rect 40776 209840 40828 209846
rect 40776 209782 40828 209788
rect 40788 209409 40816 209782
rect 40774 209400 40830 209409
rect 40774 209335 40830 209344
rect 40960 208616 41012 208622
rect 40960 208558 41012 208564
rect 40130 207360 40186 207369
rect 40130 207295 40186 207304
rect 35808 207256 35860 207262
rect 35808 207198 35860 207204
rect 40776 207256 40828 207262
rect 40776 207198 40828 207204
rect 40788 205737 40816 207198
rect 40972 206553 41000 208558
rect 41524 208185 41552 211414
rect 41696 211336 41748 211342
rect 41696 211278 41748 211284
rect 41510 208176 41566 208185
rect 41510 208111 41566 208120
rect 40958 206544 41014 206553
rect 40958 206479 41014 206488
rect 40774 205728 40830 205737
rect 40774 205663 40830 205672
rect 41708 205634 41736 211278
rect 42982 209400 43038 209409
rect 42982 209335 43038 209344
rect 42798 205728 42854 205737
rect 42798 205663 42854 205672
rect 41708 205606 41920 205634
rect 35622 205320 35678 205329
rect 35622 205255 35678 205264
rect 35636 204338 35664 205255
rect 35806 204504 35862 204513
rect 35806 204439 35808 204448
rect 35860 204439 35862 204448
rect 41694 204504 41750 204513
rect 41694 204439 41696 204448
rect 35808 204410 35860 204416
rect 41748 204439 41750 204448
rect 41696 204410 41748 204416
rect 35624 204332 35676 204338
rect 35624 204274 35676 204280
rect 41696 204332 41748 204338
rect 41696 204274 41748 204280
rect 41708 204105 41736 204274
rect 41694 204096 41750 204105
rect 41694 204031 41750 204040
rect 35806 203688 35862 203697
rect 35806 203623 35862 203632
rect 33046 202192 33102 202201
rect 33046 202127 33102 202136
rect 35820 200705 35848 203623
rect 41892 202201 41920 205606
rect 41878 202192 41934 202201
rect 41878 202127 41934 202136
rect 35806 200696 35862 200705
rect 35806 200631 35862 200640
rect 42430 197296 42486 197305
rect 42430 197231 42486 197240
rect 42444 196670 42472 197231
rect 42182 196642 42472 196670
rect 41786 195800 41842 195809
rect 41786 195735 41842 195744
rect 41800 195432 41828 195735
rect 41970 195120 42026 195129
rect 41970 195055 42026 195064
rect 41984 194820 42012 195055
rect 42430 193216 42486 193225
rect 42430 193151 42486 193160
rect 42444 192998 42472 193151
rect 42168 192930 42196 192984
rect 42260 192970 42472 192998
rect 42260 192930 42288 192970
rect 42168 192902 42288 192930
rect 42168 191706 42196 191760
rect 42338 191720 42394 191729
rect 42168 191678 42338 191706
rect 42338 191655 42394 191664
rect 41786 191584 41842 191593
rect 41786 191519 41842 191528
rect 41800 191148 41828 191519
rect 42430 190496 42486 190505
rect 42182 190454 42430 190482
rect 42430 190431 42486 190440
rect 42430 189952 42486 189961
rect 42182 189910 42430 189938
rect 42430 189887 42486 189896
rect 42430 187640 42486 187649
rect 42430 187575 42486 187584
rect 42444 187459 42472 187575
rect 42182 187431 42472 187459
rect 41786 187232 41842 187241
rect 41786 187167 41842 187176
rect 41800 186796 41828 187167
rect 41786 186416 41842 186425
rect 41786 186351 41842 186360
rect 41800 186184 41828 186351
rect 41786 186008 41842 186017
rect 41786 185943 41842 185952
rect 41800 185605 41828 185943
rect 42168 183530 42196 183765
rect 42156 183524 42208 183530
rect 42156 183466 42208 183472
rect 42812 183274 42840 205663
rect 42996 183530 43024 209335
rect 43166 206544 43222 206553
rect 43166 206479 43222 206488
rect 42984 183524 43036 183530
rect 42984 183466 43036 183472
rect 42536 183246 42840 183274
rect 42536 183138 42564 183246
rect 42182 183110 42564 183138
rect 42182 182463 42472 182491
rect 42444 182170 42472 182463
rect 43180 182170 43208 206479
rect 42432 182164 42484 182170
rect 42432 182106 42484 182112
rect 43168 182164 43220 182170
rect 43168 182106 43220 182112
rect 42076 179353 42104 181900
rect 42062 179344 42118 179353
rect 42062 179279 42118 179288
rect 43456 44198 43484 230423
rect 43640 44334 43668 230446
rect 43824 214305 43852 237895
rect 44008 230625 44036 240106
rect 43994 230616 44050 230625
rect 43994 230551 44050 230560
rect 43810 214296 43866 214305
rect 43810 214231 43866 214240
rect 44192 212129 44220 254759
rect 44376 213761 44404 256391
rect 44652 255241 44680 298007
rect 44822 293992 44878 294001
rect 44822 293927 44878 293936
rect 44836 272921 44864 293927
rect 46216 292466 46244 300455
rect 46204 292460 46256 292466
rect 46204 292402 46256 292408
rect 45006 291544 45062 291553
rect 45006 291479 45062 291488
rect 45020 278497 45048 291479
rect 46204 285728 46256 285734
rect 46204 285670 46256 285676
rect 45006 278488 45062 278497
rect 45006 278423 45062 278432
rect 44822 272912 44878 272921
rect 44822 272847 44878 272856
rect 46216 258097 46244 285670
rect 47584 284368 47636 284374
rect 47584 284310 47636 284316
rect 46202 258088 46258 258097
rect 46202 258023 46258 258032
rect 47596 257689 47624 284310
rect 47780 278730 47808 419863
rect 47964 400110 47992 430879
rect 54482 430536 54538 430545
rect 54482 430471 54538 430480
rect 51080 400240 51132 400246
rect 51080 400182 51132 400188
rect 47952 400104 48004 400110
rect 47952 400046 48004 400052
rect 50712 397452 50764 397458
rect 50712 397394 50764 397400
rect 47950 387696 48006 387705
rect 47950 387631 48006 387640
rect 47964 356046 47992 387631
rect 47952 356040 48004 356046
rect 47952 355982 48004 355988
rect 50342 331800 50398 331809
rect 50342 331735 50398 331744
rect 48962 289912 49018 289921
rect 48962 289847 49018 289856
rect 47952 280220 48004 280226
rect 47952 280162 48004 280168
rect 47768 278724 47820 278730
rect 47768 278666 47820 278672
rect 47582 257680 47638 257689
rect 47582 257615 47638 257624
rect 44914 255640 44970 255649
rect 44914 255575 44970 255584
rect 44638 255232 44694 255241
rect 44638 255167 44694 255176
rect 44546 251560 44602 251569
rect 44546 251495 44602 251504
rect 44560 240145 44588 251495
rect 44730 248296 44786 248305
rect 44730 248231 44786 248240
rect 44546 240136 44602 240145
rect 44546 240071 44602 240080
rect 44744 235929 44772 248231
rect 44730 235920 44786 235929
rect 44730 235855 44786 235864
rect 44928 234614 44956 255575
rect 45558 253600 45614 253609
rect 45558 253535 45614 253544
rect 44836 234586 44956 234614
rect 44362 213752 44418 213761
rect 44362 213687 44418 213696
rect 44836 212945 44864 234586
rect 45572 227633 45600 253535
rect 47214 252376 47270 252385
rect 47214 252311 47270 252320
rect 45926 251968 45982 251977
rect 45926 251903 45982 251912
rect 45742 249112 45798 249121
rect 45742 249047 45798 249056
rect 45756 228993 45784 249047
rect 45940 231985 45968 251903
rect 47030 251152 47086 251161
rect 47030 251087 47086 251096
rect 46110 249520 46166 249529
rect 46110 249455 46166 249464
rect 46124 233345 46152 249455
rect 46110 233336 46166 233345
rect 46110 233271 46166 233280
rect 45926 231976 45982 231985
rect 45926 231911 45982 231920
rect 45742 228984 45798 228993
rect 45742 228919 45798 228928
rect 45558 227624 45614 227633
rect 45558 227559 45614 227568
rect 47044 224913 47072 251087
rect 47228 226273 47256 252311
rect 47582 246664 47638 246673
rect 47582 246599 47638 246608
rect 47214 226264 47270 226273
rect 47214 226199 47270 226208
rect 47030 224904 47086 224913
rect 47030 224839 47086 224848
rect 44822 212936 44878 212945
rect 44822 212871 44878 212880
rect 44178 212120 44234 212129
rect 44178 212055 44234 212064
rect 46938 208856 46994 208865
rect 46938 208791 46994 208800
rect 44362 206816 44418 206825
rect 44362 206751 44418 206760
rect 44178 206000 44234 206009
rect 44178 205935 44234 205944
rect 43810 204504 43866 204513
rect 43810 204439 43866 204448
rect 43824 45218 43852 204439
rect 43994 204096 44050 204105
rect 43994 204031 44050 204040
rect 44008 190505 44036 204031
rect 43994 190496 44050 190505
rect 43994 190431 44050 190440
rect 44192 187649 44220 205935
rect 44376 193225 44404 206751
rect 44546 205184 44602 205193
rect 44546 205119 44602 205128
rect 44362 193216 44418 193225
rect 44362 193151 44418 193160
rect 44560 191729 44588 205119
rect 44822 204776 44878 204785
rect 44822 204711 44878 204720
rect 44546 191720 44602 191729
rect 44546 191655 44602 191664
rect 44178 187640 44234 187649
rect 44178 187575 44234 187584
rect 44836 74534 44864 204711
rect 46202 203552 46258 203561
rect 46202 203487 46258 203496
rect 44836 74506 45508 74534
rect 45480 50386 45508 74506
rect 46216 53106 46244 203487
rect 46952 189961 46980 208791
rect 47122 208448 47178 208457
rect 47122 208383 47178 208392
rect 47136 197305 47164 208383
rect 47122 197296 47178 197305
rect 47122 197231 47178 197240
rect 46938 189952 46994 189961
rect 46938 189887 46994 189896
rect 46204 53100 46256 53106
rect 46204 53042 46256 53048
rect 47596 51746 47624 246599
rect 47964 214985 47992 280162
rect 47950 214976 48006 214985
rect 47950 214911 48006 214920
rect 47766 213344 47822 213353
rect 47766 213279 47822 213288
rect 47780 190505 47808 213279
rect 47950 210896 48006 210905
rect 47950 210831 48006 210840
rect 47964 195922 47992 210831
rect 48594 202192 48650 202201
rect 48594 202127 48650 202136
rect 48608 196489 48636 202127
rect 48594 196480 48650 196489
rect 48594 196415 48650 196424
rect 47964 195894 48360 195922
rect 48332 194449 48360 195894
rect 48318 194440 48374 194449
rect 48318 194375 48374 194384
rect 47766 190496 47822 190505
rect 47766 190431 47822 190440
rect 48976 53242 49004 289847
rect 49146 247480 49202 247489
rect 49146 247415 49202 247424
rect 48964 53236 49016 53242
rect 48964 53178 49016 53184
rect 47584 51740 47636 51746
rect 47584 51682 47636 51688
rect 45468 50380 45520 50386
rect 45468 50322 45520 50328
rect 49160 49026 49188 247415
rect 49606 208176 49662 208185
rect 49606 208111 49662 208120
rect 49620 192409 49648 208111
rect 49606 192400 49662 192409
rect 49606 192335 49662 192344
rect 49148 49020 49200 49026
rect 49148 48962 49200 48968
rect 43812 45212 43864 45218
rect 43812 45154 43864 45160
rect 50356 44470 50384 331735
rect 50526 290728 50582 290737
rect 50526 290663 50582 290672
rect 50540 51882 50568 290663
rect 50724 278322 50752 397394
rect 51092 395729 51120 400182
rect 54496 398818 54524 430471
rect 54484 398812 54536 398818
rect 54484 398754 54536 398760
rect 51078 395720 51134 395729
rect 51078 395655 51134 395664
rect 51724 357468 51776 357474
rect 51724 357410 51776 357416
rect 51736 353297 51764 357410
rect 51722 353288 51778 353297
rect 51722 353223 51778 353232
rect 51722 334112 51778 334121
rect 51722 334047 51778 334056
rect 50712 278316 50764 278322
rect 50712 278258 50764 278264
rect 50712 218884 50764 218890
rect 50712 218826 50764 218832
rect 50724 179353 50752 218826
rect 50710 179344 50766 179353
rect 50710 179279 50766 179288
rect 51736 52018 51764 334047
rect 53838 320784 53894 320793
rect 53838 320719 53894 320728
rect 53102 320104 53158 320113
rect 53102 320039 53158 320048
rect 53116 315994 53144 320039
rect 53852 317422 53880 320719
rect 53840 317416 53892 317422
rect 53840 317358 53892 317364
rect 53104 315988 53156 315994
rect 53104 315930 53156 315936
rect 53840 314764 53892 314770
rect 53840 314706 53892 314712
rect 53852 310457 53880 314706
rect 53838 310448 53894 310457
rect 53838 310383 53894 310392
rect 51908 301776 51960 301782
rect 51908 301718 51960 301724
rect 51920 295118 51948 301718
rect 51908 295112 51960 295118
rect 51908 295054 51960 295060
rect 53104 294024 53156 294030
rect 53104 293966 53156 293972
rect 53116 275913 53144 293966
rect 54484 292596 54536 292602
rect 54484 292538 54536 292544
rect 53102 275904 53158 275913
rect 53102 275839 53158 275848
rect 54496 266257 54524 292538
rect 54482 266248 54538 266257
rect 54482 266183 54538 266192
rect 55876 264217 55904 676194
rect 56508 295112 56560 295118
rect 56508 295054 56560 295060
rect 56520 289814 56548 295054
rect 56508 289808 56560 289814
rect 56508 289750 56560 289756
rect 55862 264208 55918 264217
rect 55862 264143 55918 264152
rect 57256 231402 57284 718966
rect 57244 231396 57296 231402
rect 57244 231338 57296 231344
rect 58636 231130 58664 763166
rect 60016 742422 60044 774182
rect 61384 772880 61436 772886
rect 61384 772822 61436 772828
rect 61396 747182 61424 772822
rect 62764 755540 62816 755546
rect 62764 755482 62816 755488
rect 62776 747697 62804 755482
rect 62762 747688 62818 747697
rect 62762 747623 62818 747632
rect 61384 747176 61436 747182
rect 61384 747118 61436 747124
rect 63040 747176 63092 747182
rect 63040 747118 63092 747124
rect 62120 746564 62172 746570
rect 62120 746506 62172 746512
rect 62132 746201 62160 746506
rect 62118 746192 62174 746201
rect 62118 746127 62174 746136
rect 62118 744152 62174 744161
rect 62118 744087 62174 744096
rect 62132 743918 62160 744087
rect 62120 743912 62172 743918
rect 62120 743854 62172 743860
rect 62120 743776 62172 743782
rect 62118 743744 62120 743753
rect 62172 743744 62174 743753
rect 62118 743679 62174 743688
rect 60004 742416 60056 742422
rect 62120 742416 62172 742422
rect 60004 742358 60056 742364
rect 62118 742384 62120 742393
rect 62172 742384 62174 742393
rect 62118 742319 62174 742328
rect 63052 741849 63080 747118
rect 63038 741840 63094 741849
rect 63038 741775 63094 741784
rect 61384 730108 61436 730114
rect 61384 730050 61436 730056
rect 61396 699689 61424 730050
rect 62764 729360 62816 729366
rect 62764 729302 62816 729308
rect 62120 705152 62172 705158
rect 62120 705094 62172 705100
rect 62132 704449 62160 705094
rect 62118 704440 62174 704449
rect 62118 704375 62174 704384
rect 62120 703792 62172 703798
rect 62120 703734 62172 703740
rect 62132 703361 62160 703734
rect 62118 703352 62174 703361
rect 62118 703287 62174 703296
rect 62210 701312 62266 701321
rect 62210 701247 62266 701256
rect 62224 701078 62252 701247
rect 62212 701072 62264 701078
rect 62212 701014 62264 701020
rect 62776 700913 62804 729302
rect 62762 700904 62818 700913
rect 62762 700839 62818 700848
rect 61382 699680 61438 699689
rect 61382 699615 61438 699624
rect 62120 698216 62172 698222
rect 62118 698184 62120 698193
rect 62172 698184 62174 698193
rect 62118 698119 62174 698128
rect 61384 687268 61436 687274
rect 61384 687210 61436 687216
rect 60004 667956 60056 667962
rect 60004 667898 60056 667904
rect 60016 659598 60044 667898
rect 60004 659592 60056 659598
rect 60004 659534 60056 659540
rect 61396 656577 61424 687210
rect 62764 686520 62816 686526
rect 62764 686462 62816 686468
rect 62120 660952 62172 660958
rect 62118 660920 62120 660929
rect 62172 660920 62174 660929
rect 62118 660855 62174 660864
rect 62120 659592 62172 659598
rect 62118 659560 62120 659569
rect 62172 659560 62174 659569
rect 62118 659495 62174 659504
rect 62118 658336 62174 658345
rect 62118 658271 62174 658280
rect 62132 657558 62160 658271
rect 62776 657665 62804 686462
rect 62762 657656 62818 657665
rect 62762 657591 62818 657600
rect 62120 657552 62172 657558
rect 62120 657494 62172 657500
rect 61382 656568 61438 656577
rect 61382 656503 61438 656512
rect 62120 655512 62172 655518
rect 62120 655454 62172 655460
rect 62132 655353 62160 655454
rect 62118 655344 62174 655353
rect 62118 655279 62174 655288
rect 61384 643136 61436 643142
rect 61384 643078 61436 643084
rect 61396 613873 61424 643078
rect 62948 642388 63000 642394
rect 62948 642330 63000 642336
rect 62120 616820 62172 616826
rect 62120 616762 62172 616768
rect 62132 616593 62160 616762
rect 62118 616584 62174 616593
rect 62118 616519 62174 616528
rect 62118 614680 62174 614689
rect 62118 614615 62174 614624
rect 62132 614174 62160 614615
rect 62120 614168 62172 614174
rect 62120 614110 62172 614116
rect 61382 613864 61438 613873
rect 61382 613799 61438 613808
rect 62120 612672 62172 612678
rect 62118 612640 62120 612649
rect 62172 612640 62174 612649
rect 62118 612575 62174 612584
rect 62960 612105 62988 642330
rect 63408 633480 63460 633486
rect 63408 633422 63460 633428
rect 63132 625864 63184 625870
rect 63132 625806 63184 625812
rect 63144 618089 63172 625806
rect 63130 618080 63186 618089
rect 63130 618015 63186 618024
rect 62946 612096 63002 612105
rect 62946 612031 63002 612040
rect 62670 595776 62726 595785
rect 62670 595711 62726 595720
rect 62396 575476 62448 575482
rect 62396 575418 62448 575424
rect 62408 574841 62436 575418
rect 62394 574832 62450 574841
rect 62394 574767 62450 574776
rect 62396 574048 62448 574054
rect 62396 573990 62448 573996
rect 62408 573617 62436 573990
rect 62394 573608 62450 573617
rect 62394 573543 62450 573552
rect 62684 573458 62712 595711
rect 63130 594144 63186 594153
rect 63130 594079 63186 594088
rect 62946 590744 63002 590753
rect 62946 590679 63002 590688
rect 62960 590594 62988 590679
rect 62960 590566 63080 590594
rect 62854 590064 62910 590073
rect 62854 589999 62910 590008
rect 62868 589914 62896 589999
rect 62408 573430 62712 573458
rect 62776 589886 62896 589914
rect 62408 571169 62436 573430
rect 62776 573322 62804 589886
rect 63052 582374 63080 590566
rect 62592 573294 62804 573322
rect 62868 582346 63080 582374
rect 62394 571160 62450 571169
rect 62394 571095 62450 571104
rect 62592 569945 62620 573294
rect 62578 569936 62634 569945
rect 62578 569871 62634 569880
rect 62210 556744 62266 556753
rect 62210 556679 62266 556688
rect 62224 538214 62252 556679
rect 62670 550216 62726 550225
rect 62670 550151 62726 550160
rect 62684 547874 62712 550151
rect 62684 547846 62804 547874
rect 62224 538186 62528 538214
rect 62304 531276 62356 531282
rect 62304 531218 62356 531224
rect 62118 531176 62174 531185
rect 62118 531111 62120 531120
rect 62172 531111 62174 531120
rect 62120 531082 62172 531088
rect 62316 530641 62344 531218
rect 62302 530632 62358 530641
rect 62302 530567 62358 530576
rect 62120 528624 62172 528630
rect 62118 528592 62120 528601
rect 62172 528592 62174 528601
rect 62118 528527 62174 528536
rect 62500 528057 62528 538186
rect 62776 528554 62804 547846
rect 62684 528526 62804 528554
rect 62486 528048 62542 528057
rect 62486 527983 62542 527992
rect 62120 527128 62172 527134
rect 62118 527096 62120 527105
rect 62172 527096 62174 527105
rect 62118 527031 62174 527040
rect 62684 525745 62712 528526
rect 62670 525736 62726 525745
rect 62670 525671 62726 525680
rect 62394 422920 62450 422929
rect 62394 422855 62450 422864
rect 62120 404320 62172 404326
rect 62120 404262 62172 404268
rect 62132 404161 62160 404262
rect 62118 404152 62174 404161
rect 62118 404087 62174 404096
rect 62120 402960 62172 402966
rect 62120 402902 62172 402908
rect 62132 402665 62160 402902
rect 62118 402656 62174 402665
rect 62118 402591 62174 402600
rect 62118 400616 62174 400625
rect 62118 400551 62174 400560
rect 62132 400246 62160 400551
rect 62120 400240 62172 400246
rect 62408 400217 62436 422855
rect 62120 400182 62172 400188
rect 62394 400208 62450 400217
rect 62394 400143 62450 400152
rect 62120 400104 62172 400110
rect 62120 400046 62172 400052
rect 62132 399401 62160 400046
rect 62118 399392 62174 399401
rect 62118 399327 62174 399336
rect 62120 398812 62172 398818
rect 62120 398754 62172 398760
rect 62132 398313 62160 398754
rect 62118 398304 62174 398313
rect 62118 398239 62174 398248
rect 62210 385928 62266 385937
rect 62210 385863 62266 385872
rect 62224 364334 62252 385863
rect 62670 381848 62726 381857
rect 62670 381783 62726 381792
rect 62684 373994 62712 381783
rect 62684 373966 62804 373994
rect 62224 364306 62344 364334
rect 62120 361548 62172 361554
rect 62120 361490 62172 361496
rect 62132 360913 62160 361490
rect 62118 360904 62174 360913
rect 62118 360839 62174 360848
rect 62120 360188 62172 360194
rect 62120 360130 62172 360136
rect 62132 359825 62160 360130
rect 62118 359816 62174 359825
rect 62118 359751 62174 359760
rect 62118 357776 62174 357785
rect 62118 357711 62174 357720
rect 62132 357474 62160 357711
rect 62120 357468 62172 357474
rect 62120 357410 62172 357416
rect 62316 357377 62344 364306
rect 62302 357368 62358 357377
rect 62302 357303 62358 357312
rect 62120 356040 62172 356046
rect 62118 356008 62120 356017
rect 62172 356008 62174 356017
rect 62118 355943 62174 355952
rect 62776 354674 62804 373966
rect 62684 354646 62804 354674
rect 62684 354521 62712 354646
rect 62670 354512 62726 354521
rect 62670 354447 62726 354456
rect 62304 342236 62356 342242
rect 62304 342178 62356 342184
rect 62120 317416 62172 317422
rect 62118 317384 62120 317393
rect 62172 317384 62174 317393
rect 62118 317319 62174 317328
rect 62118 316024 62174 316033
rect 62118 315959 62120 315968
rect 62172 315959 62174 315968
rect 62120 315930 62172 315936
rect 62118 314800 62174 314809
rect 62118 314735 62120 314744
rect 62172 314735 62174 314744
rect 62120 314706 62172 314712
rect 62316 314129 62344 342178
rect 62670 341728 62726 341737
rect 62670 341663 62726 341672
rect 62486 341456 62542 341465
rect 62486 341391 62542 341400
rect 62302 314120 62358 314129
rect 62302 314055 62358 314064
rect 62500 313041 62528 341391
rect 62486 313032 62542 313041
rect 62486 312967 62542 312976
rect 62684 311817 62712 341663
rect 62670 311808 62726 311817
rect 62670 311743 62726 311752
rect 60002 300928 60058 300937
rect 60002 300863 60058 300872
rect 60016 291174 60044 300863
rect 62670 298752 62726 298761
rect 62670 298687 62726 298696
rect 61566 295352 61622 295361
rect 61566 295287 61622 295296
rect 60004 291168 60056 291174
rect 60004 291110 60056 291116
rect 58808 289808 58860 289814
rect 58808 289750 58860 289756
rect 58820 278458 58848 289750
rect 60004 288516 60056 288522
rect 60004 288458 60056 288464
rect 58808 278452 58860 278458
rect 58808 278394 58860 278400
rect 58624 231124 58676 231130
rect 58624 231066 58676 231072
rect 57244 228404 57296 228410
rect 57244 228346 57296 228352
rect 56508 227044 56560 227050
rect 56508 226986 56560 226992
rect 56520 218210 56548 226986
rect 55680 218204 55732 218210
rect 55680 218146 55732 218152
rect 56508 218204 56560 218210
rect 56508 218146 56560 218152
rect 55692 217138 55720 218146
rect 57256 218074 57284 228346
rect 58992 225616 59044 225622
rect 58992 225558 59044 225564
rect 57428 218204 57480 218210
rect 57428 218146 57480 218152
rect 56508 218068 56560 218074
rect 56508 218010 56560 218016
rect 57244 218068 57296 218074
rect 57244 218010 57296 218016
rect 56520 217138 56548 218010
rect 57440 217274 57468 218146
rect 58164 218068 58216 218074
rect 58164 218010 58216 218016
rect 55646 217110 55720 217138
rect 56474 217110 56548 217138
rect 57302 217246 57468 217274
rect 55646 216988 55674 217110
rect 56474 216988 56502 217110
rect 57302 216988 57330 217246
rect 58176 217138 58204 218010
rect 59004 217274 59032 225558
rect 60016 223553 60044 288458
rect 61382 280392 61438 280401
rect 61382 280327 61438 280336
rect 60648 227452 60700 227458
rect 60648 227394 60700 227400
rect 60002 223544 60058 223553
rect 60002 223479 60058 223488
rect 59360 221468 59412 221474
rect 59360 221410 59412 221416
rect 59372 218074 59400 221410
rect 59820 218748 59872 218754
rect 59820 218690 59872 218696
rect 59360 218068 59412 218074
rect 59360 218010 59412 218016
rect 58130 217110 58204 217138
rect 58958 217246 59032 217274
rect 58130 216988 58158 217110
rect 58958 216988 58986 217246
rect 59832 217138 59860 218690
rect 60660 217274 60688 227394
rect 61396 219434 61424 280327
rect 61580 278769 61608 295287
rect 62210 294264 62266 294273
rect 62210 294199 62266 294208
rect 62224 294030 62252 294199
rect 62212 294024 62264 294030
rect 62212 293966 62264 293972
rect 62302 292768 62358 292777
rect 62302 292703 62358 292712
rect 62316 292602 62344 292703
rect 62304 292596 62356 292602
rect 62304 292538 62356 292544
rect 62118 292496 62174 292505
rect 62118 292431 62120 292440
rect 62172 292431 62174 292440
rect 62120 292402 62172 292408
rect 62304 291168 62356 291174
rect 62304 291110 62356 291116
rect 62316 291009 62344 291110
rect 62302 291000 62358 291009
rect 62302 290935 62358 290944
rect 62684 289785 62712 298687
rect 62670 289776 62726 289785
rect 62670 289711 62726 289720
rect 62118 288552 62174 288561
rect 62118 288487 62120 288496
rect 62172 288487 62174 288496
rect 62120 288458 62172 288464
rect 62394 287192 62450 287201
rect 62394 287127 62450 287136
rect 62118 285968 62174 285977
rect 62118 285903 62174 285912
rect 62132 285734 62160 285903
rect 62120 285728 62172 285734
rect 62120 285670 62172 285676
rect 62210 282160 62266 282169
rect 62210 282095 62266 282104
rect 62224 281514 62252 282095
rect 62224 281486 62344 281514
rect 62118 280936 62174 280945
rect 62118 280871 62174 280880
rect 62132 280226 62160 280871
rect 62120 280220 62172 280226
rect 62120 280162 62172 280168
rect 61566 278760 61622 278769
rect 61566 278695 61622 278704
rect 62316 277394 62344 281486
rect 62224 277366 62344 277394
rect 62224 237969 62252 277366
rect 62408 267073 62436 287127
rect 62868 287054 62896 582346
rect 63144 568585 63172 594079
rect 63130 568576 63186 568585
rect 63130 568511 63186 568520
rect 63222 332616 63278 332625
rect 63222 332551 63278 332560
rect 62776 287026 62896 287054
rect 62776 283878 62804 287026
rect 62946 284608 63002 284617
rect 62946 284543 63002 284552
rect 62960 284374 62988 284543
rect 62948 284368 63000 284374
rect 62948 284310 63000 284316
rect 62776 283850 62896 283878
rect 62670 283248 62726 283257
rect 62670 283183 62726 283192
rect 62394 267064 62450 267073
rect 62394 266999 62450 267008
rect 62210 237960 62266 237969
rect 62210 237895 62266 237904
rect 61660 228540 61712 228546
rect 61660 228482 61712 228488
rect 61304 219406 61424 219434
rect 61304 217977 61332 219406
rect 61672 218210 61700 228482
rect 62028 225208 62080 225214
rect 62028 225150 62080 225156
rect 61660 218204 61712 218210
rect 61660 218146 61712 218152
rect 62040 218074 62068 225150
rect 62304 219020 62356 219026
rect 62304 218962 62356 218968
rect 61476 218068 61528 218074
rect 61476 218010 61528 218016
rect 62028 218068 62080 218074
rect 62028 218010 62080 218016
rect 61290 217968 61346 217977
rect 61290 217903 61346 217912
rect 59786 217110 59860 217138
rect 60614 217246 60688 217274
rect 59786 216988 59814 217110
rect 60614 216988 60642 217246
rect 61488 217138 61516 218010
rect 62316 217138 62344 218962
rect 62684 218890 62712 283183
rect 62868 278594 62896 283850
rect 62856 278588 62908 278594
rect 62856 278530 62908 278536
rect 63236 278186 63264 332551
rect 63420 278769 63448 633422
rect 63406 278760 63462 278769
rect 63406 278695 63462 278704
rect 63224 278180 63276 278186
rect 63224 278122 63276 278128
rect 64156 231266 64184 805938
rect 653404 790832 653456 790838
rect 653404 790774 653456 790780
rect 651470 778424 651526 778433
rect 651470 778359 651526 778368
rect 651484 777646 651512 778359
rect 651472 777640 651524 777646
rect 651472 777582 651524 777588
rect 652022 777064 652078 777073
rect 652022 776999 652078 777008
rect 651470 776112 651526 776121
rect 651470 776047 651526 776056
rect 651484 775606 651512 776047
rect 651472 775600 651524 775606
rect 651472 775542 651524 775548
rect 651380 775328 651432 775334
rect 651378 775296 651380 775305
rect 651432 775296 651434 775305
rect 651378 775231 651434 775240
rect 651470 774208 651526 774217
rect 651470 774143 651472 774152
rect 651524 774143 651526 774152
rect 651472 774114 651524 774120
rect 651472 773832 651524 773838
rect 651472 773774 651524 773780
rect 651484 773401 651512 773774
rect 651470 773392 651526 773401
rect 651470 773327 651526 773336
rect 652036 736234 652064 776999
rect 653416 775334 653444 790774
rect 670608 789404 670660 789410
rect 670608 789346 670660 789352
rect 655520 781108 655572 781114
rect 655520 781050 655572 781056
rect 655060 778388 655112 778394
rect 655060 778330 655112 778336
rect 653404 775328 653456 775334
rect 653404 775270 653456 775276
rect 655072 773838 655100 778330
rect 655532 774178 655560 781050
rect 660304 777640 660356 777646
rect 660304 777582 660356 777588
rect 655520 774172 655572 774178
rect 655520 774114 655572 774120
rect 655060 773832 655112 773838
rect 655060 773774 655112 773780
rect 652024 736228 652076 736234
rect 652024 736170 652076 736176
rect 653404 736228 653456 736234
rect 653404 736170 653456 736176
rect 651470 734224 651526 734233
rect 651470 734159 651526 734168
rect 651484 733446 651512 734159
rect 651472 733440 651524 733446
rect 651472 733382 651524 733388
rect 651470 733000 651526 733009
rect 651470 732935 651526 732944
rect 651484 732834 651512 732935
rect 651472 732828 651524 732834
rect 651472 732770 651524 732776
rect 651470 731776 651526 731785
rect 651470 731711 651526 731720
rect 651484 731474 651512 731711
rect 651472 731468 651524 731474
rect 651472 731410 651524 731416
rect 651472 731332 651524 731338
rect 651472 731274 651524 731280
rect 651484 731105 651512 731274
rect 651470 731096 651526 731105
rect 651470 731031 651526 731040
rect 651472 730040 651524 730046
rect 651472 729982 651524 729988
rect 651484 729881 651512 729982
rect 651470 729872 651526 729881
rect 651470 729807 651526 729816
rect 651472 728544 651524 728550
rect 651470 728512 651472 728521
rect 651524 728512 651526 728521
rect 651470 728447 651526 728456
rect 653416 716310 653444 736170
rect 657544 735616 657596 735622
rect 657544 735558 657596 735564
rect 654784 734188 654836 734194
rect 654784 734130 654836 734136
rect 654796 728550 654824 734130
rect 657556 730046 657584 735558
rect 658924 731468 658976 731474
rect 658924 731410 658976 731416
rect 657544 730040 657596 730046
rect 657544 729982 657596 729988
rect 654784 728544 654836 728550
rect 654784 728486 654836 728492
rect 653404 716304 653456 716310
rect 653404 716246 653456 716252
rect 654784 701208 654836 701214
rect 654784 701150 654836 701156
rect 651470 689480 651526 689489
rect 651470 689415 651526 689424
rect 651484 688702 651512 689415
rect 652760 688832 652812 688838
rect 651654 688800 651710 688809
rect 652760 688774 652812 688780
rect 651654 688735 651710 688744
rect 651472 688696 651524 688702
rect 651472 688638 651524 688644
rect 651470 687440 651526 687449
rect 651470 687375 651526 687384
rect 651484 687274 651512 687375
rect 651472 687268 651524 687274
rect 651472 687210 651524 687216
rect 651472 687064 651524 687070
rect 651472 687006 651524 687012
rect 651484 686769 651512 687006
rect 651470 686760 651526 686769
rect 651470 686695 651526 686704
rect 651668 686526 651696 688735
rect 651656 686520 651708 686526
rect 651656 686462 651708 686468
rect 651472 685568 651524 685574
rect 651472 685510 651524 685516
rect 651484 685273 651512 685510
rect 651470 685264 651526 685273
rect 651470 685199 651526 685208
rect 652574 684448 652630 684457
rect 652772 684434 652800 688774
rect 654796 687070 654824 701150
rect 656808 690056 656860 690062
rect 656808 689998 656860 690004
rect 654784 687064 654836 687070
rect 654784 687006 654836 687012
rect 656820 685574 656848 689998
rect 657544 688696 657596 688702
rect 657544 688638 657596 688644
rect 656808 685568 656860 685574
rect 656808 685510 656860 685516
rect 652630 684406 652800 684434
rect 652574 684383 652630 684392
rect 653404 655580 653456 655586
rect 653404 655522 653456 655528
rect 651470 643240 651526 643249
rect 651470 643175 651526 643184
rect 651484 642394 651512 643175
rect 651472 642388 651524 642394
rect 651472 642330 651524 642336
rect 652022 641880 652078 641889
rect 652022 641815 652078 641824
rect 651470 640792 651526 640801
rect 651470 640727 651526 640736
rect 651484 640354 651512 640727
rect 651472 640348 651524 640354
rect 651472 640290 651524 640296
rect 651380 640144 651432 640150
rect 651378 640112 651380 640121
rect 651432 640112 651434 640121
rect 651378 640047 651434 640056
rect 651656 638920 651708 638926
rect 651656 638862 651708 638868
rect 651472 638784 651524 638790
rect 651472 638726 651524 638732
rect 651484 638625 651512 638726
rect 651470 638616 651526 638625
rect 651470 638551 651526 638560
rect 651668 638217 651696 638862
rect 651654 638208 651710 638217
rect 651654 638143 651710 638152
rect 651470 597952 651526 597961
rect 651470 597887 651526 597896
rect 651484 597582 651512 597887
rect 651472 597576 651524 597582
rect 651472 597518 651524 597524
rect 651470 596728 651526 596737
rect 651470 596663 651526 596672
rect 651484 596222 651512 596663
rect 651472 596216 651524 596222
rect 651472 596158 651524 596164
rect 651656 595536 651708 595542
rect 651656 595478 651708 595484
rect 651470 595368 651526 595377
rect 651470 595303 651526 595312
rect 651484 594862 651512 595303
rect 651668 595105 651696 595478
rect 651654 595096 651710 595105
rect 651654 595031 651710 595040
rect 651472 594856 651524 594862
rect 651472 594798 651524 594804
rect 651472 594720 651524 594726
rect 651472 594662 651524 594668
rect 651484 594153 651512 594662
rect 651470 594144 651526 594153
rect 651470 594079 651526 594088
rect 651472 593088 651524 593094
rect 651472 593030 651524 593036
rect 651484 592793 651512 593030
rect 651470 592784 651526 592793
rect 651470 592719 651526 592728
rect 652036 581058 652064 641815
rect 653416 640150 653444 655522
rect 655520 645924 655572 645930
rect 655520 645866 655572 645872
rect 655336 643136 655388 643142
rect 655336 643078 655388 643084
rect 653404 640144 653456 640150
rect 653404 640086 653456 640092
rect 655348 638926 655376 643078
rect 655336 638920 655388 638926
rect 655336 638862 655388 638868
rect 655532 638790 655560 645866
rect 655520 638784 655572 638790
rect 655520 638726 655572 638732
rect 657556 625326 657584 688638
rect 658936 669526 658964 731410
rect 660316 715018 660344 777582
rect 669778 775840 669834 775849
rect 669778 775775 669834 775784
rect 668398 775024 668454 775033
rect 668398 774959 668454 774968
rect 668032 733440 668084 733446
rect 668032 733382 668084 733388
rect 661684 732828 661736 732834
rect 661684 732770 661736 732776
rect 660304 715012 660356 715018
rect 660304 714954 660356 714960
rect 661696 670750 661724 732770
rect 667848 703860 667900 703866
rect 667848 703802 667900 703808
rect 666468 701072 666520 701078
rect 666468 701014 666520 701020
rect 661684 670744 661736 670750
rect 661684 670686 661736 670692
rect 658924 669520 658976 669526
rect 658924 669462 658976 669468
rect 660304 642388 660356 642394
rect 660304 642330 660356 642336
rect 657544 625320 657596 625326
rect 657544 625262 657596 625268
rect 653404 611380 653456 611386
rect 653404 611322 653456 611328
rect 653416 595542 653444 611322
rect 657544 600364 657596 600370
rect 657544 600306 657596 600312
rect 654784 599004 654836 599010
rect 654784 598946 654836 598952
rect 653404 595536 653456 595542
rect 653404 595478 653456 595484
rect 654796 593094 654824 598946
rect 657556 594726 657584 600306
rect 658924 594856 658976 594862
rect 658924 594798 658976 594804
rect 657544 594720 657596 594726
rect 657544 594662 657596 594668
rect 654784 593088 654836 593094
rect 654784 593030 654836 593036
rect 652024 581052 652076 581058
rect 652024 580994 652076 581000
rect 653404 565888 653456 565894
rect 653404 565830 653456 565836
rect 651470 553480 651526 553489
rect 651470 553415 651526 553424
rect 651484 552702 651512 553415
rect 651472 552696 651524 552702
rect 651472 552638 651524 552644
rect 652022 552120 652078 552129
rect 652022 552055 652078 552064
rect 651470 551168 651526 551177
rect 651470 551103 651526 551112
rect 651484 550662 651512 551103
rect 651472 550656 651524 550662
rect 651472 550598 651524 550604
rect 651380 550384 651432 550390
rect 651378 550352 651380 550361
rect 651432 550352 651434 550361
rect 651378 550287 651434 550296
rect 651470 549264 651526 549273
rect 651470 549199 651472 549208
rect 651524 549199 651526 549208
rect 651472 549170 651524 549176
rect 651472 548888 651524 548894
rect 651472 548830 651524 548836
rect 651484 548457 651512 548830
rect 651470 548448 651526 548457
rect 651470 548383 651526 548392
rect 652036 493338 652064 552055
rect 653416 550390 653444 565830
rect 657820 554804 657872 554810
rect 657820 554746 657872 554752
rect 655152 553444 655204 553450
rect 655152 553386 655204 553392
rect 653404 550384 653456 550390
rect 653404 550326 653456 550332
rect 655164 548894 655192 553386
rect 657832 549234 657860 554746
rect 657820 549228 657872 549234
rect 657820 549170 657872 549176
rect 655152 548888 655204 548894
rect 655152 548830 655204 548836
rect 658936 534138 658964 594798
rect 660316 579698 660344 642330
rect 666480 621178 666508 701014
rect 667204 686520 667256 686526
rect 667204 686462 667256 686468
rect 667020 647352 667072 647358
rect 667020 647294 667072 647300
rect 666468 621172 666520 621178
rect 666468 621114 666520 621120
rect 661684 596216 661736 596222
rect 661684 596158 661736 596164
rect 660304 579692 660356 579698
rect 660304 579634 660356 579640
rect 661696 535498 661724 596158
rect 667032 574122 667060 647294
rect 667216 625666 667244 686462
rect 667662 639840 667718 639849
rect 667662 639775 667718 639784
rect 667204 625660 667256 625666
rect 667204 625602 667256 625608
rect 667388 597576 667440 597582
rect 667388 597518 667440 597524
rect 667020 574116 667072 574122
rect 667020 574058 667072 574064
rect 667204 570580 667256 570586
rect 667204 570522 667256 570528
rect 667018 562184 667074 562193
rect 667018 562119 667074 562128
rect 665824 552696 665876 552702
rect 665824 552638 665876 552644
rect 661684 535492 661736 535498
rect 661684 535434 661736 535440
rect 658924 534132 658976 534138
rect 658924 534074 658976 534080
rect 652208 520940 652260 520946
rect 652208 520882 652260 520888
rect 652024 493332 652076 493338
rect 652024 493274 652076 493280
rect 652220 476134 652248 520882
rect 665836 491366 665864 552638
rect 665824 491360 665876 491366
rect 665824 491302 665876 491308
rect 667032 484430 667060 562119
rect 667020 484424 667072 484430
rect 667020 484366 667072 484372
rect 658924 480956 658976 480962
rect 658924 480898 658976 480904
rect 650644 476128 650696 476134
rect 650644 476070 650696 476076
rect 652208 476128 652260 476134
rect 652208 476070 652260 476076
rect 649264 291916 649316 291922
rect 649264 291858 649316 291864
rect 649276 278322 649304 291858
rect 650656 278458 650684 476070
rect 658936 466478 658964 480898
rect 656164 466472 656216 466478
rect 656164 466414 656216 466420
rect 658924 466472 658976 466478
rect 658924 466414 658976 466420
rect 656176 458454 656204 466414
rect 651380 458448 651432 458454
rect 651380 458390 651432 458396
rect 656164 458448 656216 458454
rect 656164 458390 656216 458396
rect 651392 454578 651420 458390
rect 650828 454572 650880 454578
rect 650828 454514 650880 454520
rect 651380 454572 651432 454578
rect 651380 454514 651432 454520
rect 650840 278730 650868 454514
rect 657542 403336 657598 403345
rect 657542 403271 657598 403280
rect 652022 400888 652078 400897
rect 652022 400823 652078 400832
rect 651472 373992 651524 373998
rect 651472 373934 651524 373940
rect 651484 373289 651512 373934
rect 651470 373280 651526 373289
rect 651470 373215 651526 373224
rect 652036 372201 652064 400823
rect 652206 396672 652262 396681
rect 652206 396607 652262 396616
rect 652220 373969 652248 396607
rect 654782 382936 654838 382945
rect 654782 382871 654838 382880
rect 652206 373960 652262 373969
rect 652206 373895 652262 373904
rect 652022 372192 652078 372201
rect 652022 372127 652078 372136
rect 654796 371006 654824 382871
rect 657556 373998 657584 403271
rect 657544 373992 657596 373998
rect 657544 373934 657596 373940
rect 651472 371000 651524 371006
rect 651472 370942 651524 370948
rect 654784 371000 654836 371006
rect 654784 370942 654836 370948
rect 651484 370705 651512 370942
rect 651470 370696 651526 370705
rect 651470 370631 651526 370640
rect 652022 356688 652078 356697
rect 652022 356623 652078 356632
rect 651472 328432 651524 328438
rect 651472 328374 651524 328380
rect 651484 328273 651512 328374
rect 651470 328264 651526 328273
rect 651470 328199 651526 328208
rect 652036 326913 652064 356623
rect 652390 351112 652446 351121
rect 652390 351047 652446 351056
rect 652404 329769 652432 351047
rect 660304 338768 660356 338774
rect 653402 338736 653458 338745
rect 660304 338710 660356 338716
rect 653402 338671 653458 338680
rect 652390 329760 652446 329769
rect 652390 329695 652446 329704
rect 652022 326904 652078 326913
rect 652022 326839 652078 326848
rect 651378 325680 651434 325689
rect 653416 325650 653444 338671
rect 651378 325615 651380 325624
rect 651432 325615 651434 325624
rect 653404 325644 653456 325650
rect 651380 325586 651432 325592
rect 653404 325586 653456 325592
rect 660316 313954 660344 338710
rect 652024 313948 652076 313954
rect 652024 313890 652076 313896
rect 660304 313948 660356 313954
rect 660304 313890 660356 313896
rect 651472 302184 651524 302190
rect 651472 302126 651524 302132
rect 651484 301889 651512 302126
rect 651470 301880 651526 301889
rect 651470 301815 651526 301824
rect 651472 300824 651524 300830
rect 651472 300766 651524 300772
rect 651484 300665 651512 300766
rect 651470 300656 651526 300665
rect 651470 300591 651526 300600
rect 651746 297528 651802 297537
rect 651802 297486 651972 297514
rect 651746 297463 651802 297472
rect 651746 296848 651802 296857
rect 651746 296783 651748 296792
rect 651800 296783 651802 296792
rect 651748 296754 651800 296760
rect 651944 296714 651972 297486
rect 651852 296686 651972 296714
rect 651654 295352 651710 295361
rect 651654 295287 651710 295296
rect 651470 294264 651526 294273
rect 651470 294199 651526 294208
rect 651484 294030 651512 294199
rect 651472 294024 651524 294030
rect 651472 293966 651524 293972
rect 651668 290465 651696 295287
rect 651470 290456 651526 290465
rect 651470 290391 651526 290400
rect 651654 290456 651710 290465
rect 651654 290391 651710 290400
rect 651484 289882 651512 290391
rect 651472 289876 651524 289882
rect 651472 289818 651524 289824
rect 651654 289232 651710 289241
rect 651654 289167 651710 289176
rect 651470 288688 651526 288697
rect 651470 288623 651526 288632
rect 651484 288454 651512 288623
rect 651472 288448 651524 288454
rect 651472 288390 651524 288396
rect 651668 287706 651696 289167
rect 651656 287700 651708 287706
rect 651656 287642 651708 287648
rect 651470 285968 651526 285977
rect 651470 285903 651526 285912
rect 651484 285734 651512 285903
rect 651472 285728 651524 285734
rect 651472 285670 651524 285676
rect 651470 284744 651526 284753
rect 651470 284679 651526 284688
rect 651484 284374 651512 284679
rect 651472 284368 651524 284374
rect 651472 284310 651524 284316
rect 651470 283520 651526 283529
rect 651470 283455 651526 283464
rect 651484 282946 651512 283455
rect 651472 282940 651524 282946
rect 651472 282882 651524 282888
rect 651470 282160 651526 282169
rect 651470 282095 651526 282104
rect 651484 281586 651512 282095
rect 651472 281580 651524 281586
rect 651472 281522 651524 281528
rect 651470 280936 651526 280945
rect 651470 280871 651526 280880
rect 651484 280226 651512 280871
rect 651472 280220 651524 280226
rect 651472 280162 651524 280168
rect 651852 279449 651880 296686
rect 652036 291922 652064 313890
rect 660302 311944 660358 311953
rect 660302 311879 660358 311888
rect 652206 311128 652262 311137
rect 652206 311063 652262 311072
rect 652220 303385 652248 311063
rect 652206 303376 652262 303385
rect 652206 303311 652262 303320
rect 660316 300830 660344 311879
rect 660304 300824 660356 300830
rect 660304 300766 660356 300772
rect 652574 298616 652630 298625
rect 652630 298574 652800 298602
rect 652574 298551 652630 298560
rect 652772 296714 652800 298574
rect 665824 296744 665876 296750
rect 652772 296686 652892 296714
rect 665824 296686 665876 296692
rect 652864 293865 652892 296686
rect 664444 294024 664496 294030
rect 664444 293966 664496 293972
rect 652850 293856 652906 293865
rect 652850 293791 652906 293800
rect 652390 292768 652446 292777
rect 652390 292703 652446 292712
rect 652024 291916 652076 291922
rect 652024 291858 652076 291864
rect 652206 291544 652262 291553
rect 652206 291479 652262 291488
rect 652022 287192 652078 287201
rect 652022 287127 652078 287136
rect 651838 279440 651894 279449
rect 651838 279375 651894 279384
rect 650828 278724 650880 278730
rect 650828 278666 650880 278672
rect 650644 278452 650696 278458
rect 650644 278394 650696 278400
rect 649264 278316 649316 278322
rect 649264 278258 649316 278264
rect 65904 272542 65932 278052
rect 67100 274242 67128 278052
rect 67088 274236 67140 274242
rect 67088 274178 67140 274184
rect 65892 272536 65944 272542
rect 65892 272478 65944 272484
rect 68204 271182 68232 278052
rect 69400 273970 69428 278052
rect 69388 273964 69440 273970
rect 69388 273906 69440 273912
rect 68192 271176 68244 271182
rect 68192 271118 68244 271124
rect 70596 269822 70624 278052
rect 71792 275330 71820 278052
rect 71780 275324 71832 275330
rect 71780 275266 71832 275272
rect 72988 272678 73016 278052
rect 74184 274718 74212 278052
rect 74172 274712 74224 274718
rect 74172 274654 74224 274660
rect 72976 272672 73028 272678
rect 72976 272614 73028 272620
rect 75380 271454 75408 278052
rect 76484 275602 76512 278052
rect 76472 275596 76524 275602
rect 76472 275538 76524 275544
rect 76840 274712 76892 274718
rect 76840 274654 76892 274660
rect 75368 271448 75420 271454
rect 75368 271390 75420 271396
rect 76852 271318 76880 274654
rect 77680 274106 77708 278052
rect 77668 274100 77720 274106
rect 77668 274042 77720 274048
rect 76840 271312 76892 271318
rect 76840 271254 76892 271260
rect 78876 270366 78904 278052
rect 78864 270360 78916 270366
rect 78864 270302 78916 270308
rect 80072 269822 80100 278052
rect 81268 275058 81296 278052
rect 81256 275052 81308 275058
rect 81256 274994 81308 275000
rect 82464 272814 82492 278052
rect 83674 278038 84148 278066
rect 84778 278038 85528 278066
rect 82452 272808 82504 272814
rect 82452 272750 82504 272756
rect 84120 270502 84148 278038
rect 84108 270496 84160 270502
rect 84108 270438 84160 270444
rect 85500 269958 85528 278038
rect 85960 274718 85988 278052
rect 86224 275596 86276 275602
rect 86224 275538 86276 275544
rect 85948 274712 86000 274718
rect 85948 274654 86000 274660
rect 85488 269952 85540 269958
rect 85488 269894 85540 269900
rect 70584 269816 70636 269822
rect 70584 269758 70636 269764
rect 79324 269816 79376 269822
rect 79324 269758 79376 269764
rect 80060 269816 80112 269822
rect 80060 269758 80112 269764
rect 79336 267170 79364 269758
rect 86236 267442 86264 275538
rect 87156 271590 87184 278052
rect 88352 273834 88380 278052
rect 89562 278038 89668 278066
rect 88340 273828 88392 273834
rect 88340 273770 88392 273776
rect 87144 271584 87196 271590
rect 87144 271526 87196 271532
rect 89640 270094 89668 278038
rect 90744 275602 90772 278052
rect 91862 278038 92428 278066
rect 90732 275596 90784 275602
rect 90732 275538 90784 275544
rect 90364 274712 90416 274718
rect 90364 274654 90416 274660
rect 89628 270088 89680 270094
rect 89628 270030 89680 270036
rect 86224 267436 86276 267442
rect 86224 267378 86276 267384
rect 79324 267164 79376 267170
rect 79324 267106 79376 267112
rect 90376 267034 90404 274654
rect 92400 268394 92428 278038
rect 93044 275738 93072 278052
rect 93032 275732 93084 275738
rect 93032 275674 93084 275680
rect 94240 272950 94268 278052
rect 95436 274378 95464 278052
rect 96632 275194 96660 278052
rect 96620 275188 96672 275194
rect 96620 275130 96672 275136
rect 95424 274372 95476 274378
rect 95424 274314 95476 274320
rect 94228 272944 94280 272950
rect 94228 272886 94280 272892
rect 97828 271726 97856 278052
rect 99038 278038 99328 278066
rect 97816 271720 97868 271726
rect 97816 271662 97868 271668
rect 99300 268530 99328 278038
rect 100128 275466 100156 278052
rect 100116 275460 100168 275466
rect 100116 275402 100168 275408
rect 101324 274514 101352 278052
rect 101312 274508 101364 274514
rect 101312 274450 101364 274456
rect 102520 273086 102548 278052
rect 103716 274718 103744 278052
rect 104912 277394 104940 278052
rect 104912 277366 105032 277394
rect 103704 274712 103756 274718
rect 103704 274654 103756 274660
rect 104808 274712 104860 274718
rect 104808 274654 104860 274660
rect 102508 273080 102560 273086
rect 102508 273022 102560 273028
rect 99288 268524 99340 268530
rect 99288 268466 99340 268472
rect 92388 268388 92440 268394
rect 92388 268330 92440 268336
rect 104820 267306 104848 274654
rect 105004 268666 105032 277366
rect 106016 271862 106044 278052
rect 107212 276010 107240 278052
rect 107200 276004 107252 276010
rect 107200 275946 107252 275952
rect 108408 273222 108436 278052
rect 109618 278038 110368 278066
rect 108396 273216 108448 273222
rect 108396 273158 108448 273164
rect 106004 271856 106056 271862
rect 106004 271798 106056 271804
rect 110340 268802 110368 278038
rect 110800 274718 110828 278052
rect 110788 274712 110840 274718
rect 110788 274654 110840 274660
rect 111708 274712 111760 274718
rect 111708 274654 111760 274660
rect 110328 268796 110380 268802
rect 110328 268738 110380 268744
rect 104992 268660 105044 268666
rect 104992 268602 105044 268608
rect 111720 267578 111748 274654
rect 111996 270230 112024 278052
rect 113206 278038 113496 278066
rect 113468 271046 113496 278038
rect 114388 274650 114416 278052
rect 115506 278038 115888 278066
rect 114376 274644 114428 274650
rect 114376 274586 114428 274592
rect 113456 271040 113508 271046
rect 113456 270982 113508 270988
rect 111984 270224 112036 270230
rect 111984 270166 112036 270172
rect 115860 268938 115888 278038
rect 116688 272406 116716 278052
rect 117898 278038 118648 278066
rect 116676 272400 116728 272406
rect 116676 272342 116728 272348
rect 118620 269074 118648 278038
rect 119080 273698 119108 278052
rect 120276 273834 120304 278052
rect 119344 273828 119396 273834
rect 119344 273770 119396 273776
rect 120264 273828 120316 273834
rect 120264 273770 120316 273776
rect 119068 273692 119120 273698
rect 119068 273634 119120 273640
rect 118608 269068 118660 269074
rect 118608 269010 118660 269016
rect 115848 268932 115900 268938
rect 115848 268874 115900 268880
rect 111708 267572 111760 267578
rect 111708 267514 111760 267520
rect 104808 267300 104860 267306
rect 104808 267242 104860 267248
rect 90364 267028 90416 267034
rect 90364 266970 90416 266976
rect 119356 266898 119384 273770
rect 121472 270638 121500 278052
rect 122590 278038 122788 278066
rect 121460 270632 121512 270638
rect 121460 270574 121512 270580
rect 122760 269686 122788 278038
rect 123772 270910 123800 278052
rect 124968 271998 124996 278052
rect 126178 278038 126928 278066
rect 124956 271992 125008 271998
rect 124956 271934 125008 271940
rect 123760 270904 123812 270910
rect 123760 270846 123812 270852
rect 122748 269680 122800 269686
rect 122748 269622 122800 269628
rect 126900 269414 126928 278038
rect 127360 272270 127388 278052
rect 128556 274786 128584 278052
rect 128544 274780 128596 274786
rect 128544 274722 128596 274728
rect 127348 272264 127400 272270
rect 127348 272206 127400 272212
rect 129660 269550 129688 278052
rect 130856 274242 130884 278052
rect 130384 274236 130436 274242
rect 130384 274178 130436 274184
rect 130844 274236 130896 274242
rect 130844 274178 130896 274184
rect 129648 269544 129700 269550
rect 129648 269486 129700 269492
rect 126888 269408 126940 269414
rect 126888 269350 126940 269356
rect 130396 267714 130424 274178
rect 132052 273562 132080 278052
rect 133262 278038 133828 278066
rect 132040 273556 132092 273562
rect 132040 273498 132092 273504
rect 133800 270366 133828 278038
rect 134444 270774 134472 278052
rect 134432 270768 134484 270774
rect 134432 270710 134484 270716
rect 132500 270360 132552 270366
rect 132500 270302 132552 270308
rect 133788 270360 133840 270366
rect 133788 270302 133840 270308
rect 130384 267708 130436 267714
rect 130384 267650 130436 267656
rect 119344 266892 119396 266898
rect 119344 266834 119396 266840
rect 132512 266626 132540 270302
rect 135640 267850 135668 278052
rect 136836 274922 136864 278052
rect 136824 274916 136876 274922
rect 136824 274858 136876 274864
rect 137652 274916 137704 274922
rect 137652 274858 137704 274864
rect 136824 272536 136876 272542
rect 136824 272478 136876 272484
rect 135628 267844 135680 267850
rect 135628 267786 135680 267792
rect 132500 266620 132552 266626
rect 132500 266562 132552 266568
rect 136836 264330 136864 272478
rect 137664 270502 137692 274858
rect 137940 272542 137968 278052
rect 139136 275874 139164 278052
rect 140346 278038 140728 278066
rect 139124 275868 139176 275874
rect 139124 275810 139176 275816
rect 139400 273964 139452 273970
rect 139400 273906 139452 273912
rect 137928 272536 137980 272542
rect 137928 272478 137980 272484
rect 138480 271176 138532 271182
rect 138480 271118 138532 271124
rect 137468 270496 137520 270502
rect 137468 270438 137520 270444
rect 137652 270496 137704 270502
rect 137652 270438 137704 270444
rect 137480 266762 137508 270438
rect 138112 267708 138164 267714
rect 138112 267650 138164 267656
rect 137468 266756 137520 266762
rect 137468 266698 137520 266704
rect 136836 264302 137310 264330
rect 138124 264316 138152 267650
rect 138492 264330 138520 271118
rect 139412 264330 139440 273906
rect 140700 268258 140728 278038
rect 141056 275324 141108 275330
rect 141056 275266 141108 275272
rect 140688 268252 140740 268258
rect 140688 268194 140740 268200
rect 140596 267164 140648 267170
rect 140596 267106 140648 267112
rect 138492 264302 138966 264330
rect 139412 264302 139794 264330
rect 140608 264316 140636 267106
rect 141068 264330 141096 275266
rect 141528 271182 141556 278052
rect 142724 272678 142752 278052
rect 142160 272672 142212 272678
rect 142160 272614 142212 272620
rect 142712 272672 142764 272678
rect 142712 272614 142764 272620
rect 141516 271176 141568 271182
rect 141516 271118 141568 271124
rect 142172 264330 142200 272614
rect 142712 271448 142764 271454
rect 142712 271390 142764 271396
rect 142724 264330 142752 271390
rect 143540 271312 143592 271318
rect 143540 271254 143592 271260
rect 143552 264330 143580 271254
rect 143920 269278 143948 278052
rect 144920 274100 144972 274106
rect 144920 274042 144972 274048
rect 143908 269272 143960 269278
rect 143908 269214 143960 269220
rect 144932 267734 144960 274042
rect 145116 272134 145144 278052
rect 145288 275052 145340 275058
rect 145288 274994 145340 275000
rect 145300 273426 145328 274994
rect 146220 274922 146248 278052
rect 146208 274916 146260 274922
rect 146208 274858 146260 274864
rect 145288 273420 145340 273426
rect 145288 273362 145340 273368
rect 147416 272678 147444 278052
rect 148612 273970 148640 278052
rect 149808 275058 149836 278052
rect 151018 278038 151768 278066
rect 149980 275188 150032 275194
rect 149980 275130 150032 275136
rect 149796 275052 149848 275058
rect 149796 274994 149848 275000
rect 148600 273964 148652 273970
rect 148600 273906 148652 273912
rect 147864 273420 147916 273426
rect 147864 273362 147916 273368
rect 145564 272672 145616 272678
rect 145564 272614 145616 272620
rect 147404 272672 147456 272678
rect 147404 272614 147456 272620
rect 145104 272128 145156 272134
rect 145104 272070 145156 272076
rect 144932 267706 145144 267734
rect 144736 267436 144788 267442
rect 144736 267378 144788 267384
rect 141068 264302 141450 264330
rect 142172 264302 142278 264330
rect 142724 264302 143106 264330
rect 143552 264302 143934 264330
rect 144748 264316 144776 267378
rect 145116 264330 145144 267706
rect 145576 267170 145604 272614
rect 146392 269816 146444 269822
rect 146392 269758 146444 269764
rect 145564 267164 145616 267170
rect 145564 267106 145616 267112
rect 145116 264302 145590 264330
rect 146404 264316 146432 269758
rect 147220 266620 147272 266626
rect 147220 266562 147272 266568
rect 147232 264316 147260 266562
rect 147876 264330 147904 273362
rect 148416 272808 148468 272814
rect 148416 272750 148468 272756
rect 148428 264330 148456 272750
rect 149704 269952 149756 269958
rect 149704 269894 149756 269900
rect 147876 264302 148074 264330
rect 148428 264302 148902 264330
rect 149716 264316 149744 269894
rect 149992 266626 150020 275130
rect 151084 271992 151136 271998
rect 151084 271934 151136 271940
rect 151096 266762 151124 271934
rect 151740 268122 151768 278038
rect 152004 271584 152056 271590
rect 152004 271526 152056 271532
rect 151728 268116 151780 268122
rect 151728 268058 151780 268064
rect 151360 267028 151412 267034
rect 151360 266970 151412 266976
rect 150532 266756 150584 266762
rect 150532 266698 150584 266704
rect 151084 266756 151136 266762
rect 151084 266698 151136 266704
rect 149980 266620 150032 266626
rect 149980 266562 150032 266568
rect 150544 264316 150572 266698
rect 151372 264316 151400 266970
rect 152016 264330 152044 271526
rect 152200 271318 152228 278052
rect 152832 275732 152884 275738
rect 152832 275674 152884 275680
rect 152188 271312 152240 271318
rect 152188 271254 152240 271260
rect 152844 269958 152872 275674
rect 153396 275194 153424 278052
rect 153384 275188 153436 275194
rect 153384 275130 153436 275136
rect 154500 274106 154528 278052
rect 154764 275596 154816 275602
rect 154764 275538 154816 275544
rect 154488 274100 154540 274106
rect 154488 274042 154540 274048
rect 153844 273556 153896 273562
rect 153844 273498 153896 273504
rect 153016 270088 153068 270094
rect 153016 270030 153068 270036
rect 152832 269952 152884 269958
rect 152832 269894 152884 269900
rect 152016 264302 152214 264330
rect 153028 264316 153056 270030
rect 153856 267442 153884 273498
rect 154776 267734 154804 275538
rect 155696 272814 155724 278052
rect 156892 275466 156920 278052
rect 158102 278038 158668 278066
rect 156880 275460 156932 275466
rect 156880 275402 156932 275408
rect 157616 274372 157668 274378
rect 157616 274314 157668 274320
rect 155960 272944 156012 272950
rect 155960 272886 156012 272892
rect 155684 272808 155736 272814
rect 155684 272750 155736 272756
rect 155500 268388 155552 268394
rect 155500 268330 155552 268336
rect 154684 267706 154804 267734
rect 153844 267436 153896 267442
rect 153844 267378 153896 267384
rect 153844 266892 153896 266898
rect 153844 266834 153896 266840
rect 153856 264316 153884 266834
rect 154684 264316 154712 267706
rect 155512 264316 155540 268330
rect 155972 264330 156000 272886
rect 157156 269952 157208 269958
rect 157156 269894 157208 269900
rect 155972 264302 156354 264330
rect 157168 264316 157196 269894
rect 157628 264330 157656 274314
rect 158640 269822 158668 278038
rect 159284 274378 159312 278052
rect 160480 275738 160508 278052
rect 160468 275732 160520 275738
rect 160468 275674 160520 275680
rect 159456 275324 159508 275330
rect 159456 275266 159508 275272
rect 159272 274372 159324 274378
rect 159272 274314 159324 274320
rect 158812 271720 158864 271726
rect 158812 271662 158864 271668
rect 158628 269816 158680 269822
rect 158628 269758 158680 269764
rect 157628 264302 158010 264330
rect 158824 264316 158852 271662
rect 159468 267034 159496 275266
rect 160928 274508 160980 274514
rect 160928 274450 160980 274456
rect 160468 268524 160520 268530
rect 160468 268466 160520 268472
rect 159456 267028 159508 267034
rect 159456 266970 159508 266976
rect 159640 266620 159692 266626
rect 159640 266562 159692 266568
rect 159652 264316 159680 266562
rect 160480 264316 160508 268466
rect 160940 264330 160968 274450
rect 161584 268394 161612 278052
rect 162780 277394 162808 278052
rect 162688 277366 162808 277394
rect 162688 271454 162716 277366
rect 163504 276004 163556 276010
rect 163504 275946 163556 275952
rect 162860 273080 162912 273086
rect 162860 273022 162912 273028
rect 162676 271448 162728 271454
rect 162676 271390 162728 271396
rect 161572 268388 161624 268394
rect 161572 268330 161624 268336
rect 162124 267028 162176 267034
rect 162124 266970 162176 266976
rect 160940 264302 161322 264330
rect 162136 264316 162164 266970
rect 162872 264330 162900 273022
rect 163516 266422 163544 275946
rect 163976 275466 164004 278052
rect 163964 275460 164016 275466
rect 163964 275402 164016 275408
rect 164976 271856 165028 271862
rect 164976 271798 165028 271804
rect 163780 268660 163832 268666
rect 163780 268602 163832 268608
rect 163504 266416 163556 266422
rect 163504 266358 163556 266364
rect 162872 264302 162978 264330
rect 163792 264316 163820 268602
rect 164608 267300 164660 267306
rect 164608 267242 164660 267248
rect 164620 264316 164648 267242
rect 164988 264330 165016 271798
rect 165172 271590 165200 278052
rect 165896 273216 165948 273222
rect 165896 273158 165948 273164
rect 165160 271584 165212 271590
rect 165160 271526 165212 271532
rect 165908 264330 165936 273158
rect 166368 272950 166396 278052
rect 167564 276010 167592 278052
rect 167552 276004 167604 276010
rect 167552 275946 167604 275952
rect 167000 274780 167052 274786
rect 167000 274722 167052 274728
rect 166356 272944 166408 272950
rect 166356 272886 166408 272892
rect 167012 268802 167040 274722
rect 168760 274514 168788 278052
rect 169024 275188 169076 275194
rect 169024 275130 169076 275136
rect 168748 274508 168800 274514
rect 168748 274450 168800 274456
rect 168104 270632 168156 270638
rect 168104 270574 168156 270580
rect 167000 268796 167052 268802
rect 167000 268738 167052 268744
rect 167920 268524 167972 268530
rect 167920 268466 167972 268472
rect 167092 266416 167144 266422
rect 167092 266358 167144 266364
rect 164988 264302 165462 264330
rect 165908 264302 166290 264330
rect 167104 264316 167132 266358
rect 167932 264316 167960 268466
rect 168116 267034 168144 270574
rect 168748 270224 168800 270230
rect 168748 270166 168800 270172
rect 168104 267028 168156 267034
rect 168104 266970 168156 266976
rect 168760 264316 168788 270166
rect 169036 266898 169064 275130
rect 169864 271726 169892 278052
rect 171060 275602 171088 278052
rect 171048 275596 171100 275602
rect 171048 275538 171100 275544
rect 171600 274644 171652 274650
rect 171600 274586 171652 274592
rect 169852 271720 169904 271726
rect 169852 271662 169904 271668
rect 169944 271040 169996 271046
rect 169944 270982 169996 270988
rect 169576 267572 169628 267578
rect 169576 267514 169628 267520
rect 169024 266892 169076 266898
rect 169024 266834 169076 266840
rect 169588 264316 169616 267514
rect 169956 264330 169984 270982
rect 171232 268660 171284 268666
rect 171232 268602 171284 268608
rect 169956 264302 170430 264330
rect 171244 264316 171272 268602
rect 171612 264330 171640 274586
rect 172256 273086 172284 278052
rect 173466 278038 173848 278066
rect 174662 278038 175136 278066
rect 175858 278038 176608 278066
rect 173256 273692 173308 273698
rect 173256 273634 173308 273640
rect 172244 273080 172296 273086
rect 172244 273022 172296 273028
rect 172520 272400 172572 272406
rect 172520 272342 172572 272348
rect 172532 264330 172560 272342
rect 173268 264330 173296 273634
rect 173820 269958 173848 278038
rect 174268 275868 174320 275874
rect 174268 275810 174320 275816
rect 174280 271862 174308 275810
rect 174268 271856 174320 271862
rect 174268 271798 174320 271804
rect 173808 269952 173860 269958
rect 173808 269894 173860 269900
rect 175108 269074 175136 278038
rect 175280 273828 175332 273834
rect 175280 273770 175332 273776
rect 174544 269068 174596 269074
rect 174544 269010 174596 269016
rect 175096 269068 175148 269074
rect 175096 269010 175148 269016
rect 171612 264302 172086 264330
rect 172532 264302 172914 264330
rect 173268 264302 173742 264330
rect 174556 264316 174584 269010
rect 175292 264330 175320 273770
rect 176580 270094 176608 278038
rect 176568 270088 176620 270094
rect 176568 270030 176620 270036
rect 176200 269680 176252 269686
rect 176200 269622 176252 269628
rect 175292 264302 175398 264330
rect 176212 264316 176240 269622
rect 176948 268666 176976 278052
rect 178144 275874 178172 278052
rect 178684 276004 178736 276010
rect 178684 275946 178736 275952
rect 178132 275868 178184 275874
rect 178132 275810 178184 275816
rect 177488 270904 177540 270910
rect 177488 270846 177540 270852
rect 176936 268660 176988 268666
rect 176936 268602 176988 268608
rect 177028 267028 177080 267034
rect 177028 266970 177080 266976
rect 177040 264316 177068 266970
rect 177500 264330 177528 270846
rect 178316 269408 178368 269414
rect 178316 269350 178368 269356
rect 177672 269068 177724 269074
rect 177672 269010 177724 269016
rect 177684 267034 177712 269010
rect 177672 267028 177724 267034
rect 177672 266970 177724 266976
rect 178328 264330 178356 269350
rect 178696 267578 178724 275946
rect 179340 274650 179368 278052
rect 180536 277394 180564 278052
rect 180536 277366 180656 277394
rect 179328 274644 179380 274650
rect 179328 274586 179380 274592
rect 179880 272264 179932 272270
rect 179880 272206 179932 272212
rect 178684 267572 178736 267578
rect 178684 267514 178736 267520
rect 179512 266756 179564 266762
rect 179512 266698 179564 266704
rect 177500 264302 177882 264330
rect 178328 264302 178710 264330
rect 179524 264316 179552 266698
rect 179892 264330 179920 272206
rect 180628 268530 180656 277366
rect 181732 272542 181760 278052
rect 182942 278038 183508 278066
rect 184138 278038 184888 278066
rect 182456 274236 182508 274242
rect 182456 274178 182508 274184
rect 181720 272536 181772 272542
rect 181720 272478 181772 272484
rect 181168 269544 181220 269550
rect 181168 269486 181220 269492
rect 180616 268524 180668 268530
rect 180616 268466 180668 268472
rect 179892 264302 180366 264330
rect 181180 264316 181208 269486
rect 181996 268796 182048 268802
rect 181996 268738 182048 268744
rect 182008 264316 182036 268738
rect 182468 264330 182496 274178
rect 183480 269686 183508 278038
rect 183652 270360 183704 270366
rect 183652 270302 183704 270308
rect 183468 269680 183520 269686
rect 183468 269622 183520 269628
rect 182468 264302 182850 264330
rect 183664 264316 183692 270302
rect 184860 270230 184888 278038
rect 185228 276010 185256 278052
rect 185216 276004 185268 276010
rect 185216 275946 185268 275952
rect 185308 274916 185360 274922
rect 185308 274858 185360 274864
rect 185124 270768 185176 270774
rect 185124 270710 185176 270716
rect 184848 270224 184900 270230
rect 184848 270166 184900 270172
rect 184480 267436 184532 267442
rect 184480 267378 184532 267384
rect 184492 264316 184520 267378
rect 185136 264330 185164 270710
rect 185320 270366 185348 274858
rect 186424 273222 186452 278052
rect 187436 278038 187634 278066
rect 186412 273216 186464 273222
rect 186412 273158 186464 273164
rect 187148 272536 187200 272542
rect 187148 272478 187200 272484
rect 186136 270496 186188 270502
rect 186136 270438 186188 270444
rect 185308 270360 185360 270366
rect 185308 270302 185360 270308
rect 185136 264302 185334 264330
rect 186148 264316 186176 270438
rect 187160 267714 187188 272478
rect 187436 271046 187464 278038
rect 188816 277394 188844 278052
rect 188816 277366 188936 277394
rect 187700 272400 187752 272406
rect 187700 272342 187752 272348
rect 187424 271040 187476 271046
rect 187424 270982 187476 270988
rect 186964 267708 187016 267714
rect 186964 267650 187016 267656
rect 187148 267708 187200 267714
rect 187148 267650 187200 267656
rect 186976 264316 187004 267650
rect 187712 264330 187740 272342
rect 188908 268938 188936 277366
rect 190012 275194 190040 278052
rect 190000 275188 190052 275194
rect 190000 275130 190052 275136
rect 189080 275052 189132 275058
rect 189080 274994 189132 275000
rect 189092 272542 189120 274994
rect 189080 272536 189132 272542
rect 189080 272478 189132 272484
rect 189264 271856 189316 271862
rect 189264 271798 189316 271804
rect 189080 271176 189132 271182
rect 189080 271118 189132 271124
rect 188896 268932 188948 268938
rect 188896 268874 188948 268880
rect 188620 268252 188672 268258
rect 188620 268194 188672 268200
rect 187712 264302 187818 264330
rect 188632 264316 188660 268194
rect 189092 265674 189120 271118
rect 189080 265668 189132 265674
rect 189080 265610 189132 265616
rect 189276 264330 189304 271798
rect 191208 271182 191236 278052
rect 192404 273834 192432 278052
rect 193508 274242 193536 278052
rect 194718 278038 195008 278066
rect 193496 274236 193548 274242
rect 193496 274178 193548 274184
rect 194784 273964 194836 273970
rect 194784 273906 194836 273912
rect 192392 273828 192444 273834
rect 192392 273770 192444 273776
rect 193220 272672 193272 272678
rect 193220 272614 193272 272620
rect 192392 272128 192444 272134
rect 192392 272070 192444 272076
rect 191196 271176 191248 271182
rect 191196 271118 191248 271124
rect 191104 269272 191156 269278
rect 191104 269214 191156 269220
rect 190552 268932 190604 268938
rect 190552 268874 190604 268880
rect 190564 267442 190592 268874
rect 190552 267436 190604 267442
rect 190552 267378 190604 267384
rect 189908 265668 189960 265674
rect 189908 265610 189960 265616
rect 189920 264330 189948 265610
rect 189276 264302 189474 264330
rect 189920 264302 190302 264330
rect 191116 264316 191144 269214
rect 191932 267300 191984 267306
rect 191932 267242 191984 267248
rect 191944 264316 191972 267242
rect 192404 264330 192432 272070
rect 193232 264330 193260 272614
rect 194416 270360 194468 270366
rect 194416 270302 194468 270308
rect 192404 264302 192786 264330
rect 193232 264302 193614 264330
rect 194428 264316 194456 270302
rect 194796 264330 194824 273906
rect 194980 272406 195008 278038
rect 195900 272678 195928 278052
rect 195888 272672 195940 272678
rect 195888 272614 195940 272620
rect 197096 272542 197124 278052
rect 198096 274100 198148 274106
rect 198096 274042 198148 274048
rect 196440 272536 196492 272542
rect 196440 272478 196492 272484
rect 197084 272536 197136 272542
rect 197084 272478 197136 272484
rect 194968 272400 195020 272406
rect 194968 272342 195020 272348
rect 196072 268116 196124 268122
rect 196072 268058 196124 268064
rect 195244 267708 195296 267714
rect 195244 267650 195296 267656
rect 195256 267442 195284 267650
rect 195244 267436 195296 267442
rect 195244 267378 195296 267384
rect 194796 264302 195270 264330
rect 196084 264316 196112 268058
rect 196452 264330 196480 272478
rect 197360 271312 197412 271318
rect 197360 271254 197412 271260
rect 197372 264330 197400 271254
rect 198108 264330 198136 274042
rect 198292 271318 198320 278052
rect 199502 278038 199976 278066
rect 199384 275732 199436 275738
rect 199384 275674 199436 275680
rect 198280 271312 198332 271318
rect 198280 271254 198332 271260
rect 199396 267170 199424 275674
rect 199948 270366 199976 278038
rect 200120 272808 200172 272814
rect 200120 272750 200172 272756
rect 199936 270360 199988 270366
rect 199936 270302 199988 270308
rect 199384 267164 199436 267170
rect 199384 267106 199436 267112
rect 199384 266892 199436 266898
rect 199384 266834 199436 266840
rect 196452 264302 196926 264330
rect 197372 264302 197754 264330
rect 198108 264302 198582 264330
rect 199396 264316 199424 266834
rect 200132 264330 200160 272750
rect 200592 268802 200620 278052
rect 201788 277394 201816 278052
rect 201696 277366 201816 277394
rect 200764 275324 200816 275330
rect 200764 275266 200816 275272
rect 200776 270502 200804 275266
rect 200764 270496 200816 270502
rect 200764 270438 200816 270444
rect 201696 269822 201724 277366
rect 202328 274372 202380 274378
rect 202328 274314 202380 274320
rect 201868 270496 201920 270502
rect 201868 270438 201920 270444
rect 201040 269816 201092 269822
rect 201040 269758 201092 269764
rect 201684 269816 201736 269822
rect 201684 269758 201736 269764
rect 200580 268796 200632 268802
rect 200580 268738 200632 268744
rect 200132 264302 200238 264330
rect 201052 264316 201080 269758
rect 201880 264316 201908 270438
rect 202340 264330 202368 274314
rect 202984 271862 203012 278052
rect 202972 271856 203024 271862
rect 202972 271798 203024 271804
rect 204180 269550 204208 278052
rect 205376 272814 205404 278052
rect 206586 278038 206876 278066
rect 206376 275460 206428 275466
rect 206376 275402 206428 275408
rect 205364 272808 205416 272814
rect 205364 272750 205416 272756
rect 205640 271584 205692 271590
rect 205640 271526 205692 271532
rect 204720 271448 204772 271454
rect 204720 271390 204772 271396
rect 204168 269544 204220 269550
rect 204168 269486 204220 269492
rect 203524 268388 203576 268394
rect 203524 268330 203576 268336
rect 202340 264302 202722 264330
rect 203536 264316 203564 268330
rect 204352 267164 204404 267170
rect 204352 267106 204404 267112
rect 204364 264316 204392 267106
rect 204732 264330 204760 271390
rect 205456 269680 205508 269686
rect 205456 269622 205508 269628
rect 205468 267170 205496 269622
rect 205456 267164 205508 267170
rect 205456 267106 205508 267112
rect 205652 264330 205680 271526
rect 206388 264330 206416 275402
rect 206848 270502 206876 278038
rect 207768 274786 207796 278052
rect 207756 274780 207808 274786
rect 207756 274722 207808 274728
rect 208400 274508 208452 274514
rect 208400 274450 208452 274456
rect 207296 272944 207348 272950
rect 207296 272886 207348 272892
rect 206836 270496 206888 270502
rect 206836 270438 206888 270444
rect 207308 264330 207336 272886
rect 208412 264330 208440 274450
rect 208872 273970 208900 278052
rect 210068 274106 210096 278052
rect 210700 274780 210752 274786
rect 210700 274722 210752 274728
rect 210056 274100 210108 274106
rect 210056 274042 210108 274048
rect 208860 273964 208912 273970
rect 208860 273906 208912 273912
rect 209780 273080 209832 273086
rect 209780 273022 209832 273028
rect 209320 267572 209372 267578
rect 209320 267514 209372 267520
rect 204732 264302 205206 264330
rect 205652 264302 206034 264330
rect 206388 264302 206862 264330
rect 207308 264302 207690 264330
rect 208412 264302 208518 264330
rect 209332 264316 209360 267514
rect 209792 265674 209820 273022
rect 209964 271720 210016 271726
rect 209964 271662 210016 271668
rect 209780 265668 209832 265674
rect 209780 265610 209832 265616
rect 209976 264330 210004 271662
rect 210712 268394 210740 274722
rect 211264 272950 211292 278052
rect 211436 275596 211488 275602
rect 211436 275538 211488 275544
rect 211252 272944 211304 272950
rect 211252 272886 211304 272892
rect 211160 270088 211212 270094
rect 211160 270030 211212 270036
rect 210700 268388 210752 268394
rect 210700 268330 210752 268336
rect 211172 266422 211200 270030
rect 211160 266416 211212 266422
rect 211160 266358 211212 266364
rect 210700 265668 210752 265674
rect 210700 265610 210752 265616
rect 210712 264330 210740 265610
rect 211448 264330 211476 275538
rect 212460 270094 212488 278052
rect 213656 271454 213684 278052
rect 214852 275330 214880 278052
rect 214840 275324 214892 275330
rect 214840 275266 214892 275272
rect 214564 274644 214616 274650
rect 214564 274586 214616 274592
rect 213644 271448 213696 271454
rect 213644 271390 213696 271396
rect 212448 270088 212500 270094
rect 212448 270030 212500 270036
rect 212632 269952 212684 269958
rect 212632 269894 212684 269900
rect 209976 264302 210174 264330
rect 210712 264302 211002 264330
rect 211448 264302 211830 264330
rect 212644 264316 212672 269894
rect 214288 267028 214340 267034
rect 214288 266970 214340 266976
rect 213460 266416 213512 266422
rect 213460 266358 213512 266364
rect 213472 264316 213500 266358
rect 214300 264316 214328 266970
rect 214576 266422 214604 274586
rect 215956 271590 215984 278052
rect 216680 275868 216732 275874
rect 216680 275810 216732 275816
rect 215944 271584 215996 271590
rect 215944 271526 215996 271532
rect 216128 271040 216180 271046
rect 216128 270982 216180 270988
rect 215116 268660 215168 268666
rect 215116 268602 215168 268608
rect 214564 266416 214616 266422
rect 214564 266358 214616 266364
rect 215128 264316 215156 268602
rect 216140 266898 216168 270982
rect 216128 266892 216180 266898
rect 216128 266834 216180 266840
rect 215944 266416 215996 266422
rect 215944 266358 215996 266364
rect 215956 264316 215984 266358
rect 216692 264330 216720 275810
rect 217152 275738 217180 278052
rect 217140 275732 217192 275738
rect 217140 275674 217192 275680
rect 218348 275602 218376 278052
rect 218336 275596 218388 275602
rect 218336 275538 218388 275544
rect 218704 273216 218756 273222
rect 218704 273158 218756 273164
rect 217600 268524 217652 268530
rect 217600 268466 217652 268472
rect 216692 264302 216798 264330
rect 217612 264316 217640 268466
rect 218428 267164 218480 267170
rect 218428 267106 218480 267112
rect 218440 264316 218468 267106
rect 218716 267034 218744 273158
rect 219544 273086 219572 278052
rect 219532 273080 219584 273086
rect 219532 273022 219584 273028
rect 220740 272950 220768 278052
rect 221280 276004 221332 276010
rect 221280 275946 221332 275952
rect 220084 272944 220136 272950
rect 220084 272886 220136 272892
rect 220728 272944 220780 272950
rect 220728 272886 220780 272892
rect 219348 270224 219400 270230
rect 219348 270166 219400 270172
rect 219360 267594 219388 270166
rect 219360 267566 219664 267594
rect 219256 267436 219308 267442
rect 219256 267378 219308 267384
rect 218704 267028 218756 267034
rect 218704 266970 218756 266976
rect 219268 264316 219296 267378
rect 219636 264330 219664 267566
rect 220096 267170 220124 272886
rect 220084 267164 220136 267170
rect 220084 267106 220136 267112
rect 220912 267028 220964 267034
rect 220912 266970 220964 266976
rect 219636 264302 220110 264330
rect 220924 264316 220952 266970
rect 221292 264330 221320 275946
rect 221936 275466 221964 278052
rect 221924 275460 221976 275466
rect 221924 275402 221976 275408
rect 222936 275188 222988 275194
rect 222936 275130 222988 275136
rect 222568 266892 222620 266898
rect 222568 266834 222620 266840
rect 221292 264302 221766 264330
rect 222580 264316 222608 266834
rect 222948 264330 222976 275130
rect 223132 274378 223160 278052
rect 224236 275874 224264 278052
rect 224224 275868 224276 275874
rect 224224 275810 224276 275816
rect 224224 275732 224276 275738
rect 224224 275674 224276 275680
rect 223120 274372 223172 274378
rect 223120 274314 223172 274320
rect 223488 269544 223540 269550
rect 223488 269486 223540 269492
rect 223500 267442 223528 269486
rect 224236 268666 224264 275674
rect 224960 273828 225012 273834
rect 224960 273770 225012 273776
rect 224224 268660 224276 268666
rect 224224 268602 224276 268608
rect 223488 267436 223540 267442
rect 223488 267378 223540 267384
rect 224224 267300 224276 267306
rect 224224 267242 224276 267248
rect 222948 264302 223422 264330
rect 224236 264316 224264 267242
rect 224972 265674 225000 273770
rect 225432 271726 225460 278052
rect 226432 274236 226484 274242
rect 226432 274178 226484 274184
rect 225420 271720 225472 271726
rect 225420 271662 225472 271668
rect 225144 271176 225196 271182
rect 225144 271118 225196 271124
rect 224960 265668 225012 265674
rect 224960 265610 225012 265616
rect 225156 265554 225184 271118
rect 225604 265668 225656 265674
rect 225604 265610 225656 265616
rect 225064 265526 225184 265554
rect 225064 264316 225092 265526
rect 225616 264330 225644 265610
rect 226444 264330 226472 274178
rect 226628 269958 226656 278052
rect 227838 278038 228128 278066
rect 228100 272678 228128 278038
rect 229020 275738 229048 278052
rect 229008 275732 229060 275738
rect 229008 275674 229060 275680
rect 227904 272672 227956 272678
rect 227904 272614 227956 272620
rect 228088 272672 228140 272678
rect 228088 272614 228140 272620
rect 227168 272400 227220 272406
rect 227168 272342 227220 272348
rect 226616 269952 226668 269958
rect 226616 269894 226668 269900
rect 227180 264330 227208 272342
rect 227916 264330 227944 272614
rect 229100 272536 229152 272542
rect 229100 272478 229152 272484
rect 228364 271720 228416 271726
rect 228364 271662 228416 271668
rect 228376 267034 228404 271662
rect 228364 267028 228416 267034
rect 228364 266970 228416 266976
rect 229112 264330 229140 272478
rect 229560 271312 229612 271318
rect 229560 271254 229612 271260
rect 229572 264330 229600 271254
rect 230216 271182 230244 278052
rect 231334 278038 231716 278066
rect 230204 271176 230256 271182
rect 230204 271118 230256 271124
rect 230848 270360 230900 270366
rect 230848 270302 230900 270308
rect 225616 264302 225906 264330
rect 226444 264302 226734 264330
rect 227180 264302 227562 264330
rect 227916 264302 228390 264330
rect 229112 264302 229218 264330
rect 229572 264302 230046 264330
rect 230860 264316 230888 270302
rect 231308 268796 231360 268802
rect 231308 268738 231360 268744
rect 231320 264330 231348 268738
rect 231688 268530 231716 278038
rect 232516 275194 232544 278052
rect 233056 275868 233108 275874
rect 233056 275810 233108 275816
rect 232504 275188 232556 275194
rect 232504 275130 232556 275136
rect 233068 270366 233096 275810
rect 233712 272542 233740 278052
rect 234922 278038 235304 278066
rect 233884 275596 233936 275602
rect 233884 275538 233936 275544
rect 233700 272536 233752 272542
rect 233700 272478 233752 272484
rect 233240 271856 233292 271862
rect 233240 271798 233292 271804
rect 233056 270360 233108 270366
rect 233056 270302 233108 270308
rect 232504 269816 232556 269822
rect 232504 269758 232556 269764
rect 231676 268524 231728 268530
rect 231676 268466 231728 268472
rect 231320 264302 231702 264330
rect 232516 264316 232544 269758
rect 233252 264330 233280 271798
rect 233896 267306 233924 275538
rect 234804 272808 234856 272814
rect 234804 272750 234856 272756
rect 234160 267436 234212 267442
rect 234160 267378 234212 267384
rect 233884 267300 233936 267306
rect 233884 267242 233936 267248
rect 233252 264302 233358 264330
rect 234172 264316 234200 267378
rect 234816 264330 234844 272750
rect 235276 271318 235304 278038
rect 236104 275874 236132 278052
rect 236092 275868 236144 275874
rect 236092 275810 236144 275816
rect 235264 271312 235316 271318
rect 235264 271254 235316 271260
rect 235816 270496 235868 270502
rect 235816 270438 235868 270444
rect 234816 264302 235014 264330
rect 235828 264316 235856 270438
rect 237208 269822 237236 278052
rect 237840 274100 237892 274106
rect 237840 274042 237892 274048
rect 237380 273964 237432 273970
rect 237380 273906 237432 273912
rect 237196 269816 237248 269822
rect 237196 269758 237248 269764
rect 236644 268388 236696 268394
rect 236644 268330 236696 268336
rect 236656 264316 236684 268330
rect 237392 264330 237420 273906
rect 237852 264330 237880 274042
rect 238496 273970 238524 278052
rect 239600 275602 239628 278052
rect 239588 275596 239640 275602
rect 239588 275538 239640 275544
rect 239404 275324 239456 275330
rect 239404 275266 239456 275272
rect 238484 273964 238536 273970
rect 238484 273906 238536 273912
rect 239128 267164 239180 267170
rect 239128 267106 239180 267112
rect 237392 264302 237498 264330
rect 237852 264302 238326 264330
rect 239140 264316 239168 267106
rect 239416 266422 239444 275266
rect 240048 275188 240100 275194
rect 240048 275130 240100 275136
rect 240060 274242 240088 275130
rect 240048 274236 240100 274242
rect 240048 274178 240100 274184
rect 240796 271454 240824 278052
rect 241992 277394 242020 278052
rect 241900 277366 242020 277394
rect 240416 271448 240468 271454
rect 240416 271390 240468 271396
rect 240784 271448 240836 271454
rect 240784 271390 240836 271396
rect 239956 270088 240008 270094
rect 239956 270030 240008 270036
rect 239404 266416 239456 266422
rect 239404 266358 239456 266364
rect 239968 264316 239996 270030
rect 240428 264330 240456 271390
rect 241900 270094 241928 277366
rect 243188 275330 243216 278052
rect 243728 275732 243780 275738
rect 243728 275674 243780 275680
rect 243544 275460 243596 275466
rect 243544 275402 243596 275408
rect 243176 275324 243228 275330
rect 243176 275266 243228 275272
rect 242072 271584 242124 271590
rect 242072 271526 242124 271532
rect 241888 270088 241940 270094
rect 241888 270030 241940 270036
rect 241612 266416 241664 266422
rect 241612 266358 241664 266364
rect 240428 264302 240810 264330
rect 241624 264316 241652 266358
rect 242084 264330 242112 271526
rect 243268 268660 243320 268666
rect 243268 268602 243320 268608
rect 242084 264302 242466 264330
rect 243280 264316 243308 268602
rect 243556 266422 243584 275402
rect 243740 267442 243768 275674
rect 244384 270230 244412 278052
rect 245396 278038 245502 278066
rect 246790 278038 246988 278066
rect 244556 273080 244608 273086
rect 244556 273022 244608 273028
rect 244372 270224 244424 270230
rect 244372 270166 244424 270172
rect 243728 267436 243780 267442
rect 243728 267378 243780 267384
rect 244096 267300 244148 267306
rect 244096 267242 244148 267248
rect 243544 266416 243596 266422
rect 243544 266358 243596 266364
rect 244108 264316 244136 267242
rect 244568 264330 244596 273022
rect 245396 272814 245424 278038
rect 245752 272944 245804 272950
rect 245752 272886 245804 272892
rect 245384 272808 245436 272814
rect 245384 272750 245436 272756
rect 244568 264302 244950 264330
rect 245764 264316 245792 272886
rect 246960 267170 246988 278038
rect 247224 274372 247276 274378
rect 247224 274314 247276 274320
rect 246948 267164 247000 267170
rect 246948 267106 247000 267112
rect 246580 266416 246632 266422
rect 246580 266358 246632 266364
rect 246592 264316 246620 266358
rect 247236 264330 247264 274314
rect 247880 272950 247908 278052
rect 249076 274106 249104 278052
rect 250272 275738 250300 278052
rect 250444 275868 250496 275874
rect 250444 275810 250496 275816
rect 250260 275732 250312 275738
rect 250260 275674 250312 275680
rect 249064 274100 249116 274106
rect 249064 274042 249116 274048
rect 247868 272944 247920 272950
rect 247868 272886 247920 272892
rect 249064 272672 249116 272678
rect 249064 272614 249116 272620
rect 248236 270360 248288 270366
rect 248236 270302 248288 270308
rect 247236 264302 247434 264330
rect 248248 264316 248276 270302
rect 249076 267306 249104 272614
rect 249892 269952 249944 269958
rect 249892 269894 249944 269900
rect 249064 267300 249116 267306
rect 249064 267242 249116 267248
rect 249064 267028 249116 267034
rect 249064 266970 249116 266976
rect 249076 264316 249104 266970
rect 249904 264316 249932 269894
rect 250456 266422 250484 275810
rect 251468 271046 251496 278052
rect 252008 271176 252060 271182
rect 252008 271118 252060 271124
rect 251456 271040 251508 271046
rect 251456 270982 251508 270988
rect 251548 267436 251600 267442
rect 251548 267378 251600 267384
rect 250720 267300 250772 267306
rect 250720 267242 250772 267248
rect 250444 266416 250496 266422
rect 250444 266358 250496 266364
rect 250732 264316 250760 267242
rect 251560 264316 251588 267378
rect 252020 264330 252048 271118
rect 252664 268394 252692 278052
rect 253860 274718 253888 278052
rect 253848 274712 253900 274718
rect 253848 274654 253900 274660
rect 253940 274236 253992 274242
rect 253940 274178 253992 274184
rect 253204 268524 253256 268530
rect 253204 268466 253256 268472
rect 252652 268388 252704 268394
rect 252652 268330 252704 268336
rect 252020 264302 252402 264330
rect 253216 264316 253244 268466
rect 253952 264330 253980 274178
rect 254964 272542 254992 278052
rect 255964 275596 256016 275602
rect 255964 275538 256016 275544
rect 254400 272536 254452 272542
rect 254400 272478 254452 272484
rect 254952 272536 255004 272542
rect 254952 272478 255004 272484
rect 254412 264330 254440 272478
rect 255320 271312 255372 271318
rect 255320 271254 255372 271260
rect 255332 264330 255360 271254
rect 255976 267034 256004 275538
rect 256160 275466 256188 278052
rect 257356 275602 257384 278052
rect 257344 275596 257396 275602
rect 257344 275538 257396 275544
rect 256148 275460 256200 275466
rect 256148 275402 256200 275408
rect 256700 275324 256752 275330
rect 256700 275266 256752 275272
rect 256712 271318 256740 275266
rect 256884 274712 256936 274718
rect 256884 274654 256936 274660
rect 256700 271312 256752 271318
rect 256700 271254 256752 271260
rect 256896 269958 256924 274654
rect 258080 273828 258132 273834
rect 258080 273770 258132 273776
rect 256884 269952 256936 269958
rect 256884 269894 256936 269900
rect 257344 269816 257396 269822
rect 257344 269758 257396 269764
rect 255964 267028 256016 267034
rect 255964 266970 256016 266976
rect 256516 266416 256568 266422
rect 256516 266358 256568 266364
rect 253952 264302 254058 264330
rect 254412 264302 254886 264330
rect 255332 264302 255714 264330
rect 256528 264316 256556 266358
rect 257356 264316 257384 269758
rect 258092 264330 258120 273770
rect 258552 269822 258580 278052
rect 259748 277394 259776 278052
rect 259748 277366 259868 277394
rect 259368 275732 259420 275738
rect 259368 275674 259420 275680
rect 259380 273562 259408 275674
rect 259368 273556 259420 273562
rect 259368 273498 259420 273504
rect 259840 271454 259868 277366
rect 260944 275806 260972 278052
rect 260932 275800 260984 275806
rect 260932 275742 260984 275748
rect 259644 271448 259696 271454
rect 259644 271390 259696 271396
rect 259828 271448 259880 271454
rect 259828 271390 259880 271396
rect 258540 269816 258592 269822
rect 258540 269758 258592 269764
rect 259000 267028 259052 267034
rect 259000 266970 259052 266976
rect 258092 264302 258198 264330
rect 259012 264316 259040 266970
rect 259656 264330 259684 271390
rect 262048 271318 262076 278052
rect 262312 275596 262364 275602
rect 262312 275538 262364 275544
rect 262324 272814 262352 275538
rect 263244 275330 263272 278052
rect 263232 275324 263284 275330
rect 263232 275266 263284 275272
rect 264244 272944 264296 272950
rect 264244 272886 264296 272892
rect 262312 272808 262364 272814
rect 262312 272750 262364 272756
rect 262680 272672 262732 272678
rect 262680 272614 262732 272620
rect 261024 271312 261076 271318
rect 261024 271254 261076 271260
rect 262036 271312 262088 271318
rect 262036 271254 262088 271260
rect 260656 270088 260708 270094
rect 260656 270030 260708 270036
rect 259656 264302 259854 264330
rect 260668 264316 260696 270030
rect 261036 264330 261064 271254
rect 262312 270224 262364 270230
rect 262312 270166 262364 270172
rect 261036 264302 261510 264330
rect 262324 264316 262352 270166
rect 262692 264330 262720 272614
rect 264256 267734 264284 272886
rect 264440 272678 264468 278052
rect 265650 278038 266216 278066
rect 265256 274100 265308 274106
rect 265256 274042 265308 274048
rect 264428 272672 264480 272678
rect 264428 272614 264480 272620
rect 264256 267706 264376 267734
rect 263968 267164 264020 267170
rect 263968 267106 264020 267112
rect 262692 264302 263166 264330
rect 263980 264316 264008 267106
rect 264348 264330 264376 267706
rect 265268 264330 265296 274042
rect 266188 270094 266216 278038
rect 266360 275800 266412 275806
rect 266360 275742 266412 275748
rect 266372 274106 266400 275742
rect 266832 275602 266860 278052
rect 266820 275596 266872 275602
rect 266820 275538 266872 275544
rect 266360 274100 266412 274106
rect 266360 274042 266412 274048
rect 266360 273556 266412 273562
rect 266360 273498 266412 273504
rect 266176 270088 266228 270094
rect 266176 270030 266228 270036
rect 266372 264330 266400 273498
rect 268028 271182 268056 278052
rect 269224 275126 269252 278052
rect 269396 275460 269448 275466
rect 269396 275402 269448 275408
rect 269212 275120 269264 275126
rect 269212 275062 269264 275068
rect 269408 272678 269436 275402
rect 269120 272672 269172 272678
rect 269120 272614 269172 272620
rect 269396 272672 269448 272678
rect 269396 272614 269448 272620
rect 269132 272406 269160 272614
rect 270328 272542 270356 278052
rect 271524 273970 271552 278052
rect 272734 278038 273116 278066
rect 271512 273964 271564 273970
rect 271512 273906 271564 273912
rect 270960 272808 271012 272814
rect 270960 272750 271012 272756
rect 270592 272672 270644 272678
rect 270592 272614 270644 272620
rect 269304 272536 269356 272542
rect 269304 272478 269356 272484
rect 270316 272536 270368 272542
rect 270316 272478 270368 272484
rect 269120 272400 269172 272406
rect 269120 272342 269172 272348
rect 268016 271176 268068 271182
rect 268016 271118 268068 271124
rect 266912 271040 266964 271046
rect 266912 270982 266964 270988
rect 266924 264330 266952 270982
rect 268936 269952 268988 269958
rect 268936 269894 268988 269900
rect 268108 268388 268160 268394
rect 268108 268330 268160 268336
rect 264348 264302 264822 264330
rect 265268 264302 265650 264330
rect 266372 264302 266478 264330
rect 266924 264302 267306 264330
rect 268120 264316 268148 268330
rect 268948 264316 268976 269894
rect 269316 264330 269344 272478
rect 269316 264302 269790 264330
rect 270604 264316 270632 272614
rect 270972 264330 271000 272750
rect 272616 271448 272668 271454
rect 272616 271390 272668 271396
rect 272248 269816 272300 269822
rect 272248 269758 272300 269764
rect 270972 264302 271446 264330
rect 272260 264316 272288 269758
rect 272628 264330 272656 271390
rect 273088 269822 273116 278038
rect 273260 275324 273312 275330
rect 273260 275266 273312 275272
rect 273076 269816 273128 269822
rect 273076 269758 273128 269764
rect 273272 269074 273300 275266
rect 273536 274100 273588 274106
rect 273536 274042 273588 274048
rect 273260 269068 273312 269074
rect 273260 269010 273312 269016
rect 273548 264330 273576 274042
rect 273916 272814 273944 278052
rect 274640 275120 274692 275126
rect 274640 275062 274692 275068
rect 273904 272808 273956 272814
rect 273904 272750 273956 272756
rect 274652 271862 274680 275062
rect 275112 274718 275140 278052
rect 276308 275330 276336 278052
rect 276480 275596 276532 275602
rect 276480 275538 276532 275544
rect 276296 275324 276348 275330
rect 276296 275266 276348 275272
rect 275100 274712 275152 274718
rect 275100 274654 275152 274660
rect 276020 272400 276072 272406
rect 276020 272342 276072 272348
rect 274640 271856 274692 271862
rect 274640 271798 274692 271804
rect 274640 271312 274692 271318
rect 274640 271254 274692 271260
rect 274652 264330 274680 271254
rect 275560 269068 275612 269074
rect 275560 269010 275612 269016
rect 272628 264302 273102 264330
rect 273548 264302 273930 264330
rect 274652 264302 274758 264330
rect 275572 264316 275600 269010
rect 276032 264330 276060 272342
rect 276492 267782 276520 275538
rect 277504 275534 277532 278052
rect 277492 275528 277544 275534
rect 277492 275470 277544 275476
rect 278412 274712 278464 274718
rect 278412 274654 278464 274660
rect 278424 270502 278452 274654
rect 278608 274106 278636 278052
rect 278596 274100 278648 274106
rect 278596 274042 278648 274048
rect 279240 271856 279292 271862
rect 279240 271798 279292 271804
rect 278872 271176 278924 271182
rect 278872 271118 278924 271124
rect 278412 270496 278464 270502
rect 278412 270438 278464 270444
rect 277216 270088 277268 270094
rect 277216 270030 277268 270036
rect 276480 267776 276532 267782
rect 276480 267718 276532 267724
rect 276032 264302 276414 264330
rect 277228 264316 277256 270030
rect 278044 267776 278096 267782
rect 278044 267718 278096 267724
rect 278056 264316 278084 267718
rect 278884 264316 278912 271118
rect 279252 264330 279280 271798
rect 279804 271182 279832 278052
rect 280344 273964 280396 273970
rect 280344 273906 280396 273912
rect 279792 271176 279844 271182
rect 279792 271118 279844 271124
rect 280356 265674 280384 273906
rect 281000 273086 281028 278052
rect 282210 278038 282776 278066
rect 280988 273080 281040 273086
rect 280988 273022 281040 273028
rect 280528 272536 280580 272542
rect 280528 272478 280580 272484
rect 280344 265668 280396 265674
rect 280344 265610 280396 265616
rect 279252 264302 279726 264330
rect 280540 264316 280568 272478
rect 282184 269816 282236 269822
rect 282184 269758 282236 269764
rect 280988 265668 281040 265674
rect 280988 265610 281040 265616
rect 281000 264330 281028 265610
rect 281000 264302 281382 264330
rect 282196 264316 282224 269758
rect 282748 269278 282776 278038
rect 283104 275324 283156 275330
rect 283104 275266 283156 275272
rect 282920 272808 282972 272814
rect 282920 272750 282972 272756
rect 282736 269272 282788 269278
rect 282736 269214 282788 269220
rect 282932 264330 282960 272750
rect 283116 270366 283144 275266
rect 283392 274718 283420 278052
rect 284588 275874 284616 278052
rect 284576 275868 284628 275874
rect 284576 275810 284628 275816
rect 285128 275528 285180 275534
rect 285128 275470 285180 275476
rect 283380 274712 283432 274718
rect 283380 274654 283432 274660
rect 283840 270496 283892 270502
rect 283840 270438 283892 270444
rect 283104 270360 283156 270366
rect 283104 270302 283156 270308
rect 282932 264302 283038 264330
rect 283852 264316 283880 270438
rect 284668 270360 284720 270366
rect 284668 270302 284720 270308
rect 284680 264316 284708 270302
rect 285140 264330 285168 275470
rect 285692 275466 285720 278052
rect 286888 275738 286916 278052
rect 286876 275732 286928 275738
rect 286876 275674 286928 275680
rect 285680 275460 285732 275466
rect 285680 275402 285732 275408
rect 288084 275058 288112 278052
rect 288072 275052 288124 275058
rect 288072 274994 288124 275000
rect 289280 274922 289308 278052
rect 290096 275868 290148 275874
rect 290096 275810 290148 275816
rect 289268 274916 289320 274922
rect 289268 274858 289320 274864
rect 289176 274712 289228 274718
rect 289176 274654 289228 274660
rect 285864 274100 285916 274106
rect 285864 274042 285916 274048
rect 285876 264330 285904 274042
rect 286324 273080 286376 273086
rect 286324 273022 286376 273028
rect 286336 267034 286364 273022
rect 287060 271176 287112 271182
rect 287060 271118 287112 271124
rect 286324 267028 286376 267034
rect 286324 266970 286376 266976
rect 287072 264330 287100 271118
rect 288808 269272 288860 269278
rect 288808 269214 288860 269220
rect 287980 267028 288032 267034
rect 287980 266970 288032 266976
rect 285140 264302 285522 264330
rect 285876 264302 286350 264330
rect 287072 264302 287178 264330
rect 287992 264316 288020 266970
rect 288820 264316 288848 269214
rect 289188 264330 289216 274654
rect 290108 264330 290136 275810
rect 290476 274718 290504 278052
rect 291200 275460 291252 275466
rect 291200 275402 291252 275408
rect 290464 274712 290516 274718
rect 290464 274654 290516 274660
rect 291212 264330 291240 275402
rect 291672 275330 291700 278052
rect 291844 275732 291896 275738
rect 291844 275674 291896 275680
rect 291660 275324 291712 275330
rect 291660 275266 291712 275272
rect 291856 264330 291884 275674
rect 292868 275194 292896 278052
rect 292856 275188 292908 275194
rect 292856 275130 292908 275136
rect 292856 275052 292908 275058
rect 292856 274994 292908 275000
rect 292672 274916 292724 274922
rect 292672 274858 292724 274864
rect 292684 265674 292712 274858
rect 292672 265668 292724 265674
rect 292672 265610 292724 265616
rect 292868 264330 292896 274994
rect 293972 274990 294000 278052
rect 293960 274984 294012 274990
rect 293960 274926 294012 274932
rect 295168 274718 295196 278052
rect 295340 275324 295392 275330
rect 295340 275266 295392 275272
rect 294144 274712 294196 274718
rect 294144 274654 294196 274660
rect 295156 274712 295208 274718
rect 295156 274654 295208 274660
rect 293500 265668 293552 265674
rect 293500 265610 293552 265616
rect 293512 264330 293540 265610
rect 294156 264330 294184 274654
rect 295352 264330 295380 275266
rect 295800 275188 295852 275194
rect 295800 275130 295852 275136
rect 295812 264330 295840 275130
rect 296364 274854 296392 278052
rect 297180 274984 297232 274990
rect 297180 274926 297232 274932
rect 296352 274848 296404 274854
rect 296352 274790 296404 274796
rect 296812 274712 296864 274718
rect 296812 274654 296864 274660
rect 296824 265674 296852 274654
rect 297192 267734 297220 274926
rect 297560 274718 297588 278052
rect 298756 275262 298784 278052
rect 299952 275398 299980 278052
rect 300964 278038 301070 278066
rect 302266 278038 302464 278066
rect 299940 275392 299992 275398
rect 299940 275334 299992 275340
rect 298744 275256 298796 275262
rect 298744 275198 298796 275204
rect 300032 275256 300084 275262
rect 300032 275198 300084 275204
rect 298376 274848 298428 274854
rect 298376 274790 298428 274796
rect 297548 274712 297600 274718
rect 297548 274654 297600 274660
rect 297100 267706 297220 267734
rect 296812 265668 296864 265674
rect 296812 265610 296864 265616
rect 289188 264302 289662 264330
rect 290108 264302 290490 264330
rect 291212 264302 291318 264330
rect 291856 264302 292146 264330
rect 292868 264302 292974 264330
rect 293512 264302 293802 264330
rect 294156 264302 294630 264330
rect 295352 264302 295458 264330
rect 295812 264302 296286 264330
rect 297100 264316 297128 267706
rect 297548 265668 297600 265674
rect 297548 265610 297600 265616
rect 297560 264330 297588 265610
rect 298388 264330 298416 274790
rect 299480 274712 299532 274718
rect 299480 274654 299532 274660
rect 299492 264330 299520 274654
rect 300044 264330 300072 275198
rect 300964 266422 300992 278038
rect 301136 275392 301188 275398
rect 301136 275334 301188 275340
rect 300952 266416 301004 266422
rect 300952 266358 301004 266364
rect 301148 264330 301176 275334
rect 302056 266416 302108 266422
rect 302056 266358 302108 266364
rect 297560 264302 297942 264330
rect 298388 264302 298770 264330
rect 299492 264302 299598 264330
rect 300044 264302 300426 264330
rect 301148 264302 301254 264330
rect 302068 264316 302096 266358
rect 302436 264330 302464 278038
rect 303448 274718 303476 278052
rect 303724 278038 304658 278066
rect 305012 278038 305854 278066
rect 306392 278038 307050 278066
rect 307772 278038 308154 278066
rect 309152 278038 309350 278066
rect 303436 274712 303488 274718
rect 303436 274654 303488 274660
rect 303724 266422 303752 278038
rect 303988 274712 304040 274718
rect 303988 274654 304040 274660
rect 303712 266416 303764 266422
rect 303712 266358 303764 266364
rect 304000 264330 304028 274654
rect 304540 266416 304592 266422
rect 304540 266358 304592 266364
rect 302436 264302 302910 264330
rect 303738 264302 304028 264330
rect 304552 264316 304580 266358
rect 305012 264330 305040 278038
rect 306392 266370 306420 278038
rect 307772 267734 307800 278038
rect 306208 266342 306420 266370
rect 307496 267706 307800 267734
rect 305012 264302 305394 264330
rect 306208 264316 306236 266342
rect 307496 264330 307524 267706
rect 308680 266688 308732 266694
rect 308680 266630 308732 266636
rect 307852 266416 307904 266422
rect 307852 266358 307904 266364
rect 307050 264302 307524 264330
rect 307864 264316 307892 266358
rect 308692 264316 308720 266630
rect 309152 266422 309180 278038
rect 310532 277394 310560 278052
rect 310992 278038 311742 278066
rect 311912 278038 312938 278066
rect 313292 278038 314134 278066
rect 314672 278038 315238 278066
rect 316052 278038 316434 278066
rect 317432 278038 317630 278066
rect 318826 278038 319300 278066
rect 310532 277366 310652 277394
rect 310624 266694 310652 277366
rect 310612 266688 310664 266694
rect 310612 266630 310664 266636
rect 310336 266552 310388 266558
rect 310336 266494 310388 266500
rect 309140 266416 309192 266422
rect 309140 266358 309192 266364
rect 309508 266416 309560 266422
rect 309508 266358 309560 266364
rect 309520 264316 309548 266358
rect 310348 264316 310376 266494
rect 310992 266422 311020 278038
rect 311912 266558 311940 278038
rect 312820 267028 312872 267034
rect 312820 266970 312872 266976
rect 311900 266552 311952 266558
rect 311900 266494 311952 266500
rect 312360 266552 312412 266558
rect 312360 266494 312412 266500
rect 310980 266416 311032 266422
rect 310980 266358 311032 266364
rect 311164 266416 311216 266422
rect 311164 266358 311216 266364
rect 311176 264316 311204 266358
rect 312372 264330 312400 266494
rect 312018 264302 312400 264330
rect 312832 264316 312860 266970
rect 313292 266422 313320 278038
rect 313648 267164 313700 267170
rect 313648 267106 313700 267112
rect 313280 266416 313332 266422
rect 313280 266358 313332 266364
rect 313660 264316 313688 267106
rect 314476 266892 314528 266898
rect 314476 266834 314528 266840
rect 314488 264316 314516 266834
rect 314672 266558 314700 278038
rect 315304 267436 315356 267442
rect 315304 267378 315356 267384
rect 314660 266552 314712 266558
rect 314660 266494 314712 266500
rect 315316 264316 315344 267378
rect 316052 267034 316080 278038
rect 317432 267170 317460 278038
rect 319076 272604 319128 272610
rect 319076 272546 319128 272552
rect 318708 272468 318760 272474
rect 318708 272410 318760 272416
rect 318720 267734 318748 272410
rect 318628 267706 318748 267734
rect 317420 267164 317472 267170
rect 317420 267106 317472 267112
rect 316040 267028 316092 267034
rect 316040 266970 316092 266976
rect 317788 267028 317840 267034
rect 317788 266970 317840 266976
rect 316960 266688 317012 266694
rect 316960 266630 317012 266636
rect 316132 266552 316184 266558
rect 316132 266494 316184 266500
rect 316144 264316 316172 266494
rect 316972 264316 317000 266630
rect 317800 264316 317828 266970
rect 318628 264316 318656 267706
rect 319088 267442 319116 272546
rect 319076 267436 319128 267442
rect 319076 267378 319128 267384
rect 319272 266898 319300 278038
rect 319640 278038 320022 278066
rect 320192 278038 321218 278066
rect 321572 278038 322414 278066
rect 322952 278038 323518 278066
rect 319640 272610 319668 278038
rect 319628 272604 319680 272610
rect 319628 272546 319680 272552
rect 319444 269136 319496 269142
rect 319444 269078 319496 269084
rect 319260 266892 319312 266898
rect 319260 266834 319312 266840
rect 319456 264316 319484 269078
rect 320192 266558 320220 278038
rect 321192 274712 321244 274718
rect 321192 274654 321244 274660
rect 321204 267734 321232 274654
rect 321376 270768 321428 270774
rect 321376 270710 321428 270716
rect 321112 267706 321232 267734
rect 320180 266552 320232 266558
rect 320180 266494 320232 266500
rect 320272 266416 320324 266422
rect 320272 266358 320324 266364
rect 320284 264316 320312 266358
rect 321112 264316 321140 267706
rect 321388 266422 321416 270710
rect 321572 266694 321600 278038
rect 322756 273964 322808 273970
rect 322756 273906 322808 273912
rect 321928 267300 321980 267306
rect 321928 267242 321980 267248
rect 321560 266688 321612 266694
rect 321560 266630 321612 266636
rect 321376 266416 321428 266422
rect 321376 266358 321428 266364
rect 321940 264316 321968 267242
rect 322768 264316 322796 273906
rect 322952 267034 322980 278038
rect 324044 272672 324096 272678
rect 324044 272614 324096 272620
rect 322940 267028 322992 267034
rect 322940 266970 322992 266976
rect 324056 264330 324084 272614
rect 324700 272474 324728 278052
rect 325712 278038 325910 278066
rect 325332 272808 325384 272814
rect 325332 272750 325384 272756
rect 324688 272468 324740 272474
rect 324688 272410 324740 272416
rect 325344 266422 325372 272750
rect 325516 271448 325568 271454
rect 325516 271390 325568 271396
rect 324412 266416 324464 266422
rect 324412 266358 324464 266364
rect 325332 266416 325384 266422
rect 325332 266358 325384 266364
rect 323610 264302 324084 264330
rect 324424 264316 324452 266358
rect 325528 264330 325556 271390
rect 325712 269142 325740 278038
rect 326436 275324 326488 275330
rect 326436 275266 326488 275272
rect 325700 269136 325752 269142
rect 325700 269078 325752 269084
rect 326448 264330 326476 275266
rect 327092 270774 327120 278052
rect 328288 274718 328316 278052
rect 328276 274712 328328 274718
rect 328276 274654 328328 274660
rect 329484 273290 329512 278052
rect 330588 273970 330616 278052
rect 330576 273964 330628 273970
rect 330576 273906 330628 273912
rect 327724 273284 327776 273290
rect 327724 273226 327776 273232
rect 329472 273284 329524 273290
rect 329472 273226 329524 273232
rect 327080 270768 327132 270774
rect 327080 270710 327132 270716
rect 326896 269816 326948 269822
rect 326896 269758 326948 269764
rect 325266 264302 325556 264330
rect 326094 264302 326476 264330
rect 326908 264316 326936 269758
rect 327736 267306 327764 273226
rect 331784 272678 331812 278052
rect 331956 274304 332008 274310
rect 331956 274246 332008 274252
rect 331772 272672 331824 272678
rect 331772 272614 331824 272620
rect 329748 272536 329800 272542
rect 329748 272478 329800 272484
rect 329564 271312 329616 271318
rect 329564 271254 329616 271260
rect 327724 267300 327776 267306
rect 327724 267242 327776 267248
rect 327724 266552 327776 266558
rect 327724 266494 327776 266500
rect 327736 264316 327764 266494
rect 328552 266416 328604 266422
rect 328552 266358 328604 266364
rect 328564 264316 328592 266358
rect 329576 264330 329604 271254
rect 329760 266422 329788 272478
rect 331128 271176 331180 271182
rect 331128 271118 331180 271124
rect 330208 269952 330260 269958
rect 330208 269894 330260 269900
rect 329748 266416 329800 266422
rect 329748 266358 329800 266364
rect 329406 264302 329604 264330
rect 330220 264316 330248 269894
rect 331140 267734 331168 271118
rect 331048 267706 331168 267734
rect 331048 264316 331076 267706
rect 331968 266558 331996 274246
rect 332980 272814 333008 278052
rect 333796 272944 333848 272950
rect 333796 272886 333848 272892
rect 332968 272808 333020 272814
rect 332968 272750 333020 272756
rect 332324 272672 332376 272678
rect 332324 272614 332376 272620
rect 331956 266552 332008 266558
rect 331956 266494 332008 266500
rect 332336 264330 332364 272614
rect 332692 266892 332744 266898
rect 332692 266834 332744 266840
rect 331890 264302 332364 264330
rect 332704 264316 332732 266834
rect 333808 264330 333836 272886
rect 334176 271454 334204 278052
rect 335372 275330 335400 278052
rect 335556 278038 336582 278066
rect 335360 275324 335412 275330
rect 335360 275266 335412 275272
rect 335268 273964 335320 273970
rect 335268 273906 335320 273912
rect 334164 271448 334216 271454
rect 334164 271390 334216 271396
rect 334348 270224 334400 270230
rect 334348 270166 334400 270172
rect 333546 264302 333836 264330
rect 334360 264316 334388 270166
rect 335280 267734 335308 273906
rect 335556 269822 335584 278038
rect 337764 274310 337792 278052
rect 337752 274304 337804 274310
rect 337752 274246 337804 274252
rect 337752 274100 337804 274106
rect 337752 274042 337804 274048
rect 335544 269816 335596 269822
rect 335544 269758 335596 269764
rect 336004 269816 336056 269822
rect 336004 269758 336056 269764
rect 335188 267706 335308 267734
rect 335188 264316 335216 267706
rect 336016 264316 336044 269758
rect 337764 267734 337792 274042
rect 338868 272542 338896 278052
rect 338856 272536 338908 272542
rect 338856 272478 338908 272484
rect 339224 272536 339276 272542
rect 339224 272478 339276 272484
rect 337936 271584 337988 271590
rect 337936 271526 337988 271532
rect 337672 267706 337792 267734
rect 336832 266416 336884 266422
rect 336832 266358 336884 266364
rect 336844 264316 336872 266358
rect 337672 264316 337700 267706
rect 337948 266422 337976 271526
rect 338488 268524 338540 268530
rect 338488 268466 338540 268472
rect 337936 266416 337988 266422
rect 337936 266358 337988 266364
rect 338500 264316 338528 268466
rect 339236 264330 339264 272478
rect 340064 271318 340092 278052
rect 340892 278038 341274 278066
rect 340052 271312 340104 271318
rect 340052 271254 340104 271260
rect 340604 271312 340656 271318
rect 340604 271254 340656 271260
rect 340616 264330 340644 271254
rect 340892 269958 340920 278038
rect 342456 271182 342484 278052
rect 343652 272678 343680 278052
rect 343836 278038 344862 278066
rect 343640 272672 343692 272678
rect 343640 272614 343692 272620
rect 342444 271176 342496 271182
rect 342444 271118 342496 271124
rect 343548 271176 343600 271182
rect 343548 271118 343600 271124
rect 340880 269952 340932 269958
rect 340880 269894 340932 269900
rect 341800 269952 341852 269958
rect 341800 269894 341852 269900
rect 340972 267436 341024 267442
rect 340972 267378 341024 267384
rect 339236 264302 339342 264330
rect 340170 264302 340644 264330
rect 340984 264316 341012 267378
rect 341812 264316 341840 269894
rect 343560 267734 343588 271118
rect 343468 267706 343588 267734
rect 342628 266484 342680 266490
rect 342628 266426 342680 266432
rect 342640 264316 342668 266426
rect 343468 264316 343496 267706
rect 343836 266898 343864 278038
rect 345952 272950 345980 278052
rect 346412 278038 347162 278066
rect 345940 272944 345992 272950
rect 345940 272886 345992 272892
rect 344652 272808 344704 272814
rect 344652 272750 344704 272756
rect 343824 266892 343876 266898
rect 343824 266834 343876 266840
rect 344664 264330 344692 272750
rect 346216 272672 346268 272678
rect 346216 272614 346268 272620
rect 345296 270088 345348 270094
rect 345296 270030 345348 270036
rect 345112 266620 345164 266626
rect 345112 266562 345164 266568
rect 344310 264302 344692 264330
rect 345124 264316 345152 266562
rect 345308 266490 345336 270030
rect 345296 266484 345348 266490
rect 345296 266426 345348 266432
rect 346228 264330 346256 272614
rect 346412 270230 346440 278038
rect 348344 273970 348372 278052
rect 349172 278038 349554 278066
rect 348332 273964 348384 273970
rect 348332 273906 348384 273912
rect 348424 272944 348476 272950
rect 348424 272886 348476 272892
rect 347688 271448 347740 271454
rect 347688 271390 347740 271396
rect 346400 270224 346452 270230
rect 346400 270166 346452 270172
rect 347504 266756 347556 266762
rect 347504 266698 347556 266704
rect 346768 266416 346820 266422
rect 346768 266358 346820 266364
rect 345966 264302 346256 264330
rect 346780 264316 346808 266358
rect 347516 264330 347544 266698
rect 347700 266422 347728 271390
rect 348436 266626 348464 272886
rect 349172 269822 349200 278038
rect 350356 273964 350408 273970
rect 350356 273906 350408 273912
rect 349160 269816 349212 269822
rect 349160 269758 349212 269764
rect 348792 268388 348844 268394
rect 348792 268330 348844 268336
rect 348424 266620 348476 266626
rect 348424 266562 348476 266568
rect 347688 266416 347740 266422
rect 347688 266358 347740 266364
rect 348804 264330 348832 268330
rect 350080 266552 350132 266558
rect 350080 266494 350132 266500
rect 349252 266416 349304 266422
rect 349252 266358 349304 266364
rect 347516 264302 347622 264330
rect 348450 264302 348832 264330
rect 349264 264316 349292 266358
rect 350092 264316 350120 266494
rect 350368 266422 350396 273906
rect 350736 271590 350764 278052
rect 351932 274106 351960 278052
rect 352116 278038 353142 278066
rect 351920 274100 351972 274106
rect 351920 274042 351972 274048
rect 351184 271720 351236 271726
rect 351184 271662 351236 271668
rect 350724 271584 350776 271590
rect 350724 271526 350776 271532
rect 350908 267300 350960 267306
rect 350908 267242 350960 267248
rect 350356 266416 350408 266422
rect 350356 266358 350408 266364
rect 350920 264316 350948 267242
rect 351196 266762 351224 271662
rect 351736 269816 351788 269822
rect 351736 269758 351788 269764
rect 351184 266756 351236 266762
rect 351184 266698 351236 266704
rect 351748 264316 351776 269758
rect 352116 268530 352144 278038
rect 353944 274100 353996 274106
rect 353944 274042 353996 274048
rect 352564 268660 352616 268666
rect 352564 268602 352616 268608
rect 352104 268524 352156 268530
rect 352104 268466 352156 268472
rect 352576 264316 352604 268602
rect 353392 267708 353444 267714
rect 353392 267650 353444 267656
rect 353404 264316 353432 267650
rect 353956 266558 353984 274042
rect 354232 272542 354260 278052
rect 355152 278038 355442 278066
rect 354220 272536 354272 272542
rect 354220 272478 354272 272484
rect 354496 272536 354548 272542
rect 354496 272478 354548 272484
rect 353944 266552 353996 266558
rect 353944 266494 353996 266500
rect 354508 264330 354536 272478
rect 355152 271318 355180 278038
rect 356624 271862 356652 278052
rect 357452 278038 357834 278066
rect 358832 278038 359030 278066
rect 355324 271856 355376 271862
rect 355324 271798 355376 271804
rect 356612 271856 356664 271862
rect 356612 271798 356664 271804
rect 355140 271312 355192 271318
rect 355140 271254 355192 271260
rect 355048 270360 355100 270366
rect 355048 270302 355100 270308
rect 354246 264302 354536 264330
rect 355060 264316 355088 270302
rect 355336 267442 355364 271798
rect 357164 271312 357216 271318
rect 357164 271254 357216 271260
rect 355324 267436 355376 267442
rect 355324 267378 355376 267384
rect 355876 266552 355928 266558
rect 355876 266494 355928 266500
rect 355888 264316 355916 266494
rect 357176 264330 357204 271254
rect 357452 269958 357480 278038
rect 358636 275460 358688 275466
rect 358636 275402 358688 275408
rect 357440 269952 357492 269958
rect 357440 269894 357492 269900
rect 357532 266416 357584 266422
rect 357532 266358 357584 266364
rect 356730 264302 357204 264330
rect 357544 264316 357572 266358
rect 358648 264330 358676 275402
rect 358832 270094 358860 278038
rect 359464 274236 359516 274242
rect 359464 274178 359516 274184
rect 358820 270088 358872 270094
rect 358820 270030 358872 270036
rect 359188 269952 359240 269958
rect 359188 269894 359240 269900
rect 358386 264302 358676 264330
rect 359200 264316 359228 269894
rect 359476 266422 359504 274178
rect 360212 271182 360240 278052
rect 361212 273080 361264 273086
rect 361212 273022 361264 273028
rect 360844 271584 360896 271590
rect 360844 271526 360896 271532
rect 360200 271176 360252 271182
rect 360200 271118 360252 271124
rect 360016 266756 360068 266762
rect 360016 266698 360068 266704
rect 359464 266416 359516 266422
rect 359464 266358 359516 266364
rect 360028 264316 360056 266698
rect 360856 266558 360884 271526
rect 360844 266552 360896 266558
rect 360844 266494 360896 266500
rect 361224 264330 361252 273022
rect 361408 272814 361436 278052
rect 362512 272950 362540 278052
rect 362776 273216 362828 273222
rect 362776 273158 362828 273164
rect 362500 272944 362552 272950
rect 362500 272886 362552 272892
rect 361396 272808 361448 272814
rect 361396 272750 361448 272756
rect 362224 272808 362276 272814
rect 362224 272750 362276 272756
rect 362236 267306 362264 272750
rect 362224 267300 362276 267306
rect 362224 267242 362276 267248
rect 362500 266892 362552 266898
rect 362500 266834 362552 266840
rect 361672 266416 361724 266422
rect 361672 266358 361724 266364
rect 360870 264302 361252 264330
rect 361684 264316 361712 266358
rect 362512 264316 362540 266834
rect 362788 266422 362816 273158
rect 363708 272678 363736 278052
rect 363880 275596 363932 275602
rect 363880 275538 363932 275544
rect 363696 272672 363748 272678
rect 363696 272614 363748 272620
rect 363892 267734 363920 275538
rect 364904 271454 364932 278052
rect 365444 272944 365496 272950
rect 365444 272886 365496 272892
rect 364892 271448 364944 271454
rect 364892 271390 364944 271396
rect 364156 271176 364208 271182
rect 364156 271118 364208 271124
rect 363800 267706 363920 267734
rect 362776 266416 362828 266422
rect 362776 266358 362828 266364
rect 363800 264330 363828 267706
rect 363354 264302 363828 264330
rect 364168 264316 364196 271118
rect 365456 264330 365484 272886
rect 366100 271726 366128 278052
rect 367112 278038 367310 278066
rect 366088 271720 366140 271726
rect 366088 271662 366140 271668
rect 366364 271448 366416 271454
rect 366364 271390 366416 271396
rect 365812 267164 365864 267170
rect 365812 267106 365864 267112
rect 365010 264302 365484 264330
rect 365824 264316 365852 267106
rect 366376 266762 366404 271390
rect 366640 270088 366692 270094
rect 366640 270030 366692 270036
rect 366364 266756 366416 266762
rect 366364 266698 366416 266704
rect 366652 264316 366680 270030
rect 367112 268394 367140 278038
rect 368492 273970 368520 278052
rect 368940 274372 368992 274378
rect 368940 274314 368992 274320
rect 368480 273964 368532 273970
rect 368480 273906 368532 273912
rect 367468 268524 367520 268530
rect 367468 268466 367520 268472
rect 367100 268388 367152 268394
rect 367100 268330 367152 268336
rect 367480 264316 367508 268466
rect 368296 267572 368348 267578
rect 368296 267514 368348 267520
rect 368308 264316 368336 267514
rect 368952 266898 368980 274314
rect 369596 274106 369624 278052
rect 369584 274100 369636 274106
rect 369584 274042 369636 274048
rect 370792 272814 370820 278052
rect 371252 278038 372002 278066
rect 372632 278038 373198 278066
rect 371056 275324 371108 275330
rect 371056 275266 371108 275272
rect 370780 272808 370832 272814
rect 370780 272750 370832 272756
rect 370504 272672 370556 272678
rect 370504 272614 370556 272620
rect 368940 266892 368992 266898
rect 368940 266834 368992 266840
rect 369952 266552 370004 266558
rect 369952 266494 370004 266500
rect 369124 266416 369176 266422
rect 369124 266358 369176 266364
rect 369136 264316 369164 266358
rect 369964 264316 369992 266494
rect 370516 266422 370544 272614
rect 370504 266416 370556 266422
rect 370504 266358 370556 266364
rect 371068 264330 371096 275266
rect 371252 269822 371280 278038
rect 372252 270224 372304 270230
rect 372252 270166 372304 270172
rect 371240 269816 371292 269822
rect 371240 269758 371292 269764
rect 371608 267436 371660 267442
rect 371608 267378 371660 267384
rect 370806 264302 371096 264330
rect 371620 264316 371648 267378
rect 372264 266558 372292 270166
rect 372632 268666 372660 278038
rect 374380 277394 374408 278052
rect 374380 277366 374500 277394
rect 373264 274100 373316 274106
rect 373264 274042 373316 274048
rect 372620 268660 372672 268666
rect 372620 268602 372672 268608
rect 372436 268388 372488 268394
rect 372436 268330 372488 268336
rect 372252 266552 372304 266558
rect 372252 266494 372304 266500
rect 372448 264316 372476 268330
rect 373276 267442 373304 274042
rect 374472 267714 374500 277366
rect 375576 272542 375604 278052
rect 376786 278038 376984 278066
rect 376116 272672 376168 272678
rect 376116 272614 376168 272620
rect 375564 272536 375616 272542
rect 375564 272478 375616 272484
rect 375288 271856 375340 271862
rect 375288 271798 375340 271804
rect 374460 267708 374512 267714
rect 374460 267650 374512 267656
rect 373264 267436 373316 267442
rect 373264 267378 373316 267384
rect 373264 267300 373316 267306
rect 373264 267242 373316 267248
rect 373276 264316 373304 267242
rect 374920 266552 374972 266558
rect 374920 266494 374972 266500
rect 374092 266416 374144 266422
rect 374092 266358 374144 266364
rect 374104 264316 374132 266358
rect 374932 264316 374960 266494
rect 375300 266422 375328 271798
rect 375288 266416 375340 266422
rect 375288 266358 375340 266364
rect 376128 264330 376156 272614
rect 376956 270366 376984 278038
rect 377680 273964 377732 273970
rect 377680 273906 377732 273912
rect 376944 270360 376996 270366
rect 376944 270302 376996 270308
rect 376576 269816 376628 269822
rect 376576 269758 376628 269764
rect 375774 264302 376156 264330
rect 376588 264316 376616 269758
rect 377692 264330 377720 273906
rect 377876 271590 377904 278052
rect 377864 271584 377916 271590
rect 377864 271526 377916 271532
rect 379072 271318 379100 278052
rect 380268 274242 380296 278052
rect 381464 275466 381492 278052
rect 382292 278038 382674 278066
rect 381452 275460 381504 275466
rect 381452 275402 381504 275408
rect 381544 274508 381596 274514
rect 381544 274450 381596 274456
rect 380256 274236 380308 274242
rect 380256 274178 380308 274184
rect 379428 272536 379480 272542
rect 379428 272478 379480 272484
rect 379060 271312 379112 271318
rect 379060 271254 379112 271260
rect 378232 267708 378284 267714
rect 378232 267650 378284 267656
rect 377430 264302 377720 264330
rect 378244 264316 378272 267650
rect 379440 264330 379468 272478
rect 380532 270360 380584 270366
rect 380532 270302 380584 270308
rect 380544 266558 380572 270302
rect 380716 267436 380768 267442
rect 380716 267378 380768 267384
rect 380532 266552 380584 266558
rect 380532 266494 380584 266500
rect 379888 266416 379940 266422
rect 379888 266358 379940 266364
rect 379086 264302 379468 264330
rect 379900 264316 379928 266358
rect 380728 264316 380756 267378
rect 381556 267170 381584 274450
rect 382004 271720 382056 271726
rect 382004 271662 382056 271668
rect 381544 267164 381596 267170
rect 381544 267106 381596 267112
rect 382016 264330 382044 271662
rect 382292 269958 382320 278038
rect 383856 271454 383884 278052
rect 385052 274666 385080 278052
rect 385960 275460 386012 275466
rect 385960 275402 386012 275408
rect 384960 274638 385080 274666
rect 384960 273086 384988 274638
rect 384948 273080 385000 273086
rect 384948 273022 385000 273028
rect 385684 273080 385736 273086
rect 385684 273022 385736 273028
rect 384948 272128 385000 272134
rect 384948 272070 385000 272076
rect 383844 271448 383896 271454
rect 383844 271390 383896 271396
rect 384764 271448 384816 271454
rect 384764 271390 384816 271396
rect 382280 269952 382332 269958
rect 382280 269894 382332 269900
rect 383016 269952 383068 269958
rect 383016 269894 383068 269900
rect 382372 268932 382424 268938
rect 382372 268874 382424 268880
rect 381570 264302 382044 264330
rect 382384 264316 382412 268874
rect 383028 266422 383056 269894
rect 383200 267164 383252 267170
rect 383200 267106 383252 267112
rect 383016 266416 383068 266422
rect 383016 266358 383068 266364
rect 383212 264316 383240 267106
rect 384028 266416 384080 266422
rect 384028 266358 384080 266364
rect 384040 264316 384068 266358
rect 384776 264330 384804 271390
rect 384960 266422 384988 272070
rect 385696 267578 385724 273022
rect 385684 267572 385736 267578
rect 385684 267514 385736 267520
rect 384948 266416 385000 266422
rect 384948 266358 385000 266364
rect 385972 264330 386000 275402
rect 386156 273222 386184 278052
rect 387352 274378 387380 278052
rect 388548 275602 388576 278052
rect 388536 275596 388588 275602
rect 388536 275538 388588 275544
rect 387340 274372 387392 274378
rect 387340 274314 387392 274320
rect 388996 274236 389048 274242
rect 388996 274178 389048 274184
rect 386144 273216 386196 273222
rect 386144 273158 386196 273164
rect 387708 271584 387760 271590
rect 387708 271526 387760 271532
rect 387340 268796 387392 268802
rect 387340 268738 387392 268744
rect 386512 266416 386564 266422
rect 386512 266358 386564 266364
rect 384776 264302 384882 264330
rect 385710 264302 386000 264330
rect 386524 264316 386552 266358
rect 387352 264316 387380 268738
rect 387720 266422 387748 271526
rect 388168 266756 388220 266762
rect 388168 266698 388220 266704
rect 387708 266416 387760 266422
rect 387708 266358 387760 266364
rect 388180 264316 388208 266698
rect 389008 264316 389036 274178
rect 389744 271182 389772 278052
rect 390940 272950 390968 278052
rect 392136 274514 392164 278052
rect 392124 274508 392176 274514
rect 392124 274450 392176 274456
rect 390928 272944 390980 272950
rect 390928 272886 390980 272892
rect 391848 272264 391900 272270
rect 391848 272206 391900 272212
rect 390284 271312 390336 271318
rect 390284 271254 390336 271260
rect 389732 271176 389784 271182
rect 389732 271118 389784 271124
rect 390296 264330 390324 271254
rect 390652 266892 390704 266898
rect 390652 266834 390704 266840
rect 389850 264302 390324 264330
rect 390664 264316 390692 266834
rect 391860 264330 391888 272206
rect 393332 270094 393360 278052
rect 393516 278038 394450 278066
rect 393320 270088 393372 270094
rect 393320 270030 393372 270036
rect 392032 269680 392084 269686
rect 392032 269622 392084 269628
rect 392044 267306 392072 269622
rect 393320 268660 393372 268666
rect 393320 268602 393372 268608
rect 392032 267300 392084 267306
rect 392032 267242 392084 267248
rect 393136 267028 393188 267034
rect 393136 266970 393188 266976
rect 392308 266416 392360 266422
rect 392308 266358 392360 266364
rect 391506 264302 391888 264330
rect 392320 264316 392348 266358
rect 393148 264316 393176 266970
rect 393332 266422 393360 268602
rect 393516 268530 393544 278038
rect 395632 273086 395660 278052
rect 395620 273080 395672 273086
rect 395620 273022 395672 273028
rect 396828 272814 396856 278052
rect 397472 278038 398038 278066
rect 397000 273828 397052 273834
rect 397000 273770 397052 273776
rect 396816 272808 396868 272814
rect 396816 272750 396868 272756
rect 395988 272400 396040 272406
rect 395988 272342 396040 272348
rect 394332 271176 394384 271182
rect 394332 271118 394384 271124
rect 393504 268524 393556 268530
rect 393504 268466 393556 268472
rect 393320 266416 393372 266422
rect 393320 266358 393372 266364
rect 394344 264330 394372 271118
rect 394700 270088 394752 270094
rect 394700 270030 394752 270036
rect 394712 267714 394740 270030
rect 394700 267708 394752 267714
rect 394700 267650 394752 267656
rect 394792 266416 394844 266422
rect 394792 266358 394844 266364
rect 393990 264302 394372 264330
rect 394804 264316 394832 266358
rect 396000 264330 396028 272342
rect 397012 267734 397040 273770
rect 397472 270230 397500 278038
rect 399220 275330 399248 278052
rect 399208 275324 399260 275330
rect 399208 275266 399260 275272
rect 400324 274106 400352 278052
rect 400508 278038 401534 278066
rect 401704 278038 402730 278066
rect 400312 274100 400364 274106
rect 400312 274042 400364 274048
rect 400036 273216 400088 273222
rect 400036 273158 400088 273164
rect 397460 270224 397512 270230
rect 397460 270166 397512 270172
rect 397920 270224 397972 270230
rect 397920 270166 397972 270172
rect 397276 268524 397328 268530
rect 397276 268466 397328 268472
rect 396920 267706 397040 267734
rect 396920 264330 396948 267706
rect 395646 264302 396028 264330
rect 396474 264302 396948 264330
rect 397288 264316 397316 268466
rect 397932 267442 397960 270166
rect 397920 267436 397972 267442
rect 397920 267378 397972 267384
rect 398104 267300 398156 267306
rect 398104 267242 398156 267248
rect 398116 264316 398144 267242
rect 399760 266620 399812 266626
rect 399760 266562 399812 266568
rect 398932 266416 398984 266422
rect 398932 266358 398984 266364
rect 398944 264316 398972 266358
rect 399772 264316 399800 266562
rect 400048 266422 400076 273158
rect 400508 268394 400536 278038
rect 401508 274100 401560 274106
rect 401508 274042 401560 274048
rect 400864 270496 400916 270502
rect 400864 270438 400916 270444
rect 400496 268388 400548 268394
rect 400496 268330 400548 268336
rect 400036 266416 400088 266422
rect 400036 266358 400088 266364
rect 400876 264330 400904 270438
rect 401520 267734 401548 274042
rect 401704 269686 401732 278038
rect 403912 271862 403940 278052
rect 404372 278038 405122 278066
rect 404176 273080 404228 273086
rect 404176 273022 404228 273028
rect 403900 271856 403952 271862
rect 403900 271798 403952 271804
rect 403624 270632 403676 270638
rect 403624 270574 403676 270580
rect 401692 269680 401744 269686
rect 401692 269622 401744 269628
rect 401692 269544 401744 269550
rect 401692 269486 401744 269492
rect 400614 264302 400904 264330
rect 401428 267706 401548 267734
rect 401428 264316 401456 267706
rect 401704 267170 401732 269486
rect 402244 268388 402296 268394
rect 402244 268330 402296 268336
rect 401692 267164 401744 267170
rect 401692 267106 401744 267112
rect 402256 264316 402284 268330
rect 403072 267572 403124 267578
rect 403072 267514 403124 267520
rect 403084 264316 403112 267514
rect 403636 266490 403664 270574
rect 403624 266484 403676 266490
rect 403624 266426 403676 266432
rect 404188 264330 404216 273022
rect 404372 270366 404400 278038
rect 405556 272944 405608 272950
rect 405556 272886 405608 272892
rect 404360 270360 404412 270366
rect 404360 270302 404412 270308
rect 404360 269680 404412 269686
rect 404360 269622 404412 269628
rect 404372 266762 404400 269622
rect 404728 267436 404780 267442
rect 404728 267378 404780 267384
rect 404360 266756 404412 266762
rect 404360 266698 404412 266704
rect 403926 264302 404216 264330
rect 404740 264316 404768 267378
rect 405568 264316 405596 272886
rect 406304 272678 406332 278052
rect 407132 278038 407514 278066
rect 406844 272808 406896 272814
rect 406844 272750 406896 272756
rect 406292 272672 406344 272678
rect 406292 272614 406344 272620
rect 406856 264330 406884 272750
rect 407132 269822 407160 278038
rect 408604 273970 408632 278052
rect 408788 278038 409814 278066
rect 408592 273964 408644 273970
rect 408592 273906 408644 273912
rect 407764 270904 407816 270910
rect 407764 270846 407816 270852
rect 407120 269816 407172 269822
rect 407120 269758 407172 269764
rect 407212 266756 407264 266762
rect 407212 266698 407264 266704
rect 406410 264302 406884 264330
rect 407224 264316 407252 266698
rect 407776 266626 407804 270846
rect 408788 270094 408816 278038
rect 410800 276004 410852 276010
rect 410800 275946 410852 275952
rect 409788 274644 409840 274650
rect 409788 274586 409840 274592
rect 409604 270360 409656 270366
rect 409604 270302 409656 270308
rect 408776 270088 408828 270094
rect 408776 270030 408828 270036
rect 408316 269408 408368 269414
rect 408316 269350 408368 269356
rect 408040 267708 408092 267714
rect 408040 267650 408092 267656
rect 407764 266620 407816 266626
rect 407764 266562 407816 266568
rect 408052 264316 408080 267650
rect 408328 266898 408356 269350
rect 408316 266892 408368 266898
rect 408316 266834 408368 266840
rect 408868 266416 408920 266422
rect 408868 266358 408920 266364
rect 408880 264316 408908 266358
rect 409616 264330 409644 270302
rect 409800 266422 409828 274586
rect 409788 266416 409840 266422
rect 409788 266358 409840 266364
rect 410812 264330 410840 275946
rect 410996 272542 411024 278052
rect 411272 278038 412206 278066
rect 412652 278038 413402 278066
rect 410984 272536 411036 272542
rect 410984 272478 411036 272484
rect 411272 269958 411300 278038
rect 412272 272672 412324 272678
rect 412272 272614 412324 272620
rect 411260 269952 411312 269958
rect 411260 269894 411312 269900
rect 412284 266422 412312 272614
rect 412652 270230 412680 278038
rect 413836 274508 413888 274514
rect 413836 274450 413888 274456
rect 412640 270224 412692 270230
rect 412640 270166 412692 270172
rect 412456 270088 412508 270094
rect 412456 270030 412508 270036
rect 411352 266416 411404 266422
rect 411352 266358 411404 266364
rect 412272 266416 412324 266422
rect 412272 266358 412324 266364
rect 409616 264302 409722 264330
rect 410550 264302 410840 264330
rect 411364 264316 411392 266358
rect 412468 264330 412496 270030
rect 413008 267164 413060 267170
rect 413008 267106 413060 267112
rect 412206 264302 412496 264330
rect 413020 264316 413048 267106
rect 413848 264316 413876 274450
rect 414584 271726 414612 278052
rect 415412 278038 415794 278066
rect 416792 278038 416898 278066
rect 414572 271720 414624 271726
rect 414572 271662 414624 271668
rect 414480 270768 414532 270774
rect 414480 270710 414532 270716
rect 414492 266762 414520 270710
rect 414664 270224 414716 270230
rect 414664 270166 414716 270172
rect 414480 266756 414532 266762
rect 414480 266698 414532 266704
rect 414676 264316 414704 270166
rect 415412 268938 415440 278038
rect 416412 275732 416464 275738
rect 416412 275674 416464 275680
rect 415400 268932 415452 268938
rect 415400 268874 415452 268880
rect 416228 268252 416280 268258
rect 416228 268194 416280 268200
rect 416240 267442 416268 268194
rect 416228 267436 416280 267442
rect 416228 267378 416280 267384
rect 416424 266422 416452 275674
rect 416596 272536 416648 272542
rect 416596 272478 416648 272484
rect 415492 266416 415544 266422
rect 415492 266358 415544 266364
rect 416412 266416 416464 266422
rect 416412 266358 416464 266364
rect 415504 264316 415532 266358
rect 416608 264330 416636 272478
rect 416792 269550 416820 278038
rect 418080 272134 418108 278052
rect 418804 275324 418856 275330
rect 418804 275266 418856 275272
rect 418068 272128 418120 272134
rect 418068 272070 418120 272076
rect 417424 271040 417476 271046
rect 417424 270982 417476 270988
rect 417148 269816 417200 269822
rect 417148 269758 417200 269764
rect 416780 269544 416832 269550
rect 416780 269486 416832 269492
rect 416346 264302 416636 264330
rect 417160 264316 417188 269758
rect 417436 267306 417464 270982
rect 417424 267300 417476 267306
rect 417424 267242 417476 267248
rect 418816 266422 418844 275266
rect 419080 274372 419132 274378
rect 419080 274314 419132 274320
rect 417976 266416 418028 266422
rect 417976 266358 418028 266364
rect 418804 266416 418856 266422
rect 418804 266358 418856 266364
rect 417988 264316 418016 266358
rect 419092 264330 419120 274314
rect 419276 271454 419304 278052
rect 420472 275466 420500 278052
rect 420460 275460 420512 275466
rect 420460 275402 420512 275408
rect 420552 275052 420604 275058
rect 420552 274994 420604 275000
rect 420184 271584 420236 271590
rect 420184 271526 420236 271532
rect 419264 271448 419316 271454
rect 419264 271390 419316 271396
rect 419632 269952 419684 269958
rect 419632 269894 419684 269900
rect 418830 264302 419120 264330
rect 419644 264316 419672 269894
rect 420196 267034 420224 271526
rect 420564 267734 420592 274994
rect 421668 271726 421696 278052
rect 422312 278038 422878 278066
rect 423692 278038 423982 278066
rect 422116 273964 422168 273970
rect 422116 273906 422168 273912
rect 421656 271720 421708 271726
rect 421656 271662 421708 271668
rect 420472 267706 420592 267734
rect 420184 267028 420236 267034
rect 420184 266970 420236 266976
rect 420472 264316 420500 267706
rect 421288 267436 421340 267442
rect 421288 267378 421340 267384
rect 421300 264316 421328 267378
rect 422128 264316 422156 273906
rect 422312 268802 422340 278038
rect 423692 269686 423720 278038
rect 425164 274242 425192 278052
rect 425152 274236 425204 274242
rect 425152 274178 425204 274184
rect 425704 274236 425756 274242
rect 425704 274178 425756 274184
rect 423680 269680 423732 269686
rect 423680 269622 423732 269628
rect 423864 269680 423916 269686
rect 423864 269622 423916 269628
rect 422300 268796 422352 268802
rect 422300 268738 422352 268744
rect 422300 268116 422352 268122
rect 422300 268058 422352 268064
rect 422312 267578 422340 268058
rect 423876 267714 423904 269622
rect 424600 269544 424652 269550
rect 424600 269486 424652 269492
rect 423864 267708 423916 267714
rect 423864 267650 423916 267656
rect 422300 267572 422352 267578
rect 422300 267514 422352 267520
rect 422944 266892 422996 266898
rect 422944 266834 422996 266840
rect 422956 264316 422984 266834
rect 423772 266552 423824 266558
rect 423772 266494 423824 266500
rect 423784 264316 423812 266494
rect 424612 264316 424640 269486
rect 425716 266558 425744 274178
rect 426360 271454 426388 278052
rect 426544 278038 427570 278066
rect 426348 271448 426400 271454
rect 426348 271390 426400 271396
rect 426544 269414 426572 278038
rect 427084 275188 427136 275194
rect 427084 275130 427136 275136
rect 426532 269408 426584 269414
rect 426532 269350 426584 269356
rect 425704 266552 425756 266558
rect 425704 266494 425756 266500
rect 426256 266552 426308 266558
rect 426256 266494 426308 266500
rect 425428 266416 425480 266422
rect 425428 266358 425480 266364
rect 425440 264316 425468 266358
rect 426268 264316 426296 266494
rect 427096 266422 427124 275130
rect 428752 272270 428780 278052
rect 429212 278038 429962 278066
rect 428740 272264 428792 272270
rect 428740 272206 428792 272212
rect 428464 271992 428516 271998
rect 428464 271934 428516 271940
rect 427452 271040 427504 271046
rect 427452 270982 427504 270988
rect 427084 266416 427136 266422
rect 427084 266358 427136 266364
rect 427464 264330 427492 270982
rect 427912 266688 427964 266694
rect 427912 266630 427964 266636
rect 427110 264302 427492 264330
rect 427924 264316 427952 266630
rect 428476 266558 428504 271934
rect 429212 268666 429240 278038
rect 430212 275868 430264 275874
rect 430212 275810 430264 275816
rect 429200 268660 429252 268666
rect 429200 268602 429252 268608
rect 428740 267572 428792 267578
rect 428740 267514 428792 267520
rect 428464 266552 428516 266558
rect 428464 266494 428516 266500
rect 428752 264316 428780 267514
rect 429568 266416 429620 266422
rect 429568 266358 429620 266364
rect 429580 264316 429608 266358
rect 430224 264330 430252 275810
rect 430396 271720 430448 271726
rect 430396 271662 430448 271668
rect 430408 266422 430436 271662
rect 431144 271590 431172 278052
rect 431684 272128 431736 272134
rect 431684 272070 431736 272076
rect 431132 271584 431184 271590
rect 431132 271526 431184 271532
rect 430396 266416 430448 266422
rect 430396 266358 430448 266364
rect 431696 264330 431724 272070
rect 432248 271318 432276 278052
rect 433156 271856 433208 271862
rect 433156 271798 433208 271804
rect 432236 271312 432288 271318
rect 432236 271254 432288 271260
rect 432880 267300 432932 267306
rect 432880 267242 432932 267248
rect 432052 266416 432104 266422
rect 432052 266358 432104 266364
rect 430224 264302 430422 264330
rect 431250 264302 431724 264330
rect 432064 264316 432092 266358
rect 432892 264316 432920 267242
rect 433168 266422 433196 271798
rect 433444 270638 433472 278052
rect 434640 272406 434668 278052
rect 435640 275460 435692 275466
rect 435640 275402 435692 275408
rect 434628 272400 434680 272406
rect 434628 272342 434680 272348
rect 433432 270632 433484 270638
rect 433432 270574 433484 270580
rect 433708 268932 433760 268938
rect 433708 268874 433760 268880
rect 433156 266416 433208 266422
rect 433156 266358 433208 266364
rect 433720 264316 433748 268874
rect 434352 267028 434404 267034
rect 434352 266970 434404 266976
rect 434364 266694 434392 266970
rect 434536 266756 434588 266762
rect 434536 266698 434588 266704
rect 434352 266688 434404 266694
rect 434352 266630 434404 266636
rect 434548 264316 434576 266698
rect 435652 264330 435680 275402
rect 435836 273834 435864 278052
rect 436112 278038 437046 278066
rect 437952 278038 438242 278066
rect 435824 273828 435876 273834
rect 435824 273770 435876 273776
rect 436112 268530 436140 278038
rect 437204 271584 437256 271590
rect 437204 271526 437256 271532
rect 436560 269068 436612 269074
rect 436560 269010 436612 269016
rect 436100 268524 436152 268530
rect 436100 268466 436152 268472
rect 436572 264330 436600 269010
rect 437216 264330 437244 271526
rect 437952 271182 437980 278038
rect 438124 273828 438176 273834
rect 438124 273770 438176 273776
rect 437940 271176 437992 271182
rect 437940 271118 437992 271124
rect 438136 266898 438164 273770
rect 439332 273222 439360 278052
rect 439320 273216 439372 273222
rect 439320 273158 439372 273164
rect 439964 271448 440016 271454
rect 439964 271390 440016 271396
rect 438676 268796 438728 268802
rect 438676 268738 438728 268744
rect 438124 266892 438176 266898
rect 438124 266834 438176 266840
rect 437848 266620 437900 266626
rect 437848 266562 437900 266568
rect 435390 264302 435680 264330
rect 436218 264302 436600 264330
rect 437046 264302 437244 264330
rect 437860 264316 437888 266562
rect 438688 264316 438716 268738
rect 439976 264330 440004 271390
rect 440528 270910 440556 278052
rect 441724 277394 441752 278052
rect 441632 277366 441752 277394
rect 440884 273692 440936 273698
rect 440884 273634 440936 273640
rect 440516 270904 440568 270910
rect 440516 270846 440568 270852
rect 440896 267442 440924 273634
rect 441344 271176 441396 271182
rect 441344 271118 441396 271124
rect 441160 268660 441212 268666
rect 441160 268602 441212 268608
rect 440884 267436 440936 267442
rect 440884 267378 440936 267384
rect 440332 266416 440384 266422
rect 440332 266358 440384 266364
rect 439530 264302 440004 264330
rect 440344 264316 440372 266358
rect 441172 264316 441200 268602
rect 441356 266422 441384 271118
rect 441632 270502 441660 277366
rect 442920 274106 442948 278052
rect 443104 278038 444130 278066
rect 444392 278038 445326 278066
rect 442908 274100 442960 274106
rect 442908 274042 442960 274048
rect 442908 271312 442960 271318
rect 442908 271254 442960 271260
rect 441620 270496 441672 270502
rect 441620 270438 441672 270444
rect 441620 269408 441672 269414
rect 441620 269350 441672 269356
rect 441632 267170 441660 269350
rect 441620 267164 441672 267170
rect 441620 267106 441672 267112
rect 442724 266892 442776 266898
rect 442724 266834 442776 266840
rect 441344 266416 441396 266422
rect 441344 266358 441396 266364
rect 441988 266416 442040 266422
rect 441988 266358 442040 266364
rect 442000 264316 442028 266358
rect 442736 264330 442764 266834
rect 442920 266422 442948 271254
rect 443104 268394 443132 278038
rect 444012 273216 444064 273222
rect 444012 273158 444064 273164
rect 443092 268388 443144 268394
rect 443092 268330 443144 268336
rect 442908 266416 442960 266422
rect 442908 266358 442960 266364
rect 444024 264330 444052 273158
rect 444392 268122 444420 278038
rect 445024 275596 445076 275602
rect 445024 275538 445076 275544
rect 445036 271182 445064 275538
rect 446508 273086 446536 278052
rect 447152 278038 447626 278066
rect 446496 273080 446548 273086
rect 446496 273022 446548 273028
rect 446864 273080 446916 273086
rect 446864 273022 446916 273028
rect 445024 271176 445076 271182
rect 445024 271118 445076 271124
rect 445668 271176 445720 271182
rect 445668 271118 445720 271124
rect 444380 268116 444432 268122
rect 444380 268058 444432 268064
rect 445300 267708 445352 267714
rect 445300 267650 445352 267656
rect 444472 266416 444524 266422
rect 444472 266358 444524 266364
rect 442736 264302 442842 264330
rect 443670 264302 444052 264330
rect 444484 264316 444512 266358
rect 445312 264316 445340 267650
rect 445680 266422 445708 271118
rect 446128 268524 446180 268530
rect 446128 268466 446180 268472
rect 445668 266416 445720 266422
rect 445668 266358 445720 266364
rect 446140 264316 446168 268466
rect 446876 264330 446904 273022
rect 447152 268258 447180 278038
rect 447784 273556 447836 273562
rect 447784 273498 447836 273504
rect 447140 268252 447192 268258
rect 447140 268194 447192 268200
rect 447796 267578 447824 273498
rect 448808 272950 448836 278052
rect 448796 272944 448848 272950
rect 448796 272886 448848 272892
rect 450004 272814 450032 278052
rect 450832 278038 451214 278066
rect 451384 278038 452410 278066
rect 449992 272808 450044 272814
rect 449992 272750 450044 272756
rect 449716 272400 449768 272406
rect 449716 272342 449768 272348
rect 449164 270904 449216 270910
rect 449164 270846 449216 270852
rect 448428 268252 448480 268258
rect 448428 268194 448480 268200
rect 447784 267572 447836 267578
rect 447784 267514 447836 267520
rect 447784 267436 447836 267442
rect 447784 267378 447836 267384
rect 446876 264302 446982 264330
rect 447796 264316 447824 267378
rect 448440 266626 448468 268194
rect 449176 266762 449204 270846
rect 449164 266756 449216 266762
rect 449164 266698 449216 266704
rect 448428 266620 448480 266626
rect 448428 266562 448480 266568
rect 448612 266416 448664 266422
rect 448612 266358 448664 266364
rect 448624 264316 448652 266358
rect 449728 264330 449756 272342
rect 450544 272264 450596 272270
rect 450544 272206 450596 272212
rect 450268 267572 450320 267578
rect 450268 267514 450320 267520
rect 449466 264302 449756 264330
rect 450280 264316 450308 267514
rect 450556 266422 450584 272206
rect 450832 270774 450860 278038
rect 451188 274100 451240 274106
rect 451188 274042 451240 274048
rect 450820 270768 450872 270774
rect 450820 270710 450872 270716
rect 451200 267734 451228 274042
rect 451384 269686 451412 278038
rect 453592 274650 453620 278052
rect 454052 278038 454710 278066
rect 453580 274644 453632 274650
rect 453580 274586 453632 274592
rect 452292 272808 452344 272814
rect 452292 272750 452344 272756
rect 451372 269680 451424 269686
rect 451372 269622 451424 269628
rect 451108 267706 451228 267734
rect 450544 266416 450596 266422
rect 450544 266358 450596 266364
rect 451108 264316 451136 267706
rect 452304 264330 452332 272750
rect 453304 270632 453356 270638
rect 453304 270574 453356 270580
rect 453316 267306 453344 270574
rect 454052 270366 454080 278038
rect 455892 276010 455920 278052
rect 455880 276004 455932 276010
rect 455880 275946 455932 275952
rect 456432 276004 456484 276010
rect 456432 275946 456484 275952
rect 456064 274508 456116 274514
rect 456064 274450 456116 274456
rect 456076 274106 456104 274450
rect 456064 274100 456116 274106
rect 456064 274042 456116 274048
rect 456248 274100 456300 274106
rect 456248 274042 456300 274048
rect 456260 273562 456288 274042
rect 456248 273556 456300 273562
rect 456248 273498 456300 273504
rect 455328 272944 455380 272950
rect 455328 272886 455380 272892
rect 454040 270360 454092 270366
rect 454040 270302 454092 270308
rect 453580 269680 453632 269686
rect 453580 269622 453632 269628
rect 453304 267300 453356 267306
rect 453304 267242 453356 267248
rect 452752 266552 452804 266558
rect 452752 266494 452804 266500
rect 451950 264302 452332 264330
rect 452764 264316 452792 266494
rect 453592 264316 453620 269622
rect 455144 267164 455196 267170
rect 455144 267106 455196 267112
rect 454408 266416 454460 266422
rect 454408 266358 454460 266364
rect 454420 264316 454448 266358
rect 455156 264330 455184 267106
rect 455340 266422 455368 272886
rect 456444 271810 456472 275946
rect 457088 272678 457116 278052
rect 458284 277394 458312 278052
rect 458192 277366 458312 277394
rect 458468 278038 459494 278066
rect 457444 273556 457496 273562
rect 457444 273498 457496 273504
rect 457076 272672 457128 272678
rect 457076 272614 457128 272620
rect 457260 272672 457312 272678
rect 457260 272614 457312 272620
rect 456076 271782 456472 271810
rect 456076 267442 456104 271782
rect 456432 270496 456484 270502
rect 456432 270438 456484 270444
rect 456064 267436 456116 267442
rect 456064 267378 456116 267384
rect 455328 266416 455380 266422
rect 455328 266358 455380 266364
rect 456444 264330 456472 270438
rect 457272 264330 457300 272614
rect 457456 267034 457484 273498
rect 458192 270094 458220 277366
rect 458180 270088 458232 270094
rect 458180 270030 458232 270036
rect 458468 269414 458496 278038
rect 460676 274650 460704 278052
rect 461228 278038 461886 278066
rect 460664 274644 460716 274650
rect 460664 274586 460716 274592
rect 461030 272912 461086 272921
rect 461030 272847 461086 272856
rect 461044 272678 461072 272847
rect 461032 272672 461084 272678
rect 460846 272640 460902 272649
rect 461032 272614 461084 272620
rect 460846 272575 460902 272584
rect 458824 270360 458876 270366
rect 458824 270302 458876 270308
rect 458456 269408 458508 269414
rect 458456 269350 458508 269356
rect 457444 267028 457496 267034
rect 457444 266970 457496 266976
rect 457720 266756 457772 266762
rect 457720 266698 457772 266704
rect 455156 264302 455262 264330
rect 456090 264302 456472 264330
rect 456918 264302 457300 264330
rect 457732 264316 457760 266698
rect 458836 264330 458864 270302
rect 460204 267436 460256 267442
rect 460204 267378 460256 267384
rect 459376 267300 459428 267306
rect 459376 267242 459428 267248
rect 458574 264302 458864 264330
rect 459388 264316 459416 267242
rect 460216 264316 460244 267378
rect 460860 267306 460888 272575
rect 461228 270230 461256 278038
rect 462976 275738 463004 278052
rect 463712 278038 464186 278066
rect 465092 278038 465382 278066
rect 462964 275732 463016 275738
rect 462964 275674 463016 275680
rect 463148 275732 463200 275738
rect 463148 275674 463200 275680
rect 463160 273578 463188 275674
rect 462976 273550 463188 273578
rect 461400 272944 461452 272950
rect 461400 272886 461452 272892
rect 461412 272678 461440 272886
rect 461400 272672 461452 272678
rect 461860 272672 461912 272678
rect 461400 272614 461452 272620
rect 461858 272640 461860 272649
rect 461912 272640 461914 272649
rect 461858 272575 461914 272584
rect 461216 270224 461268 270230
rect 461216 270166 461268 270172
rect 461400 270224 461452 270230
rect 461400 270166 461452 270172
rect 460848 267300 460900 267306
rect 460848 267242 460900 267248
rect 461412 264330 461440 270166
rect 461860 268388 461912 268394
rect 461860 268330 461912 268336
rect 461058 264302 461440 264330
rect 461872 264316 461900 268330
rect 462976 266558 463004 273550
rect 463240 273420 463292 273426
rect 463240 273362 463292 273368
rect 463252 273254 463280 273362
rect 463160 273226 463280 273254
rect 462964 266552 463016 266558
rect 462964 266494 463016 266500
rect 463160 264330 463188 273226
rect 463712 272542 463740 278038
rect 464436 274644 464488 274650
rect 464436 274586 464488 274592
rect 464448 273562 464476 274586
rect 464436 273556 464488 273562
rect 464436 273498 464488 273504
rect 463700 272536 463752 272542
rect 463700 272478 463752 272484
rect 464710 272504 464766 272513
rect 464710 272439 464766 272448
rect 463516 270088 463568 270094
rect 463516 270030 463568 270036
rect 462714 264302 463188 264330
rect 463528 264316 463556 270030
rect 464724 264330 464752 272439
rect 465092 269822 465120 278038
rect 466564 275330 466592 278052
rect 466552 275324 466604 275330
rect 466552 275266 466604 275272
rect 467564 275324 467616 275330
rect 467564 275266 467616 275272
rect 465908 274508 465960 274514
rect 465908 274450 465960 274456
rect 466092 274508 466144 274514
rect 466092 274450 466144 274456
rect 465920 273970 465948 274450
rect 465724 273964 465776 273970
rect 465724 273906 465776 273912
rect 465908 273964 465960 273970
rect 465908 273906 465960 273912
rect 465736 273698 465764 273906
rect 465724 273692 465776 273698
rect 465724 273634 465776 273640
rect 466104 273426 466132 274450
rect 466092 273420 466144 273426
rect 466092 273362 466144 273368
rect 466274 272912 466330 272921
rect 466274 272847 466330 272856
rect 466288 272626 466316 272847
rect 466414 272672 466466 272678
rect 466288 272620 466414 272626
rect 466288 272614 466466 272620
rect 466288 272598 466454 272614
rect 465080 269816 465132 269822
rect 465080 269758 465132 269764
rect 466000 269816 466052 269822
rect 466000 269758 466052 269764
rect 465172 267300 465224 267306
rect 465172 267242 465224 267248
rect 464370 264302 464752 264330
rect 465184 264316 465212 267242
rect 466012 264316 466040 269758
rect 466828 265124 466880 265130
rect 466828 265066 466880 265072
rect 466840 264316 466868 265066
rect 467576 264330 467604 275266
rect 467760 274378 467788 278052
rect 467944 278038 468970 278066
rect 467748 274372 467800 274378
rect 467748 274314 467800 274320
rect 467944 269958 467972 278038
rect 470152 275058 470180 278052
rect 470416 276276 470468 276282
rect 470416 276218 470468 276224
rect 470140 275052 470192 275058
rect 470140 274994 470192 275000
rect 467932 269952 467984 269958
rect 467932 269894 467984 269900
rect 468484 269952 468536 269958
rect 468484 269894 468536 269900
rect 467576 264302 467682 264330
rect 468496 264316 468524 269894
rect 470428 267034 470456 276218
rect 471256 273562 471284 278052
rect 472256 274236 472308 274242
rect 472256 274178 472308 274184
rect 472268 273970 472296 274178
rect 472256 273964 472308 273970
rect 472256 273906 472308 273912
rect 472452 273698 472480 278052
rect 473084 274916 473136 274922
rect 473084 274858 473136 274864
rect 472440 273692 472492 273698
rect 472440 273634 472492 273640
rect 471244 273556 471296 273562
rect 471244 273498 471296 273504
rect 470554 272536 470606 272542
rect 470692 272536 470744 272542
rect 470554 272478 470606 272484
rect 470690 272504 470692 272513
rect 470744 272504 470746 272513
rect 470566 272354 470594 272478
rect 470690 272439 470746 272448
rect 470566 272326 470732 272354
rect 470704 271998 470732 272326
rect 470554 271992 470606 271998
rect 470552 271960 470554 271969
rect 470692 271992 470744 271998
rect 470606 271960 470608 271969
rect 470692 271934 470744 271940
rect 470552 271895 470608 271904
rect 470968 269408 471020 269414
rect 470968 269350 471020 269356
rect 469312 267028 469364 267034
rect 469312 266970 469364 266976
rect 470416 267028 470468 267034
rect 470416 266970 470468 266976
rect 470600 267028 470652 267034
rect 470600 266970 470652 266976
rect 469324 264316 469352 266970
rect 470612 266914 470640 266970
rect 470520 266886 470640 266914
rect 470520 264330 470548 266886
rect 470166 264302 470548 264330
rect 470980 264316 471008 269350
rect 471796 265260 471848 265266
rect 471796 265202 471848 265208
rect 471808 264316 471836 265202
rect 473096 264330 473124 274858
rect 473648 273834 473676 278052
rect 474844 274378 474872 278052
rect 475028 278038 476054 278066
rect 474832 274372 474884 274378
rect 474832 274314 474884 274320
rect 473636 273828 473688 273834
rect 473636 273770 473688 273776
rect 474648 273828 474700 273834
rect 474648 273770 474700 273776
rect 474280 269272 474332 269278
rect 474280 269214 474332 269220
rect 473452 266416 473504 266422
rect 473452 266358 473504 266364
rect 472650 264302 473124 264330
rect 473464 264316 473492 266358
rect 474292 264316 474320 269214
rect 474660 266422 474688 273770
rect 475028 269550 475056 278038
rect 477236 275194 477264 278052
rect 478064 278038 478354 278066
rect 479168 278038 479550 278066
rect 477224 275188 477276 275194
rect 477224 275130 477276 275136
rect 476764 274780 476816 274786
rect 476764 274722 476816 274728
rect 476028 273556 476080 273562
rect 476028 273498 476080 273504
rect 475016 269544 475068 269550
rect 475016 269486 475068 269492
rect 476040 267734 476068 273498
rect 475948 267706 476068 267734
rect 475108 266552 475160 266558
rect 475108 266494 475160 266500
rect 474648 266416 474700 266422
rect 474648 266358 474700 266364
rect 475120 264316 475148 266494
rect 475948 264316 475976 267706
rect 476776 266762 476804 274722
rect 478064 271969 478092 278038
rect 478512 276412 478564 276418
rect 478512 276354 478564 276360
rect 478050 271960 478106 271969
rect 478050 271895 478106 271904
rect 476764 266756 476816 266762
rect 476764 266698 476816 266704
rect 478524 266422 478552 276354
rect 478696 273420 478748 273426
rect 478696 273362 478748 273368
rect 477592 266416 477644 266422
rect 477592 266358 477644 266364
rect 478512 266416 478564 266422
rect 478512 266358 478564 266364
rect 476764 265396 476816 265402
rect 476764 265338 476816 265344
rect 476776 264316 476804 265338
rect 477604 264316 477632 266358
rect 478708 264330 478736 273362
rect 479168 271046 479196 278038
rect 479984 276548 480036 276554
rect 479984 276490 480036 276496
rect 479522 271824 479578 271833
rect 479522 271759 479578 271768
rect 479156 271040 479208 271046
rect 479156 270982 479208 270988
rect 479536 266558 479564 271759
rect 479996 267734 480024 276490
rect 480732 274650 480760 278052
rect 480720 274644 480772 274650
rect 480720 274586 480772 274592
rect 481364 274236 481416 274242
rect 481364 274178 481416 274184
rect 480258 272368 480314 272377
rect 480258 272303 480314 272312
rect 480272 272218 480300 272303
rect 480180 272190 480300 272218
rect 480180 272134 480208 272190
rect 480168 272128 480220 272134
rect 480168 272070 480220 272076
rect 479720 267706 480024 267734
rect 479524 266552 479576 266558
rect 479524 266494 479576 266500
rect 479720 264330 479748 267706
rect 480076 266348 480128 266354
rect 480076 266290 480128 266296
rect 478446 264302 478736 264330
rect 479274 264302 479748 264330
rect 480088 264316 480116 266290
rect 481376 264330 481404 274178
rect 481928 273970 481956 278052
rect 483124 277394 483152 278052
rect 483032 277366 483152 277394
rect 481916 273964 481968 273970
rect 481916 273906 481968 273912
rect 483032 271726 483060 277366
rect 484032 277228 484084 277234
rect 484032 277170 484084 277176
rect 483204 271992 483256 271998
rect 483204 271934 483256 271940
rect 483216 271833 483244 271934
rect 483202 271824 483258 271833
rect 483202 271759 483258 271768
rect 483020 271720 483072 271726
rect 483020 271662 483072 271668
rect 482284 271040 482336 271046
rect 482284 270982 482336 270988
rect 482296 266626 482324 270982
rect 482284 266620 482336 266626
rect 482284 266562 482336 266568
rect 482560 266620 482612 266626
rect 482560 266562 482612 266568
rect 481732 265532 481784 265538
rect 481732 265474 481784 265480
rect 480930 264302 481404 264330
rect 481744 264316 481772 265474
rect 482572 264316 482600 266562
rect 483388 266484 483440 266490
rect 483388 266426 483440 266432
rect 483400 264316 483428 266426
rect 484044 264330 484072 277170
rect 484320 275874 484348 278052
rect 484872 278038 485530 278066
rect 484308 275868 484360 275874
rect 484308 275810 484360 275816
rect 484216 273692 484268 273698
rect 484216 273634 484268 273640
rect 484228 266490 484256 273634
rect 484872 272377 484900 278038
rect 485504 277092 485556 277098
rect 485504 277034 485556 277040
rect 485044 275868 485096 275874
rect 485044 275810 485096 275816
rect 485056 275466 485084 275810
rect 485044 275460 485096 275466
rect 485044 275402 485096 275408
rect 485320 274236 485372 274242
rect 485320 274178 485372 274184
rect 485332 273698 485360 274178
rect 485320 273692 485372 273698
rect 485320 273634 485372 273640
rect 484858 272368 484914 272377
rect 484858 272303 484914 272312
rect 485044 271856 485096 271862
rect 485044 271798 485096 271804
rect 485056 266626 485084 271798
rect 485516 267734 485544 277034
rect 485780 275460 485832 275466
rect 485780 275402 485832 275408
rect 485792 274514 485820 275402
rect 485780 274508 485832 274514
rect 485780 274450 485832 274456
rect 486620 271726 486648 278052
rect 486792 274644 486844 274650
rect 486792 274586 486844 274592
rect 486608 271720 486660 271726
rect 486608 271662 486660 271668
rect 485424 267706 485544 267734
rect 485044 266620 485096 266626
rect 485044 266562 485096 266568
rect 484216 266484 484268 266490
rect 484216 266426 484268 266432
rect 485424 264330 485452 267706
rect 486804 266490 486832 274586
rect 486976 270768 487028 270774
rect 486976 270710 487028 270716
rect 485872 266484 485924 266490
rect 485872 266426 485924 266432
rect 486792 266484 486844 266490
rect 486792 266426 486844 266432
rect 484044 264302 484242 264330
rect 485070 264302 485452 264330
rect 485884 264316 485912 266426
rect 486988 264330 487016 270710
rect 487816 270638 487844 278052
rect 488552 278038 489026 278066
rect 488356 274508 488408 274514
rect 488356 274450 488408 274456
rect 487804 270632 487856 270638
rect 487804 270574 487856 270580
rect 487528 266212 487580 266218
rect 487528 266154 487580 266160
rect 486726 264302 487016 264330
rect 487540 264316 487568 266154
rect 488368 264316 488396 274450
rect 488552 268938 488580 278038
rect 489918 272640 489974 272649
rect 489918 272575 489974 272584
rect 489932 272218 489960 272575
rect 489886 272190 489960 272218
rect 489886 272134 489914 272190
rect 489874 272128 489926 272134
rect 489874 272070 489926 272076
rect 490012 272128 490064 272134
rect 490012 272070 490064 272076
rect 490024 271862 490052 272070
rect 490012 271856 490064 271862
rect 490012 271798 490064 271804
rect 490208 270910 490236 278052
rect 491404 275874 491432 278052
rect 491680 278038 492614 278066
rect 491392 275868 491444 275874
rect 491392 275810 491444 275816
rect 490196 270904 490248 270910
rect 490196 270846 490248 270852
rect 489644 270632 489696 270638
rect 489644 270574 489696 270580
rect 488540 268932 488592 268938
rect 488540 268874 488592 268880
rect 489656 264330 489684 270574
rect 491680 269074 491708 278038
rect 493704 271590 493732 278052
rect 494072 278038 494914 278066
rect 495452 278038 496110 278066
rect 493692 271584 493744 271590
rect 493692 271526 493744 271532
rect 492496 270904 492548 270910
rect 492496 270846 492548 270852
rect 491668 269068 491720 269074
rect 491668 269010 491720 269016
rect 490840 267980 490892 267986
rect 490840 267922 490892 267928
rect 490012 266756 490064 266762
rect 490012 266698 490064 266704
rect 489210 264302 489684 264330
rect 490024 264316 490052 266698
rect 490852 264316 490880 267922
rect 492508 267734 492536 270846
rect 492772 269544 492824 269550
rect 492772 269486 492824 269492
rect 492784 267734 492812 269486
rect 493324 269068 493376 269074
rect 493324 269010 493376 269016
rect 492416 267706 492536 267734
rect 492600 267706 492812 267734
rect 492416 266490 492444 267706
rect 491668 266484 491720 266490
rect 491668 266426 491720 266432
rect 492404 266484 492456 266490
rect 492404 266426 492456 266432
rect 491680 264316 491708 266426
rect 492600 265690 492628 267706
rect 492508 265662 492628 265690
rect 492508 264316 492536 265662
rect 493336 264316 493364 269010
rect 494072 268258 494100 278038
rect 495072 276956 495124 276962
rect 495072 276898 495124 276904
rect 494704 271720 494756 271726
rect 494704 271662 494756 271668
rect 494716 271046 494744 271662
rect 494704 271040 494756 271046
rect 494704 270982 494756 270988
rect 494060 268252 494112 268258
rect 494060 268194 494112 268200
rect 495084 267734 495112 276898
rect 495256 271040 495308 271046
rect 495256 270982 495308 270988
rect 494992 267706 495112 267734
rect 494152 266484 494204 266490
rect 494152 266426 494204 266432
rect 494164 264316 494192 266426
rect 494992 264316 495020 267706
rect 495268 266490 495296 270982
rect 495452 268802 495480 278038
rect 496544 271856 496596 271862
rect 496544 271798 496596 271804
rect 495440 268796 495492 268802
rect 495440 268738 495492 268744
rect 495808 268252 495860 268258
rect 495808 268194 495860 268200
rect 495256 266484 495308 266490
rect 495256 266426 495308 266432
rect 495820 264316 495848 268194
rect 496556 264330 496584 271798
rect 497292 271454 497320 278052
rect 498488 275602 498516 278052
rect 499698 278038 500172 278066
rect 498476 275596 498528 275602
rect 498476 275538 498528 275544
rect 498844 275596 498896 275602
rect 498844 275538 498896 275544
rect 497924 275052 497976 275058
rect 497924 274994 497976 275000
rect 497280 271448 497332 271454
rect 497280 271390 497332 271396
rect 497936 264330 497964 274994
rect 498292 268932 498344 268938
rect 498292 268874 498344 268880
rect 496556 264302 496662 264330
rect 497490 264302 497964 264330
rect 498304 264316 498332 268874
rect 498856 267714 498884 275538
rect 499948 273216 500000 273222
rect 499948 273158 500000 273164
rect 499488 273080 499540 273086
rect 499486 273048 499488 273057
rect 499540 273048 499542 273057
rect 499960 273034 499988 273158
rect 499486 272983 499542 272992
rect 499684 273006 499988 273034
rect 499684 272898 499712 273006
rect 499592 272870 499712 272898
rect 499592 272762 499620 272870
rect 499500 272734 499620 272762
rect 499500 272406 499528 272734
rect 499670 272640 499726 272649
rect 499670 272575 499726 272584
rect 499684 272406 499712 272575
rect 499488 272400 499540 272406
rect 499488 272342 499540 272348
rect 499672 272400 499724 272406
rect 499672 272342 499724 272348
rect 499304 271584 499356 271590
rect 499304 271526 499356 271532
rect 498844 267708 498896 267714
rect 498844 267650 498896 267656
rect 499316 264330 499344 271526
rect 500144 268666 500172 278038
rect 500880 271318 500908 278052
rect 501800 278038 501998 278066
rect 501800 271726 501828 278038
rect 503180 273086 503208 278052
rect 503536 277432 503588 277438
rect 503536 277374 503588 277380
rect 503168 273080 503220 273086
rect 503352 273080 503404 273086
rect 503168 273022 503220 273028
rect 503350 273048 503352 273057
rect 503404 273048 503406 273057
rect 503350 272983 503406 272992
rect 501788 271720 501840 271726
rect 501788 271662 501840 271668
rect 501972 271720 502024 271726
rect 501972 271662 502024 271668
rect 500868 271312 500920 271318
rect 500868 271254 500920 271260
rect 500776 268796 500828 268802
rect 500776 268738 500828 268744
rect 500132 268660 500184 268666
rect 500132 268602 500184 268608
rect 499948 266892 500000 266898
rect 499948 266834 500000 266840
rect 499146 264302 499344 264330
rect 499960 264316 499988 266834
rect 500788 264316 500816 268738
rect 501984 264330 502012 271662
rect 503260 268660 503312 268666
rect 503260 268602 503312 268608
rect 502432 266484 502484 266490
rect 502432 266426 502484 266432
rect 501630 264302 502012 264330
rect 502444 264316 502472 266426
rect 503272 264316 503300 268602
rect 503548 266490 503576 277374
rect 504376 271182 504404 278052
rect 505572 275602 505600 278052
rect 506492 278038 506782 278066
rect 505560 275596 505612 275602
rect 505560 275538 505612 275544
rect 505744 275596 505796 275602
rect 505744 275538 505796 275544
rect 505008 271448 505060 271454
rect 505008 271390 505060 271396
rect 504364 271176 504416 271182
rect 504364 271118 504416 271124
rect 504824 266620 504876 266626
rect 504824 266562 504876 266568
rect 503536 266484 503588 266490
rect 503536 266426 503588 266432
rect 504088 266484 504140 266490
rect 504088 266426 504140 266432
rect 504100 264316 504128 266426
rect 504836 264330 504864 266562
rect 505020 266490 505048 271390
rect 505756 267578 505784 275538
rect 506204 274372 506256 274378
rect 506204 274314 506256 274320
rect 505744 267572 505796 267578
rect 505744 267514 505796 267520
rect 505008 266484 505060 266490
rect 505008 266426 505060 266432
rect 506216 264330 506244 274314
rect 506492 268530 506520 278038
rect 507492 275188 507544 275194
rect 507492 275130 507544 275136
rect 506480 268524 506532 268530
rect 506480 268466 506532 268472
rect 507504 267734 507532 275130
rect 507964 273086 507992 278052
rect 509068 276010 509096 278052
rect 509056 276004 509108 276010
rect 509056 275946 509108 275952
rect 507952 273080 508004 273086
rect 507952 273022 508004 273028
rect 509700 273080 509752 273086
rect 509700 273022 509752 273028
rect 507676 271312 507728 271318
rect 507676 271254 507728 271260
rect 507412 267706 507532 267734
rect 506572 266484 506624 266490
rect 506572 266426 506624 266432
rect 504836 264302 504942 264330
rect 505770 264302 506244 264330
rect 506584 264316 506612 266426
rect 507412 264316 507440 267706
rect 507688 266490 507716 271254
rect 509238 269920 509294 269929
rect 509238 269855 509294 269864
rect 509252 269686 509280 269855
rect 509240 269680 509292 269686
rect 509240 269622 509292 269628
rect 509146 269512 509202 269521
rect 509146 269447 509202 269456
rect 508228 268524 508280 268530
rect 508228 268466 508280 268472
rect 507860 266892 507912 266898
rect 507860 266834 507912 266840
rect 507872 266490 507900 266834
rect 507676 266484 507728 266490
rect 507676 266426 507728 266432
rect 507860 266484 507912 266490
rect 507860 266426 507912 266432
rect 508240 264316 508268 268466
rect 509160 267734 509188 269447
rect 509068 267706 509188 267734
rect 509068 264316 509096 267706
rect 509712 266762 509740 273022
rect 510264 272270 510292 278052
rect 511460 273222 511488 278052
rect 512656 275602 512684 278052
rect 513196 276004 513248 276010
rect 513196 275946 513248 275952
rect 512644 275596 512696 275602
rect 512644 275538 512696 275544
rect 511632 274236 511684 274242
rect 511632 274178 511684 274184
rect 511448 273216 511500 273222
rect 511448 273158 511500 273164
rect 510252 272264 510304 272270
rect 510252 272206 510304 272212
rect 509884 269544 509936 269550
rect 509882 269512 509884 269521
rect 509936 269512 509938 269521
rect 509882 269447 509938 269456
rect 509884 267708 509936 267714
rect 509884 267650 509936 267656
rect 509700 266756 509752 266762
rect 509700 266698 509752 266704
rect 509896 264316 509924 267650
rect 511644 266762 511672 274178
rect 513208 266762 513236 275946
rect 513852 274106 513880 278052
rect 514484 276820 514536 276826
rect 514484 276762 514536 276768
rect 513840 274100 513892 274106
rect 513840 274042 513892 274048
rect 513564 273080 513616 273086
rect 513564 273022 513616 273028
rect 513576 272814 513604 273022
rect 513564 272808 513616 272814
rect 513564 272750 513616 272756
rect 513748 272808 513800 272814
rect 513748 272750 513800 272756
rect 513760 272406 513788 272750
rect 513748 272400 513800 272406
rect 513748 272342 513800 272348
rect 510712 266756 510764 266762
rect 510712 266698 510764 266704
rect 511632 266756 511684 266762
rect 511632 266698 511684 266704
rect 512368 266756 512420 266762
rect 512368 266698 512420 266704
rect 513196 266756 513248 266762
rect 513196 266698 513248 266704
rect 510724 264316 510752 266698
rect 511540 266076 511592 266082
rect 511540 266018 511592 266024
rect 511552 264316 511580 266018
rect 512380 264316 512408 266698
rect 513196 265940 513248 265946
rect 513196 265882 513248 265888
rect 513208 264316 513236 265882
rect 514496 264330 514524 276762
rect 515048 272950 515076 278052
rect 516244 275738 516272 278052
rect 516520 278038 517362 278066
rect 516232 275732 516284 275738
rect 516232 275674 516284 275680
rect 515220 273216 515272 273222
rect 515220 273158 515272 273164
rect 515404 273216 515456 273222
rect 515404 273158 515456 273164
rect 515232 272950 515260 273158
rect 515036 272944 515088 272950
rect 515036 272886 515088 272892
rect 515220 272944 515272 272950
rect 515220 272886 515272 272892
rect 514852 267572 514904 267578
rect 514852 267514 514904 267520
rect 514050 264302 514524 264330
rect 514864 264316 514892 267514
rect 515416 267170 515444 273158
rect 516520 269929 516548 278038
rect 516784 275596 516836 275602
rect 516784 275538 516836 275544
rect 516506 269920 516562 269929
rect 516506 269855 516562 269864
rect 516796 267442 516824 275538
rect 518544 273086 518572 278052
rect 519740 273222 519768 278052
rect 520292 278038 520950 278066
rect 519728 273216 519780 273222
rect 519728 273158 519780 273164
rect 518532 273080 518584 273086
rect 518532 273022 518584 273028
rect 517428 272400 517480 272406
rect 517428 272342 517480 272348
rect 516784 267436 516836 267442
rect 516784 267378 516836 267384
rect 515404 267164 515456 267170
rect 515404 267106 515456 267112
rect 517244 267164 517296 267170
rect 517244 267106 517296 267112
rect 516508 266756 516560 266762
rect 516508 266698 516560 266704
rect 515680 265804 515732 265810
rect 515680 265746 515732 265752
rect 515692 264316 515720 265746
rect 516520 264316 516548 266698
rect 517256 264330 517284 267106
rect 517440 266762 517468 272342
rect 520096 272264 520148 272270
rect 520096 272206 520148 272212
rect 519820 267436 519872 267442
rect 519820 267378 519872 267384
rect 517428 266756 517480 266762
rect 517428 266698 517480 266704
rect 518992 266756 519044 266762
rect 518992 266698 519044 266704
rect 518164 265668 518216 265674
rect 518164 265610 518216 265616
rect 517256 264302 517362 264330
rect 518176 264316 518204 265610
rect 519004 264316 519032 266698
rect 519832 264316 519860 267378
rect 520108 266762 520136 272206
rect 520292 270502 520320 278038
rect 521108 276684 521160 276690
rect 521108 276626 521160 276632
rect 520280 270496 520332 270502
rect 520280 270438 520332 270444
rect 520096 266756 520148 266762
rect 520096 266698 520148 266704
rect 521120 264330 521148 276626
rect 521476 273216 521528 273222
rect 521476 273158 521528 273164
rect 520674 264302 521148 264330
rect 521488 264316 521516 273158
rect 522132 272678 522160 278052
rect 522764 275868 522816 275874
rect 522764 275810 522816 275816
rect 522120 272672 522172 272678
rect 522120 272614 522172 272620
rect 522776 264330 522804 275810
rect 523328 274786 523356 278052
rect 524432 278038 524538 278066
rect 523316 274780 523368 274786
rect 523316 274722 523368 274728
rect 523684 274780 523736 274786
rect 523684 274722 523736 274728
rect 523132 270496 523184 270502
rect 523132 270438 523184 270444
rect 522330 264302 522804 264330
rect 523144 264316 523172 270438
rect 523696 267306 523724 274722
rect 524052 271176 524104 271182
rect 524052 271118 524104 271124
rect 524064 267734 524092 271118
rect 524432 270366 524460 278038
rect 525628 272814 525656 278052
rect 526824 275602 526852 278052
rect 527192 278038 528034 278066
rect 528572 278038 529230 278066
rect 526812 275596 526864 275602
rect 526812 275538 526864 275544
rect 525616 272808 525668 272814
rect 525616 272750 525668 272756
rect 526812 272672 526864 272678
rect 526812 272614 526864 272620
rect 524420 270360 524472 270366
rect 524420 270302 524472 270308
rect 525616 270360 525668 270366
rect 525616 270302 525668 270308
rect 523972 267706 524092 267734
rect 523684 267300 523736 267306
rect 523684 267242 523736 267248
rect 523972 264316 524000 267706
rect 524788 267300 524840 267306
rect 524788 267242 524840 267248
rect 524800 264316 524828 267242
rect 525628 264316 525656 270302
rect 526824 264330 526852 272614
rect 527192 270230 527220 278038
rect 528192 275732 528244 275738
rect 528192 275674 528244 275680
rect 527180 270224 527232 270230
rect 527180 270166 527232 270172
rect 527180 268116 527232 268122
rect 527180 268058 527232 268064
rect 527192 267170 527220 268058
rect 527180 267164 527232 267170
rect 527180 267106 527232 267112
rect 528204 266762 528232 275674
rect 528376 270224 528428 270230
rect 528376 270166 528428 270172
rect 527272 266756 527324 266762
rect 527272 266698 527324 266704
rect 528192 266756 528244 266762
rect 528192 266698 528244 266704
rect 526470 264302 526852 264330
rect 527284 264316 527312 266698
rect 528388 264330 528416 270166
rect 528572 268394 528600 278038
rect 530412 275466 530440 278052
rect 531332 278038 531622 278066
rect 530400 275460 530452 275466
rect 530400 275402 530452 275408
rect 529848 272808 529900 272814
rect 529848 272750 529900 272756
rect 528560 268388 528612 268394
rect 528560 268330 528612 268336
rect 529664 267164 529716 267170
rect 529664 267106 529716 267112
rect 528928 266756 528980 266762
rect 528928 266698 528980 266704
rect 528126 264302 528416 264330
rect 528940 264316 528968 266698
rect 529676 264330 529704 267106
rect 529860 266762 529888 272750
rect 531332 270178 531360 278038
rect 532332 275596 532384 275602
rect 532332 275538 532384 275544
rect 532344 270314 532372 275538
rect 532516 272944 532568 272950
rect 532516 272886 532568 272892
rect 532344 270286 532464 270314
rect 530780 270150 531360 270178
rect 532238 270192 532294 270201
rect 530780 270094 530808 270150
rect 532238 270127 532294 270136
rect 530768 270088 530820 270094
rect 530768 270030 530820 270036
rect 530952 270088 531004 270094
rect 530952 270030 531004 270036
rect 529848 266756 529900 266762
rect 529848 266698 529900 266704
rect 530964 264330 530992 270030
rect 532252 269822 532280 270127
rect 532240 269816 532292 269822
rect 532240 269758 532292 269764
rect 531412 266756 531464 266762
rect 531412 266698 531464 266704
rect 529676 264302 529782 264330
rect 530610 264302 530992 264330
rect 531424 264316 531452 266698
rect 532436 264330 532464 270286
rect 532528 267734 532556 272886
rect 532712 272542 532740 278052
rect 533908 274786 533936 278052
rect 534092 278038 535118 278066
rect 535748 278038 536314 278066
rect 533896 274780 533948 274786
rect 533896 274722 533948 274728
rect 532884 272808 532936 272814
rect 532884 272750 532936 272756
rect 533712 272808 533764 272814
rect 533712 272750 533764 272756
rect 532896 272542 532924 272750
rect 532700 272536 532752 272542
rect 532700 272478 532752 272484
rect 532884 272536 532936 272542
rect 532884 272478 532936 272484
rect 532988 270558 533384 270586
rect 532792 270496 532844 270502
rect 532792 270438 532844 270444
rect 532804 269686 532832 270438
rect 532988 270094 533016 270558
rect 533356 270450 533384 270558
rect 533356 270422 533568 270450
rect 533540 270366 533568 270422
rect 533528 270360 533580 270366
rect 533528 270302 533580 270308
rect 533252 270224 533304 270230
rect 533528 270224 533580 270230
rect 533304 270184 533528 270212
rect 533252 270166 533304 270172
rect 533528 270166 533580 270172
rect 532976 270088 533028 270094
rect 532976 270030 533028 270036
rect 532792 269680 532844 269686
rect 532792 269622 532844 269628
rect 532528 267706 532648 267734
rect 532620 266762 532648 267706
rect 532608 266756 532660 266762
rect 532608 266698 532660 266704
rect 533068 266756 533120 266762
rect 533068 266698 533120 266704
rect 532266 264302 532464 264330
rect 533080 264316 533108 266698
rect 533724 264330 533752 272750
rect 534092 270201 534120 278038
rect 534724 274780 534776 274786
rect 534724 274722 534776 274728
rect 534078 270192 534134 270201
rect 534078 270127 534134 270136
rect 533988 269952 534040 269958
rect 533988 269894 534040 269900
rect 534000 266762 534028 269894
rect 534736 267034 534764 274722
rect 534724 267028 534776 267034
rect 534724 266970 534776 266976
rect 535552 267028 535604 267034
rect 535552 266970 535604 266976
rect 534724 266892 534776 266898
rect 534724 266834 534776 266840
rect 533988 266756 534040 266762
rect 533988 266698 534040 266704
rect 533724 264302 533922 264330
rect 534736 264316 534764 266834
rect 535564 264316 535592 266970
rect 535748 265130 535776 278038
rect 537496 275330 537524 278052
rect 538508 278038 538706 278066
rect 537668 275460 537720 275466
rect 537668 275402 537720 275408
rect 537484 275324 537536 275330
rect 537484 275266 537536 275272
rect 536748 274100 536800 274106
rect 536748 274042 536800 274048
rect 536562 272504 536618 272513
rect 536562 272439 536618 272448
rect 535736 265124 535788 265130
rect 535736 265066 535788 265072
rect 536576 264330 536604 272439
rect 536760 267034 536788 274042
rect 536748 267028 536800 267034
rect 536748 266970 536800 266976
rect 537680 264330 537708 275402
rect 538508 273254 538536 278038
rect 539888 276282 539916 278052
rect 539876 276276 539928 276282
rect 539876 276218 539928 276224
rect 540992 274786 541020 278052
rect 541636 278038 542202 278066
rect 542372 278038 543398 278066
rect 540980 274780 541032 274786
rect 540980 274722 541032 274728
rect 539322 274000 539378 274009
rect 539322 273935 539378 273944
rect 538324 273226 538536 273254
rect 538324 270094 538352 273226
rect 539048 272944 539100 272950
rect 538508 272892 539048 272898
rect 538508 272886 539100 272892
rect 538508 272870 539088 272886
rect 538508 272542 538536 272870
rect 538680 272808 538732 272814
rect 538680 272750 538732 272756
rect 538692 272542 538720 272750
rect 538496 272536 538548 272542
rect 538496 272478 538548 272484
rect 538680 272536 538732 272542
rect 538680 272478 538732 272484
rect 538312 270088 538364 270094
rect 538312 270030 538364 270036
rect 538692 269878 539088 269906
rect 538034 269784 538090 269793
rect 538034 269719 538090 269728
rect 536406 264302 536604 264330
rect 537234 264302 537708 264330
rect 538048 264316 538076 269719
rect 538692 269414 538720 269878
rect 539060 269822 539088 269878
rect 538864 269816 538916 269822
rect 538864 269758 538916 269764
rect 539048 269816 539100 269822
rect 539048 269758 539100 269764
rect 538876 269414 538904 269758
rect 538680 269408 538732 269414
rect 538680 269350 538732 269356
rect 538864 269408 538916 269414
rect 538864 269350 538916 269356
rect 539336 264330 539364 273935
rect 540520 269952 540572 269958
rect 540520 269894 540572 269900
rect 539692 267028 539744 267034
rect 539692 266970 539744 266976
rect 538890 264302 539364 264330
rect 539704 264316 539732 266970
rect 540532 264316 540560 269894
rect 541636 269822 541664 278038
rect 542084 275324 542136 275330
rect 542084 275266 542136 275272
rect 541624 269816 541676 269822
rect 541808 269816 541860 269822
rect 541624 269758 541676 269764
rect 541806 269784 541808 269793
rect 541860 269784 541862 269793
rect 541806 269719 541862 269728
rect 541348 268388 541400 268394
rect 541348 268330 541400 268336
rect 541360 264316 541388 268330
rect 542096 264330 542124 275266
rect 542372 265266 542400 278038
rect 544580 274922 544608 278052
rect 544568 274916 544620 274922
rect 544568 274858 544620 274864
rect 545776 273970 545804 278052
rect 546512 278038 546986 278066
rect 547892 278038 548090 278066
rect 545946 274000 546002 274009
rect 545764 273964 545816 273970
rect 545946 273935 545948 273944
rect 545764 273906 545816 273912
rect 546000 273935 546002 273944
rect 545948 273906 546000 273912
rect 546512 269278 546540 278038
rect 547694 272504 547750 272513
rect 547694 272439 547750 272448
rect 547708 271998 547736 272439
rect 547512 271992 547564 271998
rect 547510 271960 547512 271969
rect 547696 271992 547748 271998
rect 547564 271960 547566 271969
rect 547892 271969 547920 278038
rect 549272 273562 549300 278052
rect 549456 278038 550482 278066
rect 549260 273556 549312 273562
rect 549260 273498 549312 273504
rect 547696 271934 547748 271940
rect 547878 271960 547934 271969
rect 547510 271895 547566 271904
rect 547878 271895 547934 271904
rect 546500 269272 546552 269278
rect 546500 269214 546552 269220
rect 543004 266756 543056 266762
rect 543004 266698 543056 266704
rect 542360 265260 542412 265266
rect 542360 265202 542412 265208
rect 542096 264302 542202 264330
rect 543016 264316 543044 266698
rect 549456 265402 549484 278038
rect 551664 276418 551692 278052
rect 551652 276412 551704 276418
rect 551652 276354 551704 276360
rect 551284 273556 551336 273562
rect 551284 273498 551336 273504
rect 551296 266490 551324 273498
rect 552860 273426 552888 278052
rect 554056 276554 554084 278052
rect 554792 278038 555266 278066
rect 554044 276548 554096 276554
rect 554044 276490 554096 276496
rect 552848 273420 552900 273426
rect 552848 273362 552900 273368
rect 552296 272128 552348 272134
rect 552296 272070 552348 272076
rect 552308 271980 552336 272070
rect 552848 271992 552900 271998
rect 552308 271952 552848 271980
rect 552848 271934 552900 271940
rect 551284 266484 551336 266490
rect 551284 266426 551336 266432
rect 554792 266354 554820 278038
rect 556356 273698 556384 278052
rect 556344 273692 556396 273698
rect 556344 273634 556396 273640
rect 556804 273692 556856 273698
rect 556804 273634 556856 273640
rect 556816 266626 556844 273634
rect 556804 266620 556856 266626
rect 556804 266562 556856 266568
rect 554780 266348 554832 266354
rect 554780 266290 554832 266296
rect 557552 265538 557580 278052
rect 558748 271998 558776 278052
rect 559944 273834 559972 278052
rect 561140 277234 561168 278052
rect 561128 277228 561180 277234
rect 561128 277170 561180 277176
rect 562336 277098 562364 278052
rect 562324 277092 562376 277098
rect 562324 277034 562376 277040
rect 563440 274650 563468 278052
rect 563428 274644 563480 274650
rect 563428 274586 563480 274592
rect 559932 273828 559984 273834
rect 559932 273770 559984 273776
rect 562140 273080 562192 273086
rect 562140 273022 562192 273028
rect 562324 273080 562376 273086
rect 562324 273022 562376 273028
rect 562152 271998 562180 273022
rect 562336 272134 562364 273022
rect 562324 272128 562376 272134
rect 562324 272070 562376 272076
rect 558736 271992 558788 271998
rect 558736 271934 558788 271940
rect 562140 271992 562192 271998
rect 562140 271934 562192 271940
rect 564636 270774 564664 278052
rect 564624 270768 564676 270774
rect 564624 270710 564676 270716
rect 565832 266218 565860 278052
rect 567028 274514 567056 278052
rect 567016 274508 567068 274514
rect 567016 274450 567068 274456
rect 567844 270768 567896 270774
rect 567844 270710 567896 270716
rect 567856 267714 567884 270710
rect 568224 270638 568252 278052
rect 569420 271998 569448 278052
rect 569972 278038 570630 278066
rect 569408 271992 569460 271998
rect 569408 271934 569460 271940
rect 568212 270632 568264 270638
rect 568212 270574 568264 270580
rect 569972 267986 570000 278038
rect 571720 270910 571748 278052
rect 572732 278038 572930 278066
rect 571708 270904 571760 270910
rect 571708 270846 571760 270852
rect 572732 269414 572760 278038
rect 572720 269408 572772 269414
rect 572720 269350 572772 269356
rect 574112 269074 574140 278052
rect 575308 271046 575336 278052
rect 576504 276962 576532 278052
rect 576872 278038 577714 278066
rect 576492 276956 576544 276962
rect 576492 276898 576544 276904
rect 575296 271040 575348 271046
rect 575296 270982 575348 270988
rect 576124 271040 576176 271046
rect 576124 270982 576176 270988
rect 574100 269068 574152 269074
rect 574100 269010 574152 269016
rect 569960 267980 570012 267986
rect 569960 267922 570012 267928
rect 567844 267708 567896 267714
rect 567844 267650 567896 267656
rect 576136 267578 576164 270982
rect 576872 268258 576900 278038
rect 578896 271862 578924 278052
rect 580000 275058 580028 278052
rect 581012 278038 581210 278066
rect 579988 275052 580040 275058
rect 579988 274994 580040 275000
rect 578884 271856 578936 271862
rect 578884 271798 578936 271804
rect 581012 268938 581040 278038
rect 582392 271590 582420 278052
rect 583588 273562 583616 278052
rect 583772 278038 584798 278066
rect 583576 273556 583628 273562
rect 583576 273498 583628 273504
rect 582380 271584 582432 271590
rect 582380 271526 582432 271532
rect 583024 271584 583076 271590
rect 583024 271526 583076 271532
rect 581000 268932 581052 268938
rect 581000 268874 581052 268880
rect 576860 268252 576912 268258
rect 576860 268194 576912 268200
rect 576124 267572 576176 267578
rect 576124 267514 576176 267520
rect 583036 267442 583064 271526
rect 583772 268802 583800 278038
rect 585980 271726 586008 278052
rect 587084 277438 587112 278052
rect 587912 278038 588294 278066
rect 587072 277432 587124 277438
rect 587072 277374 587124 277380
rect 585968 271720 586020 271726
rect 585968 271662 586020 271668
rect 583760 268796 583812 268802
rect 583760 268738 583812 268744
rect 587912 268666 587940 278038
rect 589476 271454 589504 278052
rect 590672 273698 590700 278052
rect 591868 274378 591896 278052
rect 591856 274372 591908 274378
rect 591856 274314 591908 274320
rect 590660 273692 590712 273698
rect 590660 273634 590712 273640
rect 589464 271448 589516 271454
rect 589464 271390 589516 271396
rect 589924 271448 589976 271454
rect 589924 271390 589976 271396
rect 587900 268660 587952 268666
rect 587900 268602 587952 268608
rect 583024 267436 583076 267442
rect 583024 267378 583076 267384
rect 589936 266898 589964 271390
rect 593064 271318 593092 278052
rect 594260 275194 594288 278052
rect 594812 278038 595378 278066
rect 596192 278038 596574 278066
rect 594248 275188 594300 275194
rect 594248 275130 594300 275136
rect 593052 271312 593104 271318
rect 593052 271254 593104 271260
rect 594812 268530 594840 278038
rect 596192 269550 596220 278038
rect 597756 270774 597784 278052
rect 598952 274242 598980 278052
rect 599136 278038 600162 278066
rect 598940 274236 598992 274242
rect 598940 274178 598992 274184
rect 598204 271312 598256 271318
rect 598204 271254 598256 271260
rect 597744 270768 597796 270774
rect 597744 270710 597796 270716
rect 596180 269544 596232 269550
rect 596180 269486 596232 269492
rect 594800 268524 594852 268530
rect 594800 268466 594852 268472
rect 589924 266892 589976 266898
rect 589924 266834 589976 266840
rect 598216 266762 598244 271254
rect 598204 266756 598256 266762
rect 598204 266698 598256 266704
rect 565820 266212 565872 266218
rect 565820 266154 565872 266160
rect 599136 266082 599164 278038
rect 601344 276010 601372 278052
rect 601712 278038 602462 278066
rect 601332 276004 601384 276010
rect 601332 275946 601384 275952
rect 601148 273080 601200 273086
rect 601148 273022 601200 273028
rect 601160 272406 601188 273022
rect 600964 272400 601016 272406
rect 600964 272342 601016 272348
rect 601148 272400 601200 272406
rect 601148 272342 601200 272348
rect 600976 272134 601004 272342
rect 600964 272128 601016 272134
rect 600964 272070 601016 272076
rect 599124 266076 599176 266082
rect 599124 266018 599176 266024
rect 601712 265946 601740 278038
rect 603644 276826 603672 278052
rect 603632 276820 603684 276826
rect 603632 276762 603684 276768
rect 604840 271046 604868 278052
rect 605852 278038 606050 278066
rect 604828 271040 604880 271046
rect 604828 270982 604880 270988
rect 601700 265940 601752 265946
rect 601700 265882 601752 265888
rect 605852 265810 605880 278038
rect 607232 272134 607260 278052
rect 607416 278038 608442 278066
rect 608612 278038 609638 278066
rect 607220 272128 607272 272134
rect 607220 272070 607272 272076
rect 607416 268122 607444 278038
rect 607404 268116 607456 268122
rect 607404 268058 607456 268064
rect 605840 265804 605892 265810
rect 605840 265746 605892 265752
rect 608612 265674 608640 278038
rect 610728 272270 610756 278052
rect 611648 278038 611938 278066
rect 610716 272264 610768 272270
rect 610716 272206 610768 272212
rect 611648 271590 611676 278038
rect 613120 276690 613148 278052
rect 613108 276684 613160 276690
rect 613108 276626 613160 276632
rect 614316 273222 614344 278052
rect 615512 275874 615540 278052
rect 615696 278038 616722 278066
rect 617352 278038 617826 278066
rect 615500 275868 615552 275874
rect 615500 275810 615552 275816
rect 614304 273216 614356 273222
rect 614304 273158 614356 273164
rect 611636 271584 611688 271590
rect 611636 271526 611688 271532
rect 612004 271584 612056 271590
rect 612004 271526 612056 271532
rect 612016 267306 612044 271526
rect 615696 269686 615724 278038
rect 617352 271182 617380 278038
rect 618444 272944 618496 272950
rect 618444 272886 618496 272892
rect 618456 272678 618484 272886
rect 618444 272672 618496 272678
rect 618444 272614 618496 272620
rect 619008 271590 619036 278052
rect 619652 278038 620218 278066
rect 618996 271584 619048 271590
rect 618996 271526 619048 271532
rect 617340 271176 617392 271182
rect 617340 271118 617392 271124
rect 617524 271176 617576 271182
rect 617524 271118 617576 271124
rect 615684 269680 615736 269686
rect 615684 269622 615736 269628
rect 612004 267300 612056 267306
rect 612004 267242 612056 267248
rect 617536 267170 617564 271118
rect 619652 270502 619680 278038
rect 621400 272950 621428 278052
rect 622596 275738 622624 278052
rect 623806 278038 624004 278066
rect 622584 275732 622636 275738
rect 622584 275674 622636 275680
rect 621388 272944 621440 272950
rect 621388 272886 621440 272892
rect 620284 272672 620336 272678
rect 620284 272614 620336 272620
rect 620296 272406 620324 272614
rect 620284 272400 620336 272406
rect 620284 272342 620336 272348
rect 619640 270496 619692 270502
rect 619640 270438 619692 270444
rect 623976 270230 624004 278038
rect 624988 273086 625016 278052
rect 624976 273080 625028 273086
rect 624976 273022 625028 273028
rect 626092 271182 626120 278052
rect 626552 278038 627302 278066
rect 626080 271176 626132 271182
rect 626080 271118 626132 271124
rect 626552 270366 626580 278038
rect 628484 272814 628512 278052
rect 629680 275602 629708 278052
rect 630692 278038 630890 278066
rect 629668 275596 629720 275602
rect 629668 275538 629720 275544
rect 628472 272808 628524 272814
rect 628472 272750 628524 272756
rect 626540 270360 626592 270366
rect 626540 270302 626592 270308
rect 623964 270224 624016 270230
rect 623964 270166 624016 270172
rect 630692 270094 630720 278038
rect 632072 272542 632100 278052
rect 632060 272536 632112 272542
rect 632060 272478 632112 272484
rect 633268 271454 633296 278052
rect 634372 274106 634400 278052
rect 634360 274100 634412 274106
rect 634360 274042 634412 274048
rect 635568 272678 635596 278052
rect 636764 275466 636792 278052
rect 637592 278038 637974 278066
rect 636752 275460 636804 275466
rect 636752 275402 636804 275408
rect 635556 272672 635608 272678
rect 635556 272614 635608 272620
rect 634084 272536 634136 272542
rect 634084 272478 634136 272484
rect 633256 271448 633308 271454
rect 633256 271390 633308 271396
rect 630680 270088 630732 270094
rect 630680 270030 630732 270036
rect 617524 267164 617576 267170
rect 617524 267106 617576 267112
rect 634096 267034 634124 272478
rect 637592 269822 637620 278038
rect 639156 273970 639184 278052
rect 639144 273964 639196 273970
rect 639144 273906 639196 273912
rect 640352 272542 640380 278052
rect 640536 278038 641470 278066
rect 641732 278038 642666 278066
rect 640340 272536 640392 272542
rect 640340 272478 640392 272484
rect 640536 269958 640564 278038
rect 640524 269952 640576 269958
rect 640524 269894 640576 269900
rect 637580 269816 637632 269822
rect 637580 269758 637632 269764
rect 641732 268394 641760 278038
rect 643848 275330 643876 278052
rect 643836 275324 643888 275330
rect 643836 275266 643888 275272
rect 645044 271318 645072 278052
rect 645872 278038 646254 278066
rect 647252 278038 647450 278066
rect 645032 271312 645084 271318
rect 645032 271254 645084 271260
rect 641720 268388 641772 268394
rect 641720 268330 641772 268336
rect 634084 267028 634136 267034
rect 634084 266970 634136 266976
rect 608600 265668 608652 265674
rect 608600 265610 608652 265616
rect 557540 265532 557592 265538
rect 557540 265474 557592 265480
rect 549444 265396 549496 265402
rect 549444 265338 549496 265344
rect 554410 262168 554466 262177
rect 554410 262103 554466 262112
rect 554424 260914 554452 262103
rect 645872 261526 645900 278038
rect 570604 261520 570656 261526
rect 570604 261462 570656 261468
rect 645860 261520 645912 261526
rect 645860 261462 645912 261468
rect 554412 260908 554464 260914
rect 554412 260850 554464 260856
rect 568580 260908 568632 260914
rect 568580 260850 568632 260856
rect 554318 259992 554374 260001
rect 554318 259927 554374 259936
rect 554332 259486 554360 259927
rect 554320 259480 554372 259486
rect 554320 259422 554372 259428
rect 560944 259480 560996 259486
rect 560944 259422 560996 259428
rect 553950 257816 554006 257825
rect 553950 257751 554006 257760
rect 553964 256766 553992 257751
rect 553952 256760 554004 256766
rect 553952 256702 554004 256708
rect 553490 255640 553546 255649
rect 553490 255575 553492 255584
rect 553544 255575 553546 255584
rect 555424 255604 555476 255610
rect 553492 255546 553544 255552
rect 555424 255546 555476 255552
rect 554410 253464 554466 253473
rect 554410 253399 554466 253408
rect 554424 252618 554452 253399
rect 554412 252612 554464 252618
rect 554412 252554 554464 252560
rect 554134 251288 554190 251297
rect 554134 251223 554136 251232
rect 554188 251223 554190 251232
rect 554136 251194 554188 251200
rect 554042 249112 554098 249121
rect 554042 249047 554098 249056
rect 553858 246936 553914 246945
rect 553858 246871 553914 246880
rect 553872 245682 553900 246871
rect 553860 245676 553912 245682
rect 553860 245618 553912 245624
rect 553674 242584 553730 242593
rect 553674 242519 553730 242528
rect 553688 241534 553716 242519
rect 553676 241528 553728 241534
rect 553676 241470 553728 241476
rect 137928 231804 137980 231810
rect 137928 231746 137980 231752
rect 152372 231804 152424 231810
rect 152372 231746 152424 231752
rect 91744 231668 91796 231674
rect 91744 231610 91796 231616
rect 64144 231260 64196 231266
rect 64144 231202 64196 231208
rect 86224 229900 86276 229906
rect 86224 229842 86276 229848
rect 68284 229764 68336 229770
rect 68284 229706 68336 229712
rect 67548 228676 67600 228682
rect 67548 228618 67600 228624
rect 64788 227724 64840 227730
rect 64788 227666 64840 227672
rect 64604 220380 64656 220386
rect 64604 220322 64656 220328
rect 64616 219434 64644 220322
rect 64800 219434 64828 227666
rect 66168 225752 66220 225758
rect 66168 225694 66220 225700
rect 63960 219428 64012 219434
rect 64616 219406 64736 219434
rect 64800 219428 64932 219434
rect 64800 219406 64880 219428
rect 63960 219370 64012 219376
rect 63132 219156 63184 219162
rect 63132 219098 63184 219104
rect 62672 218884 62724 218890
rect 62672 218826 62724 218832
rect 63144 217138 63172 219098
rect 63972 217138 64000 219370
rect 64708 217274 64736 219406
rect 64880 219370 64932 219376
rect 66180 218074 66208 225694
rect 67272 218204 67324 218210
rect 67272 218146 67324 218152
rect 65616 218068 65668 218074
rect 65616 218010 65668 218016
rect 66168 218068 66220 218074
rect 66168 218010 66220 218016
rect 66444 218068 66496 218074
rect 66444 218010 66496 218016
rect 64708 217246 64782 217274
rect 61442 217110 61516 217138
rect 62270 217110 62344 217138
rect 63098 217110 63172 217138
rect 63926 217110 64000 217138
rect 61442 216988 61470 217110
rect 62270 216988 62298 217110
rect 63098 216988 63126 217110
rect 63926 216988 63954 217110
rect 64754 216988 64782 217246
rect 65628 217138 65656 218010
rect 66456 217138 66484 218010
rect 67284 217138 67312 218146
rect 67560 218074 67588 228618
rect 68296 218210 68324 229706
rect 82084 229628 82136 229634
rect 82084 229570 82136 229576
rect 72424 226160 72476 226166
rect 72424 226102 72476 226108
rect 68928 224256 68980 224262
rect 68928 224198 68980 224204
rect 68744 223168 68796 223174
rect 68744 223110 68796 223116
rect 68284 218204 68336 218210
rect 68284 218146 68336 218152
rect 68756 218074 68784 223110
rect 67548 218068 67600 218074
rect 67548 218010 67600 218016
rect 68100 218068 68152 218074
rect 68100 218010 68152 218016
rect 68744 218068 68796 218074
rect 68744 218010 68796 218016
rect 68112 217138 68140 218010
rect 68940 217274 68968 224198
rect 71412 222896 71464 222902
rect 71412 222838 71464 222844
rect 69756 219564 69808 219570
rect 69756 219506 69808 219512
rect 69768 217274 69796 219506
rect 70584 219156 70636 219162
rect 70584 219098 70636 219104
rect 65582 217110 65656 217138
rect 66410 217110 66484 217138
rect 67238 217110 67312 217138
rect 68066 217110 68140 217138
rect 68894 217246 68968 217274
rect 69722 217246 69796 217274
rect 65582 216988 65610 217110
rect 66410 216988 66438 217110
rect 67238 216988 67266 217110
rect 68066 216988 68094 217110
rect 68894 216988 68922 217246
rect 69722 216988 69750 217246
rect 70596 217138 70624 219098
rect 71424 217274 71452 222838
rect 72436 219026 72464 226102
rect 76564 225888 76616 225894
rect 76564 225830 76616 225836
rect 73712 224392 73764 224398
rect 73712 224334 73764 224340
rect 73068 220244 73120 220250
rect 73068 220186 73120 220192
rect 72424 219020 72476 219026
rect 72424 218962 72476 218968
rect 72240 218068 72292 218074
rect 72240 218010 72292 218016
rect 70550 217110 70624 217138
rect 71378 217246 71452 217274
rect 70550 216988 70578 217110
rect 71378 216988 71406 217246
rect 72252 217138 72280 218010
rect 73080 217274 73108 220186
rect 73724 218074 73752 224334
rect 75828 223032 75880 223038
rect 75828 222974 75880 222980
rect 73896 221604 73948 221610
rect 73896 221546 73948 221552
rect 73712 218068 73764 218074
rect 73712 218010 73764 218016
rect 73908 217274 73936 221546
rect 75552 218204 75604 218210
rect 75552 218146 75604 218152
rect 74724 218068 74776 218074
rect 74724 218010 74776 218016
rect 72206 217110 72280 217138
rect 73034 217246 73108 217274
rect 73862 217246 73936 217274
rect 72206 216988 72234 217110
rect 73034 216988 73062 217246
rect 73862 216988 73890 217246
rect 74736 217138 74764 218010
rect 75564 217138 75592 218146
rect 75840 218074 75868 222974
rect 76380 220516 76432 220522
rect 76380 220458 76432 220464
rect 75828 218068 75880 218074
rect 75828 218010 75880 218016
rect 76392 217274 76420 220458
rect 76576 218210 76604 225830
rect 79968 224528 80020 224534
rect 79968 224470 80020 224476
rect 78588 222760 78640 222766
rect 78588 222702 78640 222708
rect 77208 219020 77260 219026
rect 77208 218962 77260 218968
rect 76564 218204 76616 218210
rect 76564 218146 76616 218152
rect 74690 217110 74764 217138
rect 75518 217110 75592 217138
rect 76346 217246 76420 217274
rect 74690 216988 74718 217110
rect 75518 216988 75546 217110
rect 76346 216988 76374 217246
rect 77220 217138 77248 218962
rect 78600 218074 78628 222702
rect 79692 220652 79744 220658
rect 79692 220594 79744 220600
rect 78036 218068 78088 218074
rect 78036 218010 78088 218016
rect 78588 218068 78640 218074
rect 78588 218010 78640 218016
rect 78864 218068 78916 218074
rect 78864 218010 78916 218016
rect 78048 217138 78076 218010
rect 78876 217138 78904 218010
rect 79704 217274 79732 220594
rect 79980 218074 80008 224470
rect 81348 223304 81400 223310
rect 81348 223246 81400 223252
rect 80520 220856 80572 220862
rect 80520 220798 80572 220804
rect 79968 218068 80020 218074
rect 79968 218010 80020 218016
rect 80532 217274 80560 220798
rect 81360 217274 81388 223246
rect 82096 221610 82124 229570
rect 86236 229094 86264 229842
rect 86144 229066 86264 229094
rect 83464 226024 83516 226030
rect 83464 225966 83516 225972
rect 82084 221604 82136 221610
rect 82084 221546 82136 221552
rect 83004 220992 83056 220998
rect 83004 220934 83056 220940
rect 82176 218068 82228 218074
rect 82176 218010 82228 218016
rect 77174 217110 77248 217138
rect 78002 217110 78076 217138
rect 78830 217110 78904 217138
rect 79658 217246 79732 217274
rect 80486 217246 80560 217274
rect 81314 217246 81388 217274
rect 77174 216988 77202 217110
rect 78002 216988 78030 217110
rect 78830 216988 78858 217110
rect 79658 216988 79686 217246
rect 80486 216988 80514 217246
rect 81314 216988 81342 217246
rect 82188 217138 82216 218010
rect 83016 217274 83044 220934
rect 83476 218074 83504 225966
rect 85488 224664 85540 224670
rect 85488 224606 85540 224612
rect 85304 222624 85356 222630
rect 85304 222566 85356 222572
rect 83832 218884 83884 218890
rect 83832 218826 83884 218832
rect 83464 218068 83516 218074
rect 83464 218010 83516 218016
rect 82142 217110 82216 217138
rect 82970 217246 83044 217274
rect 82142 216988 82170 217110
rect 82970 216988 82998 217246
rect 83844 217138 83872 218826
rect 85316 218074 85344 222566
rect 84660 218068 84712 218074
rect 84660 218010 84712 218016
rect 85304 218068 85356 218074
rect 85304 218010 85356 218016
rect 84672 217138 84700 218010
rect 85500 217274 85528 224606
rect 86144 220862 86172 229066
rect 88248 227860 88300 227866
rect 88248 227802 88300 227808
rect 87972 223576 88024 223582
rect 87972 223518 88024 223524
rect 86316 221604 86368 221610
rect 86316 221546 86368 221552
rect 86132 220856 86184 220862
rect 86132 220798 86184 220804
rect 86328 217274 86356 221546
rect 87144 218068 87196 218074
rect 87144 218010 87196 218016
rect 83798 217110 83872 217138
rect 84626 217110 84700 217138
rect 85454 217246 85528 217274
rect 86282 217246 86356 217274
rect 83798 216988 83826 217110
rect 84626 216988 84654 217110
rect 85454 216988 85482 217246
rect 86282 216988 86310 217246
rect 87156 217138 87184 218010
rect 87984 217274 88012 223518
rect 88260 218074 88288 227802
rect 89628 227180 89680 227186
rect 89628 227122 89680 227128
rect 89444 224800 89496 224806
rect 89444 224742 89496 224748
rect 89456 218074 89484 224742
rect 88248 218068 88300 218074
rect 88248 218010 88300 218016
rect 88800 218068 88852 218074
rect 88800 218010 88852 218016
rect 89444 218068 89496 218074
rect 89444 218010 89496 218016
rect 87110 217110 87184 217138
rect 87938 217246 88012 217274
rect 87110 216988 87138 217110
rect 87938 216988 87966 217246
rect 88812 217138 88840 218010
rect 89640 217274 89668 227122
rect 91284 222012 91336 222018
rect 91284 221954 91336 221960
rect 90456 218068 90508 218074
rect 90456 218010 90508 218016
rect 88766 217110 88840 217138
rect 89594 217246 89668 217274
rect 88766 216988 88794 217110
rect 89594 216988 89622 217246
rect 90468 217138 90496 218010
rect 91296 217274 91324 221954
rect 91756 218074 91784 231610
rect 128268 231532 128320 231538
rect 128268 231474 128320 231480
rect 97908 230920 97960 230926
rect 97908 230862 97960 230868
rect 95240 230172 95292 230178
rect 95240 230114 95292 230120
rect 93768 228812 93820 228818
rect 93768 228754 93820 228760
rect 93780 218074 93808 228754
rect 95252 227866 95280 230114
rect 95240 227860 95292 227866
rect 95240 227802 95292 227808
rect 96436 227316 96488 227322
rect 96436 227258 96488 227264
rect 96252 224936 96304 224942
rect 96252 224878 96304 224884
rect 94596 221876 94648 221882
rect 94596 221818 94648 221824
rect 91744 218068 91796 218074
rect 91744 218010 91796 218016
rect 92940 218068 92992 218074
rect 92940 218010 92992 218016
rect 93768 218068 93820 218074
rect 93768 218010 93820 218016
rect 92112 217456 92164 217462
rect 92112 217398 92164 217404
rect 90422 217110 90496 217138
rect 91250 217246 91324 217274
rect 90422 216988 90450 217110
rect 91250 216988 91278 217246
rect 92124 217138 92152 217398
rect 92952 217138 92980 218010
rect 93768 217320 93820 217326
rect 94608 217308 94636 221818
rect 96264 218074 96292 224878
rect 95424 218068 95476 218074
rect 95424 218010 95476 218016
rect 96252 218068 96304 218074
rect 96252 218010 96304 218016
rect 93768 217262 93820 217268
rect 94562 217280 94636 217308
rect 93780 217138 93808 217262
rect 92078 217110 92152 217138
rect 92906 217110 92980 217138
rect 93734 217110 93808 217138
rect 92078 216988 92106 217110
rect 92906 216988 92934 217110
rect 93734 216988 93762 217110
rect 94562 216988 94590 217280
rect 95436 217138 95464 218010
rect 96448 217138 96476 227258
rect 97724 221740 97776 221746
rect 97724 221682 97776 221688
rect 97736 219434 97764 221682
rect 97736 219406 97856 219434
rect 97080 218068 97132 218074
rect 97080 218010 97132 218016
rect 97092 217138 97120 218010
rect 97828 217308 97856 219406
rect 97920 218090 97948 230862
rect 110328 230784 110380 230790
rect 110328 230726 110380 230732
rect 102140 229492 102192 229498
rect 102140 229434 102192 229440
rect 100668 229084 100720 229090
rect 100668 229026 100720 229032
rect 99288 223440 99340 223446
rect 99288 223382 99340 223388
rect 97920 218074 98040 218090
rect 99300 218074 99328 223382
rect 100392 218612 100444 218618
rect 100392 218554 100444 218560
rect 97920 218068 98052 218074
rect 97920 218062 98000 218068
rect 98000 218010 98052 218016
rect 98736 218068 98788 218074
rect 98736 218010 98788 218016
rect 99288 218068 99340 218074
rect 99288 218010 99340 218016
rect 99564 218068 99616 218074
rect 99564 218010 99616 218016
rect 97828 217280 97902 217308
rect 95390 217110 95464 217138
rect 96218 217110 96476 217138
rect 97046 217110 97120 217138
rect 95390 216988 95418 217110
rect 96218 216988 96246 217110
rect 97046 216988 97074 217110
rect 97874 216988 97902 217280
rect 98748 217138 98776 218010
rect 99576 217138 99604 218010
rect 100404 217138 100432 218554
rect 100680 218074 100708 229026
rect 102152 227458 102180 229434
rect 106188 229084 106240 229090
rect 106188 229026 106240 229032
rect 102140 227452 102192 227458
rect 102140 227394 102192 227400
rect 103428 227452 103480 227458
rect 103428 227394 103480 227400
rect 102048 224120 102100 224126
rect 102048 224062 102100 224068
rect 101220 220108 101272 220114
rect 101220 220050 101272 220056
rect 100668 218068 100720 218074
rect 100668 218010 100720 218016
rect 101232 217308 101260 220050
rect 102060 217308 102088 224062
rect 103440 218074 103468 227394
rect 106004 223984 106056 223990
rect 106004 223926 106056 223932
rect 104532 221332 104584 221338
rect 104532 221274 104584 221280
rect 102876 218068 102928 218074
rect 102876 218010 102928 218016
rect 103428 218068 103480 218074
rect 103428 218010 103480 218016
rect 98702 217110 98776 217138
rect 99530 217110 99604 217138
rect 100358 217110 100432 217138
rect 101186 217280 101260 217308
rect 102014 217280 102088 217308
rect 98702 216988 98730 217110
rect 99530 216988 99558 217110
rect 100358 216988 100386 217110
rect 101186 216988 101214 217280
rect 102014 216988 102042 217280
rect 102888 217138 102916 218010
rect 103704 217592 103756 217598
rect 103704 217534 103756 217540
rect 103716 217138 103744 217534
rect 104544 217274 104572 221274
rect 105820 219446 105872 219452
rect 105820 219388 105872 219394
rect 105832 218618 105860 219388
rect 105820 218612 105872 218618
rect 105820 218554 105872 218560
rect 106016 218074 106044 223926
rect 105360 218068 105412 218074
rect 105360 218010 105412 218016
rect 106004 218068 106056 218074
rect 106004 218010 106056 218016
rect 102842 217110 102916 217138
rect 103670 217110 103744 217138
rect 104498 217246 104572 217274
rect 102842 216988 102870 217110
rect 103670 216988 103698 217110
rect 104498 216988 104526 217246
rect 105372 217138 105400 218010
rect 106200 217274 106228 229026
rect 110144 227588 110196 227594
rect 110144 227530 110196 227536
rect 106924 226500 106976 226506
rect 106924 226442 106976 226448
rect 106936 219298 106964 226442
rect 108672 223848 108724 223854
rect 108672 223790 108724 223796
rect 107844 220788 107896 220794
rect 107844 220730 107896 220736
rect 106924 219292 106976 219298
rect 106924 219234 106976 219240
rect 107016 218612 107068 218618
rect 107016 218554 107068 218560
rect 105326 217110 105400 217138
rect 106154 217246 106228 217274
rect 105326 216988 105354 217110
rect 106154 216988 106182 217246
rect 107028 217138 107056 218554
rect 107856 217274 107884 220730
rect 108684 217274 108712 223790
rect 110156 218074 110184 227530
rect 109500 218068 109552 218074
rect 109500 218010 109552 218016
rect 110144 218068 110196 218074
rect 110144 218010 110196 218016
rect 106982 217110 107056 217138
rect 107810 217246 107884 217274
rect 108638 217246 108712 217274
rect 106982 216988 107010 217110
rect 107810 216988 107838 217246
rect 108638 216988 108666 217246
rect 109512 217138 109540 218010
rect 110340 217274 110368 230726
rect 118608 230648 118660 230654
rect 118608 230590 118660 230596
rect 111064 229356 111116 229362
rect 111064 229298 111116 229304
rect 111076 227730 111104 229298
rect 112812 228268 112864 228274
rect 112812 228210 112864 228216
rect 111064 227724 111116 227730
rect 111064 227666 111116 227672
rect 111984 222148 112036 222154
rect 111984 222090 112036 222096
rect 111156 221196 111208 221202
rect 111156 221138 111208 221144
rect 111168 217274 111196 221138
rect 111996 217274 112024 222090
rect 112824 217274 112852 228210
rect 117228 227724 117280 227730
rect 117228 227666 117280 227672
rect 115296 223712 115348 223718
rect 115296 223654 115348 223660
rect 114468 219972 114520 219978
rect 114468 219914 114520 219920
rect 113640 219292 113692 219298
rect 113640 219234 113692 219240
rect 109466 217110 109540 217138
rect 110294 217246 110368 217274
rect 111122 217246 111196 217274
rect 111950 217246 112024 217274
rect 112778 217246 112852 217274
rect 109466 216988 109494 217110
rect 110294 216988 110322 217246
rect 111122 216988 111150 217246
rect 111950 216988 111978 217246
rect 112778 216988 112806 217246
rect 113652 217138 113680 219234
rect 114480 217274 114508 219914
rect 115308 217274 115336 223654
rect 117240 218074 117268 227666
rect 118424 222488 118476 222494
rect 118424 222430 118476 222436
rect 118436 219434 118464 222430
rect 118436 219406 118556 219434
rect 117964 219156 118016 219162
rect 117964 219098 118016 219104
rect 117976 218346 118004 219098
rect 117964 218340 118016 218346
rect 117964 218282 118016 218288
rect 116124 218068 116176 218074
rect 116124 218010 116176 218016
rect 117228 218068 117280 218074
rect 117228 218010 117280 218016
rect 117780 218068 117832 218074
rect 117780 218010 117832 218016
rect 113606 217110 113680 217138
rect 114434 217246 114508 217274
rect 115262 217246 115336 217274
rect 113606 216988 113634 217110
rect 114434 216988 114462 217246
rect 115262 216988 115290 217246
rect 116136 217138 116164 218010
rect 116952 217728 117004 217734
rect 116952 217670 117004 217676
rect 116964 217138 116992 217670
rect 117792 217138 117820 218010
rect 118528 217274 118556 219406
rect 118620 218090 118648 230590
rect 126888 230036 126940 230042
rect 126888 229978 126940 229984
rect 123484 229220 123536 229226
rect 123484 229162 123536 229168
rect 119988 228132 120040 228138
rect 119988 228074 120040 228080
rect 118620 218074 118740 218090
rect 120000 218074 120028 228074
rect 122748 226908 122800 226914
rect 122748 226850 122800 226856
rect 122564 226296 122616 226302
rect 122564 226238 122616 226244
rect 121092 219836 121144 219842
rect 121092 219778 121144 219784
rect 120264 218476 120316 218482
rect 120264 218418 120316 218424
rect 118620 218068 118752 218074
rect 118620 218062 118700 218068
rect 118700 218010 118752 218016
rect 119436 218068 119488 218074
rect 119436 218010 119488 218016
rect 119988 218068 120040 218074
rect 119988 218010 120040 218016
rect 118528 217246 118602 217274
rect 116090 217110 116164 217138
rect 116918 217110 116992 217138
rect 117746 217110 117820 217138
rect 116090 216988 116118 217110
rect 116918 216988 116946 217110
rect 117746 216988 117774 217110
rect 118574 216988 118602 217246
rect 119448 217138 119476 218010
rect 120276 217138 120304 218418
rect 121104 217274 121132 219778
rect 122576 218074 122604 226238
rect 121920 218068 121972 218074
rect 121920 218010 121972 218016
rect 122564 218068 122616 218074
rect 122564 218010 122616 218016
rect 119402 217110 119476 217138
rect 120230 217110 120304 217138
rect 121058 217246 121132 217274
rect 119402 216988 119430 217110
rect 120230 216988 120258 217110
rect 121058 216988 121086 217246
rect 121932 217138 121960 218010
rect 122760 217274 122788 226850
rect 123496 218346 123524 229162
rect 126704 227996 126756 228002
rect 126704 227938 126756 227944
rect 125232 225480 125284 225486
rect 125232 225422 125284 225428
rect 124404 221060 124456 221066
rect 124404 221002 124456 221008
rect 123484 218340 123536 218346
rect 123484 218282 123536 218288
rect 123576 218204 123628 218210
rect 123576 218146 123628 218152
rect 121886 217110 121960 217138
rect 122714 217246 122788 217274
rect 121886 216988 121914 217110
rect 122714 216988 122742 217246
rect 123588 217138 123616 218146
rect 124416 217274 124444 221002
rect 125244 217274 125272 225422
rect 126716 218074 126744 227938
rect 126060 218068 126112 218074
rect 126060 218010 126112 218016
rect 126704 218068 126756 218074
rect 126704 218010 126756 218016
rect 123542 217110 123616 217138
rect 124370 217246 124444 217274
rect 125198 217246 125272 217274
rect 123542 216988 123570 217110
rect 124370 216988 124398 217246
rect 125198 216988 125226 217246
rect 126072 217138 126100 218010
rect 126900 217274 126928 229978
rect 127624 222760 127676 222766
rect 127624 222702 127676 222708
rect 127808 222760 127860 222766
rect 127808 222702 127860 222708
rect 127636 222494 127664 222702
rect 127624 222488 127676 222494
rect 127624 222430 127676 222436
rect 127820 222358 127848 222702
rect 127808 222352 127860 222358
rect 127808 222294 127860 222300
rect 128280 218074 128308 231474
rect 130384 230444 130436 230450
rect 130384 230386 130436 230392
rect 129556 226772 129608 226778
rect 129556 226714 129608 226720
rect 129372 225344 129424 225350
rect 129372 225286 129424 225292
rect 129384 218074 129412 225286
rect 127716 218068 127768 218074
rect 127716 218010 127768 218016
rect 128268 218068 128320 218074
rect 128268 218010 128320 218016
rect 128544 218068 128596 218074
rect 128544 218010 128596 218016
rect 129372 218068 129424 218074
rect 129372 218010 129424 218016
rect 126026 217110 126100 217138
rect 126854 217246 126928 217274
rect 126026 216988 126054 217110
rect 126854 216988 126882 217246
rect 127728 217138 127756 218010
rect 128556 217138 128584 218010
rect 129568 217274 129596 226714
rect 130396 225214 130424 230386
rect 133788 230308 133840 230314
rect 133788 230250 133840 230256
rect 133512 227860 133564 227866
rect 133512 227802 133564 227808
rect 130384 225208 130436 225214
rect 130384 225150 130436 225156
rect 132408 225208 132460 225214
rect 132408 225150 132460 225156
rect 132420 218346 132448 225150
rect 132592 219156 132644 219162
rect 132592 219098 132644 219104
rect 131856 218340 131908 218346
rect 131856 218282 131908 218288
rect 132408 218340 132460 218346
rect 132408 218282 132460 218288
rect 130200 218068 130252 218074
rect 130200 218010 130252 218016
rect 127682 217110 127756 217138
rect 128510 217110 128584 217138
rect 129338 217246 129596 217274
rect 127682 216988 127710 217110
rect 128510 216988 128538 217110
rect 129338 216988 129366 217246
rect 130212 217138 130240 218010
rect 131028 217864 131080 217870
rect 131028 217806 131080 217812
rect 131040 217138 131068 217806
rect 131868 217138 131896 218282
rect 132604 218226 132632 219098
rect 132512 218198 132632 218226
rect 132512 218074 132540 218198
rect 133524 218074 133552 227802
rect 133800 219434 133828 230250
rect 136548 226636 136600 226642
rect 136548 226578 136600 226584
rect 135168 225072 135220 225078
rect 135168 225014 135220 225020
rect 134340 219836 134392 219842
rect 134340 219778 134392 219784
rect 133708 219406 133828 219434
rect 132500 218068 132552 218074
rect 132500 218010 132552 218016
rect 132684 218068 132736 218074
rect 132684 218010 132736 218016
rect 133512 218068 133564 218074
rect 133512 218010 133564 218016
rect 132696 217138 132724 218010
rect 133708 217274 133736 219406
rect 134352 217274 134380 219778
rect 135180 217274 135208 225014
rect 136560 218074 136588 226578
rect 137940 219434 137968 231746
rect 139860 229492 139912 229498
rect 139860 229434 139912 229440
rect 139872 229378 139900 229434
rect 139872 229362 140360 229378
rect 139872 229356 140372 229362
rect 139872 229350 140320 229356
rect 140320 229298 140372 229304
rect 140042 229256 140098 229265
rect 140042 229191 140098 229200
rect 139306 228712 139362 228721
rect 139306 228647 139362 228656
rect 139124 222352 139176 222358
rect 139124 222294 139176 222300
rect 137664 219406 137968 219434
rect 136824 218340 136876 218346
rect 136824 218282 136876 218288
rect 135996 218068 136048 218074
rect 135996 218010 136048 218016
rect 136548 218068 136600 218074
rect 136548 218010 136600 218016
rect 130166 217110 130240 217138
rect 130994 217110 131068 217138
rect 131822 217110 131896 217138
rect 132650 217110 132724 217138
rect 133478 217246 133736 217274
rect 134306 217246 134380 217274
rect 135134 217246 135208 217274
rect 130166 216988 130194 217110
rect 130994 216988 131022 217110
rect 131822 216988 131850 217110
rect 132650 216988 132678 217110
rect 133478 216988 133506 217246
rect 134306 216988 134334 217246
rect 135134 216988 135162 217246
rect 136008 217138 136036 218010
rect 136836 217138 136864 218282
rect 137664 217274 137692 219406
rect 139136 218074 139164 222294
rect 138480 218068 138532 218074
rect 138480 218010 138532 218016
rect 139124 218068 139176 218074
rect 139124 218010 139176 218016
rect 135962 217110 136036 217138
rect 136790 217110 136864 217138
rect 137618 217246 137692 217274
rect 135962 216988 135990 217110
rect 136790 216988 136818 217110
rect 137618 216988 137646 217246
rect 138492 217138 138520 218010
rect 139320 217274 139348 228647
rect 140056 219026 140084 229191
rect 141160 228410 141188 231676
rect 141344 231662 141818 231690
rect 142172 231662 142462 231690
rect 142632 231662 143106 231690
rect 141148 228404 141200 228410
rect 141148 228346 141200 228352
rect 141148 226160 141200 226166
rect 141146 226128 141148 226137
rect 141200 226128 141202 226137
rect 141146 226063 141202 226072
rect 141344 221474 141372 231662
rect 142172 227050 142200 231662
rect 142632 230602 142660 231662
rect 142448 230574 142660 230602
rect 142448 228546 142476 230574
rect 142618 230480 142674 230489
rect 142618 230415 142620 230424
rect 142672 230415 142674 230424
rect 142804 230444 142856 230450
rect 142620 230386 142672 230392
rect 142804 230386 142856 230392
rect 142816 229770 142844 230386
rect 142804 229764 142856 229770
rect 142804 229706 142856 229712
rect 142988 229764 143040 229770
rect 142988 229706 143040 229712
rect 143000 229362 143028 229706
rect 142988 229356 143040 229362
rect 142988 229298 143040 229304
rect 142988 229084 143040 229090
rect 142988 229026 143040 229032
rect 143448 229084 143500 229090
rect 143448 229026 143500 229032
rect 143000 228682 143028 229026
rect 142988 228676 143040 228682
rect 142988 228618 143040 228624
rect 142436 228540 142488 228546
rect 142436 228482 142488 228488
rect 142160 227044 142212 227050
rect 142160 226986 142212 226992
rect 143264 227044 143316 227050
rect 143264 226986 143316 226992
rect 141516 226160 141568 226166
rect 141516 226102 141568 226108
rect 141528 225622 141556 226102
rect 141516 225616 141568 225622
rect 141516 225558 141568 225564
rect 141792 225616 141844 225622
rect 141792 225558 141844 225564
rect 141332 221468 141384 221474
rect 141332 221410 141384 221416
rect 140778 219872 140834 219881
rect 140778 219807 140780 219816
rect 140832 219807 140834 219816
rect 140964 219836 141016 219842
rect 140780 219778 140832 219784
rect 140964 219778 141016 219784
rect 140044 219020 140096 219026
rect 140044 218962 140096 218968
rect 139492 218340 139544 218346
rect 139492 218282 139544 218288
rect 140136 218340 140188 218346
rect 140136 218282 140188 218288
rect 139504 218074 139532 218282
rect 139492 218068 139544 218074
rect 139492 218010 139544 218016
rect 138446 217110 138520 217138
rect 139274 217246 139348 217274
rect 138446 216988 138474 217110
rect 139274 216988 139302 217246
rect 140148 217138 140176 218282
rect 140976 217274 141004 219778
rect 141804 217274 141832 225558
rect 141974 220416 142030 220425
rect 141974 220351 141976 220360
rect 142028 220351 142030 220360
rect 141976 220322 142028 220328
rect 141988 220238 142384 220266
rect 141988 219842 142016 220238
rect 142158 219872 142214 219881
rect 141976 219836 142028 219842
rect 142158 219807 142160 219816
rect 141976 219778 142028 219784
rect 142212 219807 142214 219816
rect 142160 219778 142212 219784
rect 142158 219600 142214 219609
rect 142356 219570 142384 220238
rect 142158 219535 142160 219544
rect 142212 219535 142214 219544
rect 142344 219564 142396 219570
rect 142160 219506 142212 219512
rect 142344 219506 142396 219512
rect 142436 219020 142488 219026
rect 142436 218962 142488 218968
rect 142448 218754 142476 218962
rect 143276 218754 143304 226986
rect 142436 218748 142488 218754
rect 142436 218690 142488 218696
rect 142620 218748 142672 218754
rect 142620 218690 142672 218696
rect 143264 218748 143316 218754
rect 143264 218690 143316 218696
rect 140102 217110 140176 217138
rect 140930 217246 141004 217274
rect 141758 217246 141832 217274
rect 140102 216988 140130 217110
rect 140930 216988 140958 217246
rect 141758 216988 141786 217246
rect 142632 217138 142660 218690
rect 143460 217274 143488 229026
rect 143736 219026 143764 231676
rect 144104 231662 144394 231690
rect 144104 230489 144132 231662
rect 144090 230480 144146 230489
rect 144090 230415 144146 230424
rect 144184 229356 144236 229362
rect 144184 229298 144236 229304
rect 144196 220425 144224 229298
rect 145024 226166 145052 231676
rect 145668 229770 145696 231676
rect 145656 229764 145708 229770
rect 145656 229706 145708 229712
rect 145840 229764 145892 229770
rect 145840 229706 145892 229712
rect 145852 229265 145880 229706
rect 145838 229256 145894 229265
rect 145838 229191 145894 229200
rect 146116 228540 146168 228546
rect 146116 228482 146168 228488
rect 145012 226160 145064 226166
rect 145196 226160 145248 226166
rect 145012 226102 145064 226108
rect 145194 226128 145196 226137
rect 145248 226128 145250 226137
rect 145194 226063 145250 226072
rect 145930 222320 145986 222329
rect 145930 222255 145986 222264
rect 144182 220416 144238 220425
rect 144182 220351 144238 220360
rect 144276 220244 144328 220250
rect 144276 220186 144328 220192
rect 143724 219020 143776 219026
rect 143724 218962 143776 218968
rect 144288 217274 144316 220186
rect 145944 218754 145972 222255
rect 145104 218748 145156 218754
rect 145104 218690 145156 218696
rect 145932 218748 145984 218754
rect 145932 218690 145984 218696
rect 142586 217110 142660 217138
rect 143414 217246 143488 217274
rect 144242 217246 144316 217274
rect 142586 216988 142614 217110
rect 143414 216988 143442 217246
rect 144242 216988 144270 217246
rect 145116 217138 145144 218690
rect 146128 217274 146156 228482
rect 146312 226506 146340 231676
rect 146956 229362 146984 231676
rect 147508 231662 147614 231690
rect 147968 231662 148258 231690
rect 146944 229356 146996 229362
rect 146944 229298 146996 229304
rect 147126 229256 147182 229265
rect 147126 229191 147182 229200
rect 147140 229090 147168 229191
rect 147128 229084 147180 229090
rect 147128 229026 147180 229032
rect 147312 229084 147364 229090
rect 147312 229026 147364 229032
rect 146482 228984 146538 228993
rect 146482 228919 146538 228928
rect 146300 226500 146352 226506
rect 146300 226442 146352 226448
rect 146496 223174 146524 228919
rect 147324 228721 147352 229026
rect 147310 228712 147366 228721
rect 147310 228647 147366 228656
rect 147508 226166 147536 231662
rect 147968 229378 147996 231662
rect 147876 229362 147996 229378
rect 147864 229356 147996 229362
rect 147916 229350 147996 229356
rect 147864 229298 147916 229304
rect 148888 228410 148916 231676
rect 149256 231662 149546 231690
rect 149808 231662 150190 231690
rect 149060 229628 149112 229634
rect 149060 229570 149112 229576
rect 149072 229226 149100 229570
rect 149060 229220 149112 229226
rect 149060 229162 149112 229168
rect 149256 228993 149284 231662
rect 149612 229492 149664 229498
rect 149612 229434 149664 229440
rect 149624 229226 149652 229434
rect 149612 229220 149664 229226
rect 149612 229162 149664 229168
rect 149242 228984 149298 228993
rect 149242 228919 149298 228928
rect 148876 228404 148928 228410
rect 148876 228346 148928 228352
rect 147496 226160 147548 226166
rect 147496 226102 147548 226108
rect 148968 226160 149020 226166
rect 148968 226102 149020 226108
rect 146484 223168 146536 223174
rect 146484 223110 146536 223116
rect 146668 223168 146720 223174
rect 146668 223110 146720 223116
rect 146680 222494 146708 223110
rect 147310 223000 147366 223009
rect 147310 222935 147366 222944
rect 146668 222488 146720 222494
rect 146668 222430 146720 222436
rect 147128 222352 147180 222358
rect 147126 222320 147128 222329
rect 147180 222320 147182 222329
rect 147126 222255 147182 222264
rect 146758 220416 146814 220425
rect 146758 220351 146814 220360
rect 146772 220250 146800 220351
rect 146760 220244 146812 220250
rect 146760 220186 146812 220192
rect 146944 220244 146996 220250
rect 146944 220186 146996 220192
rect 146956 219706 146984 220186
rect 146944 219700 146996 219706
rect 146944 219642 146996 219648
rect 147324 219434 147352 222935
rect 147588 221468 147640 221474
rect 147588 221410 147640 221416
rect 147128 219428 147352 219434
rect 147180 219406 147352 219428
rect 147128 219370 147180 219376
rect 146760 219020 146812 219026
rect 146760 218962 146812 218968
rect 145070 217110 145144 217138
rect 145898 217246 146156 217274
rect 145070 216988 145098 217110
rect 145898 216988 145926 217246
rect 146772 217138 146800 218962
rect 147600 217274 147628 221410
rect 147770 219600 147826 219609
rect 147770 219535 147772 219544
rect 147824 219535 147826 219544
rect 147772 219506 147824 219512
rect 148980 218754 149008 226102
rect 149808 225758 149836 231662
rect 150820 230450 150848 231676
rect 151004 231662 151478 231690
rect 150808 230444 150860 230450
rect 150808 230386 150860 230392
rect 149980 229492 150032 229498
rect 149980 229434 150032 229440
rect 149992 229265 150020 229434
rect 150346 229392 150402 229401
rect 150346 229327 150402 229336
rect 149978 229256 150034 229265
rect 149978 229191 150034 229200
rect 150072 226500 150124 226506
rect 150072 226442 150124 226448
rect 149796 225752 149848 225758
rect 149796 225694 149848 225700
rect 150084 218754 150112 226442
rect 150360 219434 150388 229327
rect 151004 224954 151032 231662
rect 151176 229356 151228 229362
rect 151176 229298 151228 229304
rect 151188 225842 151216 229298
rect 150728 224926 151032 224954
rect 151096 225814 151216 225842
rect 150728 219570 150756 224926
rect 151096 220930 151124 225814
rect 151268 225752 151320 225758
rect 151268 225694 151320 225700
rect 151084 220924 151136 220930
rect 151084 220866 151136 220872
rect 150716 219564 150768 219570
rect 150716 219506 150768 219512
rect 150900 219564 150952 219570
rect 150900 219506 150952 219512
rect 150268 219406 150388 219434
rect 148416 218748 148468 218754
rect 148416 218690 148468 218696
rect 148968 218748 149020 218754
rect 148968 218690 149020 218696
rect 149244 218748 149296 218754
rect 149244 218690 149296 218696
rect 150072 218748 150124 218754
rect 150072 218690 150124 218696
rect 146726 217110 146800 217138
rect 147554 217246 147628 217274
rect 146726 216988 146754 217110
rect 147554 216988 147582 217246
rect 148428 217138 148456 218690
rect 149256 217138 149284 218690
rect 150268 217274 150296 219406
rect 150440 219020 150492 219026
rect 150440 218962 150492 218968
rect 150452 218754 150480 218962
rect 150440 218748 150492 218754
rect 150440 218690 150492 218696
rect 150912 217274 150940 219506
rect 151280 219434 151308 225694
rect 151912 223304 151964 223310
rect 151910 223272 151912 223281
rect 151964 223272 151966 223281
rect 151910 223207 151966 223216
rect 151450 223000 151506 223009
rect 151506 222958 151814 222986
rect 151450 222935 151506 222944
rect 151786 222902 151814 222958
rect 151636 222896 151688 222902
rect 151636 222838 151688 222844
rect 151774 222896 151826 222902
rect 151774 222838 151826 222844
rect 151648 222737 151676 222838
rect 152108 222737 152136 231676
rect 152384 230518 152412 231746
rect 152372 230512 152424 230518
rect 152372 230454 152424 230460
rect 152464 228676 152516 228682
rect 152464 228618 152516 228624
rect 152476 228410 152504 228618
rect 152464 228404 152516 228410
rect 152464 228346 152516 228352
rect 152752 224262 152780 231676
rect 153396 229634 153424 231676
rect 153672 231662 154054 231690
rect 154698 231662 154988 231690
rect 153384 229628 153436 229634
rect 153384 229570 153436 229576
rect 153108 228676 153160 228682
rect 153108 228618 153160 228624
rect 152740 224256 152792 224262
rect 152740 224198 152792 224204
rect 152372 223032 152424 223038
rect 152372 222974 152424 222980
rect 151634 222728 151690 222737
rect 151634 222663 151690 222672
rect 152094 222728 152150 222737
rect 152094 222663 152150 222672
rect 151636 220380 151688 220386
rect 151636 220322 151688 220328
rect 151772 220382 151828 220391
rect 151648 219609 151676 220322
rect 151772 220317 151828 220326
rect 151634 219600 151690 219609
rect 151634 219535 151690 219544
rect 151280 219406 151676 219434
rect 148382 217110 148456 217138
rect 149210 217110 149284 217138
rect 150038 217246 150296 217274
rect 150866 217246 150940 217274
rect 151648 217274 151676 219406
rect 152384 218618 152412 222974
rect 153120 218618 153148 228618
rect 153672 219609 153700 231662
rect 153844 229628 153896 229634
rect 153844 229570 153896 229576
rect 153658 219600 153714 219609
rect 153658 219535 153714 219544
rect 153384 219020 153436 219026
rect 153384 218962 153436 218968
rect 152372 218612 152424 218618
rect 152372 218554 152424 218560
rect 152556 218612 152608 218618
rect 152556 218554 152608 218560
rect 153108 218612 153160 218618
rect 153108 218554 153160 218560
rect 151648 217246 151722 217274
rect 148382 216988 148410 217110
rect 149210 216988 149238 217110
rect 150038 216988 150066 217246
rect 150866 216988 150894 217246
rect 151694 216988 151722 217246
rect 152568 217138 152596 218554
rect 153396 217138 153424 218962
rect 153856 218890 153884 229570
rect 154960 223174 154988 231662
rect 155328 224398 155356 231676
rect 155972 229226 156000 231676
rect 156156 231662 156630 231690
rect 156892 231662 157274 231690
rect 157918 231662 158300 231690
rect 155960 229220 156012 229226
rect 155960 229162 156012 229168
rect 155316 224392 155368 224398
rect 155316 224334 155368 224340
rect 155868 224256 155920 224262
rect 155868 224198 155920 224204
rect 154948 223168 155000 223174
rect 154948 223110 155000 223116
rect 155040 220924 155092 220930
rect 155040 220866 155092 220872
rect 154026 220688 154082 220697
rect 154026 220623 154028 220632
rect 154080 220623 154082 220632
rect 154212 220652 154264 220658
rect 154028 220594 154080 220600
rect 154212 220594 154264 220600
rect 153844 218884 153896 218890
rect 153844 218826 153896 218832
rect 154224 217274 154252 220594
rect 155052 217274 155080 220866
rect 155880 217274 155908 224198
rect 156156 220522 156184 231662
rect 156694 229936 156750 229945
rect 156694 229871 156696 229880
rect 156748 229871 156750 229880
rect 156696 229842 156748 229848
rect 156326 229392 156382 229401
rect 156326 229327 156328 229336
rect 156380 229327 156382 229336
rect 156328 229298 156380 229304
rect 156694 227488 156750 227497
rect 156694 227423 156750 227432
rect 156708 227186 156736 227423
rect 156696 227180 156748 227186
rect 156696 227122 156748 227128
rect 156892 224954 156920 231662
rect 157294 230172 157346 230178
rect 157294 230114 157346 230120
rect 157432 230172 157484 230178
rect 157432 230114 157484 230120
rect 157306 229770 157334 230114
rect 157444 229945 157472 230114
rect 157430 229936 157486 229945
rect 157430 229871 157486 229880
rect 157294 229764 157346 229770
rect 157294 229706 157346 229712
rect 157706 229664 157762 229673
rect 157706 229599 157708 229608
rect 157760 229599 157762 229608
rect 157984 229628 158036 229634
rect 157708 229570 157760 229576
rect 157984 229570 158036 229576
rect 156432 224926 156920 224954
rect 156432 223310 156460 224926
rect 157996 224398 158024 229570
rect 158272 225894 158300 231662
rect 158548 229906 158576 231676
rect 158916 231662 159206 231690
rect 158536 229900 158588 229906
rect 158536 229842 158588 229848
rect 158720 229900 158772 229906
rect 158720 229842 158772 229848
rect 158732 229673 158760 229842
rect 158718 229664 158774 229673
rect 158718 229599 158774 229608
rect 158260 225888 158312 225894
rect 158260 225830 158312 225836
rect 157248 224392 157300 224398
rect 157248 224334 157300 224340
rect 157984 224392 158036 224398
rect 157984 224334 158036 224340
rect 156420 223304 156472 223310
rect 156420 223246 156472 223252
rect 156604 223304 156656 223310
rect 156604 223246 156656 223252
rect 156420 223168 156472 223174
rect 156420 223110 156472 223116
rect 156432 222902 156460 223110
rect 156420 222896 156472 222902
rect 156420 222838 156472 222844
rect 156616 222630 156644 223246
rect 156604 222624 156656 222630
rect 156604 222566 156656 222572
rect 156970 220688 157026 220697
rect 156788 220652 156840 220658
rect 156970 220623 156972 220632
rect 156788 220594 156840 220600
rect 157024 220623 157026 220632
rect 156972 220594 157024 220600
rect 156144 220516 156196 220522
rect 156144 220458 156196 220464
rect 156604 220516 156656 220522
rect 156604 220458 156656 220464
rect 156616 220250 156644 220458
rect 156800 220250 156828 220594
rect 156604 220244 156656 220250
rect 156604 220186 156656 220192
rect 156788 220244 156840 220250
rect 156788 220186 156840 220192
rect 156236 219292 156288 219298
rect 156236 219234 156288 219240
rect 156248 218890 156276 219234
rect 156236 218884 156288 218890
rect 156236 218826 156288 218832
rect 157260 218618 157288 224334
rect 158076 223032 158128 223038
rect 158076 222974 158128 222980
rect 158088 219434 158116 222974
rect 158258 221504 158314 221513
rect 158258 221439 158314 221448
rect 158272 220930 158300 221439
rect 158260 220924 158312 220930
rect 158260 220866 158312 220872
rect 158444 220924 158496 220930
rect 158444 220866 158496 220872
rect 158088 219406 158300 219434
rect 158272 218618 158300 219406
rect 156696 218612 156748 218618
rect 156696 218554 156748 218560
rect 157248 218612 157300 218618
rect 157248 218554 157300 218560
rect 157524 218612 157576 218618
rect 157524 218554 157576 218560
rect 158260 218612 158312 218618
rect 158260 218554 158312 218560
rect 152522 217110 152596 217138
rect 153350 217110 153424 217138
rect 154178 217246 154252 217274
rect 155006 217246 155080 217274
rect 155834 217246 155908 217274
rect 152522 216988 152550 217110
rect 153350 216988 153378 217110
rect 154178 216988 154206 217246
rect 155006 216988 155034 217246
rect 155834 216988 155862 217246
rect 156708 217138 156736 218554
rect 157536 217138 157564 218554
rect 158456 217274 158484 220866
rect 158916 220658 158944 231662
rect 159836 223281 159864 231676
rect 160006 228168 160062 228177
rect 160006 228103 160062 228112
rect 159822 223272 159878 223281
rect 159822 223207 159878 223216
rect 158904 220652 158956 220658
rect 158904 220594 158956 220600
rect 159824 219428 159876 219434
rect 159824 219370 159876 219376
rect 159180 218612 159232 218618
rect 159180 218554 159232 218560
rect 156662 217110 156736 217138
rect 157490 217110 157564 217138
rect 158318 217246 158484 217274
rect 156662 216988 156690 217110
rect 157490 216988 157518 217110
rect 158318 216988 158346 217246
rect 159192 217138 159220 218554
rect 159836 217274 159864 219370
rect 160020 218618 160048 228103
rect 160192 227180 160244 227186
rect 160192 227122 160244 227128
rect 160204 224262 160232 227122
rect 160480 224534 160508 231676
rect 161124 230178 161152 231676
rect 161112 230172 161164 230178
rect 161112 230114 161164 230120
rect 161768 229226 161796 231676
rect 161952 231662 162426 231690
rect 161756 229220 161808 229226
rect 161756 229162 161808 229168
rect 160468 224528 160520 224534
rect 160468 224470 160520 224476
rect 160192 224256 160244 224262
rect 160192 224198 160244 224204
rect 161952 223310 161980 231662
rect 163056 226030 163084 231676
rect 163700 229906 163728 231676
rect 163688 229900 163740 229906
rect 163688 229842 163740 229848
rect 163964 229900 164016 229906
rect 163964 229842 164016 229848
rect 163044 226024 163096 226030
rect 163044 225966 163096 225972
rect 162768 224392 162820 224398
rect 162768 224334 162820 224340
rect 161940 223304 161992 223310
rect 161940 223246 161992 223252
rect 162124 223304 162176 223310
rect 162124 223246 162176 223252
rect 161432 221912 161488 221921
rect 161432 221847 161434 221856
rect 161486 221847 161488 221856
rect 161572 221876 161624 221882
rect 161434 221818 161486 221824
rect 161572 221818 161624 221824
rect 161584 221762 161612 221818
rect 161492 221734 161612 221762
rect 161492 221610 161520 221734
rect 161662 221640 161718 221649
rect 161480 221604 161532 221610
rect 161662 221575 161664 221584
rect 161480 221546 161532 221552
rect 161716 221575 161718 221584
rect 161664 221546 161716 221552
rect 160836 220652 160888 220658
rect 160836 220594 160888 220600
rect 160008 218612 160060 218618
rect 160008 218554 160060 218560
rect 160848 217274 160876 220594
rect 162136 218890 162164 223246
rect 162492 219292 162544 219298
rect 162492 219234 162544 219240
rect 162124 218884 162176 218890
rect 162124 218826 162176 218832
rect 161480 218612 161532 218618
rect 161480 218554 161532 218560
rect 161492 218210 161520 218554
rect 161480 218204 161532 218210
rect 161480 218146 161532 218152
rect 161664 218204 161716 218210
rect 161664 218146 161716 218152
rect 159836 217246 160002 217274
rect 159146 217110 159220 217138
rect 159146 216988 159174 217110
rect 159974 216988 160002 217246
rect 160802 217246 160876 217274
rect 160802 216988 160830 217246
rect 161676 217138 161704 218146
rect 162504 217138 162532 219234
rect 162780 218210 162808 224334
rect 163976 218210 164004 229842
rect 164344 224954 164372 231676
rect 164608 229220 164660 229226
rect 164608 229162 164660 229168
rect 164620 228954 164648 229162
rect 164608 228948 164660 228954
rect 164608 228890 164660 228896
rect 164344 224926 164464 224954
rect 164436 222034 164464 224926
rect 164988 223582 165016 231676
rect 165632 224670 165660 231676
rect 166276 229770 166304 231676
rect 166552 231662 166934 231690
rect 167196 231662 167578 231690
rect 166264 229764 166316 229770
rect 166264 229706 166316 229712
rect 166552 227497 166580 231662
rect 166814 228984 166870 228993
rect 166814 228919 166870 228928
rect 166828 228818 166856 228919
rect 166816 228812 166868 228818
rect 166816 228754 166868 228760
rect 166954 228812 167006 228818
rect 166954 228754 167006 228760
rect 166966 228698 166994 228754
rect 166828 228670 166994 228698
rect 166828 228410 166856 228670
rect 166816 228404 166868 228410
rect 166816 228346 166868 228352
rect 166954 228404 167006 228410
rect 166954 228346 167006 228352
rect 166966 228290 166994 228346
rect 166828 228262 166994 228290
rect 166828 228177 166856 228262
rect 166814 228168 166870 228177
rect 166814 228103 166870 228112
rect 166538 227488 166594 227497
rect 166538 227423 166594 227432
rect 165620 224664 165672 224670
rect 165620 224606 165672 224612
rect 165528 224528 165580 224534
rect 165528 224470 165580 224476
rect 164976 223576 165028 223582
rect 164976 223518 165028 223524
rect 164344 222006 164464 222034
rect 164344 221882 164372 222006
rect 164514 221912 164570 221921
rect 164332 221876 164384 221882
rect 164514 221847 164516 221856
rect 164332 221818 164384 221824
rect 164568 221847 164570 221856
rect 164516 221818 164568 221824
rect 164146 220688 164202 220697
rect 164146 220623 164202 220632
rect 162768 218204 162820 218210
rect 162768 218146 162820 218152
rect 163320 218204 163372 218210
rect 163320 218146 163372 218152
rect 163964 218204 164016 218210
rect 163964 218146 164016 218152
rect 163332 217138 163360 218146
rect 164160 217308 164188 220623
rect 165540 218210 165568 224470
rect 166172 224392 166224 224398
rect 166172 224334 166224 224340
rect 166184 219434 166212 224334
rect 166356 222624 166408 222630
rect 166356 222566 166408 222572
rect 166092 219406 166212 219434
rect 165804 218884 165856 218890
rect 165804 218826 165856 218832
rect 164976 218204 165028 218210
rect 164976 218146 165028 218152
rect 165528 218204 165580 218210
rect 165528 218146 165580 218152
rect 161630 217110 161704 217138
rect 162458 217110 162532 217138
rect 163286 217110 163360 217138
rect 164114 217280 164188 217308
rect 161630 216988 161658 217110
rect 162458 216988 162486 217110
rect 163286 216988 163314 217110
rect 164114 216988 164142 217280
rect 164988 217138 165016 218146
rect 165816 217138 165844 218826
rect 166092 218618 166120 219406
rect 166080 218612 166132 218618
rect 166080 218554 166132 218560
rect 166368 218498 166396 222566
rect 167196 222018 167224 231662
rect 167366 228984 167422 228993
rect 167366 228919 167368 228928
rect 167420 228919 167422 228928
rect 167368 228890 167420 228896
rect 168208 224806 168236 231676
rect 168576 231674 168866 231690
rect 168564 231668 168866 231674
rect 168616 231662 168866 231668
rect 168564 231610 168616 231616
rect 169496 228954 169524 231676
rect 169864 231662 170154 231690
rect 170324 231662 170798 231690
rect 169484 228948 169536 228954
rect 169484 228890 169536 228896
rect 169482 227352 169538 227361
rect 169482 227287 169484 227296
rect 169536 227287 169538 227296
rect 169484 227258 169536 227264
rect 169668 225888 169720 225894
rect 169668 225830 169720 225836
rect 168196 224800 168248 224806
rect 168196 224742 168248 224748
rect 168012 224392 168064 224398
rect 168012 224334 168064 224340
rect 167184 222012 167236 222018
rect 167184 221954 167236 221960
rect 167460 222012 167512 222018
rect 167460 221954 167512 221960
rect 167472 221746 167500 221954
rect 167460 221740 167512 221746
rect 167460 221682 167512 221688
rect 167644 221740 167696 221746
rect 167644 221682 167696 221688
rect 167656 221202 167684 221682
rect 167828 221604 167880 221610
rect 167828 221546 167880 221552
rect 167840 221202 167868 221546
rect 167644 221196 167696 221202
rect 167644 221138 167696 221144
rect 167828 221196 167880 221202
rect 167828 221138 167880 221144
rect 167090 220688 167146 220697
rect 167090 220623 167146 220632
rect 167104 220522 167132 220623
rect 166954 220516 167006 220522
rect 166954 220458 167006 220464
rect 167092 220516 167144 220522
rect 167092 220458 167144 220464
rect 166966 220402 166994 220458
rect 166966 220374 167132 220402
rect 166952 220144 167008 220153
rect 167104 220114 167132 220374
rect 166952 220079 166954 220088
rect 167006 220079 167008 220088
rect 167092 220108 167144 220114
rect 166954 220050 167006 220056
rect 167092 220050 167144 220056
rect 166540 219292 166592 219298
rect 166540 219234 166592 219240
rect 167460 219292 167512 219298
rect 167460 219234 167512 219240
rect 166552 218890 166580 219234
rect 166540 218884 166592 218890
rect 166540 218826 166592 218832
rect 166632 218612 166684 218618
rect 166632 218554 166684 218560
rect 166092 218482 166396 218498
rect 166080 218476 166396 218482
rect 166132 218470 166396 218476
rect 166080 218418 166132 218424
rect 166644 217138 166672 218554
rect 167472 217138 167500 219234
rect 168024 217274 168052 224334
rect 168196 221740 168248 221746
rect 168196 221682 168248 221688
rect 168208 219298 168236 221682
rect 169680 219298 169708 225830
rect 169864 221882 169892 231662
rect 169852 221876 169904 221882
rect 169852 221818 169904 221824
rect 168196 219292 168248 219298
rect 168196 219234 168248 219240
rect 169116 219292 169168 219298
rect 169116 219234 169168 219240
rect 169668 219292 169720 219298
rect 169668 219234 169720 219240
rect 169944 219292 169996 219298
rect 169944 219234 169996 219240
rect 168024 217246 168282 217274
rect 164942 217110 165016 217138
rect 165770 217110 165844 217138
rect 166598 217110 166672 217138
rect 167426 217110 167500 217138
rect 164942 216988 164970 217110
rect 165770 216988 165798 217110
rect 166598 216988 166626 217110
rect 167426 216988 167454 217110
rect 168254 216988 168282 217246
rect 169128 217138 169156 219234
rect 169956 217138 169984 219234
rect 170324 217462 170352 231662
rect 171048 229764 171100 229770
rect 171048 229706 171100 229712
rect 170864 224800 170916 224806
rect 170864 224742 170916 224748
rect 170876 224126 170904 224742
rect 170864 224120 170916 224126
rect 170864 224062 170916 224068
rect 171060 219298 171088 229706
rect 171230 227624 171286 227633
rect 171230 227559 171286 227568
rect 171244 227458 171272 227559
rect 171232 227452 171284 227458
rect 171232 227394 171284 227400
rect 171428 226930 171456 231676
rect 171704 231662 172086 231690
rect 171704 227361 171732 231662
rect 172150 227624 172206 227633
rect 172150 227559 172206 227568
rect 172164 227458 172192 227559
rect 172152 227452 172204 227458
rect 172152 227394 172204 227400
rect 171690 227352 171746 227361
rect 171690 227287 171746 227296
rect 171600 227180 171652 227186
rect 171600 227122 171652 227128
rect 171336 226902 171456 226930
rect 171048 219292 171100 219298
rect 171048 219234 171100 219240
rect 171140 218884 171192 218890
rect 171140 218826 171192 218832
rect 170954 218512 171010 218521
rect 171152 218482 171180 218826
rect 170954 218447 170956 218456
rect 171008 218447 171010 218456
rect 171140 218476 171192 218482
rect 170956 218418 171008 218424
rect 171140 218418 171192 218424
rect 171336 218362 171364 226902
rect 171612 225894 171640 227122
rect 171600 225888 171652 225894
rect 171600 225830 171652 225836
rect 171784 225888 171836 225894
rect 171784 225830 171836 225836
rect 171796 224954 171824 225830
rect 171244 218334 171364 218362
rect 171428 224926 171824 224954
rect 170772 218068 170824 218074
rect 170772 218010 170824 218016
rect 170312 217456 170364 217462
rect 170312 217398 170364 217404
rect 170784 217138 170812 218010
rect 171244 217326 171272 218334
rect 171428 218210 171456 224926
rect 171796 224726 172192 224754
rect 171796 224670 171824 224726
rect 171784 224664 171836 224670
rect 171784 224606 171836 224612
rect 171968 224664 172020 224670
rect 171968 224606 172020 224612
rect 171554 224392 171606 224398
rect 171606 224340 171824 224346
rect 171554 224334 171824 224340
rect 171566 224318 171824 224334
rect 171796 224126 171824 224318
rect 171980 224262 172008 224606
rect 172164 224398 172192 224726
rect 172152 224392 172204 224398
rect 172152 224334 172204 224340
rect 171968 224256 172020 224262
rect 171968 224198 172020 224204
rect 172152 224256 172204 224262
rect 172152 224198 172204 224204
rect 171784 224120 171836 224126
rect 171784 224062 171836 224068
rect 171784 223576 171836 223582
rect 171784 223518 171836 223524
rect 171796 222902 171824 223518
rect 171784 222896 171836 222902
rect 171784 222838 171836 222844
rect 172164 219298 172192 224198
rect 172716 222018 172744 231676
rect 172992 231662 173374 231690
rect 172992 224942 173020 231662
rect 174004 230926 174032 231676
rect 174280 231662 174662 231690
rect 175306 231662 175596 231690
rect 175950 231662 176148 231690
rect 173992 230920 174044 230926
rect 173992 230862 174044 230868
rect 174280 229226 174308 231662
rect 174268 229220 174320 229226
rect 174268 229162 174320 229168
rect 173162 228848 173218 228857
rect 173162 228783 173218 228792
rect 174818 228848 174874 228857
rect 174818 228783 174820 228792
rect 172980 224936 173032 224942
rect 172980 224878 173032 224884
rect 172888 222896 172940 222902
rect 172888 222838 172940 222844
rect 172704 222012 172756 222018
rect 172704 221954 172756 221960
rect 171600 219292 171652 219298
rect 171600 219234 171652 219240
rect 172152 219292 172204 219298
rect 172152 219234 172204 219240
rect 172428 219292 172480 219298
rect 172428 219234 172480 219240
rect 171416 218204 171468 218210
rect 171416 218146 171468 218152
rect 171232 217320 171284 217326
rect 171232 217262 171284 217268
rect 171612 217138 171640 219234
rect 172440 217138 172468 219234
rect 172900 218521 172928 222838
rect 173176 219298 173204 228783
rect 174872 228783 174874 228792
rect 174820 228754 174872 228760
rect 174084 221876 174136 221882
rect 174084 221818 174136 221824
rect 173164 219292 173216 219298
rect 173164 219234 173216 219240
rect 172886 218512 172942 218521
rect 172886 218447 172942 218456
rect 173256 218204 173308 218210
rect 173256 218146 173308 218152
rect 173268 217138 173296 218146
rect 174096 217138 174124 221818
rect 174912 221740 174964 221746
rect 174912 221682 174964 221688
rect 174924 217138 174952 221682
rect 175568 220153 175596 231662
rect 176120 224954 176148 231662
rect 176028 224926 176148 224954
rect 176488 231662 176594 231690
rect 176028 223446 176056 224926
rect 176290 224904 176346 224913
rect 176290 224839 176346 224848
rect 176304 224262 176332 224839
rect 176292 224256 176344 224262
rect 176292 224198 176344 224204
rect 176488 223938 176516 231662
rect 176752 230172 176804 230178
rect 176752 230114 176804 230120
rect 176764 229094 176792 230114
rect 176304 223910 176516 223938
rect 176672 229066 176792 229094
rect 176016 223440 176068 223446
rect 176304 223394 176332 223910
rect 176672 223530 176700 229066
rect 177224 227458 177252 231676
rect 177408 231662 177882 231690
rect 177212 227452 177264 227458
rect 177212 227394 177264 227400
rect 176844 224936 176896 224942
rect 176842 224904 176844 224913
rect 176896 224904 176898 224913
rect 176842 224839 176898 224848
rect 177408 224210 177436 231662
rect 178512 224806 178540 231676
rect 178788 231662 179170 231690
rect 178500 224800 178552 224806
rect 178500 224742 178552 224748
rect 176016 223382 176068 223388
rect 176212 223366 176332 223394
rect 176580 223502 176700 223530
rect 177316 224182 177436 224210
rect 176212 223258 176240 223366
rect 176120 223230 176240 223258
rect 176120 223174 176148 223230
rect 176108 223168 176160 223174
rect 176108 223110 176160 223116
rect 176580 221626 176608 223502
rect 176304 221598 176608 221626
rect 175554 220144 175610 220153
rect 175554 220079 175610 220088
rect 175740 218748 175792 218754
rect 175740 218690 175792 218696
rect 175752 217138 175780 218690
rect 176304 217274 176332 221598
rect 177316 221377 177344 224182
rect 177488 224120 177540 224126
rect 177488 224062 177540 224068
rect 176474 221368 176530 221377
rect 176474 221303 176476 221312
rect 176528 221303 176530 221312
rect 177302 221368 177358 221377
rect 177302 221303 177358 221312
rect 176476 221274 176528 221280
rect 177304 221196 177356 221202
rect 177304 221138 177356 221144
rect 176474 220824 176530 220833
rect 176474 220759 176476 220768
rect 176528 220759 176530 220768
rect 176614 220788 176666 220794
rect 176476 220730 176528 220736
rect 176614 220730 176666 220736
rect 176626 220674 176654 220730
rect 176488 220646 176654 220674
rect 176488 218074 176516 220646
rect 176476 218068 176528 218074
rect 176476 218010 176528 218016
rect 177316 217274 177344 221138
rect 177500 219162 177528 224062
rect 178788 219434 178816 231662
rect 179800 228954 179828 231676
rect 179984 231662 180458 231690
rect 179788 228948 179840 228954
rect 179788 228890 179840 228896
rect 179328 224936 179380 224942
rect 179328 224878 179380 224884
rect 178420 219406 178816 219434
rect 177488 219156 177540 219162
rect 177488 219098 177540 219104
rect 178224 218068 178276 218074
rect 178224 218010 178276 218016
rect 176304 217246 176562 217274
rect 177316 217246 177390 217274
rect 169082 217110 169156 217138
rect 169910 217110 169984 217138
rect 170738 217110 170812 217138
rect 171566 217110 171640 217138
rect 172394 217110 172468 217138
rect 173222 217110 173296 217138
rect 174050 217110 174124 217138
rect 174878 217110 174952 217138
rect 175706 217110 175780 217138
rect 169082 216988 169110 217110
rect 169910 216988 169938 217110
rect 170738 216988 170766 217110
rect 171566 216988 171594 217110
rect 172394 216988 172422 217110
rect 173222 216988 173250 217110
rect 174050 216988 174078 217110
rect 174878 216988 174906 217110
rect 175706 216988 175734 217110
rect 176534 216988 176562 217246
rect 177362 216988 177390 217246
rect 178236 217138 178264 218010
rect 178420 217598 178448 219406
rect 179052 219156 179104 219162
rect 179052 219098 179104 219104
rect 178408 217592 178460 217598
rect 178408 217534 178460 217540
rect 179064 217138 179092 219098
rect 179340 218074 179368 224878
rect 179786 220824 179842 220833
rect 179984 220810 180012 231662
rect 180156 228948 180208 228954
rect 180156 228890 180208 228896
rect 179842 220782 180012 220810
rect 179786 220759 179842 220768
rect 180168 219434 180196 228890
rect 181088 223990 181116 231676
rect 181352 227452 181404 227458
rect 181352 227394 181404 227400
rect 181076 223984 181128 223990
rect 181076 223926 181128 223932
rect 180524 220788 180576 220794
rect 180524 220730 180576 220736
rect 180708 220788 180760 220794
rect 180708 220730 180760 220736
rect 180536 220153 180564 220730
rect 180522 220144 180578 220153
rect 180522 220079 180578 220088
rect 180076 219406 180196 219434
rect 180076 218890 180104 219406
rect 180064 218884 180116 218890
rect 180064 218826 180116 218832
rect 179880 218204 179932 218210
rect 179880 218146 179932 218152
rect 179328 218068 179380 218074
rect 179328 218010 179380 218016
rect 179892 217138 179920 218146
rect 180720 217274 180748 220730
rect 180890 220008 180946 220017
rect 180890 219943 180892 219952
rect 180944 219943 180946 219952
rect 180892 219914 180944 219920
rect 181168 218748 181220 218754
rect 181168 218690 181220 218696
rect 181180 218346 181208 218690
rect 181364 218482 181392 227394
rect 181732 223582 181760 231676
rect 182376 227594 182404 231676
rect 182652 231662 183034 231690
rect 183678 231662 183876 231690
rect 182364 227588 182416 227594
rect 182364 227530 182416 227536
rect 181720 223576 181772 223582
rect 181720 223518 181772 223524
rect 181996 223168 182048 223174
rect 181996 223110 182048 223116
rect 181534 220280 181590 220289
rect 181534 220215 181590 220224
rect 181548 220114 181576 220215
rect 181536 220108 181588 220114
rect 181536 220050 181588 220056
rect 181352 218476 181404 218482
rect 181352 218418 181404 218424
rect 182008 218346 182036 223110
rect 182652 221610 182680 231662
rect 183848 223854 183876 231662
rect 184308 230790 184336 231676
rect 184296 230784 184348 230790
rect 184296 230726 184348 230732
rect 184664 229220 184716 229226
rect 184664 229162 184716 229168
rect 183836 223848 183888 223854
rect 183836 223790 183888 223796
rect 184388 223848 184440 223854
rect 184388 223790 184440 223796
rect 183192 223576 183244 223582
rect 183192 223518 183244 223524
rect 182640 221604 182692 221610
rect 182640 221546 182692 221552
rect 182364 219292 182416 219298
rect 182364 219234 182416 219240
rect 181168 218340 181220 218346
rect 181168 218282 181220 218288
rect 181536 218340 181588 218346
rect 181536 218282 181588 218288
rect 181996 218340 182048 218346
rect 181996 218282 182048 218288
rect 178190 217110 178264 217138
rect 179018 217110 179092 217138
rect 179846 217110 179920 217138
rect 180674 217246 180748 217274
rect 178190 216988 178218 217110
rect 179018 216988 179046 217110
rect 179846 216988 179874 217110
rect 180674 216988 180702 217246
rect 181548 217138 181576 218282
rect 182376 217138 182404 219234
rect 183204 217274 183232 223518
rect 184400 218754 184428 223790
rect 184676 223582 184704 229162
rect 184952 228274 184980 231676
rect 185136 231662 185610 231690
rect 185872 231662 186254 231690
rect 184940 228268 184992 228274
rect 184940 228210 184992 228216
rect 184664 223576 184716 223582
rect 184664 223518 184716 223524
rect 184848 223576 184900 223582
rect 184848 223518 184900 223524
rect 184662 221776 184718 221785
rect 184662 221711 184718 221720
rect 184676 219434 184704 221711
rect 184676 219406 184796 219434
rect 184388 218748 184440 218754
rect 184388 218690 184440 218696
rect 184020 218340 184072 218346
rect 184020 218282 184072 218288
rect 181502 217110 181576 217138
rect 182330 217110 182404 217138
rect 183158 217246 183232 217274
rect 181502 216988 181530 217110
rect 182330 216988 182358 217110
rect 183158 216988 183186 217246
rect 184032 217138 184060 218282
rect 184768 217274 184796 219406
rect 184860 218362 184888 223518
rect 185136 220017 185164 231662
rect 185872 229094 185900 231662
rect 185872 229066 185992 229094
rect 185400 227724 185452 227730
rect 185400 227666 185452 227672
rect 185412 226914 185440 227666
rect 185584 227316 185636 227322
rect 185584 227258 185636 227264
rect 185596 226914 185624 227258
rect 185400 226908 185452 226914
rect 185400 226850 185452 226856
rect 185584 226908 185636 226914
rect 185584 226850 185636 226856
rect 185584 224936 185636 224942
rect 185584 224878 185636 224884
rect 185768 224936 185820 224942
rect 185768 224878 185820 224884
rect 185596 224670 185624 224878
rect 185400 224664 185452 224670
rect 185400 224606 185452 224612
rect 185584 224664 185636 224670
rect 185584 224606 185636 224612
rect 185412 224126 185440 224606
rect 185400 224120 185452 224126
rect 185400 224062 185452 224068
rect 185780 223990 185808 224878
rect 185768 223984 185820 223990
rect 185768 223926 185820 223932
rect 185964 222154 185992 229066
rect 186136 227452 186188 227458
rect 186136 227394 186188 227400
rect 185952 222148 186004 222154
rect 185952 222090 186004 222096
rect 185766 221776 185822 221785
rect 185766 221711 185768 221720
rect 185820 221711 185822 221720
rect 185768 221682 185820 221688
rect 185860 221332 185912 221338
rect 185860 221274 185912 221280
rect 185872 221218 185900 221274
rect 185320 221202 185900 221218
rect 185308 221196 185900 221202
rect 185360 221190 185900 221196
rect 185308 221138 185360 221144
rect 185122 220008 185178 220017
rect 185122 219943 185178 219952
rect 184860 218346 184980 218362
rect 186148 218346 186176 227394
rect 186884 223310 186912 231676
rect 187528 227594 187556 231676
rect 188172 230654 188200 231676
rect 188160 230648 188212 230654
rect 188160 230590 188212 230596
rect 187516 227588 187568 227594
rect 187516 227530 187568 227536
rect 188816 223718 188844 231676
rect 189092 231662 189474 231690
rect 189092 229094 189120 231662
rect 189092 229066 189304 229094
rect 188804 223712 188856 223718
rect 188804 223654 188856 223660
rect 187332 223440 187384 223446
rect 187332 223382 187384 223388
rect 186872 223304 186924 223310
rect 186872 223246 186924 223252
rect 186504 218884 186556 218890
rect 186504 218826 186556 218832
rect 184860 218340 184992 218346
rect 184860 218334 184940 218340
rect 184940 218282 184992 218288
rect 185676 218340 185728 218346
rect 185676 218282 185728 218288
rect 186136 218340 186188 218346
rect 186136 218282 186188 218288
rect 184768 217246 184842 217274
rect 183986 217110 184060 217138
rect 183986 216988 184014 217110
rect 184814 216988 184842 217246
rect 185688 217138 185716 218282
rect 186516 217138 186544 218826
rect 187344 217274 187372 223382
rect 188896 223304 188948 223310
rect 188896 223246 188948 223252
rect 188908 218346 188936 223246
rect 188160 218340 188212 218346
rect 188160 218282 188212 218288
rect 188896 218340 188948 218346
rect 188896 218282 188948 218288
rect 189080 218340 189132 218346
rect 189080 218282 189132 218288
rect 185642 217110 185716 217138
rect 186470 217110 186544 217138
rect 187298 217246 187372 217274
rect 185642 216988 185670 217110
rect 186470 216988 186498 217110
rect 187298 216988 187326 217246
rect 188172 217138 188200 218282
rect 189092 218226 189120 218282
rect 188908 218198 189120 218226
rect 188908 217274 188936 218198
rect 189276 217734 189304 229066
rect 189724 228268 189776 228274
rect 189724 228210 189776 228216
rect 189736 219298 189764 228210
rect 190104 228138 190132 231676
rect 190656 231662 190762 231690
rect 190656 229094 190684 231662
rect 190472 229066 190684 229094
rect 190092 228132 190144 228138
rect 190092 228074 190144 228080
rect 189908 227452 189960 227458
rect 189908 227394 189960 227400
rect 189724 219292 189776 219298
rect 189724 219234 189776 219240
rect 189920 218754 189948 227394
rect 190472 219978 190500 229066
rect 191392 222766 191420 231676
rect 191564 223984 191616 223990
rect 191564 223926 191616 223932
rect 191380 222760 191432 222766
rect 191380 222702 191432 222708
rect 190460 219972 190512 219978
rect 190460 219914 190512 219920
rect 190644 219972 190696 219978
rect 190644 219914 190696 219920
rect 189908 218748 189960 218754
rect 189908 218690 189960 218696
rect 189816 218476 189868 218482
rect 189816 218418 189868 218424
rect 189264 217728 189316 217734
rect 189264 217670 189316 217676
rect 188908 217246 188982 217274
rect 188126 217110 188200 217138
rect 188126 216988 188154 217110
rect 188954 216988 188982 217246
rect 189828 217138 189856 218418
rect 190656 217274 190684 219914
rect 191576 219434 191604 223926
rect 192036 222630 192064 231676
rect 192680 227730 192708 231676
rect 193036 228132 193088 228138
rect 193036 228074 193088 228080
rect 192668 227724 192720 227730
rect 192668 227666 192720 227672
rect 192024 222624 192076 222630
rect 192024 222566 192076 222572
rect 191484 219406 191604 219434
rect 191484 217274 191512 219406
rect 192852 219292 192904 219298
rect 192852 219234 192904 219240
rect 191932 218748 191984 218754
rect 191932 218690 191984 218696
rect 191944 218482 191972 218690
rect 191932 218476 191984 218482
rect 191932 218418 191984 218424
rect 192300 218340 192352 218346
rect 192300 218282 192352 218288
rect 189782 217110 189856 217138
rect 190610 217246 190684 217274
rect 191438 217246 191512 217274
rect 189782 216988 189810 217110
rect 190610 216988 190638 217246
rect 191438 216988 191466 217246
rect 192312 217138 192340 218282
rect 192864 217274 192892 219234
rect 193048 218346 193076 228074
rect 193324 221066 193352 231676
rect 193968 226302 193996 231676
rect 193956 226296 194008 226302
rect 193956 226238 194008 226244
rect 193772 226024 193824 226030
rect 193772 225966 193824 225972
rect 193312 221060 193364 221066
rect 193312 221002 193364 221008
rect 193784 218482 193812 225966
rect 194612 224126 194640 231676
rect 195060 230648 195112 230654
rect 195060 230590 195112 230596
rect 195072 230042 195100 230590
rect 195060 230036 195112 230042
rect 195060 229978 195112 229984
rect 195256 228002 195284 231676
rect 195900 231538 195928 231676
rect 196176 231662 196558 231690
rect 196912 231662 197202 231690
rect 197464 231662 197846 231690
rect 198016 231662 198490 231690
rect 195888 231532 195940 231538
rect 195888 231474 195940 231480
rect 195428 230036 195480 230042
rect 195428 229978 195480 229984
rect 195244 227996 195296 228002
rect 195244 227938 195296 227944
rect 195244 226296 195296 226302
rect 195244 226238 195296 226244
rect 195256 225214 195284 226238
rect 195244 225208 195296 225214
rect 195244 225150 195296 225156
rect 194600 224120 194652 224126
rect 194600 224062 194652 224068
rect 194508 222624 194560 222630
rect 194508 222566 194560 222572
rect 193772 218476 193824 218482
rect 193772 218418 193824 218424
rect 194520 218346 194548 222566
rect 195440 219434 195468 229978
rect 196176 225486 196204 231662
rect 196912 230654 196940 231662
rect 196900 230648 196952 230654
rect 196900 230590 196952 230596
rect 197464 226778 197492 231662
rect 198016 229094 198044 231662
rect 197740 229066 198044 229094
rect 197452 226772 197504 226778
rect 197452 226714 197504 226720
rect 196164 225480 196216 225486
rect 196164 225422 196216 225428
rect 196624 225208 196676 225214
rect 196624 225150 196676 225156
rect 195888 224120 195940 224126
rect 195888 224062 195940 224068
rect 195256 219406 195468 219434
rect 195256 218754 195284 219406
rect 195244 218748 195296 218754
rect 195244 218690 195296 218696
rect 195612 218748 195664 218754
rect 195612 218690 195664 218696
rect 193036 218340 193088 218346
rect 193036 218282 193088 218288
rect 193956 218340 194008 218346
rect 193956 218282 194008 218288
rect 194508 218340 194560 218346
rect 194508 218282 194560 218288
rect 194784 218340 194836 218346
rect 194784 218282 194836 218288
rect 192864 217246 193122 217274
rect 192266 217110 192340 217138
rect 192266 216988 192294 217110
rect 193094 216988 193122 217246
rect 193968 217138 193996 218282
rect 194796 217138 194824 218282
rect 195624 217138 195652 218690
rect 195900 218346 195928 224062
rect 196636 219162 196664 225150
rect 197176 222760 197228 222766
rect 197176 222702 197228 222708
rect 196624 219156 196676 219162
rect 196624 219098 196676 219104
rect 195888 218340 195940 218346
rect 195888 218282 195940 218288
rect 196440 218340 196492 218346
rect 196440 218282 196492 218288
rect 196452 217138 196480 218282
rect 197188 217274 197216 222702
rect 197740 217870 197768 229066
rect 198004 225480 198056 225486
rect 198004 225422 198056 225428
rect 198016 218754 198044 225422
rect 199120 225350 199148 231676
rect 199292 226024 199344 226030
rect 199292 225966 199344 225972
rect 199476 226024 199528 226030
rect 199476 225966 199528 225972
rect 199304 225350 199332 225966
rect 199108 225344 199160 225350
rect 199108 225286 199160 225292
rect 199292 225344 199344 225350
rect 199292 225286 199344 225292
rect 199488 225214 199516 225966
rect 199476 225208 199528 225214
rect 199476 225150 199528 225156
rect 199764 224942 199792 231676
rect 200408 227866 200436 231676
rect 200592 231662 201066 231690
rect 200396 227860 200448 227866
rect 200396 227802 200448 227808
rect 200028 227724 200080 227730
rect 200028 227666 200080 227672
rect 200040 225026 200068 227666
rect 200040 224998 200160 225026
rect 199752 224936 199804 224942
rect 199752 224878 199804 224884
rect 199936 224936 199988 224942
rect 199936 224878 199988 224884
rect 199948 224074 199976 224878
rect 200132 224754 200160 224998
rect 199856 224046 199976 224074
rect 200040 224726 200160 224754
rect 199856 223990 199884 224046
rect 199844 223984 199896 223990
rect 199844 223926 199896 223932
rect 200040 219298 200068 224726
rect 200592 222306 200620 231662
rect 201696 226302 201724 231676
rect 202340 230314 202368 231676
rect 202998 231662 203196 231690
rect 202328 230308 202380 230314
rect 202328 230250 202380 230256
rect 202878 229120 202934 229129
rect 202878 229055 202880 229064
rect 202932 229055 202934 229064
rect 202880 229026 202932 229032
rect 203168 226642 203196 231662
rect 203628 230518 203656 231676
rect 203616 230512 203668 230518
rect 203616 230454 203668 230460
rect 203524 227860 203576 227866
rect 203524 227802 203576 227808
rect 203156 226636 203208 226642
rect 203156 226578 203208 226584
rect 201684 226296 201736 226302
rect 201684 226238 201736 226244
rect 203156 226296 203208 226302
rect 203156 226238 203208 226244
rect 203168 225622 203196 226238
rect 203156 225616 203208 225622
rect 203156 225558 203208 225564
rect 202788 225208 202840 225214
rect 202788 225150 202840 225156
rect 201408 223984 201460 223990
rect 201408 223926 201460 223932
rect 200224 222278 200620 222306
rect 200224 219842 200252 222278
rect 200396 222148 200448 222154
rect 200396 222090 200448 222096
rect 200212 219836 200264 219842
rect 200212 219778 200264 219784
rect 198188 219292 198240 219298
rect 198188 219234 198240 219240
rect 198924 219292 198976 219298
rect 198924 219234 198976 219240
rect 200028 219292 200080 219298
rect 200028 219234 200080 219240
rect 198200 218754 198228 219234
rect 198004 218748 198056 218754
rect 198004 218690 198056 218696
rect 198188 218748 198240 218754
rect 198188 218690 198240 218696
rect 198096 218476 198148 218482
rect 198096 218418 198148 218424
rect 197728 217864 197780 217870
rect 197728 217806 197780 217812
rect 197188 217246 197262 217274
rect 193922 217110 193996 217138
rect 194750 217110 194824 217138
rect 195578 217110 195652 217138
rect 196406 217110 196480 217138
rect 193922 216988 193950 217110
rect 194750 216988 194778 217110
rect 195578 216988 195606 217110
rect 196406 216988 196434 217110
rect 197234 216988 197262 217246
rect 198108 217138 198136 218418
rect 198936 217138 198964 219234
rect 199752 219156 199804 219162
rect 199752 219098 199804 219104
rect 199764 217138 199792 219098
rect 200408 218482 200436 222090
rect 200580 219836 200632 219842
rect 200580 219778 200632 219784
rect 200396 218476 200448 218482
rect 200396 218418 200448 218424
rect 200592 217274 200620 219778
rect 201420 217274 201448 223926
rect 202604 219292 202656 219298
rect 202604 219234 202656 219240
rect 202616 218618 202644 219234
rect 202604 218612 202656 218618
rect 202604 218554 202656 218560
rect 202800 218482 202828 225150
rect 203536 219026 203564 227802
rect 204076 227044 204128 227050
rect 204076 226986 204128 226992
rect 204088 226642 204116 226986
rect 204076 226636 204128 226642
rect 204076 226578 204128 226584
rect 203890 225448 203946 225457
rect 203890 225383 203946 225392
rect 203524 219020 203576 219026
rect 203524 218962 203576 218968
rect 203064 218612 203116 218618
rect 203064 218554 203116 218560
rect 202236 218476 202288 218482
rect 202236 218418 202288 218424
rect 202788 218476 202840 218482
rect 202788 218418 202840 218424
rect 198062 217110 198136 217138
rect 198890 217110 198964 217138
rect 199718 217110 199792 217138
rect 200546 217246 200620 217274
rect 201374 217246 201448 217274
rect 198062 216988 198090 217110
rect 198890 216988 198918 217110
rect 199718 216988 199746 217110
rect 200546 216988 200574 217246
rect 201374 216988 201402 217246
rect 202248 217138 202276 218418
rect 203076 217138 203104 218554
rect 203904 217274 203932 225383
rect 204272 225078 204300 231676
rect 204720 229084 204772 229090
rect 204720 229026 204772 229032
rect 204732 228138 204760 229026
rect 204720 228132 204772 228138
rect 204720 228074 204772 228080
rect 204916 227882 204944 231676
rect 205192 231662 205574 231690
rect 205836 231662 206218 231690
rect 205192 229129 205220 231662
rect 205178 229120 205234 229129
rect 205178 229055 205234 229064
rect 205456 227996 205508 228002
rect 205456 227938 205508 227944
rect 204548 227854 204944 227882
rect 204548 225894 204576 227854
rect 204904 227724 204956 227730
rect 204904 227666 204956 227672
rect 204916 227458 204944 227666
rect 204720 227452 204772 227458
rect 204720 227394 204772 227400
rect 204904 227452 204956 227458
rect 204904 227394 204956 227400
rect 204732 226778 204760 227394
rect 204720 226772 204772 226778
rect 204720 226714 204772 226720
rect 204536 225888 204588 225894
rect 204536 225830 204588 225836
rect 204720 225888 204772 225894
rect 204720 225830 204772 225836
rect 204732 225486 204760 225830
rect 204904 225752 204956 225758
rect 204904 225694 204956 225700
rect 204720 225480 204772 225486
rect 204720 225422 204772 225428
rect 204916 225350 204944 225694
rect 205088 225480 205140 225486
rect 205086 225448 205088 225457
rect 205140 225448 205142 225457
rect 205086 225383 205142 225392
rect 204904 225344 204956 225350
rect 204904 225286 204956 225292
rect 204628 225208 204680 225214
rect 204628 225150 204680 225156
rect 204260 225072 204312 225078
rect 204260 225014 204312 225020
rect 204640 219434 204668 225150
rect 204904 221468 204956 221474
rect 204904 221410 204956 221416
rect 205088 221468 205140 221474
rect 205088 221410 205140 221416
rect 204916 221202 204944 221410
rect 204904 221196 204956 221202
rect 204904 221138 204956 221144
rect 205100 221066 205128 221410
rect 205088 221060 205140 221066
rect 205088 221002 205140 221008
rect 204536 219428 204668 219434
rect 204588 219406 204668 219428
rect 204536 219370 204588 219376
rect 204720 218476 204772 218482
rect 204720 218418 204772 218424
rect 202202 217110 202276 217138
rect 203030 217110 203104 217138
rect 203858 217246 203932 217274
rect 202202 216988 202230 217110
rect 203030 216988 203058 217110
rect 203858 216988 203886 217246
rect 204732 217138 204760 218418
rect 205468 217274 205496 227938
rect 205836 219706 205864 231662
rect 206284 230444 206336 230450
rect 206284 230386 206336 230392
rect 205824 219700 205876 219706
rect 205824 219642 205876 219648
rect 206296 219434 206324 230386
rect 206848 222494 206876 231676
rect 207492 223854 207520 231676
rect 208136 226642 208164 231676
rect 208596 231662 208794 231690
rect 208124 226636 208176 226642
rect 208124 226578 208176 226584
rect 207480 223848 207532 223854
rect 207480 223790 207532 223796
rect 207664 223712 207716 223718
rect 207664 223654 207716 223660
rect 206836 222488 206888 222494
rect 206836 222430 206888 222436
rect 207204 219700 207256 219706
rect 207204 219642 207256 219648
rect 206204 219406 206324 219434
rect 206204 218618 206232 219406
rect 206376 219020 206428 219026
rect 206376 218962 206428 218968
rect 206192 218612 206244 218618
rect 206192 218554 206244 218560
rect 205468 217246 205542 217274
rect 204686 217110 204760 217138
rect 204686 216988 204714 217110
rect 205514 216988 205542 217246
rect 206388 217138 206416 218962
rect 207216 217274 207244 219642
rect 207676 219298 207704 223654
rect 207848 222488 207900 222494
rect 207848 222430 207900 222436
rect 207664 219292 207716 219298
rect 207664 219234 207716 219240
rect 207860 218482 207888 222430
rect 208596 220386 208624 231662
rect 209424 226302 209452 231676
rect 210068 229498 210096 231676
rect 210424 230308 210476 230314
rect 210424 230250 210476 230256
rect 210056 229492 210108 229498
rect 210056 229434 210108 229440
rect 209412 226296 209464 226302
rect 209412 226238 209464 226244
rect 209596 226296 209648 226302
rect 209596 226238 209648 226244
rect 209608 225706 209636 226238
rect 209332 225678 209636 225706
rect 209332 225486 209360 225678
rect 209320 225480 209372 225486
rect 209320 225422 209372 225428
rect 209504 225480 209556 225486
rect 209504 225422 209556 225428
rect 208584 220380 208636 220386
rect 208584 220322 208636 220328
rect 208032 218612 208084 218618
rect 208032 218554 208084 218560
rect 207848 218476 207900 218482
rect 207848 218418 207900 218424
rect 206342 217110 206416 217138
rect 207170 217246 207244 217274
rect 206342 216988 206370 217110
rect 207170 216988 207198 217246
rect 208044 217138 208072 218554
rect 209516 218482 209544 225422
rect 210436 219434 210464 230250
rect 210712 228546 210740 231676
rect 211172 231662 211370 231690
rect 210700 228540 210752 228546
rect 210700 228482 210752 228488
rect 210976 227860 211028 227866
rect 210976 227802 211028 227808
rect 209688 219428 209740 219434
rect 209688 219370 209740 219376
rect 210424 219428 210476 219434
rect 210424 219370 210476 219376
rect 208860 218476 208912 218482
rect 208860 218418 208912 218424
rect 209504 218476 209556 218482
rect 209504 218418 209556 218424
rect 208872 217138 208900 218418
rect 209700 217138 209728 219370
rect 210148 218612 210200 218618
rect 210148 218554 210200 218560
rect 210160 218346 210188 218554
rect 210148 218340 210200 218346
rect 210148 218282 210200 218288
rect 210332 218340 210384 218346
rect 210332 218282 210384 218288
rect 210344 218074 210372 218282
rect 210988 218074 211016 227802
rect 211172 221202 211200 231662
rect 212000 222358 212028 231676
rect 212356 229084 212408 229090
rect 212356 229026 212408 229032
rect 212368 228682 212396 229026
rect 212356 228676 212408 228682
rect 212356 228618 212408 228624
rect 212172 226636 212224 226642
rect 212172 226578 212224 226584
rect 211988 222352 212040 222358
rect 211988 222294 212040 222300
rect 211160 221196 211212 221202
rect 211160 221138 211212 221144
rect 211528 221196 211580 221202
rect 211528 221138 211580 221144
rect 211344 219292 211396 219298
rect 211344 219234 211396 219240
rect 210332 218068 210384 218074
rect 210332 218010 210384 218016
rect 210516 218068 210568 218074
rect 210516 218010 210568 218016
rect 210976 218068 211028 218074
rect 210976 218010 211028 218016
rect 210528 217138 210556 218010
rect 211356 217138 211384 219234
rect 211540 218482 211568 221138
rect 211528 218476 211580 218482
rect 211528 218418 211580 218424
rect 212184 217274 212212 226578
rect 212644 222902 212672 231676
rect 213288 226506 213316 231676
rect 213946 231662 214144 231690
rect 214116 229094 214144 231662
rect 213932 229066 214144 229094
rect 214576 229094 214604 231676
rect 214748 230036 214800 230042
rect 214748 229978 214800 229984
rect 214760 229634 214788 229978
rect 214748 229628 214800 229634
rect 214748 229570 214800 229576
rect 215220 229362 215248 231676
rect 215208 229356 215260 229362
rect 215208 229298 215260 229304
rect 214380 229084 214432 229090
rect 213276 226500 213328 226506
rect 213276 226442 213328 226448
rect 212632 222896 212684 222902
rect 212632 222838 212684 222844
rect 213184 222896 213236 222902
rect 213184 222838 213236 222844
rect 213000 219428 213052 219434
rect 213000 219370 213052 219376
rect 207998 217110 208072 217138
rect 208826 217110 208900 217138
rect 209654 217110 209728 217138
rect 210482 217110 210556 217138
rect 211310 217110 211384 217138
rect 212138 217246 212212 217274
rect 207998 216988 208026 217110
rect 208826 216988 208854 217110
rect 209654 216988 209682 217110
rect 210482 216988 210510 217110
rect 211310 216988 211338 217110
rect 212138 216988 212166 217246
rect 213012 217138 213040 219370
rect 213196 218346 213224 222838
rect 213932 220810 213960 229066
rect 214576 229066 214788 229094
rect 214380 229026 214432 229032
rect 214392 228002 214420 229026
rect 214564 228404 214616 228410
rect 214564 228346 214616 228352
rect 214576 228138 214604 228346
rect 214564 228132 214616 228138
rect 214564 228074 214616 228080
rect 214380 227996 214432 228002
rect 214380 227938 214432 227944
rect 214760 227746 214788 229066
rect 215864 228546 215892 231676
rect 216048 231662 216522 231690
rect 215852 228540 215904 228546
rect 215852 228482 215904 228488
rect 214576 227718 214788 227746
rect 214104 227044 214156 227050
rect 214104 226986 214156 226992
rect 214116 226778 214144 226986
rect 214104 226772 214156 226778
rect 214104 226714 214156 226720
rect 214576 226166 214604 227718
rect 214748 227588 214800 227594
rect 214748 227530 214800 227536
rect 214932 227588 214984 227594
rect 214932 227530 214984 227536
rect 214760 226914 214788 227530
rect 214748 226908 214800 226914
rect 214748 226850 214800 226856
rect 214944 226642 214972 227530
rect 214932 226636 214984 226642
rect 214932 226578 214984 226584
rect 214564 226160 214616 226166
rect 214564 226102 214616 226108
rect 215208 225072 215260 225078
rect 215208 225014 215260 225020
rect 213932 220782 214052 220810
rect 213828 220380 213880 220386
rect 213828 220322 213880 220328
rect 213184 218340 213236 218346
rect 213184 218282 213236 218288
rect 213840 217274 213868 220322
rect 214024 219570 214052 220782
rect 214012 219564 214064 219570
rect 214012 219506 214064 219512
rect 215220 218074 215248 225014
rect 216048 224954 216076 231662
rect 216220 228540 216272 228546
rect 216220 228482 216272 228488
rect 216232 224954 216260 228482
rect 216404 226500 216456 226506
rect 216404 226442 216456 226448
rect 216416 224954 216444 226442
rect 217152 225622 217180 231676
rect 217508 228404 217560 228410
rect 217508 228346 217560 228352
rect 217140 225616 217192 225622
rect 217140 225558 217192 225564
rect 215956 224926 216076 224954
rect 216140 224926 216260 224954
rect 216324 224926 216444 224954
rect 215956 220250 215984 224926
rect 215944 220244 215996 220250
rect 215944 220186 215996 220192
rect 216140 218074 216168 224926
rect 214656 218068 214708 218074
rect 214656 218010 214708 218016
rect 215208 218068 215260 218074
rect 215208 218010 215260 218016
rect 215484 218068 215536 218074
rect 215484 218010 215536 218016
rect 216128 218068 216180 218074
rect 216128 218010 216180 218016
rect 212966 217110 213040 217138
rect 213794 217246 213868 217274
rect 212966 216988 212994 217110
rect 213794 216988 213822 217246
rect 214668 217138 214696 218010
rect 215496 217138 215524 218010
rect 216324 217274 216352 224926
rect 217140 220244 217192 220250
rect 217140 220186 217192 220192
rect 217152 217274 217180 220186
rect 217520 219434 217548 228346
rect 217796 227730 217824 231676
rect 217784 227724 217836 227730
rect 217784 227666 217836 227672
rect 218440 226778 218468 231676
rect 218428 226772 218480 226778
rect 218428 226714 218480 226720
rect 219084 223038 219112 231676
rect 219742 231662 220216 231690
rect 219992 230036 220044 230042
rect 219992 229978 220044 229984
rect 220004 229770 220032 229978
rect 219992 229764 220044 229770
rect 219992 229706 220044 229712
rect 219808 228812 219860 228818
rect 219808 228754 219860 228760
rect 219622 228712 219678 228721
rect 219622 228647 219678 228656
rect 219636 228546 219664 228647
rect 219624 228540 219676 228546
rect 219624 228482 219676 228488
rect 219820 228138 219848 228754
rect 219992 228540 220044 228546
rect 219992 228482 220044 228488
rect 219808 228132 219860 228138
rect 219808 228074 219860 228080
rect 220004 227866 220032 228482
rect 219992 227860 220044 227866
rect 219992 227802 220044 227808
rect 219808 227724 219860 227730
rect 219808 227666 219860 227672
rect 219532 227316 219584 227322
rect 219532 227258 219584 227264
rect 219348 226772 219400 226778
rect 219348 226714 219400 226720
rect 219072 223032 219124 223038
rect 219072 222974 219124 222980
rect 218060 221060 218112 221066
rect 218060 221002 218112 221008
rect 217336 219406 217548 219434
rect 217336 218618 217364 219406
rect 218072 219298 218100 221002
rect 218060 219292 218112 219298
rect 218060 219234 218112 219240
rect 217324 218612 217376 218618
rect 217324 218554 217376 218560
rect 217968 218476 218020 218482
rect 217968 218418 218020 218424
rect 214622 217110 214696 217138
rect 215450 217110 215524 217138
rect 216278 217246 216352 217274
rect 217106 217246 217180 217274
rect 214622 216988 214650 217110
rect 215450 216988 215478 217110
rect 216278 216988 216306 217246
rect 217106 216988 217134 217246
rect 217980 217138 218008 218418
rect 219360 218074 219388 226714
rect 219544 226642 219572 227258
rect 219820 227186 219848 227666
rect 219992 227316 220044 227322
rect 219992 227258 220044 227264
rect 219808 227180 219860 227186
rect 219808 227122 219860 227128
rect 220004 226914 220032 227258
rect 219992 226908 220044 226914
rect 219992 226850 220044 226856
rect 219532 226636 219584 226642
rect 219532 226578 219584 226584
rect 219992 225616 220044 225622
rect 219992 225558 220044 225564
rect 220004 225078 220032 225558
rect 219992 225072 220044 225078
rect 219992 225014 220044 225020
rect 220188 221474 220216 231662
rect 220372 229498 220400 231676
rect 220360 229492 220412 229498
rect 220360 229434 220412 229440
rect 220728 229492 220780 229498
rect 220728 229434 220780 229440
rect 220360 228948 220412 228954
rect 220360 228890 220412 228896
rect 220372 228682 220400 228890
rect 220542 228712 220598 228721
rect 220360 228676 220412 228682
rect 220542 228647 220544 228656
rect 220360 228618 220412 228624
rect 220596 228647 220598 228656
rect 220544 228618 220596 228624
rect 220740 226624 220768 229434
rect 221016 228002 221044 231676
rect 221292 231662 221674 231690
rect 221004 227996 221056 228002
rect 221004 227938 221056 227944
rect 220556 226596 220768 226624
rect 220556 226506 220584 226596
rect 220544 226500 220596 226506
rect 220544 226442 220596 226448
rect 220728 226500 220780 226506
rect 220728 226442 220780 226448
rect 220176 221468 220228 221474
rect 220176 221410 220228 221416
rect 220740 219434 220768 226442
rect 221004 221468 221056 221474
rect 221004 221410 221056 221416
rect 221016 221066 221044 221410
rect 221004 221060 221056 221066
rect 221004 221002 221056 221008
rect 221292 220658 221320 231662
rect 221464 228404 221516 228410
rect 221464 228346 221516 228352
rect 221476 228002 221504 228346
rect 221464 227996 221516 228002
rect 221464 227938 221516 227944
rect 221832 227044 221884 227050
rect 221832 226986 221884 226992
rect 221280 220652 221332 220658
rect 221280 220594 221332 220600
rect 220464 219406 220768 219434
rect 219624 218612 219676 218618
rect 219624 218554 219676 218560
rect 218796 218068 218848 218074
rect 218796 218010 218848 218016
rect 219348 218068 219400 218074
rect 219348 218010 219400 218016
rect 218808 217138 218836 218010
rect 219636 217138 219664 218554
rect 220464 217274 220492 219406
rect 221844 218074 221872 226986
rect 222016 226160 222068 226166
rect 222016 226102 222068 226108
rect 221280 218068 221332 218074
rect 221280 218010 221332 218016
rect 221832 218068 221884 218074
rect 221832 218010 221884 218016
rect 217934 217110 218008 217138
rect 218762 217110 218836 217138
rect 219590 217110 219664 217138
rect 220418 217246 220492 217274
rect 217934 216988 217962 217110
rect 218762 216988 218790 217110
rect 219590 216988 219618 217110
rect 220418 216988 220446 217246
rect 221292 217138 221320 218010
rect 222028 217274 222056 226102
rect 222304 220930 222332 231676
rect 222948 225350 222976 231676
rect 223592 226642 223620 231676
rect 223776 231662 224250 231690
rect 223580 226636 223632 226642
rect 223580 226578 223632 226584
rect 222936 225344 222988 225350
rect 222936 225286 222988 225292
rect 222292 220924 222344 220930
rect 222292 220866 222344 220872
rect 223488 220924 223540 220930
rect 223488 220866 223540 220872
rect 223500 218482 223528 220866
rect 223776 220658 223804 231662
rect 224592 228404 224644 228410
rect 224592 228346 224644 228352
rect 223764 220652 223816 220658
rect 223764 220594 223816 220600
rect 223764 220516 223816 220522
rect 223764 220458 223816 220464
rect 223488 218476 223540 218482
rect 223488 218418 223540 218424
rect 222936 218340 222988 218346
rect 222936 218282 222988 218288
rect 222028 217246 222102 217274
rect 221246 217110 221320 217138
rect 221246 216988 221274 217110
rect 222074 216988 222102 217246
rect 222948 217138 222976 218282
rect 223776 217274 223804 220458
rect 224604 217274 224632 228346
rect 224880 224534 224908 231676
rect 225524 229906 225552 231676
rect 225512 229900 225564 229906
rect 225512 229842 225564 229848
rect 226168 228818 226196 231676
rect 226536 231662 226826 231690
rect 226156 228812 226208 228818
rect 226156 228754 226208 228760
rect 226156 227860 226208 227866
rect 226156 227802 226208 227808
rect 225604 226636 225656 226642
rect 225604 226578 225656 226584
rect 224868 224528 224920 224534
rect 224868 224470 224920 224476
rect 225616 218210 225644 226578
rect 225972 218476 226024 218482
rect 225972 218418 226024 218424
rect 225604 218204 225656 218210
rect 225604 218146 225656 218152
rect 225420 218068 225472 218074
rect 225420 218010 225472 218016
rect 222902 217110 222976 217138
rect 223730 217246 223804 217274
rect 224558 217246 224632 217274
rect 222902 216988 222930 217110
rect 223730 216988 223758 217246
rect 224558 216988 224586 217246
rect 225432 217138 225460 218010
rect 225984 217274 226012 218418
rect 226168 218074 226196 227802
rect 226536 222018 226564 231662
rect 227456 224398 227484 231676
rect 227444 224392 227496 224398
rect 227444 224334 227496 224340
rect 227536 223848 227588 223854
rect 227536 223790 227588 223796
rect 226524 222012 226576 222018
rect 226524 221954 226576 221960
rect 227548 218074 227576 223790
rect 228100 223718 228128 231676
rect 228744 227730 228772 231676
rect 229296 231662 229402 231690
rect 228732 227724 228784 227730
rect 228732 227666 228784 227672
rect 228916 227724 228968 227730
rect 228916 227666 228968 227672
rect 228928 226506 228956 227666
rect 228916 226500 228968 226506
rect 228916 226442 228968 226448
rect 228732 224528 228784 224534
rect 228732 224470 228784 224476
rect 228088 223712 228140 223718
rect 228088 223654 228140 223660
rect 227904 221060 227956 221066
rect 227904 221002 227956 221008
rect 226156 218068 226208 218074
rect 226156 218010 226208 218016
rect 227076 218068 227128 218074
rect 227076 218010 227128 218016
rect 227536 218068 227588 218074
rect 227536 218010 227588 218016
rect 225984 217246 226242 217274
rect 225386 217110 225460 217138
rect 225386 216988 225414 217110
rect 226214 216988 226242 217246
rect 227088 217138 227116 218010
rect 227916 217274 227944 221002
rect 228744 217274 228772 224470
rect 229296 220114 229324 231662
rect 230032 224262 230060 231676
rect 230676 230042 230704 231676
rect 230664 230036 230716 230042
rect 230664 229978 230716 229984
rect 230480 229900 230532 229906
rect 230480 229842 230532 229848
rect 230020 224256 230072 224262
rect 230492 224210 230520 229842
rect 231124 229492 231176 229498
rect 231124 229434 231176 229440
rect 230020 224198 230072 224204
rect 230400 224182 230520 224210
rect 229284 220108 229336 220114
rect 229284 220050 229336 220056
rect 230204 220108 230256 220114
rect 230204 220050 230256 220056
rect 230216 219434 230244 220050
rect 230216 219406 230336 219434
rect 229560 218068 229612 218074
rect 229560 218010 229612 218016
rect 227042 217110 227116 217138
rect 227870 217246 227944 217274
rect 228698 217246 228772 217274
rect 227042 216988 227070 217110
rect 227870 216988 227898 217246
rect 228698 216988 228726 217246
rect 229572 217138 229600 218010
rect 230308 217274 230336 219406
rect 230400 218090 230428 224182
rect 231136 219434 231164 229434
rect 231320 228138 231348 231676
rect 231308 228132 231360 228138
rect 231308 228074 231360 228080
rect 231676 224256 231728 224262
rect 231676 224198 231728 224204
rect 231044 219406 231164 219434
rect 231044 218346 231072 219406
rect 231032 218340 231084 218346
rect 231032 218282 231084 218288
rect 230400 218074 230520 218090
rect 231688 218074 231716 224198
rect 231964 221882 231992 231676
rect 232608 224806 232636 231676
rect 233252 229094 233280 231676
rect 233896 229094 233924 231676
rect 233252 229066 233372 229094
rect 232596 224800 232648 224806
rect 232596 224742 232648 224748
rect 233148 224392 233200 224398
rect 233148 224334 233200 224340
rect 232136 222012 232188 222018
rect 232136 221954 232188 221960
rect 231952 221876 232004 221882
rect 231952 221818 232004 221824
rect 232148 221610 232176 221954
rect 232136 221604 232188 221610
rect 232136 221546 232188 221552
rect 232872 218340 232924 218346
rect 232872 218282 232924 218288
rect 230400 218068 230532 218074
rect 230400 218062 230480 218068
rect 230480 218010 230532 218016
rect 231216 218068 231268 218074
rect 231216 218010 231268 218016
rect 231676 218068 231728 218074
rect 231676 218010 231728 218016
rect 232044 218068 232096 218074
rect 232044 218010 232096 218016
rect 230308 217246 230382 217274
rect 229526 217110 229600 217138
rect 229526 216988 229554 217110
rect 230354 216988 230382 217246
rect 231228 217138 231256 218010
rect 232056 217138 232084 218010
rect 232884 217138 232912 218282
rect 233160 218074 233188 224334
rect 233344 222902 233372 229066
rect 233712 229066 233924 229094
rect 234172 231662 234554 231690
rect 234724 231662 235198 231690
rect 234172 229094 234200 231662
rect 234172 229066 234292 229094
rect 233712 227186 233740 229066
rect 233884 228132 233936 228138
rect 233884 228074 233936 228080
rect 233896 227866 233924 228074
rect 233884 227860 233936 227866
rect 233884 227802 233936 227808
rect 233700 227180 233752 227186
rect 233700 227122 233752 227128
rect 233332 222896 233384 222902
rect 233332 222838 233384 222844
rect 233700 221876 233752 221882
rect 233700 221818 233752 221824
rect 233148 218068 233200 218074
rect 233148 218010 233200 218016
rect 233712 217274 233740 221818
rect 234068 221468 234120 221474
rect 234068 221410 234120 221416
rect 234080 221066 234108 221410
rect 234264 221338 234292 229066
rect 234528 222896 234580 222902
rect 234528 222838 234580 222844
rect 234252 221332 234304 221338
rect 234252 221274 234304 221280
rect 234068 221060 234120 221066
rect 234068 221002 234120 221008
rect 234540 217274 234568 222838
rect 234724 222018 234752 231662
rect 235828 230178 235856 231676
rect 235816 230172 235868 230178
rect 235816 230114 235868 230120
rect 235816 226772 235868 226778
rect 235816 226714 235868 226720
rect 234712 222012 234764 222018
rect 234712 221954 234764 221960
rect 235828 218074 235856 226714
rect 236472 226030 236500 231676
rect 236748 231662 237130 231690
rect 236460 226024 236512 226030
rect 236460 225966 236512 225972
rect 236748 220794 236776 231662
rect 237760 224670 237788 231676
rect 238404 226642 238432 231676
rect 238576 228812 238628 228818
rect 238576 228754 238628 228760
rect 238392 226636 238444 226642
rect 238392 226578 238444 226584
rect 237748 224664 237800 224670
rect 237748 224606 237800 224612
rect 237012 222352 237064 222358
rect 237012 222294 237064 222300
rect 236736 220788 236788 220794
rect 236736 220730 236788 220736
rect 236184 220652 236236 220658
rect 236184 220594 236236 220600
rect 235356 218068 235408 218074
rect 235356 218010 235408 218016
rect 235816 218068 235868 218074
rect 235816 218010 235868 218016
rect 231182 217110 231256 217138
rect 232010 217110 232084 217138
rect 232838 217110 232912 217138
rect 233666 217246 233740 217274
rect 234494 217246 234568 217274
rect 231182 216988 231210 217110
rect 232010 216988 232038 217110
rect 232838 216988 232866 217110
rect 233666 216988 233694 217246
rect 234494 216988 234522 217246
rect 235368 217138 235396 218010
rect 236196 217274 236224 220594
rect 237024 217274 237052 222294
rect 237840 221332 237892 221338
rect 237840 221274 237892 221280
rect 237852 217274 237880 221274
rect 235322 217110 235396 217138
rect 236150 217246 236224 217274
rect 236978 217246 237052 217274
rect 237806 217246 237880 217274
rect 238588 217274 238616 228754
rect 239048 228274 239076 231676
rect 239036 228268 239088 228274
rect 239036 228210 239088 228216
rect 239312 227860 239364 227866
rect 239312 227802 239364 227808
rect 239324 218890 239352 227802
rect 239692 223582 239720 231676
rect 239680 223576 239732 223582
rect 239680 223518 239732 223524
rect 240336 223174 240364 231676
rect 240980 229226 241008 231676
rect 240968 229220 241020 229226
rect 240968 229162 241020 229168
rect 241624 227322 241652 231676
rect 241612 227316 241664 227322
rect 241612 227258 241664 227264
rect 241152 227180 241204 227186
rect 241152 227122 241204 227128
rect 240324 223168 240376 223174
rect 240324 223110 240376 223116
rect 239496 219292 239548 219298
rect 239496 219234 239548 219240
rect 239312 218884 239364 218890
rect 239312 218826 239364 218832
rect 238588 217246 238662 217274
rect 235322 216988 235350 217110
rect 236150 216988 236178 217246
rect 236978 216988 237006 217246
rect 237806 216988 237834 217246
rect 238634 216988 238662 217246
rect 239508 217138 239536 219234
rect 240324 218068 240376 218074
rect 240324 218010 240376 218016
rect 240336 217138 240364 218010
rect 241164 217274 241192 227122
rect 242268 223446 242296 231676
rect 242926 231662 243124 231690
rect 242532 230036 242584 230042
rect 242532 229978 242584 229984
rect 242544 229094 242572 229978
rect 242544 229066 242756 229094
rect 242256 223440 242308 223446
rect 242256 223382 242308 223388
rect 241336 223168 241388 223174
rect 241336 223110 241388 223116
rect 241348 218074 241376 223110
rect 241980 218204 242032 218210
rect 241980 218146 242032 218152
rect 241336 218068 241388 218074
rect 241336 218010 241388 218016
rect 239462 217110 239536 217138
rect 240290 217110 240364 217138
rect 241118 217246 241192 217274
rect 239462 216988 239490 217110
rect 240290 216988 240318 217110
rect 241118 216988 241146 217246
rect 241992 217138 242020 218146
rect 242728 217274 242756 229066
rect 242900 225344 242952 225350
rect 242820 225292 242900 225298
rect 242820 225286 242952 225292
rect 242820 225270 242940 225286
rect 242820 218226 242848 225270
rect 243096 221746 243124 231662
rect 243556 227866 243584 231676
rect 243544 227860 243596 227866
rect 243544 227802 243596 227808
rect 244200 225758 244228 231676
rect 244476 231662 244858 231690
rect 245120 231662 245502 231690
rect 244188 225752 244240 225758
rect 244188 225694 244240 225700
rect 244096 223440 244148 223446
rect 244096 223382 244148 223388
rect 243084 221740 243136 221746
rect 243084 221682 243136 221688
rect 243728 221604 243780 221610
rect 243728 221546 243780 221552
rect 243740 221338 243768 221546
rect 243728 221332 243780 221338
rect 243728 221274 243780 221280
rect 243544 219156 243596 219162
rect 243544 219098 243596 219104
rect 242820 218210 242940 218226
rect 243556 218210 243584 219098
rect 242820 218204 242952 218210
rect 242820 218198 242900 218204
rect 242900 218146 242952 218152
rect 243544 218204 243596 218210
rect 243544 218146 243596 218152
rect 244108 218074 244136 223382
rect 244476 219978 244504 231662
rect 245120 223310 245148 231662
rect 246132 229770 246160 231676
rect 246120 229764 246172 229770
rect 246120 229706 246172 229712
rect 246488 229356 246540 229362
rect 246488 229298 246540 229304
rect 246304 227860 246356 227866
rect 246304 227802 246356 227808
rect 245476 224800 245528 224806
rect 245476 224742 245528 224748
rect 245108 223304 245160 223310
rect 245108 223246 245160 223252
rect 245292 223032 245344 223038
rect 245292 222974 245344 222980
rect 244464 219972 244516 219978
rect 244464 219914 244516 219920
rect 245304 218074 245332 222974
rect 243636 218068 243688 218074
rect 243636 218010 243688 218016
rect 244096 218068 244148 218074
rect 244096 218010 244148 218016
rect 244464 218068 244516 218074
rect 244464 218010 244516 218016
rect 245292 218068 245344 218074
rect 245292 218010 245344 218016
rect 242728 217246 242802 217274
rect 241946 217110 242020 217138
rect 241946 216988 241974 217110
rect 242774 216988 242802 217246
rect 243648 217138 243676 218010
rect 244476 217138 244504 218010
rect 245488 217274 245516 224742
rect 246120 218884 246172 218890
rect 246120 218826 246172 218832
rect 243602 217110 243676 217138
rect 244430 217110 244504 217138
rect 245258 217246 245516 217274
rect 243602 216988 243630 217110
rect 244430 216988 244458 217110
rect 245258 216988 245286 217246
rect 246132 217138 246160 218826
rect 246316 218754 246344 227802
rect 246500 220658 246528 229298
rect 246776 228954 246804 231676
rect 246764 228948 246816 228954
rect 246764 228890 246816 228896
rect 247420 222630 247448 231676
rect 248064 224942 248092 231676
rect 248708 227866 248736 231676
rect 249260 231662 249366 231690
rect 248696 227860 248748 227866
rect 248696 227802 248748 227808
rect 249064 227860 249116 227866
rect 249064 227802 249116 227808
rect 248052 224936 248104 224942
rect 248052 224878 248104 224884
rect 248328 224664 248380 224670
rect 248328 224606 248380 224612
rect 247408 222624 247460 222630
rect 247408 222566 247460 222572
rect 246948 220788 247000 220794
rect 246948 220730 247000 220736
rect 246488 220652 246540 220658
rect 246488 220594 246540 220600
rect 246304 218748 246356 218754
rect 246304 218690 246356 218696
rect 246960 217274 246988 220730
rect 248340 218074 248368 224606
rect 249076 218210 249104 227802
rect 249260 225894 249288 231662
rect 249432 227316 249484 227322
rect 249432 227258 249484 227264
rect 249248 225888 249300 225894
rect 249248 225830 249300 225836
rect 249444 223666 249472 227258
rect 249260 223638 249472 223666
rect 249064 218204 249116 218210
rect 249064 218146 249116 218152
rect 249260 218074 249288 223638
rect 249432 223576 249484 223582
rect 249432 223518 249484 223524
rect 247776 218068 247828 218074
rect 247776 218010 247828 218016
rect 248328 218068 248380 218074
rect 248328 218010 248380 218016
rect 248604 218068 248656 218074
rect 248604 218010 248656 218016
rect 249248 218068 249300 218074
rect 249248 218010 249300 218016
rect 246086 217110 246160 217138
rect 246914 217246 246988 217274
rect 246086 216988 246114 217110
rect 246914 216988 246942 217246
rect 247788 217138 247816 218010
rect 248616 217138 248644 218010
rect 249444 217274 249472 223518
rect 249996 222766 250024 231676
rect 250640 224126 250668 231676
rect 251284 228002 251312 231676
rect 251272 227996 251324 228002
rect 251272 227938 251324 227944
rect 251928 227458 251956 231676
rect 252586 231662 252784 231690
rect 251916 227452 251968 227458
rect 251916 227394 251968 227400
rect 252468 226024 252520 226030
rect 252468 225966 252520 225972
rect 251088 225752 251140 225758
rect 251088 225694 251140 225700
rect 250628 224120 250680 224126
rect 250628 224062 250680 224068
rect 250904 223304 250956 223310
rect 250904 223246 250956 223252
rect 249984 222760 250036 222766
rect 249984 222702 250036 222708
rect 250916 218074 250944 223246
rect 250260 218068 250312 218074
rect 250260 218010 250312 218016
rect 250904 218068 250956 218074
rect 250904 218010 250956 218016
rect 247742 217110 247816 217138
rect 248570 217110 248644 217138
rect 249398 217246 249472 217274
rect 247742 216988 247770 217110
rect 248570 216988 248598 217110
rect 249398 216988 249426 217246
rect 250272 217138 250300 218010
rect 251100 217274 251128 225694
rect 252480 218074 252508 225966
rect 252756 219842 252784 231662
rect 252940 231662 253230 231690
rect 252940 222154 252968 231662
rect 253860 227866 253888 231676
rect 253848 227860 253900 227866
rect 253848 227802 253900 227808
rect 254504 225214 254532 231676
rect 254952 228268 255004 228274
rect 254952 228210 255004 228216
rect 254492 225208 254544 225214
rect 254492 225150 254544 225156
rect 252928 222148 252980 222154
rect 252928 222090 252980 222096
rect 253388 220924 253440 220930
rect 253388 220866 253440 220872
rect 252744 219836 252796 219842
rect 252744 219778 252796 219784
rect 253400 219026 253428 220866
rect 254400 220652 254452 220658
rect 254400 220594 254452 220600
rect 253572 219972 253624 219978
rect 253572 219914 253624 219920
rect 253388 219020 253440 219026
rect 253388 218962 253440 218968
rect 252744 218748 252796 218754
rect 252744 218690 252796 218696
rect 251916 218068 251968 218074
rect 251916 218010 251968 218016
rect 252468 218068 252520 218074
rect 252468 218010 252520 218016
rect 250226 217110 250300 217138
rect 251054 217246 251128 217274
rect 250226 216988 250254 217110
rect 251054 216988 251082 217246
rect 251928 217138 251956 218010
rect 252756 217138 252784 218690
rect 253584 217274 253612 219914
rect 254412 217274 254440 220594
rect 254964 219434 254992 228210
rect 255148 226302 255176 231676
rect 255136 226296 255188 226302
rect 255136 226238 255188 226244
rect 255792 223990 255820 231676
rect 256436 230450 256464 231676
rect 256424 230444 256476 230450
rect 256424 230386 256476 230392
rect 256516 229764 256568 229770
rect 256516 229706 256568 229712
rect 255780 223984 255832 223990
rect 255780 223926 255832 223932
rect 254964 219406 255176 219434
rect 251882 217110 251956 217138
rect 252710 217110 252784 217138
rect 253538 217246 253612 217274
rect 254366 217246 254440 217274
rect 255148 217274 255176 219406
rect 256528 218074 256556 229706
rect 257080 229090 257108 231676
rect 257264 231662 257738 231690
rect 257068 229084 257120 229090
rect 257068 229026 257120 229032
rect 257264 219706 257292 231662
rect 257528 229084 257580 229090
rect 257528 229026 257580 229032
rect 257252 219700 257304 219706
rect 257252 219642 257304 219648
rect 257540 218074 257568 229026
rect 257712 228948 257764 228954
rect 257712 228890 257764 228896
rect 256056 218068 256108 218074
rect 256056 218010 256108 218016
rect 256516 218068 256568 218074
rect 256516 218010 256568 218016
rect 256884 218068 256936 218074
rect 256884 218010 256936 218016
rect 257528 218068 257580 218074
rect 257528 218010 257580 218016
rect 255148 217246 255222 217274
rect 251882 216988 251910 217110
rect 252710 216988 252738 217110
rect 253538 216988 253566 217246
rect 254366 216988 254394 217246
rect 255194 216988 255222 217246
rect 256068 217138 256096 218010
rect 256896 217138 256924 218010
rect 257724 217274 257752 228890
rect 258368 222494 258396 231676
rect 258644 231662 259026 231690
rect 258356 222488 258408 222494
rect 258356 222430 258408 222436
rect 258080 222148 258132 222154
rect 258080 222090 258132 222096
rect 258092 219434 258120 222090
rect 258644 220930 258672 231662
rect 259368 226636 259420 226642
rect 259368 226578 259420 226584
rect 258632 220924 258684 220930
rect 258632 220866 258684 220872
rect 258080 219428 258132 219434
rect 258080 219370 258132 219376
rect 259184 219020 259236 219026
rect 259184 218962 259236 218968
rect 258540 218068 258592 218074
rect 258540 218010 258592 218016
rect 256022 217110 256096 217138
rect 256850 217110 256924 217138
rect 257678 217246 257752 217274
rect 256022 216988 256050 217110
rect 256850 216988 256878 217110
rect 257678 216988 257706 217246
rect 258552 217138 258580 218010
rect 259196 217274 259224 218962
rect 259380 218074 259408 226578
rect 259656 225486 259684 231676
rect 260300 228546 260328 231676
rect 260944 229094 260972 231676
rect 261588 230314 261616 231676
rect 261576 230308 261628 230314
rect 261576 230250 261628 230256
rect 260852 229066 260972 229094
rect 260288 228540 260340 228546
rect 260288 228482 260340 228488
rect 260656 226296 260708 226302
rect 260656 226238 260708 226244
rect 259644 225480 259696 225486
rect 259644 225422 259696 225428
rect 260668 219434 260696 226238
rect 260852 221202 260880 229066
rect 262232 227594 262260 231676
rect 262416 231662 262890 231690
rect 263152 231662 263534 231690
rect 263888 231662 264178 231690
rect 262220 227588 262272 227594
rect 262220 227530 262272 227536
rect 261852 225888 261904 225894
rect 261852 225830 261904 225836
rect 261024 222012 261076 222018
rect 261024 221954 261076 221960
rect 260840 221196 260892 221202
rect 260840 221138 260892 221144
rect 260668 219406 260788 219434
rect 260760 218074 260788 219406
rect 259368 218068 259420 218074
rect 259368 218010 259420 218016
rect 260196 218068 260248 218074
rect 260196 218010 260248 218016
rect 260748 218068 260800 218074
rect 260748 218010 260800 218016
rect 259196 217246 259362 217274
rect 258506 217110 258580 217138
rect 258506 216988 258534 217110
rect 259334 216988 259362 217246
rect 260208 217138 260236 218010
rect 261036 217274 261064 221954
rect 261864 217274 261892 225830
rect 262416 220386 262444 231662
rect 263152 221746 263180 231662
rect 263888 222154 263916 231662
rect 264244 230172 264296 230178
rect 264244 230114 264296 230120
rect 263876 222148 263928 222154
rect 263876 222090 263928 222096
rect 263140 221740 263192 221746
rect 263140 221682 263192 221688
rect 263508 221740 263560 221746
rect 263508 221682 263560 221688
rect 262404 220380 262456 220386
rect 262404 220322 262456 220328
rect 262680 220380 262732 220386
rect 262680 220322 262732 220328
rect 262692 217274 262720 220322
rect 263520 217274 263548 221682
rect 264256 220386 264284 230114
rect 264808 228682 264836 231676
rect 265176 231662 265466 231690
rect 264796 228676 264848 228682
rect 264796 228618 264848 228624
rect 264796 227452 264848 227458
rect 264796 227394 264848 227400
rect 264244 220380 264296 220386
rect 264244 220322 264296 220328
rect 264612 220380 264664 220386
rect 264612 220322 264664 220328
rect 264624 218618 264652 220322
rect 264612 218612 264664 218618
rect 264612 218554 264664 218560
rect 264808 218074 264836 227394
rect 265176 220250 265204 231662
rect 266096 225622 266124 231676
rect 266740 229634 266768 231676
rect 266728 229628 266780 229634
rect 266728 229570 266780 229576
rect 267384 226914 267412 231676
rect 268028 227730 268056 231676
rect 268212 231662 268686 231690
rect 268016 227724 268068 227730
rect 268016 227666 268068 227672
rect 267372 226908 267424 226914
rect 267372 226850 267424 226856
rect 266084 225616 266136 225622
rect 266084 225558 266136 225564
rect 267004 225616 267056 225622
rect 267004 225558 267056 225564
rect 266268 224120 266320 224126
rect 266268 224062 266320 224068
rect 265164 220244 265216 220250
rect 265164 220186 265216 220192
rect 265992 218612 266044 218618
rect 265992 218554 266044 218560
rect 264336 218068 264388 218074
rect 264336 218010 264388 218016
rect 264796 218068 264848 218074
rect 264796 218010 264848 218016
rect 265164 218068 265216 218074
rect 265164 218010 265216 218016
rect 260162 217110 260236 217138
rect 260990 217246 261064 217274
rect 261818 217246 261892 217274
rect 262646 217246 262720 217274
rect 263474 217246 263548 217274
rect 260162 216988 260190 217110
rect 260990 216988 261018 217246
rect 261818 216988 261846 217246
rect 262646 216988 262674 217246
rect 263474 216988 263502 217246
rect 264348 217138 264376 218010
rect 265176 217138 265204 218010
rect 266004 217138 266032 218554
rect 266280 218074 266308 224062
rect 266820 221332 266872 221338
rect 266820 221274 266872 221280
rect 266268 218068 266320 218074
rect 266268 218010 266320 218016
rect 266832 217274 266860 221274
rect 267016 218482 267044 225558
rect 268212 221066 268240 231662
rect 268936 228540 268988 228546
rect 268936 228482 268988 228488
rect 268200 221060 268252 221066
rect 268200 221002 268252 221008
rect 267648 220244 267700 220250
rect 267648 220186 267700 220192
rect 267004 218476 267056 218482
rect 267004 218418 267056 218424
rect 267660 217274 267688 220186
rect 268948 218074 268976 228482
rect 269316 220386 269344 231676
rect 269960 226166 269988 231676
rect 269948 226160 270000 226166
rect 269948 226102 270000 226108
rect 270224 226160 270276 226166
rect 270224 226102 270276 226108
rect 270040 222148 270092 222154
rect 270040 222090 270092 222096
rect 269304 220380 269356 220386
rect 269304 220322 269356 220328
rect 268476 218068 268528 218074
rect 268476 218010 268528 218016
rect 268936 218068 268988 218074
rect 268936 218010 268988 218016
rect 269304 218068 269356 218074
rect 269304 218010 269356 218016
rect 264302 217110 264376 217138
rect 265130 217110 265204 217138
rect 265958 217110 266032 217138
rect 266786 217246 266860 217274
rect 267614 217246 267688 217274
rect 264302 216988 264330 217110
rect 265130 216988 265158 217110
rect 265958 216988 265986 217110
rect 266786 216988 266814 217246
rect 267614 216988 267642 217246
rect 268488 217138 268516 218010
rect 269316 217138 269344 218010
rect 270052 217274 270080 222090
rect 270236 218074 270264 226102
rect 270604 220522 270632 231676
rect 271248 227050 271276 231676
rect 271892 229498 271920 231676
rect 271880 229492 271932 229498
rect 271880 229434 271932 229440
rect 272536 228138 272564 231676
rect 272524 228132 272576 228138
rect 272524 228074 272576 228080
rect 271236 227044 271288 227050
rect 271236 226986 271288 226992
rect 271788 227044 271840 227050
rect 271788 226986 271840 226992
rect 270592 220516 270644 220522
rect 270592 220458 270644 220464
rect 270776 219564 270828 219570
rect 270776 219506 270828 219512
rect 270788 218346 270816 219506
rect 270776 218340 270828 218346
rect 270776 218282 270828 218288
rect 270224 218068 270276 218074
rect 270224 218010 270276 218016
rect 270960 218068 271012 218074
rect 270960 218010 271012 218016
rect 270052 217246 270126 217274
rect 268442 217110 268516 217138
rect 269270 217110 269344 217138
rect 268442 216988 268470 217110
rect 269270 216988 269298 217110
rect 270098 216988 270126 217246
rect 270972 217138 271000 218010
rect 271800 217274 271828 226986
rect 272524 224936 272576 224942
rect 272524 224878 272576 224884
rect 272340 219156 272392 219162
rect 272340 219098 272392 219104
rect 272352 218618 272380 219098
rect 272340 218612 272392 218618
rect 272340 218554 272392 218560
rect 272536 218074 272564 224878
rect 273180 223854 273208 231676
rect 273824 228410 273852 231676
rect 273812 228404 273864 228410
rect 273812 228346 273864 228352
rect 274272 228404 274324 228410
rect 274272 228346 274324 228352
rect 273168 223848 273220 223854
rect 273168 223790 273220 223796
rect 273444 220380 273496 220386
rect 273444 220322 273496 220328
rect 272892 219428 272944 219434
rect 272892 219370 272944 219376
rect 272708 219292 272760 219298
rect 272708 219234 272760 219240
rect 272720 218618 272748 219234
rect 272708 218612 272760 218618
rect 272708 218554 272760 218560
rect 272524 218068 272576 218074
rect 272524 218010 272576 218016
rect 272904 217274 272932 219370
rect 273456 217274 273484 220322
rect 274284 217274 274312 228346
rect 274468 225622 274496 231676
rect 275112 229094 275140 231676
rect 274928 229066 275140 229094
rect 275296 231662 275770 231690
rect 276124 231662 276414 231690
rect 274456 225616 274508 225622
rect 274456 225558 274508 225564
rect 274928 224534 274956 229066
rect 274916 224528 274968 224534
rect 274916 224470 274968 224476
rect 275100 224528 275152 224534
rect 275100 224470 275152 224476
rect 275112 217274 275140 224470
rect 275296 220114 275324 231662
rect 275652 230308 275704 230314
rect 275652 230250 275704 230256
rect 275664 229094 275692 230250
rect 275664 229066 275876 229094
rect 275284 220108 275336 220114
rect 275284 220050 275336 220056
rect 270926 217110 271000 217138
rect 271754 217246 271828 217274
rect 272582 217246 272932 217274
rect 273410 217246 273484 217274
rect 274238 217246 274312 217274
rect 275066 217246 275140 217274
rect 275848 217274 275876 229066
rect 276124 221474 276152 231662
rect 276296 230444 276348 230450
rect 276296 230386 276348 230392
rect 276308 223582 276336 230386
rect 277044 229906 277072 231676
rect 277032 229900 277084 229906
rect 277032 229842 277084 229848
rect 277688 224398 277716 231676
rect 277964 231662 278346 231690
rect 277676 224392 277728 224398
rect 277676 224334 277728 224340
rect 276296 223576 276348 223582
rect 276296 223518 276348 223524
rect 277964 221882 277992 231662
rect 278412 225616 278464 225622
rect 278412 225558 278464 225564
rect 277952 221876 278004 221882
rect 277952 221818 278004 221824
rect 276112 221468 276164 221474
rect 276112 221410 276164 221416
rect 276756 220108 276808 220114
rect 276756 220050 276808 220056
rect 276768 217274 276796 220050
rect 277584 218068 277636 218074
rect 277584 218010 277636 218016
rect 275848 217246 275922 217274
rect 270926 216988 270954 217110
rect 271754 216988 271782 217246
rect 272582 216988 272610 217246
rect 273410 216988 273438 217246
rect 274238 216988 274266 217246
rect 275066 216988 275094 217246
rect 275894 216988 275922 217246
rect 276722 217246 276796 217274
rect 276722 216988 276750 217246
rect 277596 217138 277624 218010
rect 278424 217274 278452 225558
rect 278976 224262 279004 231676
rect 279160 231662 279634 231690
rect 278964 224256 279016 224262
rect 278964 224198 279016 224204
rect 278596 223576 278648 223582
rect 278596 223518 278648 223524
rect 278608 218074 278636 223518
rect 279160 219570 279188 231662
rect 280264 226778 280292 231676
rect 280252 226772 280304 226778
rect 280252 226714 280304 226720
rect 279424 223916 279476 223922
rect 279424 223858 279476 223864
rect 279148 219564 279200 219570
rect 279148 219506 279200 219512
rect 279056 219156 279108 219162
rect 279056 219098 279108 219104
rect 279068 218890 279096 219098
rect 279056 218884 279108 218890
rect 279056 218826 279108 218832
rect 279240 218884 279292 218890
rect 279240 218826 279292 218832
rect 278596 218068 278648 218074
rect 278596 218010 278648 218016
rect 277550 217110 277624 217138
rect 278378 217246 278452 217274
rect 277550 216988 277578 217110
rect 278378 216988 278406 217246
rect 279252 217138 279280 218826
rect 279436 218618 279464 223858
rect 280908 222358 280936 231676
rect 281356 227588 281408 227594
rect 281356 227530 281408 227536
rect 280896 222352 280948 222358
rect 280896 222294 280948 222300
rect 280068 221876 280120 221882
rect 280068 221818 280120 221824
rect 279424 218612 279476 218618
rect 279424 218554 279476 218560
rect 280080 217274 280108 221818
rect 281368 219434 281396 227530
rect 281552 222902 281580 231676
rect 282196 229362 282224 231676
rect 282552 229900 282604 229906
rect 282552 229842 282604 229848
rect 282184 229356 282236 229362
rect 282184 229298 282236 229304
rect 281540 222896 281592 222902
rect 281540 222838 281592 222844
rect 281368 219406 281488 219434
rect 281460 218074 281488 219406
rect 280896 218068 280948 218074
rect 280896 218010 280948 218016
rect 281448 218068 281500 218074
rect 281448 218010 281500 218016
rect 281724 218068 281776 218074
rect 281724 218010 281776 218016
rect 279206 217110 279280 217138
rect 280034 217246 280108 217274
rect 279206 216988 279234 217110
rect 280034 216988 280062 217246
rect 280908 217138 280936 218010
rect 281736 217138 281764 218010
rect 282564 217274 282592 229842
rect 282840 228818 282868 231676
rect 282828 228812 282880 228818
rect 282828 228754 282880 228760
rect 283484 223174 283512 231676
rect 283760 231662 284142 231690
rect 283472 223168 283524 223174
rect 283472 223110 283524 223116
rect 282736 222896 282788 222902
rect 282736 222838 282788 222844
rect 282748 218074 282776 222838
rect 283760 221610 283788 231662
rect 284772 223922 284800 231676
rect 285048 231662 285430 231690
rect 285048 225350 285076 231662
rect 285496 228676 285548 228682
rect 285496 228618 285548 228624
rect 285036 225344 285088 225350
rect 285036 225286 285088 225292
rect 284760 223916 284812 223922
rect 284760 223858 284812 223864
rect 284208 222760 284260 222766
rect 284208 222702 284260 222708
rect 283748 221604 283800 221610
rect 283748 221546 283800 221552
rect 284024 221468 284076 221474
rect 284024 221410 284076 221416
rect 284036 219434 284064 221410
rect 284036 219406 284156 219434
rect 282736 218068 282788 218074
rect 282736 218010 282788 218016
rect 283380 218068 283432 218074
rect 283380 218010 283432 218016
rect 280862 217110 280936 217138
rect 281690 217110 281764 217138
rect 282518 217246 282592 217274
rect 280862 216988 280890 217110
rect 281690 216988 281718 217110
rect 282518 216988 282546 217246
rect 283392 217138 283420 218010
rect 284128 217274 284156 219406
rect 284220 218090 284248 222702
rect 284220 218074 284340 218090
rect 285508 218074 285536 228618
rect 286060 223446 286088 231676
rect 286704 227186 286732 231676
rect 287348 230042 287376 231676
rect 287716 231662 288006 231690
rect 287336 230036 287388 230042
rect 287336 229978 287388 229984
rect 287520 230036 287572 230042
rect 287520 229978 287572 229984
rect 286692 227180 286744 227186
rect 286692 227122 286744 227128
rect 287532 226166 287560 229978
rect 287520 226160 287572 226166
rect 287520 226102 287572 226108
rect 287716 224806 287744 231662
rect 288072 226160 288124 226166
rect 288072 226102 288124 226108
rect 287704 224800 287756 224806
rect 287704 224742 287756 224748
rect 286324 224392 286376 224398
rect 286324 224334 286376 224340
rect 286048 223440 286100 223446
rect 286048 223382 286100 223388
rect 286336 219162 286364 224334
rect 286692 219836 286744 219842
rect 286692 219778 286744 219784
rect 286324 219156 286376 219162
rect 286324 219098 286376 219104
rect 285864 218884 285916 218890
rect 285864 218826 285916 218832
rect 284220 218068 284352 218074
rect 284220 218062 284300 218068
rect 284300 218010 284352 218016
rect 285036 218068 285088 218074
rect 285036 218010 285088 218016
rect 285496 218068 285548 218074
rect 285496 218010 285548 218016
rect 284128 217246 284202 217274
rect 283346 217110 283420 217138
rect 283346 216988 283374 217110
rect 284174 216988 284202 217246
rect 285048 217138 285076 218010
rect 285876 217138 285904 218826
rect 286704 217274 286732 219778
rect 288084 218074 288112 226102
rect 288256 223168 288308 223174
rect 288256 223110 288308 223116
rect 287520 218068 287572 218074
rect 287520 218010 287572 218016
rect 288072 218068 288124 218074
rect 288072 218010 288124 218016
rect 285002 217110 285076 217138
rect 285830 217110 285904 217138
rect 286658 217246 286732 217274
rect 285002 216988 285030 217110
rect 285830 216988 285858 217110
rect 286658 216988 286686 217246
rect 287532 217138 287560 218010
rect 288268 217274 288296 223110
rect 288636 220794 288664 231676
rect 288992 223304 289044 223310
rect 288992 223246 289044 223252
rect 288624 220788 288676 220794
rect 288624 220730 288676 220736
rect 289004 218482 289032 223246
rect 289280 223038 289308 231676
rect 289924 224398 289952 231676
rect 290568 227322 290596 231676
rect 290556 227316 290608 227322
rect 290556 227258 290608 227264
rect 291016 227316 291068 227322
rect 291016 227258 291068 227264
rect 289912 224392 289964 224398
rect 289912 224334 289964 224340
rect 290832 224392 290884 224398
rect 290832 224334 290884 224340
rect 289636 224256 289688 224262
rect 289636 224198 289688 224204
rect 289268 223032 289320 223038
rect 289268 222974 289320 222980
rect 288992 218476 289044 218482
rect 288992 218418 289044 218424
rect 289648 218074 289676 224198
rect 289820 219564 289872 219570
rect 289820 219506 289872 219512
rect 289832 219298 289860 219506
rect 289820 219292 289872 219298
rect 289820 219234 289872 219240
rect 289176 218068 289228 218074
rect 289176 218010 289228 218016
rect 289636 218068 289688 218074
rect 289636 218010 289688 218016
rect 290004 218068 290056 218074
rect 290004 218010 290056 218016
rect 288268 217246 288342 217274
rect 287486 217110 287560 217138
rect 287486 216988 287514 217110
rect 288314 216988 288342 217246
rect 289188 217138 289216 218010
rect 290016 217138 290044 218010
rect 290844 217274 290872 224334
rect 291028 219434 291056 227258
rect 291212 223446 291240 231676
rect 291856 224670 291884 231676
rect 292500 230450 292528 231676
rect 292488 230444 292540 230450
rect 292488 230386 292540 230392
rect 293144 226030 293172 231676
rect 293328 231662 293802 231690
rect 293132 226024 293184 226030
rect 293132 225966 293184 225972
rect 291844 224664 291896 224670
rect 291844 224606 291896 224612
rect 291200 223440 291252 223446
rect 291200 223382 291252 223388
rect 291660 223032 291712 223038
rect 291660 222974 291712 222980
rect 291028 219406 291148 219434
rect 291120 218074 291148 219406
rect 291672 219026 291700 222974
rect 292488 220516 292540 220522
rect 292488 220458 292540 220464
rect 292028 219292 292080 219298
rect 292028 219234 292080 219240
rect 291660 219020 291712 219026
rect 291660 218962 291712 218968
rect 292040 218890 292068 219234
rect 292028 218884 292080 218890
rect 292028 218826 292080 218832
rect 291660 218748 291712 218754
rect 291660 218690 291712 218696
rect 291108 218068 291160 218074
rect 291108 218010 291160 218016
rect 291672 217274 291700 218690
rect 292500 217274 292528 220458
rect 293328 219978 293356 231662
rect 293776 227724 293828 227730
rect 293776 227666 293828 227672
rect 293316 219972 293368 219978
rect 293316 219914 293368 219920
rect 293788 218074 293816 227666
rect 294432 225758 294460 231676
rect 294420 225752 294472 225758
rect 294420 225694 294472 225700
rect 294880 224664 294932 224670
rect 294880 224606 294932 224612
rect 294892 219434 294920 224606
rect 295076 223310 295104 231676
rect 295720 228274 295748 231676
rect 296364 229090 296392 231676
rect 296824 231662 297022 231690
rect 296352 229084 296404 229090
rect 296352 229026 296404 229032
rect 296628 228812 296680 228818
rect 296628 228754 296680 228760
rect 295708 228268 295760 228274
rect 295708 228210 295760 228216
rect 296444 225752 296496 225758
rect 296444 225694 296496 225700
rect 295064 223304 295116 223310
rect 295064 223246 295116 223252
rect 296456 219434 296484 225694
rect 294892 219406 295012 219434
rect 296456 219406 296576 219434
rect 294144 218476 294196 218482
rect 294144 218418 294196 218424
rect 293316 218068 293368 218074
rect 293316 218010 293368 218016
rect 293776 218068 293828 218074
rect 293776 218010 293828 218016
rect 289142 217110 289216 217138
rect 289970 217110 290044 217138
rect 290798 217246 290872 217274
rect 291626 217246 291700 217274
rect 292454 217246 292528 217274
rect 289142 216988 289170 217110
rect 289970 216988 289998 217110
rect 290798 216988 290826 217246
rect 291626 216988 291654 217246
rect 292454 216988 292482 217246
rect 293328 217138 293356 218010
rect 294156 217138 294184 218418
rect 294984 217274 295012 219406
rect 295800 219156 295852 219162
rect 295800 219098 295852 219104
rect 293282 217110 293356 217138
rect 294110 217110 294184 217138
rect 294938 217246 295012 217274
rect 293282 216988 293310 217110
rect 294110 216988 294138 217110
rect 294938 216988 294966 217246
rect 295812 217138 295840 219098
rect 296548 217274 296576 219406
rect 296640 219178 296668 228754
rect 296824 220658 296852 231662
rect 297652 229770 297680 231676
rect 297640 229764 297692 229770
rect 297640 229706 297692 229712
rect 296996 229628 297048 229634
rect 296996 229570 297048 229576
rect 297008 224262 297036 229570
rect 298296 226642 298324 231676
rect 298284 226636 298336 226642
rect 298284 226578 298336 226584
rect 298940 226302 298968 231676
rect 299584 228954 299612 231676
rect 299572 228948 299624 228954
rect 299572 228890 299624 228896
rect 298928 226296 298980 226302
rect 298928 226238 298980 226244
rect 299388 226024 299440 226030
rect 299388 225966 299440 225972
rect 297364 225480 297416 225486
rect 297364 225422 297416 225428
rect 296996 224256 297048 224262
rect 296996 224198 297048 224204
rect 296812 220652 296864 220658
rect 296812 220594 296864 220600
rect 296640 219162 296760 219178
rect 296640 219156 296772 219162
rect 296640 219150 296720 219156
rect 296720 219098 296772 219104
rect 297376 219026 297404 225422
rect 299112 224256 299164 224262
rect 299112 224198 299164 224204
rect 297548 223372 297600 223378
rect 297548 223314 297600 223320
rect 297560 219434 297588 223314
rect 297548 219428 297600 219434
rect 297548 219370 297600 219376
rect 297364 219020 297416 219026
rect 297364 218962 297416 218968
rect 297456 218204 297508 218210
rect 297456 218146 297508 218152
rect 296548 217246 296622 217274
rect 295766 217110 295840 217138
rect 295766 216988 295794 217110
rect 296594 216988 296622 217246
rect 297468 217138 297496 218146
rect 298284 218068 298336 218074
rect 298284 218010 298336 218016
rect 298296 217138 298324 218010
rect 299124 217274 299152 224198
rect 299400 218074 299428 225966
rect 300228 223038 300256 231676
rect 300676 228948 300728 228954
rect 300676 228890 300728 228896
rect 300216 223032 300268 223038
rect 300216 222974 300268 222980
rect 300492 219156 300544 219162
rect 300492 219098 300544 219104
rect 299388 218068 299440 218074
rect 299388 218010 299440 218016
rect 299940 218068 299992 218074
rect 299940 218010 299992 218016
rect 297422 217110 297496 217138
rect 298250 217110 298324 217138
rect 299078 217246 299152 217274
rect 297422 216988 297450 217110
rect 298250 216988 298278 217110
rect 299078 216988 299106 217246
rect 299952 217138 299980 218010
rect 300504 217274 300532 219098
rect 300688 218074 300716 228890
rect 300872 225894 300900 231676
rect 301056 231662 301530 231690
rect 301700 231662 302174 231690
rect 300860 225888 300912 225894
rect 300860 225830 300912 225836
rect 301056 221746 301084 231662
rect 301700 222018 301728 231662
rect 302804 230178 302832 231676
rect 302792 230172 302844 230178
rect 302792 230114 302844 230120
rect 302976 230172 303028 230178
rect 302976 230114 303028 230120
rect 302148 229084 302200 229090
rect 302148 229026 302200 229032
rect 301688 222012 301740 222018
rect 301688 221954 301740 221960
rect 301044 221740 301096 221746
rect 301044 221682 301096 221688
rect 302160 218074 302188 229026
rect 302424 221604 302476 221610
rect 302424 221546 302476 221552
rect 300676 218068 300728 218074
rect 300676 218010 300728 218016
rect 301596 218068 301648 218074
rect 301596 218010 301648 218016
rect 302148 218068 302200 218074
rect 302148 218010 302200 218016
rect 300504 217246 300762 217274
rect 299906 217110 299980 217138
rect 299906 216988 299934 217110
rect 300734 216988 300762 217246
rect 301608 217138 301636 218010
rect 302436 217274 302464 221546
rect 302988 219434 303016 230114
rect 303448 224126 303476 231676
rect 303816 231662 304106 231690
rect 303436 224120 303488 224126
rect 303436 224062 303488 224068
rect 303252 221740 303304 221746
rect 303252 221682 303304 221688
rect 302896 219406 303016 219434
rect 302896 218210 302924 219406
rect 302884 218204 302936 218210
rect 302884 218146 302936 218152
rect 303264 217274 303292 221682
rect 303816 221338 303844 231662
rect 304736 227458 304764 231676
rect 304724 227452 304776 227458
rect 304724 227394 304776 227400
rect 304264 224120 304316 224126
rect 304264 224062 304316 224068
rect 303804 221332 303856 221338
rect 303804 221274 303856 221280
rect 304080 219428 304132 219434
rect 304080 219370 304132 219376
rect 301562 217110 301636 217138
rect 302390 217246 302464 217274
rect 303218 217246 303292 217274
rect 301562 216988 301590 217110
rect 302390 216988 302418 217246
rect 303218 216988 303246 217246
rect 304092 217138 304120 219370
rect 304276 218618 304304 224062
rect 305380 223378 305408 231676
rect 306024 228546 306052 231676
rect 306392 231662 306682 231690
rect 306852 231662 307326 231690
rect 306012 228540 306064 228546
rect 306012 228482 306064 228488
rect 306196 227180 306248 227186
rect 306196 227122 306248 227128
rect 305368 223372 305420 223378
rect 305368 223314 305420 223320
rect 304908 220652 304960 220658
rect 304908 220594 304960 220600
rect 304264 218612 304316 218618
rect 304264 218554 304316 218560
rect 304920 217274 304948 220594
rect 306208 218074 306236 227122
rect 306392 222154 306420 231662
rect 306380 222148 306432 222154
rect 306380 222090 306432 222096
rect 306852 220250 306880 231662
rect 307956 230042 307984 231676
rect 308404 230444 308456 230450
rect 308404 230386 308456 230392
rect 307944 230036 307996 230042
rect 307944 229978 307996 229984
rect 307668 223304 307720 223310
rect 307668 223246 307720 223252
rect 306840 220244 306892 220250
rect 306840 220186 306892 220192
rect 307392 219020 307444 219026
rect 307392 218962 307444 218968
rect 305736 218068 305788 218074
rect 305736 218010 305788 218016
rect 306196 218068 306248 218074
rect 306196 218010 306248 218016
rect 306564 218068 306616 218074
rect 306564 218010 306616 218016
rect 304046 217110 304120 217138
rect 304874 217246 304948 217274
rect 304046 216988 304074 217110
rect 304874 216988 304902 217246
rect 305748 217138 305776 218010
rect 306576 217138 306604 218010
rect 307404 217138 307432 218962
rect 307680 218074 307708 223246
rect 308416 219434 308444 230386
rect 308600 227050 308628 231676
rect 308588 227044 308640 227050
rect 308588 226986 308640 226992
rect 308864 226296 308916 226302
rect 308864 226238 308916 226244
rect 308404 219428 308456 219434
rect 308404 219370 308456 219376
rect 308876 218074 308904 226238
rect 309244 220386 309272 231676
rect 309888 224942 309916 231676
rect 310336 227044 310388 227050
rect 310336 226986 310388 226992
rect 309876 224936 309928 224942
rect 309876 224878 309928 224884
rect 309232 220380 309284 220386
rect 309232 220322 309284 220328
rect 309048 220244 309100 220250
rect 309048 220186 309100 220192
rect 307668 218068 307720 218074
rect 307668 218010 307720 218016
rect 308220 218068 308272 218074
rect 308220 218010 308272 218016
rect 308864 218068 308916 218074
rect 308864 218010 308916 218016
rect 308232 217138 308260 218010
rect 309060 217274 309088 220186
rect 310348 218074 310376 226986
rect 310532 225486 310560 231676
rect 310520 225480 310572 225486
rect 310520 225422 310572 225428
rect 311176 224534 311204 231676
rect 311360 231662 311834 231690
rect 311164 224528 311216 224534
rect 311164 224470 311216 224476
rect 310704 222148 310756 222154
rect 310704 222090 310756 222096
rect 309876 218068 309928 218074
rect 309876 218010 309928 218016
rect 310336 218068 310388 218074
rect 310336 218010 310388 218016
rect 305702 217110 305776 217138
rect 306530 217110 306604 217138
rect 307358 217110 307432 217138
rect 308186 217110 308260 217138
rect 309014 217246 309088 217274
rect 305702 216988 305730 217110
rect 306530 216988 306558 217110
rect 307358 216988 307386 217110
rect 308186 216988 308214 217110
rect 309014 216988 309042 217246
rect 309888 217138 309916 218010
rect 310716 217274 310744 222090
rect 311360 220114 311388 231662
rect 312464 228410 312492 231676
rect 313108 230314 313136 231676
rect 313292 231662 313766 231690
rect 313936 231662 314410 231690
rect 313096 230308 313148 230314
rect 313096 230250 313148 230256
rect 312636 230036 312688 230042
rect 312636 229978 312688 229984
rect 312452 228404 312504 228410
rect 312452 228346 312504 228352
rect 311532 224800 311584 224806
rect 311532 224742 311584 224748
rect 311348 220108 311400 220114
rect 311348 220050 311400 220056
rect 311544 217274 311572 224742
rect 312648 222154 312676 229978
rect 312912 225888 312964 225894
rect 312912 225830 312964 225836
rect 312636 222148 312688 222154
rect 312636 222090 312688 222096
rect 312924 218074 312952 225830
rect 313292 225622 313320 231662
rect 313936 229094 313964 231662
rect 313752 229066 313964 229094
rect 313280 225616 313332 225622
rect 313280 225558 313332 225564
rect 313188 222012 313240 222018
rect 313188 221954 313240 221960
rect 312360 218068 312412 218074
rect 312360 218010 312412 218016
rect 312912 218068 312964 218074
rect 312912 218010 312964 218016
rect 309842 217110 309916 217138
rect 310670 217246 310744 217274
rect 311498 217246 311572 217274
rect 309842 216988 309870 217110
rect 310670 216988 310698 217246
rect 311498 216988 311526 217246
rect 312372 217138 312400 218010
rect 313200 217274 313228 221954
rect 313752 221882 313780 229066
rect 313924 228540 313976 228546
rect 313924 228482 313976 228488
rect 313740 221876 313792 221882
rect 313740 221818 313792 221824
rect 313936 219298 313964 228482
rect 315040 223582 315068 231676
rect 315408 231662 315698 231690
rect 315408 229094 315436 231662
rect 315316 229066 315436 229094
rect 315316 224126 315344 229066
rect 315488 227452 315540 227458
rect 315488 227394 315540 227400
rect 315304 224120 315356 224126
rect 315304 224062 315356 224068
rect 315028 223576 315080 223582
rect 315028 223518 315080 223524
rect 313924 219292 313976 219298
rect 313924 219234 313976 219240
rect 314016 218884 314068 218890
rect 314016 218826 314068 218832
rect 312326 217110 312400 217138
rect 313154 217246 313228 217274
rect 312326 216988 312354 217110
rect 313154 216988 313182 217246
rect 314028 217138 314056 218826
rect 315500 218074 315528 227394
rect 315672 223032 315724 223038
rect 315672 222974 315724 222980
rect 314844 218068 314896 218074
rect 314844 218010 314896 218016
rect 315488 218068 315540 218074
rect 315488 218010 315540 218016
rect 314856 217138 314884 218010
rect 315684 217274 315712 222974
rect 316328 222902 316356 231676
rect 316684 223440 316736 223446
rect 316684 223382 316736 223388
rect 316316 222896 316368 222902
rect 316316 222838 316368 222844
rect 316500 220380 316552 220386
rect 316500 220322 316552 220328
rect 316512 217274 316540 220322
rect 316696 218482 316724 223382
rect 316972 222766 317000 231676
rect 317616 227594 317644 231676
rect 318260 229906 318288 231676
rect 318248 229900 318300 229906
rect 318248 229842 318300 229848
rect 318064 229764 318116 229770
rect 318064 229706 318116 229712
rect 317604 227588 317656 227594
rect 317604 227530 317656 227536
rect 316960 222760 317012 222766
rect 316960 222702 317012 222708
rect 318076 219434 318104 229706
rect 318904 228682 318932 231676
rect 319088 231662 319562 231690
rect 320206 231662 320404 231690
rect 318892 228676 318944 228682
rect 318892 228618 318944 228624
rect 318248 221876 318300 221882
rect 318248 221818 318300 221824
rect 318260 219434 318288 221818
rect 319088 219842 319116 231662
rect 320088 228404 320140 228410
rect 320088 228346 320140 228352
rect 319812 224936 319864 224942
rect 319812 224878 319864 224884
rect 319076 219836 319128 219842
rect 319076 219778 319128 219784
rect 317984 219406 318104 219434
rect 318168 219406 318288 219434
rect 316684 218476 316736 218482
rect 316684 218418 316736 218424
rect 317984 218074 318012 219406
rect 317328 218068 317380 218074
rect 317328 218010 317380 218016
rect 317972 218068 318024 218074
rect 317972 218010 318024 218016
rect 313982 217110 314056 217138
rect 314810 217110 314884 217138
rect 315638 217246 315712 217274
rect 316466 217246 316540 217274
rect 313982 216988 314010 217110
rect 314810 216988 314838 217110
rect 315638 216988 315666 217246
rect 316466 216988 316494 217246
rect 317340 217138 317368 218010
rect 318168 217274 318196 219406
rect 318984 218068 319036 218074
rect 318984 218010 319036 218016
rect 317294 217110 317368 217138
rect 318122 217246 318196 217274
rect 317294 216988 317322 217110
rect 318122 216988 318150 217246
rect 318996 217138 319024 218010
rect 319824 217274 319852 224878
rect 320100 218074 320128 228346
rect 320376 221474 320404 231662
rect 320836 228546 320864 231676
rect 320824 228540 320876 228546
rect 320824 228482 320876 228488
rect 321480 223174 321508 231676
rect 322124 227322 322152 231676
rect 322112 227316 322164 227322
rect 322112 227258 322164 227264
rect 322296 227316 322348 227322
rect 322296 227258 322348 227264
rect 321468 223168 321520 223174
rect 321468 223110 321520 223116
rect 321468 222896 321520 222902
rect 321468 222838 321520 222844
rect 320364 221468 320416 221474
rect 320364 221410 320416 221416
rect 320640 219428 320692 219434
rect 320640 219370 320692 219376
rect 320088 218068 320140 218074
rect 320088 218010 320140 218016
rect 318950 217110 319024 217138
rect 319778 217246 319852 217274
rect 318950 216988 318978 217110
rect 319778 216988 319806 217246
rect 320652 217138 320680 219370
rect 321480 217274 321508 222838
rect 322308 219434 322336 227258
rect 322768 226166 322796 231676
rect 323412 229634 323440 231676
rect 323400 229628 323452 229634
rect 323400 229570 323452 229576
rect 322756 226160 322808 226166
rect 322756 226102 322808 226108
rect 322848 224528 322900 224534
rect 322848 224470 322900 224476
rect 322124 219406 322336 219434
rect 322124 219162 322152 219406
rect 322112 219156 322164 219162
rect 322112 219098 322164 219104
rect 322860 218074 322888 224470
rect 324056 224398 324084 231676
rect 324228 229900 324280 229906
rect 324228 229842 324280 229848
rect 324044 224392 324096 224398
rect 324044 224334 324096 224340
rect 323952 223168 324004 223174
rect 323952 223110 324004 223116
rect 323964 218074 323992 223110
rect 324240 219434 324268 229842
rect 324700 219434 324728 231676
rect 325344 227730 325372 231676
rect 325516 228676 325568 228682
rect 325516 228618 325568 228624
rect 325332 227724 325384 227730
rect 325332 227666 325384 227672
rect 324148 219406 324268 219434
rect 324608 219406 324728 219434
rect 322296 218068 322348 218074
rect 322296 218010 322348 218016
rect 322848 218068 322900 218074
rect 322848 218010 322900 218016
rect 323124 218068 323176 218074
rect 323124 218010 323176 218016
rect 323952 218068 324004 218074
rect 323952 218010 324004 218016
rect 320606 217110 320680 217138
rect 321434 217246 321508 217274
rect 320606 216988 320634 217110
rect 321434 216988 321462 217246
rect 322308 217138 322336 218010
rect 323136 217138 323164 218010
rect 324148 217274 324176 219406
rect 324608 218754 324636 219406
rect 325332 219156 325384 219162
rect 325332 219098 325384 219104
rect 324596 218748 324648 218754
rect 324596 218690 324648 218696
rect 324780 218068 324832 218074
rect 324780 218010 324832 218016
rect 322262 217110 322336 217138
rect 323090 217110 323164 217138
rect 323918 217246 324176 217274
rect 322262 216988 322290 217110
rect 323090 216988 323118 217110
rect 323918 216988 323946 217246
rect 324792 217138 324820 218010
rect 325344 217274 325372 219098
rect 325528 218074 325556 228618
rect 325988 224670 326016 231676
rect 326172 231662 326646 231690
rect 325976 224664 326028 224670
rect 325976 224606 326028 224612
rect 326172 220522 326200 231662
rect 326896 228540 326948 228546
rect 326896 228482 326948 228488
rect 326160 220516 326212 220522
rect 326160 220458 326212 220464
rect 326908 218074 326936 228482
rect 327276 223446 327304 231676
rect 327920 225758 327948 231676
rect 328564 226030 328592 231676
rect 329208 228818 329236 231676
rect 329852 230178 329880 231676
rect 329840 230172 329892 230178
rect 329840 230114 329892 230120
rect 330496 228954 330524 231676
rect 331140 229090 331168 231676
rect 331128 229084 331180 229090
rect 331128 229026 331180 229032
rect 330484 228948 330536 228954
rect 330484 228890 330536 228896
rect 329196 228812 329248 228818
rect 329196 228754 329248 228760
rect 331036 227792 331088 227798
rect 331036 227734 331088 227740
rect 328552 226024 328604 226030
rect 328552 225966 328604 225972
rect 327908 225752 327960 225758
rect 327908 225694 327960 225700
rect 329748 225752 329800 225758
rect 329748 225694 329800 225700
rect 327724 225616 327776 225622
rect 327724 225558 327776 225564
rect 327264 223440 327316 223446
rect 327264 223382 327316 223388
rect 327736 219162 327764 225558
rect 328092 220516 328144 220522
rect 328092 220458 328144 220464
rect 327724 219156 327776 219162
rect 327724 219098 327776 219104
rect 327264 218748 327316 218754
rect 327264 218690 327316 218696
rect 325516 218068 325568 218074
rect 325516 218010 325568 218016
rect 326436 218068 326488 218074
rect 326436 218010 326488 218016
rect 326896 218068 326948 218074
rect 326896 218010 326948 218016
rect 325344 217246 325602 217274
rect 324746 217110 324820 217138
rect 324746 216988 324774 217110
rect 325574 216988 325602 217246
rect 326448 217138 326476 218010
rect 327276 217138 327304 218690
rect 328104 217274 328132 220458
rect 328920 220108 328972 220114
rect 328920 220050 328972 220056
rect 328932 217274 328960 220050
rect 329760 217274 329788 225694
rect 331048 218074 331076 227734
rect 331784 224262 331812 231676
rect 332428 227322 332456 231676
rect 332796 231662 333086 231690
rect 333440 231662 333730 231690
rect 334084 231662 334374 231690
rect 332416 227316 332468 227322
rect 332416 227258 332468 227264
rect 331772 224256 331824 224262
rect 331772 224198 331824 224204
rect 331864 223984 331916 223990
rect 331864 223926 331916 223932
rect 331404 222148 331456 222154
rect 331404 222090 331456 222096
rect 330576 218068 330628 218074
rect 330576 218010 330628 218016
rect 331036 218068 331088 218074
rect 331036 218010 331088 218016
rect 326402 217110 326476 217138
rect 327230 217110 327304 217138
rect 328058 217246 328132 217274
rect 328886 217246 328960 217274
rect 329714 217246 329788 217274
rect 326402 216988 326430 217110
rect 327230 216988 327258 217110
rect 328058 216988 328086 217246
rect 328886 216988 328914 217246
rect 329714 216988 329742 217246
rect 330588 217138 330616 218010
rect 331416 217274 331444 222090
rect 331876 219026 331904 223926
rect 332796 221746 332824 231662
rect 332784 221740 332836 221746
rect 332784 221682 332836 221688
rect 333440 220658 333468 231662
rect 333888 227316 333940 227322
rect 333888 227258 333940 227264
rect 333612 221468 333664 221474
rect 333612 221410 333664 221416
rect 333428 220652 333480 220658
rect 333428 220594 333480 220600
rect 331864 219020 331916 219026
rect 331864 218962 331916 218968
rect 333428 219020 333480 219026
rect 333428 218962 333480 218968
rect 333060 218204 333112 218210
rect 333060 218146 333112 218152
rect 332232 218068 332284 218074
rect 332232 218010 332284 218016
rect 330542 217110 330616 217138
rect 331370 217246 331444 217274
rect 330542 216988 330570 217110
rect 331370 216988 331398 217246
rect 332244 217138 332272 218010
rect 333072 217138 333100 218146
rect 333440 217274 333468 218962
rect 333624 218074 333652 221410
rect 333900 218210 333928 227258
rect 334084 221610 334112 231662
rect 335004 230450 335032 231676
rect 334992 230444 335044 230450
rect 334992 230386 335044 230392
rect 334256 230172 334308 230178
rect 334256 230114 334308 230120
rect 334268 227798 334296 230114
rect 334256 227792 334308 227798
rect 334256 227734 334308 227740
rect 335176 226024 335228 226030
rect 335176 225966 335228 225972
rect 334072 221604 334124 221610
rect 334072 221546 334124 221552
rect 333888 218204 333940 218210
rect 333888 218146 333940 218152
rect 335188 218074 335216 225966
rect 335648 223310 335676 231676
rect 336292 226302 336320 231676
rect 336464 228812 336516 228818
rect 336464 228754 336516 228760
rect 336280 226296 336332 226302
rect 336280 226238 336332 226244
rect 335636 223304 335688 223310
rect 335636 223246 335688 223252
rect 336476 219434 336504 228754
rect 336936 227186 336964 231676
rect 336924 227180 336976 227186
rect 336924 227122 336976 227128
rect 337580 223990 337608 231676
rect 337752 227588 337804 227594
rect 337752 227530 337804 227536
rect 337568 223984 337620 223990
rect 337568 223926 337620 223932
rect 336384 219406 336504 219434
rect 335544 218204 335596 218210
rect 335544 218146 335596 218152
rect 333612 218068 333664 218074
rect 333612 218010 333664 218016
rect 334716 218068 334768 218074
rect 334716 218010 334768 218016
rect 335176 218068 335228 218074
rect 335176 218010 335228 218016
rect 333440 217246 333882 217274
rect 332198 217110 332272 217138
rect 333026 217110 333100 217138
rect 332198 216988 332226 217110
rect 333026 216988 333054 217110
rect 333854 216988 333882 217246
rect 334728 217138 334756 218010
rect 335556 217138 335584 218146
rect 336384 217274 336412 219406
rect 337764 218074 337792 227530
rect 338224 227050 338252 231676
rect 338212 227044 338264 227050
rect 338212 226986 338264 226992
rect 338672 227044 338724 227050
rect 338672 226986 338724 226992
rect 337936 223304 337988 223310
rect 337936 223246 337988 223252
rect 337200 218068 337252 218074
rect 337200 218010 337252 218016
rect 337752 218068 337804 218074
rect 337752 218010 337804 218016
rect 334682 217110 334756 217138
rect 335510 217110 335584 217138
rect 336338 217246 336412 217274
rect 334682 216988 334710 217110
rect 335510 216988 335538 217110
rect 336338 216988 336366 217246
rect 337212 217138 337240 218010
rect 337948 217274 337976 223246
rect 338684 218210 338712 226986
rect 338868 224806 338896 231676
rect 339526 231662 339724 231690
rect 338856 224800 338908 224806
rect 338856 224742 338908 224748
rect 339408 224256 339460 224262
rect 339408 224198 339460 224204
rect 338672 218204 338724 218210
rect 338672 218146 338724 218152
rect 339420 218074 339448 224198
rect 339696 220250 339724 231662
rect 340156 230042 340184 231676
rect 340432 231662 340814 231690
rect 340144 230036 340196 230042
rect 340144 229978 340196 229984
rect 340432 222018 340460 231662
rect 341444 227458 341472 231676
rect 341720 231662 342102 231690
rect 342364 231662 342746 231690
rect 342916 231662 343390 231690
rect 343652 231662 344034 231690
rect 341432 227452 341484 227458
rect 341432 227394 341484 227400
rect 340696 227180 340748 227186
rect 340696 227122 340748 227128
rect 340420 222012 340472 222018
rect 340420 221954 340472 221960
rect 340052 220788 340104 220794
rect 340052 220730 340104 220736
rect 339684 220244 339736 220250
rect 339684 220186 339736 220192
rect 340064 218890 340092 220730
rect 340512 219156 340564 219162
rect 340512 219098 340564 219104
rect 340052 218884 340104 218890
rect 340052 218826 340104 218832
rect 338856 218068 338908 218074
rect 338856 218010 338908 218016
rect 339408 218068 339460 218074
rect 339408 218010 339460 218016
rect 339684 218068 339736 218074
rect 339684 218010 339736 218016
rect 337948 217246 338022 217274
rect 337166 217110 337240 217138
rect 337166 216988 337194 217110
rect 337994 216988 338022 217246
rect 338868 217138 338896 218010
rect 339696 217138 339724 218010
rect 340524 217138 340552 219098
rect 340708 218074 340736 227122
rect 341720 225894 341748 231662
rect 341708 225888 341760 225894
rect 341708 225830 341760 225836
rect 341984 225888 342036 225894
rect 341984 225830 342036 225836
rect 341996 219434 342024 225830
rect 342168 224392 342220 224398
rect 342168 224334 342220 224340
rect 342180 219434 342208 224334
rect 342364 220794 342392 231662
rect 342352 220788 342404 220794
rect 342352 220730 342404 220736
rect 342916 220386 342944 231662
rect 343652 221882 343680 231662
rect 344664 223038 344692 231676
rect 345020 229764 345072 229770
rect 345020 229706 345072 229712
rect 345032 227594 345060 229706
rect 345308 229634 345336 231676
rect 345296 229628 345348 229634
rect 345296 229570 345348 229576
rect 345020 227588 345072 227594
rect 345020 227530 345072 227536
rect 345952 224942 345980 231676
rect 345940 224936 345992 224942
rect 345940 224878 345992 224884
rect 346308 224664 346360 224670
rect 346308 224606 346360 224612
rect 344652 223032 344704 223038
rect 344652 222974 344704 222980
rect 345296 222896 345348 222902
rect 345296 222838 345348 222844
rect 343640 221876 343692 221882
rect 343640 221818 343692 221824
rect 344652 221740 344704 221746
rect 344652 221682 344704 221688
rect 342904 220380 342956 220386
rect 342904 220322 342956 220328
rect 342996 220244 343048 220250
rect 342996 220186 343048 220192
rect 341340 219428 341392 219434
rect 341996 219406 342116 219434
rect 342180 219428 342312 219434
rect 342180 219406 342260 219428
rect 341340 219370 341392 219376
rect 340696 218068 340748 218074
rect 340696 218010 340748 218016
rect 341352 217138 341380 219370
rect 342088 217274 342116 219406
rect 342260 219370 342312 219376
rect 343008 217274 343036 220186
rect 343824 219428 343876 219434
rect 343824 219370 343876 219376
rect 342088 217246 342162 217274
rect 338822 217110 338896 217138
rect 339650 217110 339724 217138
rect 340478 217110 340552 217138
rect 341306 217110 341380 217138
rect 338822 216988 338850 217110
rect 339650 216988 339678 217110
rect 340478 216988 340506 217110
rect 341306 216988 341334 217110
rect 342134 216988 342162 217246
rect 342962 217246 343036 217274
rect 342962 216988 342990 217246
rect 343836 217138 343864 219370
rect 344664 217274 344692 221682
rect 345308 219298 345336 222838
rect 345296 219292 345348 219298
rect 345296 219234 345348 219240
rect 345480 218068 345532 218074
rect 345480 218010 345532 218016
rect 343790 217110 343864 217138
rect 344618 217246 344692 217274
rect 343790 216988 343818 217110
rect 344618 216988 344646 217246
rect 345492 217138 345520 218010
rect 346320 217274 346348 224606
rect 346596 223038 346624 231676
rect 346872 231662 347254 231690
rect 346872 228410 346900 231662
rect 346860 228404 346912 228410
rect 346860 228346 346912 228352
rect 347044 228404 347096 228410
rect 347044 228346 347096 228352
rect 346584 223032 346636 223038
rect 346584 222974 346636 222980
rect 347056 219434 347084 228346
rect 347884 222902 347912 231676
rect 348528 223174 348556 231676
rect 349172 228682 349200 231676
rect 349160 228676 349212 228682
rect 349160 228618 349212 228624
rect 349816 224534 349844 231676
rect 350460 229906 350488 231676
rect 350448 229900 350500 229906
rect 350448 229842 350500 229848
rect 350172 228676 350224 228682
rect 350172 228618 350224 228624
rect 349804 224528 349856 224534
rect 349804 224470 349856 224476
rect 348516 223168 348568 223174
rect 348516 223110 348568 223116
rect 349068 223032 349120 223038
rect 349068 222974 349120 222980
rect 347872 222896 347924 222902
rect 347872 222838 347924 222844
rect 347228 222760 347280 222766
rect 347228 222702 347280 222708
rect 347044 219428 347096 219434
rect 347044 219370 347096 219376
rect 347044 218884 347096 218890
rect 347044 218826 347096 218832
rect 345446 217110 345520 217138
rect 346274 217246 346348 217274
rect 345446 216988 345474 217110
rect 346274 216988 346302 217246
rect 347056 217138 347084 218826
rect 347240 218074 347268 222702
rect 348792 221604 348844 221610
rect 348792 221546 348844 221552
rect 347228 218068 347280 218074
rect 347228 218010 347280 218016
rect 347964 218068 348016 218074
rect 347964 218010 348016 218016
rect 347976 217138 348004 218010
rect 348804 217274 348832 221546
rect 349080 218074 349108 222974
rect 350184 218074 350212 228618
rect 351104 228546 351132 231676
rect 351288 231662 351762 231690
rect 351092 228540 351144 228546
rect 351092 228482 351144 228488
rect 351092 227792 351144 227798
rect 351092 227734 351144 227740
rect 350356 224868 350408 224874
rect 350356 224810 350408 224816
rect 349068 218068 349120 218074
rect 349068 218010 349120 218016
rect 349620 218068 349672 218074
rect 349620 218010 349672 218016
rect 350172 218068 350224 218074
rect 350172 218010 350224 218016
rect 347056 217110 347130 217138
rect 347102 216988 347130 217110
rect 347930 217110 348004 217138
rect 348758 217246 348832 217274
rect 347930 216988 347958 217110
rect 348758 216988 348786 217246
rect 349632 217138 349660 218010
rect 350368 217274 350396 224810
rect 351104 218754 351132 227734
rect 351288 220522 351316 231662
rect 352392 225622 352420 231676
rect 353036 227798 353064 231676
rect 353024 227792 353076 227798
rect 353024 227734 353076 227740
rect 352564 227452 352616 227458
rect 352564 227394 352616 227400
rect 352380 225616 352432 225622
rect 352380 225558 352432 225564
rect 351276 220516 351328 220522
rect 351276 220458 351328 220464
rect 351276 220380 351328 220386
rect 351276 220322 351328 220328
rect 351092 218748 351144 218754
rect 351092 218690 351144 218696
rect 351288 217274 351316 220322
rect 352576 219162 352604 227394
rect 353680 225758 353708 231676
rect 353956 231662 354338 231690
rect 354784 231662 354982 231690
rect 353668 225752 353720 225758
rect 353668 225694 353720 225700
rect 352932 225616 352984 225622
rect 352932 225558 352984 225564
rect 352564 219156 352616 219162
rect 352564 219098 352616 219104
rect 352104 218068 352156 218074
rect 352104 218010 352156 218016
rect 350368 217246 350442 217274
rect 349586 217110 349660 217138
rect 349586 216988 349614 217110
rect 350414 216988 350442 217246
rect 351242 217246 351316 217274
rect 351242 216988 351270 217246
rect 352116 217138 352144 218010
rect 352944 217274 352972 225558
rect 353956 222154 353984 231662
rect 354588 228540 354640 228546
rect 354588 228482 354640 228488
rect 353944 222148 353996 222154
rect 353944 222090 353996 222096
rect 353300 221876 353352 221882
rect 353300 221818 353352 221824
rect 353312 218074 353340 221818
rect 353760 218748 353812 218754
rect 353760 218690 353812 218696
rect 353300 218068 353352 218074
rect 353300 218010 353352 218016
rect 352070 217110 352144 217138
rect 352898 217246 352972 217274
rect 352070 216988 352098 217110
rect 352898 216988 352926 217246
rect 353772 217138 353800 218690
rect 354600 217274 354628 228482
rect 354784 220114 354812 231662
rect 355612 230178 355640 231676
rect 355600 230172 355652 230178
rect 355600 230114 355652 230120
rect 354956 230036 355008 230042
rect 354956 229978 355008 229984
rect 354968 224874 354996 229978
rect 356256 227322 356284 231676
rect 356244 227316 356296 227322
rect 356244 227258 356296 227264
rect 356900 226030 356928 231676
rect 357256 227316 357308 227322
rect 357256 227258 357308 227264
rect 356888 226024 356940 226030
rect 356888 225966 356940 225972
rect 355232 225004 355284 225010
rect 355232 224946 355284 224952
rect 354956 224868 355008 224874
rect 354956 224810 355008 224816
rect 354772 220108 354824 220114
rect 354772 220050 354824 220056
rect 355244 219026 355272 224946
rect 355416 220108 355468 220114
rect 355416 220050 355468 220056
rect 355232 219020 355284 219026
rect 355232 218962 355284 218968
rect 355428 217274 355456 220050
rect 357072 219020 357124 219026
rect 357072 218962 357124 218968
rect 356244 218068 356296 218074
rect 356244 218010 356296 218016
rect 353726 217110 353800 217138
rect 354554 217246 354628 217274
rect 355382 217246 355456 217274
rect 353726 216988 353754 217110
rect 354554 216988 354582 217246
rect 355382 216988 355410 217246
rect 356256 217138 356284 218010
rect 357084 217138 357112 218962
rect 357268 218074 357296 227258
rect 357544 221474 357572 231676
rect 358188 225010 358216 231676
rect 358832 228818 358860 231676
rect 359200 231662 359490 231690
rect 358820 228812 358872 228818
rect 358820 228754 358872 228760
rect 358176 225004 358228 225010
rect 358176 224946 358228 224952
rect 359200 223310 359228 231662
rect 359924 228812 359976 228818
rect 359924 228754 359976 228760
rect 359464 224528 359516 224534
rect 359464 224470 359516 224476
rect 359188 223304 359240 223310
rect 359188 223246 359240 223252
rect 358544 223168 358596 223174
rect 358544 223110 358596 223116
rect 357532 221468 357584 221474
rect 357532 221410 357584 221416
rect 358556 218074 358584 223110
rect 359476 218210 359504 224470
rect 359936 219434 359964 228754
rect 360120 227050 360148 231676
rect 360764 229770 360792 231676
rect 360752 229764 360804 229770
rect 360752 229706 360804 229712
rect 361212 229764 361264 229770
rect 361212 229706 361264 229712
rect 361224 229094 361252 229706
rect 361040 229066 361252 229094
rect 360108 227044 360160 227050
rect 360108 226986 360160 226992
rect 359936 219406 360148 219434
rect 358728 218204 358780 218210
rect 358728 218146 358780 218152
rect 359464 218204 359516 218210
rect 359464 218146 359516 218152
rect 357256 218068 357308 218074
rect 357256 218010 357308 218016
rect 357900 218068 357952 218074
rect 357900 218010 357952 218016
rect 358544 218068 358596 218074
rect 358544 218010 358596 218016
rect 357912 217138 357940 218010
rect 358740 217138 358768 218146
rect 360120 218074 360148 219406
rect 361040 218074 361068 229066
rect 361408 227186 361436 231676
rect 361396 227180 361448 227186
rect 361396 227122 361448 227128
rect 361212 226024 361264 226030
rect 361212 225966 361264 225972
rect 359556 218068 359608 218074
rect 359556 218010 359608 218016
rect 360108 218068 360160 218074
rect 360108 218010 360160 218016
rect 360384 218068 360436 218074
rect 360384 218010 360436 218016
rect 361028 218068 361080 218074
rect 361028 218010 361080 218016
rect 359568 217138 359596 218010
rect 360396 217138 360424 218010
rect 361224 217274 361252 225966
rect 362052 224398 362080 231676
rect 362328 231662 362710 231690
rect 362040 224392 362092 224398
rect 362040 224334 362092 224340
rect 362328 224262 362356 231662
rect 363340 227458 363368 231676
rect 363524 231662 363998 231690
rect 364536 231662 364642 231690
rect 363328 227452 363380 227458
rect 363328 227394 363380 227400
rect 363524 227338 363552 231662
rect 363340 227310 363552 227338
rect 362776 227044 362828 227050
rect 362776 226986 362828 226992
rect 362316 224256 362368 224262
rect 362316 224198 362368 224204
rect 362040 219156 362092 219162
rect 362040 219098 362092 219104
rect 362052 217274 362080 219098
rect 356210 217110 356284 217138
rect 357038 217110 357112 217138
rect 357866 217110 357940 217138
rect 358694 217110 358768 217138
rect 359522 217110 359596 217138
rect 360350 217110 360424 217138
rect 361178 217246 361252 217274
rect 362006 217246 362080 217274
rect 362788 217274 362816 226986
rect 363340 220250 363368 227310
rect 363512 227180 363564 227186
rect 363512 227122 363564 227128
rect 363328 220244 363380 220250
rect 363328 220186 363380 220192
rect 363524 218890 363552 227122
rect 364536 221746 364564 231662
rect 365272 225894 365300 231676
rect 365916 228410 365944 231676
rect 365904 228404 365956 228410
rect 365904 228346 365956 228352
rect 365260 225888 365312 225894
rect 365260 225830 365312 225836
rect 365352 225752 365404 225758
rect 365352 225694 365404 225700
rect 364524 221740 364576 221746
rect 364524 221682 364576 221688
rect 364524 220516 364576 220522
rect 364524 220458 364576 220464
rect 363696 220244 363748 220250
rect 363696 220186 363748 220192
rect 363512 218884 363564 218890
rect 363512 218826 363564 218832
rect 363708 217274 363736 220186
rect 364536 217274 364564 220458
rect 365364 217274 365392 225694
rect 366560 224670 366588 231676
rect 366732 229900 366784 229906
rect 366732 229842 366784 229848
rect 366744 229094 366772 229842
rect 366744 229066 366956 229094
rect 366548 224664 366600 224670
rect 366548 224606 366600 224612
rect 366732 224392 366784 224398
rect 366732 224334 366784 224340
rect 366744 219570 366772 224334
rect 366732 219564 366784 219570
rect 366732 219506 366784 219512
rect 366180 219428 366232 219434
rect 366180 219370 366232 219376
rect 362788 217246 362862 217274
rect 356210 216988 356238 217110
rect 357038 216988 357066 217110
rect 357866 216988 357894 217110
rect 358694 216988 358722 217110
rect 359522 216988 359550 217110
rect 360350 216988 360378 217110
rect 361178 216988 361206 217246
rect 362006 216988 362034 217246
rect 362834 216988 362862 217246
rect 363662 217246 363736 217274
rect 364490 217246 364564 217274
rect 365318 217246 365392 217274
rect 363662 216988 363690 217246
rect 364490 216988 364518 217246
rect 365318 216988 365346 217246
rect 366192 217138 366220 219370
rect 366928 217274 366956 229066
rect 367204 223038 367232 231676
rect 367192 223032 367244 223038
rect 367192 222974 367244 222980
rect 367848 222902 367876 231676
rect 368492 227186 368520 231676
rect 369136 228682 369164 231676
rect 369320 231662 369794 231690
rect 370056 231662 370438 231690
rect 369124 228676 369176 228682
rect 369124 228618 369176 228624
rect 368480 227180 368532 227186
rect 368480 227122 368532 227128
rect 369124 226500 369176 226506
rect 369124 226442 369176 226448
rect 368388 223032 368440 223038
rect 368388 222974 368440 222980
rect 367836 222896 367888 222902
rect 367836 222838 367888 222844
rect 368400 218074 368428 222974
rect 369136 219026 369164 226442
rect 369320 220386 369348 231662
rect 370056 221610 370084 231662
rect 371068 230042 371096 231676
rect 371056 230036 371108 230042
rect 371056 229978 371108 229984
rect 371712 229094 371740 231676
rect 371620 229066 371740 229094
rect 371148 228404 371200 228410
rect 371148 228346 371200 228352
rect 370964 221740 371016 221746
rect 370964 221682 371016 221688
rect 370044 221604 370096 221610
rect 370044 221546 370096 221552
rect 369492 221468 369544 221474
rect 369492 221410 369544 221416
rect 369308 220380 369360 220386
rect 369308 220322 369360 220328
rect 369124 219020 369176 219026
rect 369124 218962 369176 218968
rect 368664 218884 368716 218890
rect 368664 218826 368716 218832
rect 367836 218068 367888 218074
rect 367836 218010 367888 218016
rect 368388 218068 368440 218074
rect 368388 218010 368440 218016
rect 366928 217246 367002 217274
rect 366146 217110 366220 217138
rect 366146 216988 366174 217110
rect 366974 216988 367002 217246
rect 367848 217138 367876 218010
rect 368676 217138 368704 218826
rect 369504 217274 369532 221410
rect 370976 219162 371004 221682
rect 370964 219156 371016 219162
rect 370964 219098 371016 219104
rect 370320 219020 370372 219026
rect 370320 218962 370372 218968
rect 367802 217110 367876 217138
rect 368630 217110 368704 217138
rect 369458 217246 369532 217274
rect 367802 216988 367830 217110
rect 368630 216988 368658 217110
rect 369458 216988 369486 217246
rect 370332 217138 370360 218962
rect 371160 217274 371188 228346
rect 371620 225622 371648 229066
rect 372356 228546 372384 231676
rect 372724 231662 373014 231690
rect 372344 228540 372396 228546
rect 372344 228482 372396 228488
rect 371792 227792 371844 227798
rect 371792 227734 371844 227740
rect 371608 225616 371660 225622
rect 371608 225558 371660 225564
rect 371804 218754 371832 227734
rect 372528 224256 372580 224262
rect 372528 224198 372580 224204
rect 371792 218748 371844 218754
rect 371792 218690 371844 218696
rect 372540 218074 372568 224198
rect 372724 221882 372752 231662
rect 373448 228540 373500 228546
rect 373448 228482 373500 228488
rect 372712 221876 372764 221882
rect 372712 221818 372764 221824
rect 373460 219434 373488 228482
rect 373644 227798 373672 231676
rect 373632 227792 373684 227798
rect 373632 227734 373684 227740
rect 374288 227322 374316 231676
rect 374656 231662 374946 231690
rect 374276 227316 374328 227322
rect 374276 227258 374328 227264
rect 374656 223174 374684 231662
rect 375012 225888 375064 225894
rect 375012 225830 375064 225836
rect 374644 223168 374696 223174
rect 374644 223110 374696 223116
rect 373724 221604 373776 221610
rect 373724 221546 373776 221552
rect 373460 219406 373580 219434
rect 373552 218074 373580 219406
rect 371976 218068 372028 218074
rect 371976 218010 372028 218016
rect 372528 218068 372580 218074
rect 372528 218010 372580 218016
rect 372804 218068 372856 218074
rect 372804 218010 372856 218016
rect 373540 218068 373592 218074
rect 373540 218010 373592 218016
rect 370286 217110 370360 217138
rect 371114 217246 371188 217274
rect 370286 216988 370314 217110
rect 371114 216988 371142 217246
rect 371988 217138 372016 218010
rect 372816 217138 372844 218010
rect 373736 217274 373764 221546
rect 375024 218074 375052 225830
rect 375196 222896 375248 222902
rect 375196 222838 375248 222844
rect 374460 218068 374512 218074
rect 374460 218010 374512 218016
rect 375012 218068 375064 218074
rect 375012 218010 375064 218016
rect 371942 217110 372016 217138
rect 372770 217110 372844 217138
rect 373598 217246 373764 217274
rect 371942 216988 371970 217110
rect 372770 216988 372798 217110
rect 373598 216988 373626 217246
rect 374472 217138 374500 218010
rect 375208 217274 375236 222838
rect 375576 220114 375604 231676
rect 376220 226506 376248 231676
rect 376864 228818 376892 231676
rect 376852 228812 376904 228818
rect 376852 228754 376904 228760
rect 376668 227180 376720 227186
rect 376668 227122 376720 227128
rect 376208 226500 376260 226506
rect 376208 226442 376260 226448
rect 375564 220108 375616 220114
rect 375564 220050 375616 220056
rect 376680 218074 376708 227122
rect 377508 226030 377536 231676
rect 377772 228676 377824 228682
rect 377772 228618 377824 228624
rect 377496 226024 377548 226030
rect 377496 225966 377548 225972
rect 376944 220380 376996 220386
rect 376944 220322 376996 220328
rect 376116 218068 376168 218074
rect 376116 218010 376168 218016
rect 376668 218068 376720 218074
rect 376668 218010 376720 218016
rect 375208 217246 375282 217274
rect 374426 217110 374500 217138
rect 374426 216988 374454 217110
rect 375254 216988 375282 217246
rect 376128 217138 376156 218010
rect 376956 217274 376984 220322
rect 377784 217274 377812 228618
rect 378152 224534 378180 231676
rect 378796 229770 378824 231676
rect 379072 231662 379454 231690
rect 379716 231662 380098 231690
rect 380360 231662 380742 231690
rect 381096 231662 381386 231690
rect 381648 231662 382030 231690
rect 378784 229764 378836 229770
rect 378784 229706 378836 229712
rect 379072 227050 379100 231662
rect 379060 227044 379112 227050
rect 379060 226986 379112 226992
rect 378784 226840 378836 226846
rect 378784 226782 378836 226788
rect 378140 224528 378192 224534
rect 378140 224470 378192 224476
rect 378796 218890 378824 226782
rect 379244 224528 379296 224534
rect 379244 224470 379296 224476
rect 378784 218884 378836 218890
rect 378784 218826 378836 218832
rect 379256 218074 379284 224470
rect 379716 220522 379744 231662
rect 380360 221882 380388 231662
rect 380348 221876 380400 221882
rect 380348 221818 380400 221824
rect 380072 221740 380124 221746
rect 380072 221682 380124 221688
rect 379704 220516 379756 220522
rect 379704 220458 379756 220464
rect 379428 220108 379480 220114
rect 379428 220050 379480 220056
rect 378600 218068 378652 218074
rect 378600 218010 378652 218016
rect 379244 218068 379296 218074
rect 379244 218010 379296 218016
rect 376082 217110 376156 217138
rect 376910 217246 376984 217274
rect 377738 217246 377812 217274
rect 376082 216988 376110 217110
rect 376910 216988 376938 217246
rect 377738 216988 377766 217246
rect 378612 217138 378640 218010
rect 379440 217274 379468 220050
rect 380084 219026 380112 221682
rect 381096 220250 381124 231662
rect 381648 224398 381676 231662
rect 382096 227316 382148 227322
rect 382096 227258 382148 227264
rect 381636 224392 381688 224398
rect 381636 224334 381688 224340
rect 381084 220244 381136 220250
rect 381084 220186 381136 220192
rect 380072 219020 380124 219026
rect 380072 218962 380124 218968
rect 380256 219020 380308 219026
rect 380256 218962 380308 218968
rect 378566 217110 378640 217138
rect 379394 217246 379468 217274
rect 378566 216988 378594 217110
rect 379394 216988 379422 217246
rect 380268 217138 380296 218962
rect 381912 218204 381964 218210
rect 381912 218146 381964 218152
rect 381084 218068 381136 218074
rect 381084 218010 381136 218016
rect 381096 217138 381124 218010
rect 381924 217138 381952 218146
rect 382108 218074 382136 227258
rect 382660 223038 382688 231676
rect 383304 225758 383332 231676
rect 383948 229906 383976 231676
rect 384132 231662 384606 231690
rect 383936 229900 383988 229906
rect 383936 229842 383988 229848
rect 383292 225752 383344 225758
rect 383292 225694 383344 225700
rect 382924 225616 382976 225622
rect 382924 225558 382976 225564
rect 382648 223032 382700 223038
rect 382648 222974 382700 222980
rect 382740 218884 382792 218890
rect 382740 218826 382792 218832
rect 382096 218068 382148 218074
rect 382096 218010 382148 218016
rect 382752 217138 382780 218826
rect 382936 218210 382964 225558
rect 383568 223032 383620 223038
rect 383568 222974 383620 222980
rect 383580 218890 383608 222974
rect 384132 221474 384160 231662
rect 384304 229560 384356 229566
rect 384304 229502 384356 229508
rect 384316 221610 384344 229502
rect 385236 228410 385264 231676
rect 385224 228404 385276 228410
rect 385224 228346 385276 228352
rect 385880 226846 385908 231676
rect 386236 228404 386288 228410
rect 386236 228346 386288 228352
rect 385868 226840 385920 226846
rect 385868 226782 385920 226788
rect 386052 226432 386104 226438
rect 386052 226374 386104 226380
rect 384304 221604 384356 221610
rect 384304 221546 384356 221552
rect 384120 221468 384172 221474
rect 384120 221410 384172 221416
rect 384396 221468 384448 221474
rect 384396 221410 384448 221416
rect 383568 218884 383620 218890
rect 383568 218826 383620 218832
rect 383568 218748 383620 218754
rect 383568 218690 383620 218696
rect 382924 218204 382976 218210
rect 382924 218146 382976 218152
rect 383580 217138 383608 218690
rect 384408 217274 384436 221410
rect 386064 218074 386092 226374
rect 385224 218068 385276 218074
rect 385224 218010 385276 218016
rect 386052 218068 386104 218074
rect 386052 218010 386104 218016
rect 380222 217110 380296 217138
rect 381050 217110 381124 217138
rect 381878 217110 381952 217138
rect 382706 217110 382780 217138
rect 383534 217110 383608 217138
rect 384362 217246 384436 217274
rect 380222 216988 380250 217110
rect 381050 216988 381078 217110
rect 381878 216988 381906 217110
rect 382706 216988 382734 217110
rect 383534 216988 383562 217110
rect 384362 216988 384390 217246
rect 385236 217138 385264 218010
rect 386248 217274 386276 228346
rect 386524 221746 386552 231676
rect 387168 228546 387196 231676
rect 387432 230376 387484 230382
rect 387432 230318 387484 230324
rect 387156 228540 387208 228546
rect 387156 228482 387208 228488
rect 387444 224262 387472 230318
rect 387812 225894 387840 231676
rect 388456 230382 388484 231676
rect 388444 230376 388496 230382
rect 388444 230318 388496 230324
rect 388444 230240 388496 230246
rect 388444 230182 388496 230188
rect 387800 225888 387852 225894
rect 387800 225830 387852 225836
rect 387708 225752 387760 225758
rect 387708 225694 387760 225700
rect 387432 224256 387484 224262
rect 387432 224198 387484 224204
rect 386512 221740 386564 221746
rect 386512 221682 386564 221688
rect 386880 218884 386932 218890
rect 386880 218826 386932 218832
rect 385190 217110 385264 217138
rect 386018 217246 386276 217274
rect 385190 216988 385218 217110
rect 386018 216988 386046 217246
rect 386892 217138 386920 218826
rect 387720 217274 387748 225694
rect 388456 220386 388484 230182
rect 389100 229566 389128 231676
rect 389088 229560 389140 229566
rect 389088 229502 389140 229508
rect 389744 227186 389772 231676
rect 390388 228682 390416 231676
rect 390376 228676 390428 228682
rect 390376 228618 390428 228624
rect 390468 228540 390520 228546
rect 390468 228482 390520 228488
rect 389732 227180 389784 227186
rect 389732 227122 389784 227128
rect 388628 226296 388680 226302
rect 388628 226238 388680 226244
rect 388444 220380 388496 220386
rect 388444 220322 388496 220328
rect 388444 220244 388496 220250
rect 388444 220186 388496 220192
rect 386846 217110 386920 217138
rect 387674 217246 387748 217274
rect 388456 217274 388484 220186
rect 388640 219026 388668 226238
rect 390192 224256 390244 224262
rect 390192 224198 390244 224204
rect 388628 219020 388680 219026
rect 388628 218962 388680 218968
rect 389364 218068 389416 218074
rect 389364 218010 389416 218016
rect 388456 217246 388530 217274
rect 386846 216988 386874 217110
rect 387674 216988 387702 217246
rect 388502 216988 388530 217246
rect 389376 217138 389404 218010
rect 390204 217274 390232 224198
rect 390480 218074 390508 228482
rect 391032 222902 391060 231676
rect 391676 230246 391704 231676
rect 392136 231662 392334 231690
rect 391664 230240 391716 230246
rect 391664 230182 391716 230188
rect 391204 229764 391256 229770
rect 391204 229706 391256 229712
rect 391216 226438 391244 229706
rect 391756 227044 391808 227050
rect 391756 226986 391808 226992
rect 391204 226432 391256 226438
rect 391204 226374 391256 226380
rect 391020 222896 391072 222902
rect 391020 222838 391072 222844
rect 391020 221604 391072 221610
rect 391020 221546 391072 221552
rect 390468 218068 390520 218074
rect 390468 218010 390520 218016
rect 391032 217274 391060 221546
rect 389330 217110 389404 217138
rect 390158 217246 390232 217274
rect 390986 217246 391060 217274
rect 391768 217274 391796 226986
rect 392136 220114 392164 231662
rect 392964 227322 392992 231676
rect 392952 227316 393004 227322
rect 392952 227258 393004 227264
rect 393136 227180 393188 227186
rect 393136 227122 393188 227128
rect 392124 220108 392176 220114
rect 392124 220050 392176 220056
rect 393148 218074 393176 227122
rect 393608 224534 393636 231676
rect 394252 226302 394280 231676
rect 394240 226296 394292 226302
rect 394240 226238 394292 226244
rect 394332 225888 394384 225894
rect 394332 225830 394384 225836
rect 393596 224528 393648 224534
rect 393596 224470 393648 224476
rect 392676 218068 392728 218074
rect 392676 218010 392728 218016
rect 393136 218068 393188 218074
rect 393136 218010 393188 218016
rect 393504 218068 393556 218074
rect 393504 218010 393556 218016
rect 391768 217246 391842 217274
rect 389330 216988 389358 217110
rect 390158 216988 390186 217246
rect 390986 216988 391014 217246
rect 391814 216988 391842 217246
rect 392688 217138 392716 218010
rect 393516 217138 393544 218010
rect 394344 217274 394372 225830
rect 394516 224392 394568 224398
rect 394516 224334 394568 224340
rect 394528 218074 394556 224334
rect 394896 223038 394924 231676
rect 395172 231662 395554 231690
rect 394884 223032 394936 223038
rect 394884 222974 394936 222980
rect 395172 221474 395200 231662
rect 396184 225622 396212 231676
rect 396368 231662 396842 231690
rect 396172 225616 396224 225622
rect 396172 225558 396224 225564
rect 395804 222896 395856 222902
rect 395804 222838 395856 222844
rect 395160 221468 395212 221474
rect 395160 221410 395212 221416
rect 395816 218074 395844 222838
rect 395988 220108 396040 220114
rect 395988 220050 396040 220056
rect 394516 218068 394568 218074
rect 394516 218010 394568 218016
rect 395160 218068 395212 218074
rect 395160 218010 395212 218016
rect 395804 218068 395856 218074
rect 395804 218010 395856 218016
rect 392642 217110 392716 217138
rect 393470 217110 393544 217138
rect 394298 217246 394372 217274
rect 392642 216988 392670 217110
rect 393470 216988 393498 217110
rect 394298 216988 394326 217246
rect 395172 217138 395200 218010
rect 396000 217274 396028 220050
rect 396368 219434 396396 231662
rect 397472 228410 397500 231676
rect 397840 231662 398130 231690
rect 397460 228404 397512 228410
rect 397460 228346 397512 228352
rect 397840 225758 397868 231662
rect 398104 230376 398156 230382
rect 398104 230318 398156 230324
rect 397828 225752 397880 225758
rect 397828 225694 397880 225700
rect 396816 221468 396868 221474
rect 396816 221410 396868 221416
rect 396276 219406 396396 219434
rect 396276 218754 396304 219406
rect 396264 218748 396316 218754
rect 396264 218690 396316 218696
rect 396828 217274 396856 221410
rect 398116 218890 398144 230318
rect 398760 229770 398788 231676
rect 399404 230382 399432 231676
rect 399392 230376 399444 230382
rect 399392 230318 399444 230324
rect 398748 229764 398800 229770
rect 398748 229706 398800 229712
rect 399852 229764 399904 229770
rect 399852 229706 399904 229712
rect 399864 219434 399892 229706
rect 400048 228546 400076 231676
rect 400232 231662 400706 231690
rect 400968 231662 401350 231690
rect 400232 229094 400260 231662
rect 400232 229066 400352 229094
rect 400036 228540 400088 228546
rect 400036 228482 400088 228488
rect 400128 228132 400180 228138
rect 400128 228074 400180 228080
rect 400140 219434 400168 228074
rect 400324 221610 400352 229066
rect 400312 221604 400364 221610
rect 400312 221546 400364 221552
rect 400968 220250 400996 231662
rect 401980 224262 402008 231676
rect 402624 227322 402652 231676
rect 402796 228404 402848 228410
rect 402796 228346 402848 228352
rect 402612 227316 402664 227322
rect 402612 227258 402664 227264
rect 402244 227180 402296 227186
rect 402244 227122 402296 227128
rect 401968 224256 402020 224262
rect 401968 224198 402020 224204
rect 401232 221604 401284 221610
rect 401232 221546 401284 221552
rect 400956 220244 401008 220250
rect 400956 220186 401008 220192
rect 399300 219428 399352 219434
rect 399864 219406 400076 219434
rect 400140 219428 400272 219434
rect 400140 219406 400220 219428
rect 399300 219370 399352 219376
rect 398104 218884 398156 218890
rect 398104 218826 398156 218832
rect 398472 218612 398524 218618
rect 398472 218554 398524 218560
rect 397644 218068 397696 218074
rect 397644 218010 397696 218016
rect 395126 217110 395200 217138
rect 395954 217246 396028 217274
rect 396782 217246 396856 217274
rect 395126 216988 395154 217110
rect 395954 216988 395982 217246
rect 396782 216988 396810 217246
rect 397656 217138 397684 218010
rect 398484 217138 398512 218554
rect 399312 217138 399340 219370
rect 400048 217274 400076 219406
rect 400220 219370 400272 219376
rect 400956 218204 401008 218210
rect 400956 218146 401008 218152
rect 400048 217246 400122 217274
rect 397610 217110 397684 217138
rect 398438 217110 398512 217138
rect 399266 217110 399340 217138
rect 397610 216988 397638 217110
rect 398438 216988 398466 217110
rect 399266 216988 399294 217110
rect 400094 216988 400122 217246
rect 400968 217138 400996 218146
rect 401244 218074 401272 221546
rect 402256 218210 402284 227122
rect 402612 218884 402664 218890
rect 402612 218826 402664 218832
rect 402244 218204 402296 218210
rect 402244 218146 402296 218152
rect 401232 218068 401284 218074
rect 401232 218010 401284 218016
rect 401784 218068 401836 218074
rect 401784 218010 401836 218016
rect 401796 217138 401824 218010
rect 402624 217138 402652 218826
rect 402808 218074 402836 228346
rect 403268 225894 403296 231676
rect 403544 231662 403926 231690
rect 403544 227050 403572 231662
rect 403532 227044 403584 227050
rect 403532 226986 403584 226992
rect 403992 226500 404044 226506
rect 403992 226442 404044 226448
rect 403256 225888 403308 225894
rect 403256 225830 403308 225836
rect 404004 218074 404032 226442
rect 404176 225004 404228 225010
rect 404176 224946 404228 224952
rect 402796 218068 402848 218074
rect 402796 218010 402848 218016
rect 403440 218068 403492 218074
rect 403440 218010 403492 218016
rect 403992 218068 404044 218074
rect 403992 218010 404044 218016
rect 403452 217138 403480 218010
rect 404188 217274 404216 224946
rect 404556 224398 404584 231676
rect 404740 231662 405214 231690
rect 404544 224392 404596 224398
rect 404544 224334 404596 224340
rect 404740 220114 404768 231662
rect 405556 224256 405608 224262
rect 405556 224198 405608 224204
rect 404728 220108 404780 220114
rect 404728 220050 404780 220056
rect 405568 218074 405596 224198
rect 405844 221610 405872 231676
rect 406488 222902 406516 231676
rect 407146 231662 407344 231690
rect 406752 223576 406804 223582
rect 406752 223518 406804 223524
rect 406476 222896 406528 222902
rect 406476 222838 406528 222844
rect 405832 221604 405884 221610
rect 405832 221546 405884 221552
rect 405924 219496 405976 219502
rect 405924 219438 405976 219444
rect 405096 218068 405148 218074
rect 405096 218010 405148 218016
rect 405556 218068 405608 218074
rect 405556 218010 405608 218016
rect 404188 217246 404262 217274
rect 400922 217110 400996 217138
rect 401750 217110 401824 217138
rect 402578 217110 402652 217138
rect 403406 217110 403480 217138
rect 400922 216988 400950 217110
rect 401750 216988 401778 217110
rect 402578 216988 402606 217110
rect 403406 216988 403434 217110
rect 404234 216988 404262 217246
rect 405108 217138 405136 218010
rect 405936 217274 405964 219438
rect 406764 217274 406792 223518
rect 407316 221474 407344 231662
rect 407776 228546 407804 231676
rect 407764 228540 407816 228546
rect 407764 228482 407816 228488
rect 408420 227186 408448 231676
rect 408696 231662 409078 231690
rect 408408 227180 408460 227186
rect 408408 227122 408460 227128
rect 408696 226370 408724 231662
rect 409708 229770 409736 231676
rect 409696 229764 409748 229770
rect 409696 229706 409748 229712
rect 409788 228540 409840 228546
rect 409788 228482 409840 228488
rect 409052 227792 409104 227798
rect 409052 227734 409104 227740
rect 407764 226364 407816 226370
rect 407764 226306 407816 226312
rect 408684 226364 408736 226370
rect 408684 226306 408736 226312
rect 407304 221468 407356 221474
rect 407304 221410 407356 221416
rect 407776 218618 407804 226306
rect 408408 221468 408460 221474
rect 408408 221410 408460 221416
rect 407764 218612 407816 218618
rect 407764 218554 407816 218560
rect 407580 218204 407632 218210
rect 407580 218146 407632 218152
rect 405062 217110 405136 217138
rect 405890 217246 405964 217274
rect 406718 217246 406792 217274
rect 405062 216988 405090 217110
rect 405890 216988 405918 217246
rect 406718 216988 406746 217246
rect 407592 217138 407620 218146
rect 408420 217274 408448 221410
rect 409064 218890 409092 227734
rect 409052 218884 409104 218890
rect 409052 218826 409104 218832
rect 409800 218074 409828 228482
rect 410352 227798 410380 231676
rect 410720 231662 411010 231690
rect 410720 229094 410748 231662
rect 410892 229764 410944 229770
rect 410892 229706 410944 229712
rect 410904 229094 410932 229706
rect 410628 229066 410748 229094
rect 410812 229066 410932 229094
rect 410340 227792 410392 227798
rect 410340 227734 410392 227740
rect 410628 225010 410656 229066
rect 410616 225004 410668 225010
rect 410616 224946 410668 224952
rect 410812 219434 410840 229066
rect 411640 228410 411668 231676
rect 411628 228404 411680 228410
rect 411628 228346 411680 228352
rect 411904 227792 411956 227798
rect 411904 227734 411956 227740
rect 410984 225616 411036 225622
rect 410984 225558 411036 225564
rect 410996 219434 411024 225558
rect 410720 219406 410840 219434
rect 410904 219406 411024 219434
rect 410720 218074 410748 219406
rect 409236 218068 409288 218074
rect 409236 218010 409288 218016
rect 409788 218068 409840 218074
rect 409788 218010 409840 218016
rect 410064 218068 410116 218074
rect 410064 218010 410116 218016
rect 410708 218068 410760 218074
rect 410708 218010 410760 218016
rect 407546 217110 407620 217138
rect 408374 217246 408448 217274
rect 407546 216988 407574 217110
rect 408374 216988 408402 217246
rect 409248 217138 409276 218010
rect 410076 217138 410104 218010
rect 410904 217274 410932 219406
rect 411720 218884 411772 218890
rect 411720 218826 411772 218832
rect 409202 217110 409276 217138
rect 410030 217110 410104 217138
rect 410858 217246 410932 217274
rect 409202 216988 409230 217110
rect 410030 216988 410058 217110
rect 410858 216988 410886 217246
rect 411732 217138 411760 218826
rect 411916 218210 411944 227734
rect 412284 226506 412312 231676
rect 412744 231662 412942 231690
rect 412548 227044 412600 227050
rect 412548 226986 412600 226992
rect 412272 226500 412324 226506
rect 412272 226442 412324 226448
rect 412560 218890 412588 226986
rect 412744 219502 412772 231662
rect 413572 227798 413600 231676
rect 413836 229356 413888 229362
rect 413836 229298 413888 229304
rect 413560 227792 413612 227798
rect 413560 227734 413612 227740
rect 412732 219496 412784 219502
rect 412732 219438 412784 219444
rect 412548 218884 412600 218890
rect 412548 218826 412600 218832
rect 412548 218748 412600 218754
rect 412548 218690 412600 218696
rect 411904 218204 411956 218210
rect 411904 218146 411956 218152
rect 412560 217138 412588 218690
rect 413848 218074 413876 229298
rect 414216 224262 414244 231676
rect 414204 224256 414256 224262
rect 414204 224198 414256 224204
rect 414860 223582 414888 231676
rect 415504 228546 415532 231676
rect 415492 228540 415544 228546
rect 415492 228482 415544 228488
rect 415032 228064 415084 228070
rect 415032 228006 415084 228012
rect 414848 223576 414900 223582
rect 414848 223518 414900 223524
rect 414204 220788 414256 220794
rect 414204 220730 414256 220736
rect 413376 218068 413428 218074
rect 413376 218010 413428 218016
rect 413836 218068 413888 218074
rect 413836 218010 413888 218016
rect 413388 217138 413416 218010
rect 414216 217274 414244 220730
rect 415044 217274 415072 228006
rect 416148 225622 416176 231676
rect 416792 229094 416820 231676
rect 417436 229770 417464 231676
rect 417712 231662 418094 231690
rect 418356 231662 418738 231690
rect 417424 229764 417476 229770
rect 417424 229706 417476 229712
rect 417712 229094 417740 231662
rect 416792 229066 416912 229094
rect 416688 227928 416740 227934
rect 416688 227870 416740 227876
rect 416136 225616 416188 225622
rect 416136 225558 416188 225564
rect 416504 225004 416556 225010
rect 416504 224946 416556 224952
rect 416516 219434 416544 224946
rect 416700 219434 416728 227870
rect 416884 221474 416912 229066
rect 417160 229066 417740 229094
rect 416872 221468 416924 221474
rect 416872 221410 416924 221416
rect 415860 219428 415912 219434
rect 416516 219406 416636 219434
rect 416700 219428 416832 219434
rect 416700 219406 416780 219428
rect 415860 219370 415912 219376
rect 411686 217110 411760 217138
rect 412514 217110 412588 217138
rect 413342 217110 413416 217138
rect 414170 217246 414244 217274
rect 414998 217246 415072 217274
rect 411686 216988 411714 217110
rect 412514 216988 412542 217110
rect 413342 216988 413370 217110
rect 414170 216988 414198 217246
rect 414998 216988 415026 217246
rect 415872 217138 415900 219370
rect 416608 217274 416636 219406
rect 416780 219370 416832 219376
rect 417160 218754 417188 229066
rect 418356 224954 418384 231662
rect 419368 227050 419396 231676
rect 420012 229362 420040 231676
rect 420000 229356 420052 229362
rect 420000 229298 420052 229304
rect 420656 227934 420684 231676
rect 421024 231662 421314 231690
rect 420644 227928 420696 227934
rect 420644 227870 420696 227876
rect 420644 227792 420696 227798
rect 420644 227734 420696 227740
rect 419356 227044 419408 227050
rect 419356 226986 419408 226992
rect 418172 224926 418384 224954
rect 418172 220794 418200 224926
rect 418344 220856 418396 220862
rect 418344 220798 418396 220804
rect 418160 220788 418212 220794
rect 418160 220730 418212 220736
rect 417516 219428 417568 219434
rect 417516 219370 417568 219376
rect 417148 218748 417200 218754
rect 417148 218690 417200 218696
rect 416608 217246 416682 217274
rect 415826 217110 415900 217138
rect 415826 216988 415854 217110
rect 416654 216988 416682 217246
rect 417528 217138 417556 219370
rect 418356 217274 418384 220798
rect 420656 219434 420684 227734
rect 420828 222896 420880 222902
rect 420828 222838 420880 222844
rect 420656 219406 420776 219434
rect 419172 219292 419224 219298
rect 419172 219234 419224 219240
rect 419184 217274 419212 219234
rect 420000 218068 420052 218074
rect 420000 218010 420052 218016
rect 417482 217110 417556 217138
rect 418310 217246 418384 217274
rect 419138 217246 419212 217274
rect 417482 216988 417510 217110
rect 418310 216988 418338 217246
rect 419138 216988 419166 217246
rect 420012 217138 420040 218010
rect 420748 217274 420776 219406
rect 420840 218090 420868 222838
rect 421024 219502 421052 231662
rect 421944 228070 421972 231676
rect 422312 231662 422602 231690
rect 422864 231662 423246 231690
rect 422312 229094 422340 231662
rect 422220 229066 422340 229094
rect 421932 228064 421984 228070
rect 421932 228006 421984 228012
rect 422220 225010 422248 229066
rect 422208 225004 422260 225010
rect 422208 224946 422260 224952
rect 421656 220108 421708 220114
rect 421656 220050 421708 220056
rect 421012 219496 421064 219502
rect 421012 219438 421064 219444
rect 420840 218074 420960 218090
rect 420840 218068 420972 218074
rect 420840 218062 420920 218068
rect 420920 218010 420972 218016
rect 421668 217274 421696 220050
rect 422864 219434 422892 231662
rect 423496 229152 423548 229158
rect 423496 229094 423548 229100
rect 423508 219434 423536 229094
rect 423876 227798 423904 231676
rect 424060 231662 424534 231690
rect 423864 227792 423916 227798
rect 423864 227734 423916 227740
rect 424060 220862 424088 231662
rect 425164 222902 425192 231676
rect 425440 231662 425822 231690
rect 425152 222896 425204 222902
rect 425152 222838 425204 222844
rect 424968 222148 425020 222154
rect 424968 222090 425020 222096
rect 424048 220856 424100 220862
rect 424048 220798 424100 220804
rect 422680 219406 422892 219434
rect 423324 219406 423536 219434
rect 422680 219298 422708 219406
rect 422668 219292 422720 219298
rect 422668 219234 422720 219240
rect 422484 218204 422536 218210
rect 422484 218146 422536 218152
rect 420748 217246 420822 217274
rect 419966 217110 420040 217138
rect 419966 216988 419994 217110
rect 420794 216988 420822 217246
rect 421622 217246 421696 217274
rect 421622 216988 421650 217246
rect 422496 217138 422524 218146
rect 423324 217274 423352 219406
rect 424140 218068 424192 218074
rect 424140 218010 424192 218016
rect 422450 217110 422524 217138
rect 423278 217246 423352 217274
rect 422450 216988 422478 217110
rect 423278 216988 423306 217246
rect 424152 217138 424180 218010
rect 424980 217274 425008 222090
rect 425440 218210 425468 231662
rect 426452 222698 426480 231676
rect 426728 231662 427110 231690
rect 426440 222692 426492 222698
rect 426440 222634 426492 222640
rect 426728 220114 426756 231662
rect 427740 229158 427768 231676
rect 427924 231662 428398 231690
rect 428660 231662 429042 231690
rect 429304 231662 429686 231690
rect 429948 231662 430330 231690
rect 430684 231662 430974 231690
rect 431236 231662 431618 231690
rect 432064 231662 432262 231690
rect 432708 231662 432906 231690
rect 433550 231662 433748 231690
rect 427728 229152 427780 229158
rect 427728 229094 427780 229100
rect 426992 222692 427044 222698
rect 426992 222634 427044 222640
rect 426716 220108 426768 220114
rect 426716 220050 426768 220056
rect 426624 218340 426676 218346
rect 426624 218282 426676 218288
rect 425428 218204 425480 218210
rect 425428 218146 425480 218152
rect 425796 218204 425848 218210
rect 425796 218146 425848 218152
rect 424106 217110 424180 217138
rect 424934 217246 425008 217274
rect 424106 216988 424134 217110
rect 424934 216988 424962 217246
rect 425808 217138 425836 218146
rect 426636 217138 426664 218282
rect 427004 218074 427032 222634
rect 427924 218210 427952 231662
rect 428660 219434 428688 231662
rect 429304 222154 429332 231662
rect 429292 222148 429344 222154
rect 429292 222090 429344 222096
rect 429948 219434 429976 231662
rect 430120 220244 430172 220250
rect 430120 220186 430172 220192
rect 428292 219406 428688 219434
rect 429580 219406 429976 219434
rect 427912 218204 427964 218210
rect 427912 218146 427964 218152
rect 428292 218074 428320 219406
rect 429580 218346 429608 219406
rect 429936 218748 429988 218754
rect 429936 218690 429988 218696
rect 429568 218340 429620 218346
rect 429568 218282 429620 218288
rect 428464 218204 428516 218210
rect 428464 218146 428516 218152
rect 426992 218068 427044 218074
rect 426992 218010 427044 218016
rect 427452 218068 427504 218074
rect 427452 218010 427504 218016
rect 428280 218068 428332 218074
rect 428280 218010 428332 218016
rect 427464 217138 427492 218010
rect 428476 217274 428504 218146
rect 429108 218068 429160 218074
rect 429108 218010 429160 218016
rect 425762 217110 425836 217138
rect 426590 217110 426664 217138
rect 427418 217110 427492 217138
rect 428246 217246 428504 217274
rect 425762 216988 425790 217110
rect 426590 216988 426618 217110
rect 427418 216988 427446 217110
rect 428246 216988 428274 217246
rect 429120 217138 429148 218010
rect 429948 217138 429976 218690
rect 430132 218210 430160 220186
rect 430684 219434 430712 231662
rect 431236 219434 431264 231662
rect 432064 220250 432092 231662
rect 432052 220244 432104 220250
rect 432052 220186 432104 220192
rect 431960 220108 432012 220114
rect 431960 220050 432012 220056
rect 430592 219406 430712 219434
rect 430776 219406 431264 219434
rect 430120 218204 430172 218210
rect 430120 218146 430172 218152
rect 430592 218074 430620 219406
rect 430580 218068 430632 218074
rect 430580 218010 430632 218016
rect 430776 217274 430804 219406
rect 431972 218090 432000 220050
rect 432708 218754 432736 231662
rect 433524 229832 433576 229838
rect 433524 229774 433576 229780
rect 433536 229094 433564 229774
rect 433720 229094 433748 231662
rect 434180 229838 434208 231676
rect 434168 229832 434220 229838
rect 434168 229774 434220 229780
rect 433536 229066 433656 229094
rect 433720 229066 433840 229094
rect 432696 218748 432748 218754
rect 432696 218690 432748 218696
rect 433248 218204 433300 218210
rect 433248 218146 433300 218152
rect 429074 217110 429148 217138
rect 429902 217110 429976 217138
rect 430730 217246 430804 217274
rect 431604 218062 432000 218090
rect 432420 218068 432472 218074
rect 429074 216988 429102 217110
rect 429902 216988 429930 217110
rect 430730 216988 430758 217246
rect 431604 217138 431632 218062
rect 432420 218010 432472 218016
rect 432432 217138 432460 218010
rect 433260 217138 433288 218146
rect 433628 217274 433656 229066
rect 433812 218074 433840 229066
rect 434824 220114 434852 231676
rect 435284 231662 435482 231690
rect 436126 231662 436692 231690
rect 434812 220108 434864 220114
rect 434812 220050 434864 220056
rect 435284 218210 435312 231662
rect 436100 230308 436152 230314
rect 436100 230250 436152 230256
rect 435272 218204 435324 218210
rect 435272 218146 435324 218152
rect 435732 218204 435784 218210
rect 435732 218146 435784 218152
rect 433800 218068 433852 218074
rect 433800 218010 433852 218016
rect 434904 218068 434956 218074
rect 434904 218010 434956 218016
rect 433628 217246 434070 217274
rect 431558 217110 431632 217138
rect 432386 217110 432460 217138
rect 433214 217110 433288 217138
rect 431558 216988 431586 217110
rect 432386 216988 432414 217110
rect 433214 216988 433242 217110
rect 434042 216988 434070 217246
rect 434916 217138 434944 218010
rect 435744 217138 435772 218146
rect 436112 217258 436140 230250
rect 436284 220380 436336 220386
rect 436284 220322 436336 220328
rect 436296 218074 436324 220322
rect 436664 218210 436692 231662
rect 436756 230330 436784 231676
rect 437032 231662 437414 231690
rect 437768 231662 438058 231690
rect 436756 230314 436876 230330
rect 436756 230308 436888 230314
rect 436756 230302 436836 230308
rect 436836 230250 436888 230256
rect 437032 220386 437060 231662
rect 437020 220380 437072 220386
rect 437020 220322 437072 220328
rect 437768 219434 437796 231662
rect 438688 230382 438716 231676
rect 439332 230586 439360 231676
rect 439516 231662 439990 231690
rect 440344 231662 440634 231690
rect 439320 230580 439372 230586
rect 439320 230522 439372 230528
rect 439516 230466 439544 231662
rect 438964 230438 439544 230466
rect 438676 230376 438728 230382
rect 438676 230318 438728 230324
rect 438964 219434 438992 230438
rect 439320 230376 439372 230382
rect 439320 230318 439372 230324
rect 439332 219434 439360 230318
rect 437492 219406 437796 219434
rect 438872 219406 438992 219434
rect 439056 219406 439360 219434
rect 436652 218204 436704 218210
rect 436652 218146 436704 218152
rect 437492 218074 437520 219406
rect 438872 218074 438900 219406
rect 436284 218068 436336 218074
rect 436284 218010 436336 218016
rect 436560 218068 436612 218074
rect 436560 218010 436612 218016
rect 437480 218068 437532 218074
rect 437480 218010 437532 218016
rect 438216 218068 438268 218074
rect 438216 218010 438268 218016
rect 438860 218068 438912 218074
rect 438860 218010 438912 218016
rect 436100 217252 436152 217258
rect 436100 217194 436152 217200
rect 436572 217138 436600 218010
rect 437342 217252 437394 217258
rect 437342 217194 437394 217200
rect 434870 217110 434944 217138
rect 435698 217110 435772 217138
rect 436526 217110 436600 217138
rect 434870 216988 434898 217110
rect 435698 216988 435726 217110
rect 436526 216988 436554 217110
rect 437354 216988 437382 217194
rect 438228 217138 438256 218010
rect 439056 217274 439084 219406
rect 440344 218074 440372 231662
rect 440700 230444 440752 230450
rect 440700 230386 440752 230392
rect 439872 218068 439924 218074
rect 439872 218010 439924 218016
rect 440332 218068 440384 218074
rect 440332 218010 440384 218016
rect 438182 217110 438256 217138
rect 439010 217246 439084 217274
rect 438182 216988 438210 217110
rect 439010 216988 439038 217246
rect 439884 217138 439912 218010
rect 440712 217274 440740 230386
rect 441264 229158 441292 231676
rect 441908 230450 441936 231676
rect 442092 231662 442566 231690
rect 443104 231662 443210 231690
rect 441896 230444 441948 230450
rect 441896 230386 441948 230392
rect 442092 230330 442120 231662
rect 441724 230302 442120 230330
rect 441252 229152 441304 229158
rect 441252 229094 441304 229100
rect 441724 219434 441752 230302
rect 442080 229152 442132 229158
rect 442080 229094 442132 229100
rect 442092 229066 442304 229094
rect 441632 219406 441752 219434
rect 441632 218090 441660 219406
rect 439838 217110 439912 217138
rect 440666 217246 440740 217274
rect 441540 218062 441660 218090
rect 439838 216988 439866 217110
rect 440666 216988 440694 217246
rect 441540 217138 441568 218062
rect 442276 217274 442304 229066
rect 443104 217274 443132 231662
rect 443460 230444 443512 230450
rect 443460 230386 443512 230392
rect 443472 229094 443500 230386
rect 443840 230382 443868 231676
rect 443828 230376 443880 230382
rect 443828 230318 443880 230324
rect 444484 230246 444512 231676
rect 444668 231662 445142 231690
rect 444472 230240 444524 230246
rect 444472 230182 444524 230188
rect 444668 229094 444696 231662
rect 444840 230376 444892 230382
rect 444840 230318 444892 230324
rect 444852 229094 444880 230318
rect 445772 229094 445800 231676
rect 446416 229430 446444 231676
rect 446404 229424 446456 229430
rect 446404 229366 446456 229372
rect 443472 229066 443960 229094
rect 444668 229066 444788 229094
rect 444852 229066 445616 229094
rect 445772 229066 446444 229094
rect 443932 217274 443960 229066
rect 444760 217274 444788 229066
rect 445588 217274 445616 229066
rect 446416 217274 446444 229066
rect 447060 227934 447088 231676
rect 447244 231662 447718 231690
rect 447048 227928 447100 227934
rect 447048 227870 447100 227876
rect 447244 219434 447272 231662
rect 447600 230240 447652 230246
rect 447600 230182 447652 230188
rect 447612 219434 447640 230182
rect 448348 229094 448376 231676
rect 448992 229566 449020 231676
rect 449636 230382 449664 231676
rect 449624 230376 449676 230382
rect 449624 230318 449676 230324
rect 448980 229560 449032 229566
rect 448980 229502 449032 229508
rect 448796 229424 448848 229430
rect 448796 229366 448848 229372
rect 448808 229094 448836 229366
rect 450280 229294 450308 231676
rect 450544 230376 450596 230382
rect 450544 230318 450596 230324
rect 450268 229288 450320 229294
rect 450268 229230 450320 229236
rect 450556 229094 450584 230318
rect 450924 229430 450952 231676
rect 451568 230246 451596 231676
rect 452226 231662 452608 231690
rect 451556 230240 451608 230246
rect 451556 230182 451608 230188
rect 451924 229560 451976 229566
rect 451924 229502 451976 229508
rect 450912 229424 450964 229430
rect 450912 229366 450964 229372
rect 451740 229288 451792 229294
rect 451740 229230 451792 229236
rect 448348 229066 448652 229094
rect 448808 229066 448928 229094
rect 450556 229066 450768 229094
rect 447152 219406 447272 219434
rect 447336 219406 447640 219434
rect 442276 217246 442350 217274
rect 443104 217246 443178 217274
rect 443932 217246 444006 217274
rect 444760 217246 444834 217274
rect 445588 217246 445662 217274
rect 446416 217246 446490 217274
rect 447152 217258 447180 219406
rect 447336 217274 447364 219406
rect 441494 217110 441568 217138
rect 441494 216988 441522 217110
rect 442322 216988 442350 217246
rect 443150 216988 443178 217246
rect 443978 216988 444006 217246
rect 444806 216988 444834 217246
rect 445634 216988 445662 217246
rect 446462 216988 446490 217246
rect 447140 217252 447192 217258
rect 447140 217194 447192 217200
rect 447290 217246 447364 217274
rect 448624 217258 448652 229066
rect 448900 217274 448928 229066
rect 450544 227928 450596 227934
rect 450544 227870 450596 227876
rect 450556 217274 450584 227870
rect 450740 218346 450768 229066
rect 451752 219434 451780 229230
rect 451936 229094 451964 229502
rect 451936 229066 452240 229094
rect 451476 219406 451780 219434
rect 450728 218340 450780 218346
rect 450728 218282 450780 218288
rect 451476 217274 451504 219406
rect 448106 217252 448158 217258
rect 447290 216988 447318 217246
rect 448106 217194 448158 217200
rect 448612 217252 448664 217258
rect 448900 217246 448974 217274
rect 448612 217194 448664 217200
rect 448118 216988 448146 217194
rect 448946 216988 448974 217246
rect 449762 217252 449814 217258
rect 450556 217246 450630 217274
rect 449762 217194 449814 217200
rect 449774 216988 449802 217194
rect 450602 216988 450630 217246
rect 451430 217246 451504 217274
rect 452212 217274 452240 229066
rect 452580 222154 452608 231662
rect 452856 230382 452884 231676
rect 452844 230376 452896 230382
rect 452844 230318 452896 230324
rect 453500 230246 453528 231676
rect 453304 230240 453356 230246
rect 453304 230182 453356 230188
rect 453488 230240 453540 230246
rect 453488 230182 453540 230188
rect 453028 229424 453080 229430
rect 453028 229366 453080 229372
rect 452568 222148 452620 222154
rect 452568 222090 452620 222096
rect 453040 217274 453068 229366
rect 453316 218074 453344 230182
rect 454144 230110 454172 231676
rect 454316 230376 454368 230382
rect 454316 230318 454368 230324
rect 454132 230104 454184 230110
rect 454132 230046 454184 230052
rect 454328 229094 454356 230318
rect 454788 229094 454816 231676
rect 455432 230382 455460 231676
rect 455420 230376 455472 230382
rect 455420 230318 455472 230324
rect 455788 230240 455840 230246
rect 455788 230182 455840 230188
rect 455328 230104 455380 230110
rect 455328 230046 455380 230052
rect 454328 229066 454724 229094
rect 454788 229066 454908 229094
rect 453856 218340 453908 218346
rect 453856 218282 453908 218288
rect 453304 218068 453356 218074
rect 453304 218010 453356 218016
rect 452212 217246 452286 217274
rect 453040 217246 453114 217274
rect 451430 216988 451458 217246
rect 452258 216988 452286 217246
rect 453086 216988 453114 217246
rect 453868 217138 453896 218282
rect 454696 217274 454724 229066
rect 454880 223582 454908 229066
rect 454868 223576 454920 223582
rect 454868 223518 454920 223524
rect 455340 220726 455368 230046
rect 455604 222148 455656 222154
rect 455604 222090 455656 222096
rect 455328 220720 455380 220726
rect 455328 220662 455380 220668
rect 455616 218074 455644 222090
rect 455800 219434 455828 230182
rect 456076 224534 456104 231676
rect 456064 224528 456116 224534
rect 456064 224470 456116 224476
rect 456720 220862 456748 231676
rect 457168 230376 457220 230382
rect 457168 230318 457220 230324
rect 456708 220856 456760 220862
rect 456708 220798 456760 220804
rect 457180 219434 457208 230318
rect 457364 230042 457392 231676
rect 457352 230036 457404 230042
rect 457352 229978 457404 229984
rect 458008 229094 458036 231676
rect 458008 229066 458128 229094
rect 455800 219406 456380 219434
rect 457180 219406 458036 219434
rect 455420 218068 455472 218074
rect 455420 218010 455472 218016
rect 455604 218068 455656 218074
rect 455604 218010 455656 218016
rect 455432 217274 455460 218010
rect 456352 217274 456380 219406
rect 457168 218068 457220 218074
rect 457168 218010 457220 218016
rect 454696 217246 454770 217274
rect 455432 217246 455598 217274
rect 456352 217246 456426 217274
rect 453868 217110 453942 217138
rect 453914 216988 453942 217110
rect 454742 216988 454770 217246
rect 455570 216988 455598 217246
rect 456398 216988 456426 217246
rect 457180 217138 457208 218010
rect 458008 217274 458036 219406
rect 458100 218498 458128 229066
rect 458652 226302 458680 231676
rect 459310 231662 459508 231690
rect 458640 226296 458692 226302
rect 458640 226238 458692 226244
rect 458824 220720 458876 220726
rect 458824 220662 458876 220668
rect 458100 218470 458220 218498
rect 458192 218414 458220 218470
rect 458180 218408 458232 218414
rect 458180 218350 458232 218356
rect 458836 217274 458864 220662
rect 459480 220250 459508 231662
rect 459744 224528 459796 224534
rect 459744 224470 459796 224476
rect 459468 220244 459520 220250
rect 459468 220186 459520 220192
rect 459756 217274 459784 224470
rect 459940 222902 459968 231676
rect 460584 224942 460612 231676
rect 461242 231662 461716 231690
rect 461886 231662 462176 231690
rect 461688 229094 461716 231662
rect 461688 229066 461992 229094
rect 460572 224936 460624 224942
rect 460572 224878 460624 224884
rect 460480 223576 460532 223582
rect 460480 223518 460532 223524
rect 459928 222896 459980 222902
rect 459928 222838 459980 222844
rect 458008 217246 458082 217274
rect 458836 217246 458910 217274
rect 457180 217110 457254 217138
rect 457226 216988 457254 217110
rect 458054 216988 458082 217246
rect 458882 216988 458910 217246
rect 459710 217246 459784 217274
rect 460492 217274 460520 223518
rect 461308 218340 461360 218346
rect 461308 218282 461360 218288
rect 460492 217246 460566 217274
rect 459710 216988 459738 217246
rect 460538 216988 460566 217246
rect 461320 217138 461348 218282
rect 461964 218210 461992 229066
rect 462148 222154 462176 231662
rect 462516 224806 462544 231676
rect 462964 226296 463016 226302
rect 462964 226238 463016 226244
rect 462504 224800 462556 224806
rect 462504 224742 462556 224748
rect 462136 222148 462188 222154
rect 462136 222090 462188 222096
rect 462136 220856 462188 220862
rect 462136 220798 462188 220804
rect 461952 218204 462004 218210
rect 461952 218146 462004 218152
rect 462148 217274 462176 220798
rect 462976 217274 463004 226238
rect 463160 225418 463188 231676
rect 463804 230382 463832 231676
rect 464462 231662 465028 231690
rect 465106 231662 465488 231690
rect 465750 231662 465948 231690
rect 463792 230376 463844 230382
rect 463792 230318 463844 230324
rect 463884 230036 463936 230042
rect 463884 229978 463936 229984
rect 463148 225412 463200 225418
rect 463148 225354 463200 225360
rect 463148 224936 463200 224942
rect 463148 224878 463200 224884
rect 463160 218074 463188 224878
rect 463148 218068 463200 218074
rect 463148 218010 463200 218016
rect 463896 217274 463924 229978
rect 465000 219638 465028 231662
rect 465460 229770 465488 231662
rect 465724 230376 465776 230382
rect 465724 230318 465776 230324
rect 465448 229764 465500 229770
rect 465448 229706 465500 229712
rect 465736 220726 465764 230318
rect 465920 227662 465948 231662
rect 466104 231662 466394 231690
rect 465908 227656 465960 227662
rect 465908 227598 465960 227604
rect 466104 220862 466132 231662
rect 467024 229906 467052 231676
rect 467012 229900 467064 229906
rect 467012 229842 467064 229848
rect 467472 229764 467524 229770
rect 467472 229706 467524 229712
rect 467288 225412 467340 225418
rect 467288 225354 467340 225360
rect 467104 222896 467156 222902
rect 467104 222838 467156 222844
rect 466092 220856 466144 220862
rect 466092 220798 466144 220804
rect 465724 220720 465776 220726
rect 465724 220662 465776 220668
rect 465448 220244 465500 220250
rect 465448 220186 465500 220192
rect 464988 219632 465040 219638
rect 464988 219574 465040 219580
rect 464620 218068 464672 218074
rect 464620 218010 464672 218016
rect 462148 217246 462222 217274
rect 462976 217246 463050 217274
rect 461320 217110 461394 217138
rect 461366 216988 461394 217110
rect 462194 216988 462222 217246
rect 463022 216988 463050 217246
rect 463850 217246 463924 217274
rect 463850 216988 463878 217246
rect 464632 217138 464660 218010
rect 465460 217274 465488 220186
rect 466276 218204 466328 218210
rect 466276 218146 466328 218152
rect 465460 217246 465534 217274
rect 464632 217110 464706 217138
rect 464678 216988 464706 217110
rect 465506 216988 465534 217246
rect 466288 217138 466316 218146
rect 467116 217274 467144 222838
rect 467300 218074 467328 225354
rect 467484 222902 467512 229706
rect 467668 225622 467696 231676
rect 468312 230246 468340 231676
rect 468300 230240 468352 230246
rect 468300 230182 468352 230188
rect 467656 225616 467708 225622
rect 467656 225558 467708 225564
rect 467472 222896 467524 222902
rect 467472 222838 467524 222844
rect 468760 222148 468812 222154
rect 468760 222090 468812 222096
rect 467288 218068 467340 218074
rect 467288 218010 467340 218016
rect 467932 218068 467984 218074
rect 467932 218010 467984 218016
rect 467116 217246 467190 217274
rect 466288 217110 466362 217138
rect 466334 216988 466362 217110
rect 467162 216988 467190 217246
rect 467944 217138 467972 218010
rect 468772 217274 468800 222090
rect 468956 221474 468984 231676
rect 469128 230240 469180 230246
rect 469128 230182 469180 230188
rect 468944 221468 468996 221474
rect 468944 221410 468996 221416
rect 469140 220522 469168 230182
rect 469600 229770 469628 231676
rect 469588 229764 469640 229770
rect 469588 229706 469640 229712
rect 469864 227656 469916 227662
rect 469864 227598 469916 227604
rect 469312 224800 469364 224806
rect 469312 224742 469364 224748
rect 469128 220516 469180 220522
rect 469128 220458 469180 220464
rect 468772 217246 468846 217274
rect 469324 217258 469352 224742
rect 469588 220720 469640 220726
rect 469588 220662 469640 220668
rect 469600 217274 469628 220662
rect 469876 218618 469904 227598
rect 470244 224262 470272 231676
rect 470888 230382 470916 231676
rect 470876 230376 470928 230382
rect 470876 230318 470928 230324
rect 471532 227798 471560 231676
rect 472176 230382 472204 231676
rect 472834 231662 473032 231690
rect 471888 230376 471940 230382
rect 471888 230318 471940 230324
rect 472164 230376 472216 230382
rect 472164 230318 472216 230324
rect 471520 227792 471572 227798
rect 471520 227734 471572 227740
rect 470232 224256 470284 224262
rect 470232 224198 470284 224204
rect 471900 222154 471928 230318
rect 471888 222148 471940 222154
rect 471888 222090 471940 222096
rect 471336 220856 471388 220862
rect 471336 220798 471388 220804
rect 471348 218754 471376 220798
rect 473004 220250 473032 231662
rect 473176 230376 473228 230382
rect 473176 230318 473228 230324
rect 473188 220386 473216 230318
rect 473464 223582 473492 231676
rect 474122 231662 474504 231690
rect 474004 229900 474056 229906
rect 474004 229842 474056 229848
rect 473452 223576 473504 223582
rect 473452 223518 473504 223524
rect 473728 222896 473780 222902
rect 473728 222838 473780 222844
rect 473176 220380 473228 220386
rect 473176 220322 473228 220328
rect 472992 220244 473044 220250
rect 472992 220186 473044 220192
rect 472072 219632 472124 219638
rect 472072 219574 472124 219580
rect 471336 218748 471388 218754
rect 471336 218690 471388 218696
rect 469864 218612 469916 218618
rect 469864 218554 469916 218560
rect 471244 218612 471296 218618
rect 471244 218554 471296 218560
rect 467944 217110 468018 217138
rect 467990 216988 468018 217110
rect 468818 216988 468846 217246
rect 469312 217252 469364 217258
rect 469600 217246 469674 217274
rect 469312 217194 469364 217200
rect 469646 216988 469674 217246
rect 470462 217252 470514 217258
rect 470462 217194 470514 217200
rect 470474 216988 470502 217194
rect 471256 217138 471284 218554
rect 472084 217274 472112 219574
rect 472900 218748 472952 218754
rect 472900 218690 472952 218696
rect 472912 217274 472940 218690
rect 473740 217274 473768 222838
rect 474016 220794 474044 229842
rect 474476 228410 474504 231662
rect 474464 228404 474516 228410
rect 474464 228346 474516 228352
rect 474752 226506 474780 231676
rect 475410 231662 475884 231690
rect 474740 226500 474792 226506
rect 474740 226442 474792 226448
rect 475568 223576 475620 223582
rect 475568 223518 475620 223524
rect 474004 220788 474056 220794
rect 474004 220730 474056 220736
rect 475384 220788 475436 220794
rect 475384 220730 475436 220736
rect 474556 220516 474608 220522
rect 474556 220458 474608 220464
rect 474568 217274 474596 220458
rect 475396 217274 475424 220730
rect 475580 218618 475608 223518
rect 475856 221610 475884 231662
rect 476040 229498 476068 231676
rect 476684 229906 476712 231676
rect 476672 229900 476724 229906
rect 476672 229842 476724 229848
rect 476764 229764 476816 229770
rect 476764 229706 476816 229712
rect 476028 229492 476080 229498
rect 476028 229434 476080 229440
rect 476580 225616 476632 225622
rect 476580 225558 476632 225564
rect 475844 221604 475896 221610
rect 475844 221546 475896 221552
rect 476212 221468 476264 221474
rect 476212 221410 476264 221416
rect 475568 218612 475620 218618
rect 475568 218554 475620 218560
rect 476224 217274 476252 221410
rect 476592 217274 476620 225558
rect 476776 220794 476804 229706
rect 477328 225622 477356 231676
rect 477986 231662 478368 231690
rect 478630 231662 478828 231690
rect 477316 225616 477368 225622
rect 477316 225558 477368 225564
rect 477868 222148 477920 222154
rect 477868 222090 477920 222096
rect 476764 220788 476816 220794
rect 476764 220730 476816 220736
rect 477880 217274 477908 222090
rect 478340 220114 478368 231662
rect 478604 229492 478656 229498
rect 478604 229434 478656 229440
rect 478616 227186 478644 229434
rect 478800 229094 478828 231662
rect 479260 229770 479288 231676
rect 479248 229764 479300 229770
rect 479248 229706 479300 229712
rect 478800 229066 478920 229094
rect 478892 228818 478920 229066
rect 478880 228812 478932 228818
rect 478880 228754 478932 228760
rect 479524 227792 479576 227798
rect 479524 227734 479576 227740
rect 478604 227180 478656 227186
rect 478604 227122 478656 227128
rect 478696 220788 478748 220794
rect 478696 220730 478748 220736
rect 478328 220108 478380 220114
rect 478328 220050 478380 220056
rect 478708 217274 478736 220730
rect 479536 217274 479564 227734
rect 479904 222902 479932 231676
rect 480548 224398 480576 231676
rect 481192 225758 481220 231676
rect 481836 229906 481864 231676
rect 482494 231662 482968 231690
rect 481640 229900 481692 229906
rect 481640 229842 481692 229848
rect 481824 229900 481876 229906
rect 481824 229842 481876 229848
rect 481652 226370 481680 229842
rect 482744 226500 482796 226506
rect 482744 226442 482796 226448
rect 481640 226364 481692 226370
rect 481640 226306 481692 226312
rect 481180 225752 481232 225758
rect 481180 225694 481232 225700
rect 480536 224392 480588 224398
rect 480536 224334 480588 224340
rect 480352 224256 480404 224262
rect 480352 224198 480404 224204
rect 479892 222896 479944 222902
rect 479892 222838 479944 222844
rect 480364 217274 480392 224198
rect 482756 222630 482784 226442
rect 482744 222624 482796 222630
rect 482744 222566 482796 222572
rect 481180 220380 481232 220386
rect 481180 220322 481232 220328
rect 481192 217274 481220 220322
rect 482008 220244 482060 220250
rect 482008 220186 482060 220192
rect 482020 217274 482048 220186
rect 482756 218754 482784 222566
rect 482940 220250 482968 231662
rect 483124 223174 483152 231676
rect 483768 224262 483796 231676
rect 484426 231662 484808 231690
rect 484584 228404 484636 228410
rect 484584 228346 484636 228352
rect 483756 224256 483808 224262
rect 483756 224198 483808 224204
rect 483112 223168 483164 223174
rect 483112 223110 483164 223116
rect 484596 222358 484624 228346
rect 484584 222352 484636 222358
rect 484584 222294 484636 222300
rect 483756 221468 483808 221474
rect 483756 221410 483808 221416
rect 482928 220244 482980 220250
rect 482928 220186 482980 220192
rect 482744 218748 482796 218754
rect 482744 218690 482796 218696
rect 482836 218612 482888 218618
rect 482836 218554 482888 218560
rect 472084 217246 472158 217274
rect 472912 217246 472986 217274
rect 473740 217246 473814 217274
rect 474568 217246 474642 217274
rect 475396 217246 475470 217274
rect 476224 217246 476298 217274
rect 476592 217246 477126 217274
rect 477880 217246 477954 217274
rect 478708 217246 478782 217274
rect 479536 217246 479610 217274
rect 480364 217246 480438 217274
rect 481192 217246 481266 217274
rect 482020 217246 482094 217274
rect 471256 217110 471330 217138
rect 471302 216988 471330 217110
rect 472130 216988 472158 217246
rect 472958 216988 472986 217246
rect 473786 216988 473814 217246
rect 474614 216988 474642 217246
rect 475442 216988 475470 217246
rect 476270 216988 476298 217246
rect 477098 216988 477126 217246
rect 477926 216988 477954 217246
rect 478754 216988 478782 217246
rect 479582 216988 479610 217246
rect 480410 216988 480438 217246
rect 481238 216988 481266 217246
rect 482066 216988 482094 217246
rect 482848 217138 482876 218554
rect 483768 217274 483796 221410
rect 484596 217274 484624 222294
rect 484780 221746 484808 231662
rect 485056 228410 485084 231676
rect 485700 228546 485728 231676
rect 486358 231662 486648 231690
rect 485688 228540 485740 228546
rect 485688 228482 485740 228488
rect 485044 228404 485096 228410
rect 485044 228346 485096 228352
rect 486620 223038 486648 231662
rect 486792 227180 486844 227186
rect 486792 227122 486844 227128
rect 486608 223032 486660 223038
rect 486608 222974 486660 222980
rect 484768 221740 484820 221746
rect 484768 221682 484820 221688
rect 486148 221604 486200 221610
rect 486148 221546 486200 221552
rect 485320 218748 485372 218754
rect 485320 218690 485372 218696
rect 483722 217246 483796 217274
rect 484550 217246 484624 217274
rect 485332 217274 485360 218690
rect 486160 217274 486188 221546
rect 486804 219434 486832 227122
rect 486988 227050 487016 231676
rect 487632 230382 487660 231676
rect 487620 230376 487672 230382
rect 487620 230318 487672 230324
rect 488080 229764 488132 229770
rect 488080 229706 488132 229712
rect 486976 227044 487028 227050
rect 486976 226986 487028 226992
rect 488092 226370 488120 229706
rect 488276 229294 488304 231676
rect 488934 231662 489408 231690
rect 488448 230376 488500 230382
rect 488448 230318 488500 230324
rect 488264 229288 488316 229294
rect 488264 229230 488316 229236
rect 487804 226364 487856 226370
rect 487804 226306 487856 226312
rect 488080 226364 488132 226370
rect 488080 226306 488132 226312
rect 486974 219464 487030 219473
rect 486804 219408 486974 219434
rect 486804 219406 487030 219408
rect 486974 219399 487030 219406
rect 486988 217274 487016 219399
rect 487816 218113 487844 226306
rect 488460 220522 488488 230318
rect 489380 225622 489408 231662
rect 489564 229094 489592 231676
rect 490208 230246 490236 231676
rect 490866 231662 491248 231690
rect 490196 230240 490248 230246
rect 490196 230182 490248 230188
rect 489920 229900 489972 229906
rect 489920 229842 489972 229848
rect 489564 229066 489684 229094
rect 488724 225616 488776 225622
rect 488724 225558 488776 225564
rect 489368 225616 489420 225622
rect 489368 225558 489420 225564
rect 488448 220516 488500 220522
rect 488448 220458 488500 220464
rect 487802 218104 487858 218113
rect 487802 218039 487858 218048
rect 487816 217274 487844 218039
rect 488736 217274 488764 225558
rect 489656 220114 489684 229066
rect 489932 227798 489960 229842
rect 490380 229288 490432 229294
rect 490380 229230 490432 229236
rect 490196 228812 490248 228818
rect 490196 228754 490248 228760
rect 489920 227792 489972 227798
rect 489920 227734 489972 227740
rect 490012 226364 490064 226370
rect 490012 226306 490064 226312
rect 490024 222426 490052 226306
rect 490012 222420 490064 222426
rect 490012 222362 490064 222368
rect 489460 220108 489512 220114
rect 489460 220050 489512 220056
rect 489644 220108 489696 220114
rect 489644 220050 489696 220056
rect 485332 217246 485406 217274
rect 486160 217246 486234 217274
rect 486988 217246 487062 217274
rect 487816 217246 487890 217274
rect 482848 217110 482922 217138
rect 482894 216988 482922 217110
rect 483722 216988 483750 217246
rect 484550 216988 484578 217246
rect 485378 216988 485406 217246
rect 486206 216988 486234 217246
rect 487034 216988 487062 217246
rect 487862 216988 487890 217246
rect 488690 217246 488764 217274
rect 489472 217274 489500 220050
rect 490024 219434 490052 222362
rect 489932 219406 490052 219434
rect 490208 219434 490236 228754
rect 490392 227186 490420 229230
rect 491220 229094 491248 231662
rect 491496 230110 491524 231676
rect 491484 230104 491536 230110
rect 491484 230046 491536 230052
rect 492140 229770 492168 231676
rect 492798 231662 493088 231690
rect 492496 230104 492548 230110
rect 492496 230046 492548 230052
rect 492128 229764 492180 229770
rect 492128 229706 492180 229712
rect 491220 229066 491340 229094
rect 490380 227180 490432 227186
rect 490380 227122 490432 227128
rect 491312 224534 491340 229066
rect 491300 224528 491352 224534
rect 491300 224470 491352 224476
rect 492036 222896 492088 222902
rect 492036 222838 492088 222844
rect 490208 219406 490420 219434
rect 489472 217246 489546 217274
rect 489932 217258 489960 219406
rect 490392 218657 490420 219406
rect 490378 218648 490434 218657
rect 490378 218583 490434 218592
rect 490392 217274 490420 218583
rect 492048 218074 492076 222838
rect 492508 221882 492536 230046
rect 492680 225752 492732 225758
rect 492680 225694 492732 225700
rect 492496 221876 492548 221882
rect 492496 221818 492548 221824
rect 492692 218385 492720 225694
rect 492864 224392 492916 224398
rect 492864 224334 492916 224340
rect 492678 218376 492734 218385
rect 492678 218311 492734 218320
rect 492036 218068 492088 218074
rect 492036 218010 492088 218016
rect 488690 217161 488718 217246
rect 488676 217152 488732 217161
rect 488676 217087 488732 217096
rect 488690 216988 488718 217087
rect 489518 216988 489546 217246
rect 489920 217252 489972 217258
rect 489920 217194 489972 217200
rect 490346 217246 490420 217274
rect 491162 217252 491214 217258
rect 490346 216988 490374 217246
rect 491162 217194 491214 217200
rect 491174 216988 491202 217194
rect 492048 217138 492076 218010
rect 492876 217274 492904 224334
rect 493060 223310 493088 231662
rect 493428 230382 493456 231676
rect 493416 230376 493468 230382
rect 493416 230318 493468 230324
rect 493784 230240 493836 230246
rect 493784 230182 493836 230188
rect 493796 225758 493824 230182
rect 493784 225752 493836 225758
rect 493784 225694 493836 225700
rect 494072 224670 494100 231676
rect 494730 231662 495112 231690
rect 494704 227792 494756 227798
rect 494704 227734 494756 227740
rect 494060 224664 494112 224670
rect 494060 224606 494112 224612
rect 493048 223304 493100 223310
rect 493048 223246 493100 223252
rect 494716 218929 494744 227734
rect 495084 227458 495112 231662
rect 495360 229294 495388 231676
rect 496004 229906 496032 231676
rect 496188 231662 496662 231690
rect 495992 229900 496044 229906
rect 495992 229842 496044 229848
rect 495348 229288 495400 229294
rect 495348 229230 495400 229236
rect 496188 229094 496216 231662
rect 497292 230382 497320 231676
rect 497476 231662 497950 231690
rect 496360 230376 496412 230382
rect 496360 230318 496412 230324
rect 497280 230376 497332 230382
rect 497280 230318 497332 230324
rect 496372 229094 496400 230318
rect 496188 229066 496308 229094
rect 496372 229066 496492 229094
rect 495072 227452 495124 227458
rect 495072 227394 495124 227400
rect 496084 223168 496136 223174
rect 496084 223110 496136 223116
rect 495348 220244 495400 220250
rect 495348 220186 495400 220192
rect 494702 218920 494758 218929
rect 494532 218878 494702 218906
rect 493782 218376 493838 218385
rect 493782 218311 493838 218320
rect 493796 217297 493824 218311
rect 492002 217110 492076 217138
rect 492830 217246 492904 217274
rect 493782 217288 493838 217297
rect 492002 216988 492030 217110
rect 492830 216988 492858 217246
rect 494532 217274 494560 218878
rect 494702 218855 494758 218864
rect 495360 217297 495388 220186
rect 493782 217223 493838 217232
rect 494486 217246 494560 217274
rect 495346 217288 495402 217297
rect 493796 217138 493824 217223
rect 493658 217110 493824 217138
rect 493658 216988 493686 217110
rect 494486 216988 494514 217246
rect 495346 217223 495402 217232
rect 495360 217138 495388 217223
rect 495314 217110 495388 217138
rect 496096 217138 496124 223110
rect 496280 221610 496308 229066
rect 496268 221604 496320 221610
rect 496268 221546 496320 221552
rect 496464 220386 496492 229066
rect 496912 224256 496964 224262
rect 496912 224198 496964 224204
rect 496452 220380 496504 220386
rect 496452 220322 496504 220328
rect 496924 218385 496952 224198
rect 497476 220250 497504 231662
rect 498108 230376 498160 230382
rect 498108 230318 498160 230324
rect 498120 226030 498148 230318
rect 498580 228682 498608 231676
rect 498568 228676 498620 228682
rect 498568 228618 498620 228624
rect 498292 228540 498344 228546
rect 498292 228482 498344 228488
rect 498108 226024 498160 226030
rect 498108 225966 498160 225972
rect 497740 221740 497792 221746
rect 497740 221682 497792 221688
rect 497752 220969 497780 221682
rect 497738 220960 497794 220969
rect 497738 220895 497794 220904
rect 497464 220244 497516 220250
rect 497464 220186 497516 220192
rect 496910 218376 496966 218385
rect 496910 218311 496966 218320
rect 496924 217138 496952 218311
rect 497752 217274 497780 220895
rect 497752 217246 497826 217274
rect 498304 217258 498332 228482
rect 498568 228404 498620 228410
rect 498568 228346 498620 228352
rect 498580 224954 498608 228346
rect 498488 224926 498608 224954
rect 498488 217297 498516 224926
rect 499224 224398 499252 231676
rect 499868 228818 499896 231676
rect 500526 231662 500816 231690
rect 500224 229288 500276 229294
rect 500224 229230 500276 229236
rect 499856 228812 499908 228818
rect 499856 228754 499908 228760
rect 500236 224954 500264 229230
rect 500236 224926 500448 224954
rect 499212 224392 499264 224398
rect 499212 224334 499264 224340
rect 500040 223032 500092 223038
rect 500040 222974 500092 222980
rect 500052 218482 500080 222974
rect 500224 222488 500276 222494
rect 500224 222430 500276 222436
rect 500236 222222 500264 222430
rect 500224 222216 500276 222222
rect 500224 222158 500276 222164
rect 500420 220794 500448 224926
rect 500788 222902 500816 231662
rect 500960 227044 501012 227050
rect 500960 226986 501012 226992
rect 500972 224954 501000 226986
rect 501156 225894 501184 231676
rect 501340 231662 501814 231690
rect 501144 225888 501196 225894
rect 501144 225830 501196 225836
rect 500972 224926 501092 224954
rect 500776 222896 500828 222902
rect 500776 222838 500828 222844
rect 500408 220788 500460 220794
rect 500408 220730 500460 220736
rect 501064 219502 501092 224926
rect 501340 221746 501368 231662
rect 502444 228546 502472 231676
rect 503102 231662 503392 231690
rect 502432 228540 502484 228546
rect 502432 228482 502484 228488
rect 503168 227180 503220 227186
rect 503168 227122 503220 227128
rect 502984 225616 503036 225622
rect 502984 225558 503036 225564
rect 501328 221740 501380 221746
rect 501328 221682 501380 221688
rect 501880 220516 501932 220522
rect 501880 220458 501932 220464
rect 501052 219496 501104 219502
rect 501052 219438 501104 219444
rect 500040 218476 500092 218482
rect 500040 218418 500092 218424
rect 498474 217288 498530 217297
rect 496096 217110 496170 217138
rect 496924 217110 496998 217138
rect 495314 216988 495342 217110
rect 496142 216988 496170 217110
rect 496970 216988 496998 217110
rect 497798 216988 497826 217246
rect 498292 217252 498344 217258
rect 500052 217274 500080 218418
rect 501064 217274 501092 219438
rect 498474 217223 498530 217232
rect 499442 217252 499494 217258
rect 498292 217194 498344 217200
rect 498488 217138 498516 217223
rect 500052 217246 500310 217274
rect 501064 217246 501138 217274
rect 499442 217194 499494 217200
rect 498488 217110 498654 217138
rect 498626 216988 498654 217110
rect 499454 216988 499482 217194
rect 500282 216988 500310 217246
rect 501110 216988 501138 217246
rect 501892 217138 501920 220458
rect 502996 217258 503024 225558
rect 503180 218346 503208 227122
rect 503364 223174 503392 231662
rect 503732 229158 503760 231676
rect 503720 229152 503772 229158
rect 503720 229094 503772 229100
rect 504376 224126 504404 231676
rect 504928 231662 505034 231690
rect 504928 227186 504956 231662
rect 505100 229764 505152 229770
rect 505100 229706 505152 229712
rect 504916 227180 504968 227186
rect 504916 227122 504968 227128
rect 504364 224120 504416 224126
rect 504364 224062 504416 224068
rect 505112 223786 505140 229706
rect 505664 229430 505692 231676
rect 505652 229424 505704 229430
rect 505652 229366 505704 229372
rect 506308 227050 506336 231676
rect 506296 227044 506348 227050
rect 506296 226986 506348 226992
rect 505284 225752 505336 225758
rect 505284 225694 505336 225700
rect 505100 223780 505152 223786
rect 505100 223722 505152 223728
rect 505296 223650 505324 225694
rect 506952 224806 506980 231676
rect 507124 229900 507176 229906
rect 507124 229842 507176 229848
rect 507136 228410 507164 229842
rect 507596 229770 507624 231676
rect 507584 229764 507636 229770
rect 507584 229706 507636 229712
rect 507124 228404 507176 228410
rect 507124 228346 507176 228352
rect 506940 224800 506992 224806
rect 506940 224742 506992 224748
rect 506020 224528 506072 224534
rect 506020 224470 506072 224476
rect 505284 223644 505336 223650
rect 505284 223586 505336 223592
rect 503352 223168 503404 223174
rect 503352 223110 503404 223116
rect 504364 220108 504416 220114
rect 504364 220050 504416 220056
rect 503168 218340 503220 218346
rect 503168 218282 503220 218288
rect 502984 217252 503036 217258
rect 502984 217194 503036 217200
rect 503180 217138 503208 218282
rect 503582 217252 503634 217258
rect 503582 217194 503634 217200
rect 501892 217110 501966 217138
rect 501938 216988 501966 217110
rect 502766 217110 503208 217138
rect 503594 217122 503622 217194
rect 504376 217138 504404 220050
rect 505296 217274 505324 223586
rect 506032 219638 506060 224470
rect 507676 223780 507728 223786
rect 507676 223722 507728 223728
rect 506848 221876 506900 221882
rect 506848 221818 506900 221824
rect 506020 219632 506072 219638
rect 506020 219574 506072 219580
rect 505652 218068 505704 218074
rect 505652 218010 505704 218016
rect 505664 217569 505692 218010
rect 505650 217560 505706 217569
rect 505650 217495 505706 217504
rect 505250 217246 505324 217274
rect 503582 217116 503634 217122
rect 502766 216988 502794 217110
rect 504376 217110 504450 217138
rect 503582 217058 503634 217064
rect 503594 216988 503622 217058
rect 504422 216988 504450 217110
rect 505250 216988 505278 217246
rect 506032 217138 506060 219574
rect 506860 217138 506888 221818
rect 507688 218210 507716 223722
rect 508240 223038 508268 231676
rect 508884 225758 508912 231676
rect 509528 229906 509556 231676
rect 509516 229900 509568 229906
rect 509516 229842 509568 229848
rect 509884 229152 509936 229158
rect 509884 229094 509936 229100
rect 508872 225752 508924 225758
rect 508872 225694 508924 225700
rect 508504 223304 508556 223310
rect 508504 223246 508556 223252
rect 508228 223032 508280 223038
rect 508228 222974 508280 222980
rect 507676 218204 507728 218210
rect 507676 218146 507728 218152
rect 507688 217138 507716 218146
rect 508516 217841 508544 223246
rect 509896 220658 509924 229094
rect 510172 225622 510200 231676
rect 510816 230382 510844 231676
rect 510804 230376 510856 230382
rect 510804 230318 510856 230324
rect 511460 230246 511488 231676
rect 511908 230376 511960 230382
rect 511908 230318 511960 230324
rect 511448 230240 511500 230246
rect 511448 230182 511500 230188
rect 510988 229424 511040 229430
rect 510988 229366 511040 229372
rect 511000 227322 511028 229366
rect 511920 229094 511948 230318
rect 511644 229066 511948 229094
rect 511172 227452 511224 227458
rect 511172 227394 511224 227400
rect 510988 227316 511040 227322
rect 510988 227258 511040 227264
rect 510160 225616 510212 225622
rect 510160 225558 510212 225564
rect 511184 224954 511212 227394
rect 511092 224926 511212 224954
rect 510160 224664 510212 224670
rect 510160 224606 510212 224612
rect 509884 220652 509936 220658
rect 509884 220594 509936 220600
rect 509332 220380 509384 220386
rect 509332 220322 509384 220328
rect 508502 217832 508558 217841
rect 508502 217767 508558 217776
rect 508516 217138 508544 217767
rect 509344 217274 509372 220322
rect 510172 217841 510200 224606
rect 510158 217832 510214 217841
rect 510158 217767 510214 217776
rect 509344 217246 509418 217274
rect 506032 217110 506106 217138
rect 506860 217110 506934 217138
rect 507688 217110 507762 217138
rect 508516 217110 508590 217138
rect 506078 216988 506106 217110
rect 506906 216988 506934 217110
rect 507734 216988 507762 217110
rect 508562 216988 508590 217110
rect 509390 216988 509418 217246
rect 510172 217138 510200 217767
rect 511092 217274 511120 224926
rect 511644 220522 511672 229066
rect 512104 228682 512132 231676
rect 512762 231662 513144 231690
rect 512092 228676 512144 228682
rect 512092 228618 512144 228624
rect 512736 228404 512788 228410
rect 512736 228346 512788 228352
rect 511816 220788 511868 220794
rect 511816 220730 511868 220736
rect 511632 220516 511684 220522
rect 511632 220458 511684 220464
rect 511046 217246 511120 217274
rect 511046 217190 511074 217246
rect 511034 217184 511086 217190
rect 510172 217110 510246 217138
rect 511034 217126 511086 217132
rect 511828 217138 511856 220730
rect 512748 218074 512776 228346
rect 513116 220114 513144 231662
rect 513392 229294 513420 231676
rect 513380 229288 513432 229294
rect 513380 229230 513432 229236
rect 514036 227458 514064 231676
rect 514024 227452 514076 227458
rect 514024 227394 514076 227400
rect 514300 226024 514352 226030
rect 514300 225966 514352 225972
rect 513564 221604 513616 221610
rect 513564 221546 513616 221552
rect 513576 221241 513604 221546
rect 513562 221232 513618 221241
rect 513562 221167 513618 221176
rect 513104 220108 513156 220114
rect 513104 220050 513156 220056
rect 512736 218068 512788 218074
rect 512736 218010 512788 218016
rect 512748 217274 512776 218010
rect 513576 217274 513604 221167
rect 512702 217246 512776 217274
rect 513530 217246 513604 217274
rect 514312 217274 514340 225966
rect 514680 223310 514708 231676
rect 515324 230042 515352 231676
rect 515312 230036 515364 230042
rect 515312 229978 515364 229984
rect 515404 229900 515456 229906
rect 515404 229842 515456 229848
rect 514668 223304 514720 223310
rect 514668 223246 514720 223252
rect 515416 220386 515444 229842
rect 515772 228812 515824 228818
rect 515772 228754 515824 228760
rect 515784 221882 515812 228754
rect 515968 224534 515996 231676
rect 516612 226030 516640 231676
rect 517256 229906 517284 231676
rect 517520 230240 517572 230246
rect 517520 230182 517572 230188
rect 517244 229900 517296 229906
rect 517244 229842 517296 229848
rect 516784 229764 516836 229770
rect 516784 229706 516836 229712
rect 516600 226024 516652 226030
rect 516600 225966 516652 225972
rect 515956 224528 516008 224534
rect 515956 224470 516008 224476
rect 516600 224392 516652 224398
rect 516600 224334 516652 224340
rect 515772 221876 515824 221882
rect 515772 221818 515824 221824
rect 515404 220380 515456 220386
rect 515404 220322 515456 220328
rect 515220 220244 515272 220250
rect 515220 220186 515272 220192
rect 515232 219473 515260 220186
rect 515218 219464 515274 219473
rect 515218 219399 515274 219408
rect 515784 219434 515812 221818
rect 516612 219434 516640 224334
rect 516796 222018 516824 229706
rect 517532 223446 517560 230182
rect 517704 228948 517756 228954
rect 517704 228890 517756 228896
rect 517716 223922 517744 228890
rect 517900 228682 517928 231676
rect 518544 228818 518572 231676
rect 519188 229158 519216 231676
rect 519360 229288 519412 229294
rect 519360 229230 519412 229236
rect 519176 229152 519228 229158
rect 519176 229094 519228 229100
rect 518532 228812 518584 228818
rect 518532 228754 518584 228760
rect 517888 228676 517940 228682
rect 517888 228618 517940 228624
rect 519176 225888 519228 225894
rect 519176 225830 519228 225836
rect 517704 223916 517756 223922
rect 517704 223858 517756 223864
rect 517520 223440 517572 223446
rect 517520 223382 517572 223388
rect 517520 222896 517572 222902
rect 517520 222838 517572 222844
rect 516784 222012 516836 222018
rect 516784 221954 516836 221960
rect 517532 221134 517560 222838
rect 517520 221128 517572 221134
rect 517520 221070 517572 221076
rect 517716 219434 517744 223858
rect 518440 221128 518492 221134
rect 518440 221070 518492 221076
rect 515784 219406 515996 219434
rect 516612 219406 516824 219434
rect 515232 217274 515260 219399
rect 514312 217246 514386 217274
rect 510218 216988 510246 217110
rect 511046 216988 511074 217126
rect 511828 217110 511902 217138
rect 511874 216988 511902 217110
rect 512702 216988 512730 217246
rect 513530 216988 513558 217246
rect 514358 216988 514386 217246
rect 515186 217246 515260 217274
rect 515968 217274 515996 219406
rect 516796 217274 516824 219406
rect 517624 219406 517744 219434
rect 517624 217274 517652 219406
rect 518452 217274 518480 221070
rect 519188 219434 519216 225830
rect 519372 224942 519400 229230
rect 519360 224936 519412 224942
rect 519360 224878 519412 224884
rect 519832 222902 519860 231676
rect 520476 224670 520504 231676
rect 521120 230178 521148 231676
rect 521108 230172 521160 230178
rect 521108 230114 521160 230120
rect 520924 228268 520976 228274
rect 520924 228210 520976 228216
rect 520464 224664 520516 224670
rect 520464 224606 520516 224612
rect 519820 222896 519872 222902
rect 519820 222838 519872 222844
rect 519636 221740 519688 221746
rect 519636 221682 519688 221688
rect 519648 221513 519676 221682
rect 519634 221504 519690 221513
rect 519634 221439 519690 221448
rect 520186 221504 520242 221513
rect 520186 221439 520242 221448
rect 519188 219406 519308 219434
rect 519280 217274 519308 219406
rect 520200 217274 520228 221439
rect 520936 221270 520964 228210
rect 521764 225894 521792 231676
rect 522422 231662 522712 231690
rect 521752 225888 521804 225894
rect 521752 225830 521804 225836
rect 521752 223168 521804 223174
rect 521752 223110 521804 223116
rect 520924 221264 520976 221270
rect 520924 221206 520976 221212
rect 515968 217246 516042 217274
rect 516796 217246 516870 217274
rect 517624 217246 517698 217274
rect 518452 217246 518526 217274
rect 519280 217246 519354 217274
rect 515186 216988 515214 217246
rect 516014 216988 516042 217246
rect 516842 216988 516870 217246
rect 517670 216988 517698 217246
rect 518498 216988 518526 217246
rect 519326 216988 519354 217246
rect 520154 217246 520228 217274
rect 520936 217274 520964 221206
rect 521764 217274 521792 223110
rect 522684 221746 522712 231662
rect 523052 229770 523080 231676
rect 523040 229764 523092 229770
rect 523040 229706 523092 229712
rect 523696 227186 523724 231676
rect 524248 231662 524354 231690
rect 523040 227180 523092 227186
rect 523040 227122 523092 227128
rect 523684 227180 523736 227186
rect 523684 227122 523736 227128
rect 522672 221740 522724 221746
rect 522672 221682 522724 221688
rect 522580 220652 522632 220658
rect 522580 220594 522632 220600
rect 522592 217841 522620 220594
rect 523052 217870 523080 227122
rect 523500 224256 523552 224262
rect 523500 224198 523552 224204
rect 523512 220998 523540 224198
rect 524248 221610 524276 231662
rect 524604 230036 524656 230042
rect 524604 229978 524656 229984
rect 524616 227594 524644 229978
rect 524984 229158 525012 231676
rect 524972 229152 525024 229158
rect 524972 229094 525024 229100
rect 524604 227588 524656 227594
rect 524604 227530 524656 227536
rect 524420 227316 524472 227322
rect 524420 227258 524472 227264
rect 524432 224058 524460 227258
rect 525628 224398 525656 231676
rect 526272 227322 526300 231676
rect 526916 230450 526944 231676
rect 526904 230444 526956 230450
rect 526904 230386 526956 230392
rect 526444 229900 526496 229906
rect 526444 229842 526496 229848
rect 526260 227316 526312 227322
rect 526260 227258 526312 227264
rect 526456 226166 526484 229842
rect 527560 228546 527588 231676
rect 528218 231662 528416 231690
rect 527548 228540 527600 228546
rect 527548 228482 527600 228488
rect 526628 227044 526680 227050
rect 526628 226986 526680 226992
rect 526444 226160 526496 226166
rect 526444 226102 526496 226108
rect 526352 224800 526404 224806
rect 526352 224742 526404 224748
rect 525616 224392 525668 224398
rect 525616 224334 525668 224340
rect 524420 224052 524472 224058
rect 524420 223994 524472 224000
rect 525064 224052 525116 224058
rect 525064 223994 525116 224000
rect 524236 221604 524288 221610
rect 524236 221546 524288 221552
rect 523500 220992 523552 220998
rect 523500 220934 523552 220940
rect 523040 217864 523092 217870
rect 522578 217832 522634 217841
rect 523040 217806 523092 217812
rect 522578 217767 522634 217776
rect 520936 217246 521010 217274
rect 521764 217246 521838 217274
rect 520154 216988 520182 217246
rect 520982 216988 521010 217246
rect 521810 216988 521838 217246
rect 522592 217138 522620 217767
rect 523512 217274 523540 220934
rect 524236 217864 524288 217870
rect 524236 217806 524288 217812
rect 523466 217246 523540 217274
rect 522592 217110 522666 217138
rect 522638 216988 522666 217110
rect 523466 216988 523494 217246
rect 524248 217138 524276 217806
rect 525076 217274 525104 223994
rect 525984 217728 526036 217734
rect 525984 217670 526036 217676
rect 525996 217274 526024 217670
rect 525076 217246 525150 217274
rect 524248 217110 524322 217138
rect 524294 216988 524322 217110
rect 525122 216988 525150 217246
rect 525950 217246 526024 217274
rect 526364 217274 526392 224742
rect 526640 219434 526668 226986
rect 527732 223032 527784 223038
rect 527732 222974 527784 222980
rect 527744 222018 527772 222974
rect 527548 222012 527600 222018
rect 527548 221954 527600 221960
rect 527732 222012 527784 222018
rect 527732 221954 527784 221960
rect 528192 222012 528244 222018
rect 528192 221954 528244 221960
rect 527560 219774 527588 221954
rect 527548 219768 527600 219774
rect 527548 219710 527600 219716
rect 526548 219406 526668 219434
rect 526548 217734 526576 219406
rect 526536 217728 526588 217734
rect 526536 217670 526588 217676
rect 526548 217462 526576 217670
rect 526536 217456 526588 217462
rect 526536 217398 526588 217404
rect 527560 217274 527588 219710
rect 528204 219434 528232 221954
rect 528388 220250 528416 231662
rect 528848 230314 528876 231676
rect 528836 230308 528888 230314
rect 528836 230250 528888 230256
rect 529204 230172 529256 230178
rect 529204 230114 529256 230120
rect 529216 229094 529244 230114
rect 529032 229066 529244 229094
rect 529032 220658 529060 229066
rect 529204 225752 529256 225758
rect 529204 225694 529256 225700
rect 529020 220652 529072 220658
rect 529020 220594 529072 220600
rect 528376 220244 528428 220250
rect 528376 220186 528428 220192
rect 528204 219406 528416 219434
rect 528388 217274 528416 219406
rect 529216 217274 529244 225694
rect 529492 223174 529520 231676
rect 530136 229634 530164 231676
rect 530124 229628 530176 229634
rect 530124 229570 530176 229576
rect 530780 229498 530808 231676
rect 531136 229628 531188 229634
rect 531136 229570 531188 229576
rect 530768 229492 530820 229498
rect 530768 229434 530820 229440
rect 529940 229152 529992 229158
rect 529940 229094 529992 229100
rect 529952 224806 529980 229094
rect 530952 225616 531004 225622
rect 530952 225558 531004 225564
rect 529940 224800 529992 224806
rect 529940 224742 529992 224748
rect 529480 223168 529532 223174
rect 529480 223110 529532 223116
rect 530032 220380 530084 220386
rect 530032 220322 530084 220328
rect 530044 219910 530072 220322
rect 530032 219904 530084 219910
rect 530032 219846 530084 219852
rect 530044 217274 530072 219846
rect 530964 217598 530992 225558
rect 531148 220386 531176 229570
rect 531424 225622 531452 231676
rect 531412 225616 531464 225622
rect 531412 225558 531464 225564
rect 532068 223038 532096 231676
rect 532712 230178 532740 231676
rect 533370 231662 533752 231690
rect 532700 230172 532752 230178
rect 532700 230114 532752 230120
rect 533344 228404 533396 228410
rect 533344 228346 533396 228352
rect 532516 223440 532568 223446
rect 532516 223382 532568 223388
rect 532056 223032 532108 223038
rect 532056 222974 532108 222980
rect 532528 222766 532556 223382
rect 532516 222760 532568 222766
rect 532516 222702 532568 222708
rect 531688 220516 531740 220522
rect 531688 220458 531740 220464
rect 531136 220380 531188 220386
rect 531136 220322 531188 220328
rect 530952 217592 531004 217598
rect 530952 217534 531004 217540
rect 526364 217246 526806 217274
rect 527560 217246 527634 217274
rect 528388 217246 528462 217274
rect 529216 217246 529290 217274
rect 530044 217246 530118 217274
rect 525950 216988 525978 217246
rect 526778 216988 526806 217246
rect 527606 216988 527634 217246
rect 528434 216988 528462 217246
rect 529262 216988 529290 217246
rect 530090 216988 530118 217246
rect 530964 217138 530992 217534
rect 531700 217274 531728 220458
rect 532528 217274 532556 222702
rect 533160 222148 533212 222154
rect 533160 222090 533212 222096
rect 533172 221474 533200 222090
rect 533160 221468 533212 221474
rect 533160 221410 533212 221416
rect 533356 219434 533384 228346
rect 533724 227050 533752 231662
rect 533712 227044 533764 227050
rect 533712 226986 533764 226992
rect 534000 222018 534028 231676
rect 534644 230042 534672 231676
rect 534632 230036 534684 230042
rect 534632 229978 534684 229984
rect 534816 229764 534868 229770
rect 534816 229706 534868 229712
rect 534828 223446 534856 229706
rect 535000 224936 535052 224942
rect 535000 224878 535052 224884
rect 534816 223440 534868 223446
rect 534816 223382 534868 223388
rect 533528 222012 533580 222018
rect 533528 221954 533580 221960
rect 533988 222012 534040 222018
rect 533988 221954 534040 221960
rect 533540 221610 533568 221954
rect 533528 221604 533580 221610
rect 533528 221546 533580 221552
rect 534172 220108 534224 220114
rect 534172 220050 534224 220056
rect 533356 219406 533476 219434
rect 533448 217734 533476 219406
rect 533436 217728 533488 217734
rect 533436 217670 533488 217676
rect 531700 217246 531774 217274
rect 532528 217246 532602 217274
rect 530918 217110 530992 217138
rect 530918 216988 530946 217110
rect 531746 216988 531774 217246
rect 532574 216988 532602 217246
rect 533448 217138 533476 217670
rect 534184 217274 534212 220050
rect 535012 217274 535040 224878
rect 535288 224262 535316 231676
rect 535736 227452 535788 227458
rect 535736 227394 535788 227400
rect 535276 224256 535328 224262
rect 535276 224198 535328 224204
rect 535460 223304 535512 223310
rect 535460 223246 535512 223252
rect 535472 217870 535500 223246
rect 535748 219434 535776 227394
rect 535932 225758 535960 231676
rect 536104 230444 536156 230450
rect 536104 230386 536156 230392
rect 536116 227458 536144 230386
rect 536576 229906 536604 231676
rect 536564 229900 536616 229906
rect 536564 229842 536616 229848
rect 537220 228410 537248 231676
rect 537878 231662 538168 231690
rect 537208 228404 537260 228410
rect 537208 228346 537260 228352
rect 537484 227588 537536 227594
rect 537484 227530 537536 227536
rect 536104 227452 536156 227458
rect 536104 227394 536156 227400
rect 535920 225752 535972 225758
rect 535920 225694 535972 225700
rect 535748 219406 535868 219434
rect 535460 217864 535512 217870
rect 535460 217806 535512 217812
rect 535840 217326 535868 219406
rect 537496 218618 537524 227530
rect 538140 220114 538168 231662
rect 538508 229770 538536 231676
rect 538692 231662 539166 231690
rect 538496 229764 538548 229770
rect 538496 229706 538548 229712
rect 538312 229628 538364 229634
rect 538312 229570 538364 229576
rect 538324 226030 538352 229570
rect 538496 226160 538548 226166
rect 538496 226102 538548 226108
rect 538312 226024 538364 226030
rect 538312 225966 538364 225972
rect 538508 225842 538536 226102
rect 538324 225814 538536 225842
rect 538128 220108 538180 220114
rect 538128 220050 538180 220056
rect 538324 219434 538352 225814
rect 538692 222154 538720 231662
rect 539600 230308 539652 230314
rect 539600 230250 539652 230256
rect 539612 228682 539640 230250
rect 547144 230172 547196 230178
rect 547144 230114 547196 230120
rect 543188 228948 543240 228954
rect 543188 228890 543240 228896
rect 541624 228812 541676 228818
rect 541624 228754 541676 228760
rect 539416 228676 539468 228682
rect 539416 228618 539468 228624
rect 539600 228676 539652 228682
rect 539600 228618 539652 228624
rect 539428 228274 539456 228618
rect 539416 228268 539468 228274
rect 539416 228210 539468 228216
rect 540796 228268 540848 228274
rect 540796 228210 540848 228216
rect 539968 226296 540020 226302
rect 539968 226238 540020 226244
rect 539508 224528 539560 224534
rect 539508 224470 539560 224476
rect 539520 222154 539548 224470
rect 539980 223786 540008 226238
rect 539968 223780 540020 223786
rect 539968 223722 540020 223728
rect 538680 222148 538732 222154
rect 538680 222090 538732 222096
rect 539508 222148 539560 222154
rect 539508 222090 539560 222096
rect 539520 220862 539548 222090
rect 538496 220856 538548 220862
rect 538496 220798 538548 220804
rect 539508 220856 539560 220862
rect 539508 220798 539560 220804
rect 538508 219434 538536 220798
rect 538232 219406 538352 219434
rect 538416 219406 538536 219434
rect 537484 218612 537536 218618
rect 537484 218554 537536 218560
rect 536656 217864 536708 217870
rect 536656 217806 536708 217812
rect 535828 217320 535880 217326
rect 534184 217246 534258 217274
rect 535012 217246 535086 217274
rect 535828 217262 535880 217268
rect 533402 217110 533476 217138
rect 533402 216988 533430 217110
rect 534230 216988 534258 217246
rect 535058 216988 535086 217246
rect 535840 217138 535868 217262
rect 536668 217138 536696 217806
rect 537496 217274 537524 218554
rect 538232 217598 538260 219406
rect 538220 217592 538272 217598
rect 538220 217534 538272 217540
rect 538416 217274 538444 219406
rect 539140 217592 539192 217598
rect 539140 217534 539192 217540
rect 537496 217246 537570 217274
rect 535840 217110 535914 217138
rect 536668 217110 536742 217138
rect 535886 216988 535914 217110
rect 536714 216988 536742 217110
rect 537542 216988 537570 217246
rect 538370 217246 538444 217274
rect 538370 216988 538398 217246
rect 539152 217138 539180 217534
rect 539980 217274 540008 223722
rect 540808 220522 540836 228210
rect 540796 220516 540848 220522
rect 540796 220458 540848 220464
rect 540808 217274 540836 220458
rect 541636 217274 541664 228754
rect 543200 224806 543228 228890
rect 545764 225888 545816 225894
rect 545764 225830 545816 225836
rect 543004 224800 543056 224806
rect 543004 224742 543056 224748
rect 543188 224800 543240 224806
rect 543188 224742 543240 224748
rect 543016 224534 543044 224742
rect 543004 224528 543056 224534
rect 543004 224470 543056 224476
rect 543004 222760 543056 222766
rect 543004 222702 543056 222708
rect 543016 222494 543044 222702
rect 542820 222488 542872 222494
rect 542820 222430 542872 222436
rect 543004 222488 543056 222494
rect 543004 222430 543056 222436
rect 542832 222222 542860 222430
rect 542820 222216 542872 222222
rect 542266 222184 542322 222193
rect 542820 222158 542872 222164
rect 542266 222119 542268 222128
rect 542320 222119 542322 222128
rect 542268 222090 542320 222096
rect 543004 222012 543056 222018
rect 543004 221954 543056 221960
rect 543016 221746 543044 221954
rect 542360 221740 542412 221746
rect 542360 221682 542412 221688
rect 543004 221740 543056 221746
rect 543004 221682 543056 221688
rect 542372 220862 542400 221682
rect 542360 220856 542412 220862
rect 542360 220798 542412 220804
rect 543200 219434 543228 224742
rect 544568 224664 544620 224670
rect 544568 224606 544620 224612
rect 543372 222896 543424 222902
rect 543372 222838 543424 222844
rect 543384 222018 543412 222838
rect 543692 222208 543748 222217
rect 543748 222166 543872 222194
rect 543692 222143 543748 222152
rect 543844 222086 543872 222166
rect 543832 222080 543884 222086
rect 543832 222022 543884 222028
rect 543372 222012 543424 222018
rect 543372 221954 543424 221960
rect 543694 222012 543746 222018
rect 543694 221954 543746 221960
rect 542464 219406 543228 219434
rect 542464 217274 542492 219406
rect 542820 218748 542872 218754
rect 542820 218690 542872 218696
rect 542832 218210 542860 218690
rect 543004 218612 543056 218618
rect 543004 218554 543056 218560
rect 543016 218210 543044 218554
rect 542820 218204 542872 218210
rect 542820 218146 542872 218152
rect 543004 218204 543056 218210
rect 543004 218146 543056 218152
rect 543384 217274 543412 221954
rect 543706 221898 543734 221954
rect 543706 221870 543872 221898
rect 543844 221746 543872 221870
rect 543694 221740 543746 221746
rect 543694 221682 543746 221688
rect 543832 221740 543884 221746
rect 543832 221682 543884 221688
rect 543706 221626 543734 221682
rect 543706 221598 544056 221626
rect 543740 221468 543792 221474
rect 543740 221410 543792 221416
rect 543554 220552 543610 220561
rect 543554 220487 543556 220496
rect 543608 220487 543610 220496
rect 543556 220458 543608 220464
rect 543752 219162 543780 221410
rect 544028 220844 544056 221598
rect 544384 220856 544436 220862
rect 544028 220816 544384 220844
rect 544384 220798 544436 220804
rect 543740 219156 543792 219162
rect 543740 219098 543792 219104
rect 544580 217274 544608 224606
rect 544752 221468 544804 221474
rect 544752 221410 544804 221416
rect 544764 220561 544792 221410
rect 544750 220552 544806 220561
rect 544750 220487 544806 220496
rect 544936 220516 544988 220522
rect 544936 220458 544988 220464
rect 544948 218890 544976 220458
rect 544936 218884 544988 218890
rect 544936 218826 544988 218832
rect 539980 217246 540054 217274
rect 540808 217246 540882 217274
rect 541636 217246 541710 217274
rect 542464 217246 542538 217274
rect 539152 217110 539226 217138
rect 539198 216988 539226 217110
rect 540026 216988 540054 217246
rect 540854 216988 540882 217246
rect 541682 216988 541710 217246
rect 542510 216988 542538 217246
rect 543338 217246 543412 217274
rect 544166 217246 544608 217274
rect 543338 216988 543366 217246
rect 544166 216988 544194 217246
rect 544948 217138 544976 218826
rect 545776 217598 545804 225830
rect 547156 221785 547184 230114
rect 549260 230036 549312 230042
rect 549260 229978 549312 229984
rect 548524 227180 548576 227186
rect 548524 227122 548576 227128
rect 548536 224954 548564 227122
rect 548352 224926 548564 224954
rect 548064 224664 548116 224670
rect 548064 224606 548116 224612
rect 548076 224398 548104 224606
rect 548064 224392 548116 224398
rect 548064 224334 548116 224340
rect 547420 223440 547472 223446
rect 547420 223382 547472 223388
rect 547142 221776 547198 221785
rect 547142 221711 547198 221720
rect 546592 220720 546644 220726
rect 546592 220662 546644 220668
rect 545764 217592 545816 217598
rect 545764 217534 545816 217540
rect 545776 217274 545804 217534
rect 545776 217246 545850 217274
rect 544948 217110 545022 217138
rect 544994 216988 545022 217110
rect 545822 216988 545850 217246
rect 546604 217138 546632 220662
rect 547432 218754 547460 223382
rect 548352 219586 548380 224926
rect 548616 224800 548668 224806
rect 548616 224742 548668 224748
rect 548984 224800 549036 224806
rect 548984 224742 549036 224748
rect 548628 224398 548656 224742
rect 548996 224534 549024 224742
rect 549272 224534 549300 229978
rect 553308 228540 553360 228546
rect 553308 228482 553360 228488
rect 552480 227452 552532 227458
rect 552480 227394 552532 227400
rect 551560 227316 551612 227322
rect 551560 227258 551612 227264
rect 549996 224800 550048 224806
rect 549996 224742 550048 224748
rect 548984 224528 549036 224534
rect 548984 224470 549036 224476
rect 549260 224528 549312 224534
rect 549260 224470 549312 224476
rect 548616 224392 548668 224398
rect 548616 224334 548668 224340
rect 548708 220244 548760 220250
rect 548708 220186 548760 220192
rect 548720 219774 548748 220186
rect 548708 219768 548760 219774
rect 548708 219710 548760 219716
rect 548892 219768 548944 219774
rect 548892 219710 548944 219716
rect 548904 219586 548932 219710
rect 548352 219558 548932 219586
rect 547420 218748 547472 218754
rect 547420 218690 547472 218696
rect 547432 217138 547460 218690
rect 548352 217274 548380 219558
rect 549076 219156 549128 219162
rect 549076 219098 549128 219104
rect 548306 217246 548380 217274
rect 546604 217110 546678 217138
rect 547432 217110 547506 217138
rect 546650 216988 546678 217110
rect 547478 216988 547506 217110
rect 548306 216988 548334 217246
rect 549088 217138 549116 219098
rect 550008 217138 550036 224742
rect 550640 224664 550692 224670
rect 550640 224606 550692 224612
rect 550652 222057 550680 224606
rect 550638 222048 550694 222057
rect 550638 221983 550694 221992
rect 550822 222048 550878 222057
rect 550822 221983 550878 221992
rect 550836 217138 550864 221983
rect 551572 217274 551600 227258
rect 552492 219298 552520 227394
rect 553320 224954 553348 228482
rect 553228 224926 553348 224954
rect 553032 220516 553084 220522
rect 553228 220504 553256 224926
rect 554056 222902 554084 249047
rect 554502 244760 554558 244769
rect 554502 244695 554558 244704
rect 554516 244322 554544 244695
rect 554504 244316 554556 244322
rect 554504 244258 554556 244264
rect 554502 240408 554558 240417
rect 554502 240343 554558 240352
rect 554516 240174 554544 240343
rect 554504 240168 554556 240174
rect 554504 240110 554556 240116
rect 554320 238740 554372 238746
rect 554320 238682 554372 238688
rect 554332 238241 554360 238682
rect 554318 238232 554374 238241
rect 554318 238167 554374 238176
rect 554504 236088 554556 236094
rect 554502 236056 554504 236065
rect 554556 236056 554558 236065
rect 554502 235991 554558 236000
rect 554412 234592 554464 234598
rect 554412 234534 554464 234540
rect 554424 233889 554452 234534
rect 554410 233880 554466 233889
rect 554410 233815 554466 233824
rect 555436 228546 555464 255546
rect 556804 251252 556856 251258
rect 556804 251194 556856 251200
rect 555976 228676 556028 228682
rect 555976 228618 556028 228624
rect 555424 228540 555476 228546
rect 555424 228482 555476 228488
rect 555988 224806 556016 228618
rect 556816 227186 556844 251194
rect 558184 246356 558236 246362
rect 558184 246298 558236 246304
rect 558196 236094 558224 246298
rect 558184 236088 558236 236094
rect 558184 236030 558236 236036
rect 559564 229900 559616 229906
rect 559564 229842 559616 229848
rect 556804 227180 556856 227186
rect 556804 227122 556856 227128
rect 556160 226024 556212 226030
rect 556160 225966 556212 225972
rect 557448 226024 557500 226030
rect 557448 225966 557500 225972
rect 554964 224800 555016 224806
rect 554964 224742 555016 224748
rect 555976 224800 556028 224806
rect 555976 224742 556028 224748
rect 554044 222896 554096 222902
rect 554044 222838 554096 222844
rect 553400 220856 553452 220862
rect 553400 220798 553452 220804
rect 553412 220674 553440 220798
rect 553582 220688 553638 220697
rect 553412 220646 553582 220674
rect 553582 220623 553638 220632
rect 553860 220516 553912 220522
rect 553228 220476 553860 220504
rect 553032 220458 553084 220464
rect 552480 219292 552532 219298
rect 552480 219234 552532 219240
rect 552492 217274 552520 219234
rect 553044 219162 553072 220458
rect 553032 219156 553084 219162
rect 553032 219098 553084 219104
rect 553320 217274 553348 220476
rect 553860 220458 553912 220464
rect 554044 220380 554096 220386
rect 554044 220322 554096 220328
rect 551572 217246 551646 217274
rect 549088 217110 549162 217138
rect 549134 216988 549162 217110
rect 549962 217110 550036 217138
rect 550790 217110 550864 217138
rect 549962 216988 549990 217110
rect 550790 216988 550818 217110
rect 551618 216988 551646 217246
rect 552446 217246 552520 217274
rect 553274 217246 553348 217274
rect 552446 216988 552474 217246
rect 553274 216988 553302 217246
rect 554056 217138 554084 220322
rect 554976 217274 555004 224742
rect 555792 224528 555844 224534
rect 555790 224496 555792 224505
rect 555844 224496 555846 224505
rect 555790 224431 555846 224440
rect 556172 224398 556200 225966
rect 557460 224806 557488 225966
rect 558184 225616 558236 225622
rect 558184 225558 558236 225564
rect 558196 224954 558224 225558
rect 558196 224926 558408 224954
rect 557264 224800 557316 224806
rect 557262 224768 557264 224777
rect 557448 224800 557500 224806
rect 557316 224768 557318 224777
rect 557448 224742 557500 224748
rect 557262 224703 557318 224712
rect 556160 224392 556212 224398
rect 556160 224334 556212 224340
rect 557356 224392 557408 224398
rect 557356 224334 557408 224340
rect 555700 223168 555752 223174
rect 555700 223110 555752 223116
rect 555712 217841 555740 223110
rect 556620 219156 556672 219162
rect 556620 219098 556672 219104
rect 555976 218884 556028 218890
rect 555976 218826 556028 218832
rect 555988 218618 556016 218826
rect 556436 218748 556488 218754
rect 556436 218690 556488 218696
rect 555976 218612 556028 218618
rect 555976 218554 556028 218560
rect 556448 218210 556476 218690
rect 556436 218204 556488 218210
rect 556436 218146 556488 218152
rect 555698 217832 555754 217841
rect 555698 217767 555754 217776
rect 554930 217246 555004 217274
rect 554056 217110 554130 217138
rect 554102 216988 554130 217110
rect 554930 216988 554958 217246
rect 555712 217138 555740 217767
rect 556632 217138 556660 219098
rect 555712 217110 555786 217138
rect 555758 216988 555786 217110
rect 556586 217110 556660 217138
rect 557368 217138 557396 224334
rect 558184 222760 558236 222766
rect 558184 222702 558236 222708
rect 558196 222222 558224 222702
rect 558184 222216 558236 222222
rect 558184 222158 558236 222164
rect 558000 220652 558052 220658
rect 558000 220594 558052 220600
rect 558012 220114 558040 220594
rect 558380 220425 558408 224926
rect 558552 224800 558604 224806
rect 558550 224768 558552 224777
rect 558604 224768 558606 224777
rect 558550 224703 558606 224712
rect 559012 223032 559064 223038
rect 559012 222974 559064 222980
rect 558552 222216 558604 222222
rect 558552 222158 558604 222164
rect 558564 221785 558592 222158
rect 558734 222048 558790 222057
rect 558734 221983 558790 221992
rect 558550 221776 558606 221785
rect 558550 221711 558606 221720
rect 558366 220416 558422 220425
rect 558366 220351 558422 220360
rect 558380 220266 558408 220351
rect 558196 220238 558408 220266
rect 558000 220108 558052 220114
rect 558000 220050 558052 220056
rect 558196 217274 558224 220238
rect 558368 220176 558420 220182
rect 558368 220118 558420 220124
rect 558380 219910 558408 220118
rect 558748 219910 558776 221983
rect 558368 219904 558420 219910
rect 558368 219846 558420 219852
rect 558736 219904 558788 219910
rect 558736 219846 558788 219852
rect 558196 217246 558270 217274
rect 557368 217110 557442 217138
rect 556586 216988 556614 217110
rect 557414 216988 557442 217110
rect 558242 216988 558270 217246
rect 559024 217138 559052 222974
rect 559576 220862 559604 229842
rect 560760 227044 560812 227050
rect 560760 226986 560812 226992
rect 559932 222216 559984 222222
rect 559932 222158 559984 222164
rect 559564 220856 559616 220862
rect 559564 220798 559616 220804
rect 559944 217138 559972 222158
rect 560772 220318 560800 226986
rect 560956 221785 560984 259422
rect 563704 256760 563756 256766
rect 563704 256702 563756 256708
rect 562324 252612 562376 252618
rect 562324 252554 562376 252560
rect 562336 229094 562364 252554
rect 562336 229066 562732 229094
rect 562704 224806 562732 229066
rect 563716 226302 563744 256702
rect 566464 229764 566516 229770
rect 566464 229706 566516 229712
rect 566476 229094 566504 229706
rect 566476 229066 566688 229094
rect 565636 228404 565688 228410
rect 565636 228346 565688 228352
rect 563704 226296 563756 226302
rect 563704 226238 563756 226244
rect 563060 225752 563112 225758
rect 563060 225694 563112 225700
rect 563072 224954 563100 225694
rect 563072 224926 564020 224954
rect 561404 224800 561456 224806
rect 561402 224768 561404 224777
rect 562692 224800 562744 224806
rect 561456 224768 561458 224777
rect 562692 224742 562744 224748
rect 561402 224703 561458 224712
rect 562600 224528 562652 224534
rect 561678 224496 561734 224505
rect 561678 224431 561734 224440
rect 562598 224496 562600 224505
rect 563152 224528 563204 224534
rect 562652 224496 562654 224505
rect 562598 224431 562654 224440
rect 563150 224496 563152 224505
rect 563204 224496 563206 224505
rect 563150 224431 563206 224440
rect 560942 221776 560998 221785
rect 560942 221711 560998 221720
rect 561494 220688 561550 220697
rect 561494 220623 561550 220632
rect 560760 220312 560812 220318
rect 560760 220254 560812 220260
rect 560772 217274 560800 220254
rect 559024 217110 559098 217138
rect 559070 216988 559098 217110
rect 559898 217110 559972 217138
rect 560726 217246 560800 217274
rect 559898 216988 559926 217110
rect 560726 216988 560754 217246
rect 561508 217138 561536 220623
rect 561692 219162 561720 224431
rect 562784 224392 562836 224398
rect 562836 224340 562916 224346
rect 562784 224334 562916 224340
rect 562796 224318 562916 224334
rect 562692 224256 562744 224262
rect 562692 224198 562744 224204
rect 562704 224097 562732 224198
rect 562888 224194 562916 224318
rect 562876 224188 562928 224194
rect 562876 224130 562928 224136
rect 562690 224088 562746 224097
rect 562690 224023 562746 224032
rect 563426 224088 563482 224097
rect 563426 224023 563482 224032
rect 563060 220856 563112 220862
rect 563060 220798 563112 220804
rect 563244 220856 563296 220862
rect 563244 220798 563296 220804
rect 563072 220697 563100 220798
rect 563058 220688 563114 220697
rect 563058 220623 563114 220632
rect 563256 220425 563284 220798
rect 563440 220425 563468 224023
rect 563242 220416 563298 220425
rect 563060 220380 563112 220386
rect 563242 220351 563298 220360
rect 563426 220416 563482 220425
rect 563426 220351 563482 220360
rect 563060 220322 563112 220328
rect 562876 220312 562928 220318
rect 562876 220254 562928 220260
rect 562888 220017 562916 220254
rect 563072 220017 563100 220322
rect 562874 220008 562930 220017
rect 562874 219943 562930 219952
rect 563058 220008 563114 220017
rect 563058 219943 563114 219952
rect 561680 219156 561732 219162
rect 561680 219098 561732 219104
rect 562416 219156 562468 219162
rect 562416 219098 562468 219104
rect 562232 218340 562284 218346
rect 562232 218282 562284 218288
rect 562244 217190 562272 218282
rect 562428 217274 562456 219098
rect 562876 218340 562928 218346
rect 562876 218282 562928 218288
rect 562888 218226 562916 218282
rect 562888 218198 563100 218226
rect 562690 217832 562746 217841
rect 562690 217767 562746 217776
rect 562874 217832 562930 217841
rect 562874 217767 562930 217776
rect 562382 217246 562456 217274
rect 562232 217184 562284 217190
rect 561508 217110 561582 217138
rect 562232 217126 562284 217132
rect 561554 216988 561582 217110
rect 562382 216988 562410 217246
rect 562704 217190 562732 217767
rect 562508 217184 562560 217190
rect 562508 217126 562560 217132
rect 562692 217184 562744 217190
rect 562692 217126 562744 217132
rect 562520 217036 562548 217126
rect 562888 217036 562916 217767
rect 563072 217190 563100 218198
rect 563440 217274 563468 220351
rect 563612 218000 563664 218006
rect 563612 217942 563664 217948
rect 563624 217841 563652 217942
rect 563610 217832 563666 217841
rect 563610 217767 563666 217776
rect 563210 217246 563468 217274
rect 563992 217274 564020 224926
rect 565174 224768 565230 224777
rect 565174 224703 565230 224712
rect 565188 224330 565216 224703
rect 565176 224324 565228 224330
rect 565176 224266 565228 224272
rect 564806 220688 564862 220697
rect 564806 220623 564862 220632
rect 564820 220017 564848 220623
rect 565648 220425 565676 228346
rect 566660 220658 566688 229066
rect 568120 226296 568172 226302
rect 568120 226238 568172 226244
rect 568132 224954 568160 226238
rect 568132 224926 568252 224954
rect 568224 222194 568252 224926
rect 568224 222166 568436 222194
rect 566464 220652 566516 220658
rect 566464 220594 566516 220600
rect 566648 220652 566700 220658
rect 566648 220594 566700 220600
rect 567292 220652 567344 220658
rect 567292 220594 567344 220600
rect 565634 220416 565690 220425
rect 565634 220351 565690 220360
rect 564806 220008 564862 220017
rect 564806 219943 564862 219952
rect 563992 217246 564066 217274
rect 563060 217184 563112 217190
rect 563060 217126 563112 217132
rect 562520 217008 562916 217036
rect 563210 216988 563238 217246
rect 564038 216988 564066 217246
rect 564820 217138 564848 219943
rect 565648 217274 565676 220351
rect 565648 217246 565722 217274
rect 564820 217110 564894 217138
rect 564866 216988 564894 217110
rect 565694 216988 565722 217246
rect 566476 217138 566504 220594
rect 567304 219201 567332 220594
rect 567290 219192 567346 219201
rect 567290 219127 567346 219136
rect 567304 217138 567332 219127
rect 567660 218884 567712 218890
rect 568212 218884 568264 218890
rect 567660 218826 567712 218832
rect 567856 218844 568212 218872
rect 567672 218634 567700 218826
rect 567856 218754 567884 218844
rect 568212 218826 568264 218832
rect 567844 218748 567896 218754
rect 567844 218690 567896 218696
rect 568028 218748 568080 218754
rect 568028 218690 568080 218696
rect 568040 218634 568068 218690
rect 567672 218606 568068 218634
rect 568408 217274 568436 222166
rect 568592 220658 568620 260850
rect 570616 234598 570644 261462
rect 647252 246362 647280 278038
rect 647240 246356 647292 246362
rect 647240 246298 647292 246304
rect 596824 245676 596876 245682
rect 596824 245618 596876 245624
rect 573364 244316 573416 244322
rect 573364 244258 573416 244264
rect 570604 234592 570656 234598
rect 570604 234534 570656 234540
rect 571340 228540 571392 228546
rect 571340 228482 571392 228488
rect 570604 227180 570656 227186
rect 570604 227122 570656 227128
rect 568946 221776 569002 221785
rect 568946 221711 569002 221720
rect 568580 220652 568632 220658
rect 568580 220594 568632 220600
rect 568178 217246 568436 217274
rect 566476 217110 566550 217138
rect 567304 217110 567378 217138
rect 566522 216988 566550 217110
rect 567350 216988 567378 217110
rect 568178 216988 568206 217246
rect 568960 217138 568988 221711
rect 569958 220688 570014 220697
rect 569776 220652 569828 220658
rect 569958 220623 569960 220632
rect 569776 220594 569828 220600
rect 570012 220623 570014 220632
rect 569960 220594 570012 220600
rect 569788 217138 569816 220594
rect 570616 217274 570644 227122
rect 571352 224954 571380 228482
rect 571352 224926 571932 224954
rect 571708 224800 571760 224806
rect 571708 224742 571760 224748
rect 571522 219192 571578 219201
rect 571340 219156 571392 219162
rect 571522 219127 571524 219136
rect 571340 219098 571392 219104
rect 571576 219127 571578 219136
rect 571524 219098 571576 219104
rect 570972 218748 571024 218754
rect 570972 218690 571024 218696
rect 570984 217841 571012 218690
rect 571352 217841 571380 219098
rect 570970 217832 571026 217841
rect 570970 217767 571026 217776
rect 571338 217832 571394 217841
rect 571338 217767 571394 217776
rect 571720 217274 571748 224742
rect 570616 217246 570690 217274
rect 568960 217110 569034 217138
rect 569788 217110 569862 217138
rect 569006 216988 569034 217110
rect 569834 216988 569862 217110
rect 570662 216988 570690 217246
rect 571490 217246 571748 217274
rect 571904 217274 571932 224926
rect 573376 220697 573404 244258
rect 576124 242208 576176 242214
rect 576124 242150 576176 242156
rect 576136 238746 576164 242150
rect 577504 240168 577556 240174
rect 577504 240110 577556 240116
rect 576124 238740 576176 238746
rect 576124 238682 576176 238688
rect 573362 220688 573418 220697
rect 573362 220623 573418 220632
rect 576582 220416 576638 220425
rect 576638 220374 576808 220402
rect 576582 220351 576638 220360
rect 576780 220250 576808 220374
rect 576768 220244 576820 220250
rect 576768 220186 576820 220192
rect 576584 220176 576636 220182
rect 576584 220118 576636 220124
rect 576596 220017 576624 220118
rect 576780 220102 577176 220130
rect 576780 220046 576808 220102
rect 576768 220040 576820 220046
rect 572534 220008 572590 220017
rect 572534 219943 572590 219952
rect 576582 220008 576638 220017
rect 576768 219982 576820 219988
rect 576952 220040 577004 220046
rect 576952 219982 577004 219988
rect 576582 219943 576638 219952
rect 572076 219020 572128 219026
rect 572076 218962 572128 218968
rect 572088 218906 572116 218962
rect 572088 218878 572208 218906
rect 572180 218226 572208 218878
rect 572548 218754 572576 219943
rect 576768 219632 576820 219638
rect 576964 219586 576992 219982
rect 576820 219580 576992 219586
rect 576768 219574 576992 219580
rect 576780 219558 576992 219574
rect 577148 219452 577176 220102
rect 577136 219446 577188 219452
rect 577136 219388 577188 219394
rect 574744 219292 574796 219298
rect 574744 219234 574796 219240
rect 572536 218748 572588 218754
rect 572536 218690 572588 218696
rect 572180 218210 572714 218226
rect 572180 218204 572726 218210
rect 572180 218198 572674 218204
rect 572674 218146 572726 218152
rect 572444 218136 572496 218142
rect 572496 218084 572668 218090
rect 572444 218078 572668 218084
rect 572456 218074 572668 218078
rect 572456 218068 572680 218074
rect 572456 218062 572628 218068
rect 572628 218010 572680 218016
rect 572444 218000 572496 218006
rect 572444 217942 572496 217948
rect 572456 217841 572484 217942
rect 572442 217832 572498 217841
rect 572442 217767 572498 217776
rect 574098 217832 574154 217841
rect 574098 217767 574154 217776
rect 574558 217832 574614 217841
rect 574558 217767 574614 217776
rect 571904 217246 572346 217274
rect 571490 216988 571518 217246
rect 572318 216988 572346 217246
rect 574112 216918 574140 217767
rect 574100 216912 574152 216918
rect 574100 216854 574152 216860
rect 574098 216744 574154 216753
rect 574098 216679 574154 216688
rect 574374 216744 574430 216753
rect 574374 216679 574430 216688
rect 574112 213518 574140 216679
rect 574100 213512 574152 213518
rect 574100 213454 574152 213460
rect 574388 213382 574416 216679
rect 574376 213376 574428 213382
rect 574376 213318 574428 213324
rect 574572 213246 574600 217767
rect 574756 214606 574784 219234
rect 575480 219020 575532 219026
rect 575480 218962 575532 218968
rect 574926 216472 574982 216481
rect 574926 216407 574982 216416
rect 574940 214742 574968 216407
rect 575492 214878 575520 218962
rect 575480 214872 575532 214878
rect 575480 214814 575532 214820
rect 574928 214736 574980 214742
rect 574928 214678 574980 214684
rect 574744 214600 574796 214606
rect 574744 214542 574796 214548
rect 574560 213240 574612 213246
rect 574560 213182 574612 213188
rect 577516 99142 577544 240110
rect 596836 231538 596864 245618
rect 648632 242214 648660 278052
rect 648620 242208 648672 242214
rect 648620 242150 648672 242156
rect 629944 241528 629996 241534
rect 629944 241470 629996 241476
rect 596824 231532 596876 231538
rect 596824 231474 596876 231480
rect 629956 229094 629984 241470
rect 633624 231532 633676 231538
rect 633624 231474 633676 231480
rect 629956 229066 630076 229094
rect 621020 224936 621072 224942
rect 621020 224878 621072 224884
rect 610440 224188 610492 224194
rect 610440 224130 610492 224136
rect 610624 224188 610676 224194
rect 610624 224130 610676 224136
rect 617064 224188 617116 224194
rect 617064 224130 617116 224136
rect 610452 223802 610480 224130
rect 610636 223922 610664 224130
rect 610624 223916 610676 223922
rect 610624 223858 610676 223864
rect 610808 223916 610860 223922
rect 610808 223858 610860 223864
rect 610820 223802 610848 223858
rect 610452 223774 610848 223802
rect 614948 223644 615000 223650
rect 614948 223586 615000 223592
rect 593972 222624 594024 222630
rect 593972 222566 594024 222572
rect 582470 220280 582526 220289
rect 582470 220215 582526 220224
rect 582484 220114 582512 220215
rect 582472 220108 582524 220114
rect 582472 220050 582524 220056
rect 581644 220040 581696 220046
rect 581828 220040 581880 220046
rect 581644 219982 581696 219988
rect 581826 220008 581828 220017
rect 582334 220040 582386 220046
rect 581880 220008 581882 220017
rect 581656 219638 581684 219982
rect 582654 220008 582710 220017
rect 582386 219988 582654 219994
rect 582334 219982 582654 219988
rect 582346 219966 582654 219982
rect 581826 219943 581882 219952
rect 582654 219943 582710 219952
rect 591946 220008 592002 220017
rect 591946 219943 592002 219952
rect 581644 219632 581696 219638
rect 581644 219574 581696 219580
rect 582380 219632 582432 219638
rect 582656 219632 582708 219638
rect 582432 219580 582512 219586
rect 582380 219574 582512 219580
rect 582656 219574 582708 219580
rect 582392 219558 582512 219574
rect 582484 219230 582512 219558
rect 582668 219366 582696 219574
rect 591960 219502 591988 219943
rect 591948 219496 592000 219502
rect 591948 219438 592000 219444
rect 582656 219360 582708 219366
rect 582656 219302 582708 219308
rect 582472 219224 582524 219230
rect 582472 219166 582524 219172
rect 578882 214024 578938 214033
rect 578882 213959 578938 213968
rect 578330 211712 578386 211721
rect 578330 211647 578386 211656
rect 578344 211206 578372 211647
rect 578332 211200 578384 211206
rect 578332 211142 578384 211148
rect 578896 208350 578924 213959
rect 580908 211200 580960 211206
rect 580908 211142 580960 211148
rect 579528 209840 579580 209846
rect 579526 209808 579528 209817
rect 579580 209808 579582 209817
rect 579526 209743 579582 209752
rect 578884 208344 578936 208350
rect 578884 208286 578936 208292
rect 579526 207496 579582 207505
rect 579582 207454 579752 207482
rect 579526 207431 579582 207440
rect 579526 205864 579582 205873
rect 579526 205799 579528 205808
rect 579580 205799 579582 205808
rect 579528 205770 579580 205776
rect 579724 204270 579752 207454
rect 580920 206922 580948 211142
rect 593984 210202 594012 222566
rect 605012 222080 605064 222086
rect 605012 222022 605064 222028
rect 600320 221876 600372 221882
rect 600320 221818 600372 221824
rect 599490 221232 599546 221241
rect 599490 221167 599546 221176
rect 596824 219360 596876 219366
rect 596824 219302 596876 219308
rect 594798 218648 594854 218657
rect 594798 218583 594854 218592
rect 594812 216782 594840 218583
rect 595166 217560 595222 217569
rect 595166 217495 595222 217504
rect 594800 216776 594852 216782
rect 594800 216718 594852 216724
rect 594800 213512 594852 213518
rect 594800 213454 594852 213460
rect 594812 210202 594840 213454
rect 595180 210202 595208 217495
rect 596362 217288 596418 217297
rect 596362 217223 596418 217232
rect 595718 217016 595774 217025
rect 595718 216951 595774 216960
rect 595732 210202 595760 216951
rect 596376 210202 596404 217223
rect 596836 210202 596864 219302
rect 597928 219224 597980 219230
rect 597928 219166 597980 219172
rect 597560 216912 597612 216918
rect 597560 216854 597612 216860
rect 597572 210202 597600 216854
rect 597940 210202 597968 219166
rect 598848 218612 598900 218618
rect 598848 218554 598900 218560
rect 598296 217864 598348 217870
rect 598296 217806 598348 217812
rect 598308 216918 598336 217806
rect 598664 217728 598716 217734
rect 598664 217670 598716 217676
rect 598676 217326 598704 217670
rect 598860 217326 598888 218554
rect 598664 217320 598716 217326
rect 598664 217262 598716 217268
rect 598848 217320 598900 217326
rect 598848 217262 598900 217268
rect 599032 217184 599084 217190
rect 599032 217126 599084 217132
rect 598296 216912 598348 216918
rect 598296 216854 598348 216860
rect 598478 215928 598534 215937
rect 598478 215863 598534 215872
rect 598492 210202 598520 215863
rect 599044 210202 599072 217126
rect 599504 210202 599532 221167
rect 600134 220144 600190 220153
rect 600134 220079 600190 220088
rect 600148 219502 600176 220079
rect 600136 219496 600188 219502
rect 600136 219438 600188 219444
rect 600136 217184 600188 217190
rect 600136 217126 600188 217132
rect 600148 216918 600176 217126
rect 600136 216912 600188 216918
rect 600136 216854 600188 216860
rect 600332 210202 600360 221818
rect 601148 221740 601200 221746
rect 601148 221682 601200 221688
rect 600688 221604 600740 221610
rect 600688 221546 600740 221552
rect 600700 221338 600728 221546
rect 601160 221474 601188 221682
rect 601148 221468 601200 221474
rect 601148 221410 601200 221416
rect 600688 221332 600740 221338
rect 600688 221274 600740 221280
rect 603172 221332 603224 221338
rect 603172 221274 603224 221280
rect 600504 221264 600556 221270
rect 600504 221206 600556 221212
rect 600516 214470 600544 221206
rect 600688 221128 600740 221134
rect 600688 221070 600740 221076
rect 600504 214464 600556 214470
rect 600504 214406 600556 214412
rect 600700 210202 600728 221070
rect 601700 220992 601752 220998
rect 601700 220934 601752 220940
rect 601146 220144 601202 220153
rect 601146 220079 601202 220088
rect 601160 219910 601188 220079
rect 600964 219904 601016 219910
rect 600964 219846 601016 219852
rect 601148 219904 601200 219910
rect 601148 219846 601200 219852
rect 600976 219502 601004 219846
rect 601516 219768 601568 219774
rect 601160 219716 601516 219722
rect 601160 219710 601568 219716
rect 601160 219694 601556 219710
rect 601160 219638 601188 219694
rect 601148 219632 601200 219638
rect 601148 219574 601200 219580
rect 600964 219496 601016 219502
rect 600964 219438 601016 219444
rect 601148 217320 601200 217326
rect 601148 217262 601200 217268
rect 601160 216782 601188 217262
rect 601148 216776 601200 216782
rect 601148 216718 601200 216724
rect 601240 214464 601292 214470
rect 601240 214406 601292 214412
rect 601252 210202 601280 214406
rect 601712 210202 601740 220934
rect 601884 218748 601936 218754
rect 601884 218690 601936 218696
rect 601896 217462 601924 218690
rect 602988 217864 603040 217870
rect 602988 217806 603040 217812
rect 601884 217456 601936 217462
rect 601884 217398 601936 217404
rect 603000 217326 603028 217806
rect 602344 217320 602396 217326
rect 602344 217262 602396 217268
rect 602988 217320 603040 217326
rect 602988 217262 603040 217268
rect 602356 210202 602384 217262
rect 603184 210202 603212 221274
rect 603354 218376 603410 218385
rect 603354 218311 603410 218320
rect 603368 217870 603396 218311
rect 604644 218068 604696 218074
rect 604644 218010 604696 218016
rect 603356 217864 603408 217870
rect 603356 217806 603408 217812
rect 604656 217734 604684 218010
rect 604276 217728 604328 217734
rect 604644 217728 604696 217734
rect 604328 217676 604500 217682
rect 604276 217670 604500 217676
rect 604644 217670 604696 217676
rect 604288 217654 604500 217670
rect 603448 217320 603500 217326
rect 603448 217262 603500 217268
rect 603460 210202 603488 217262
rect 604000 217184 604052 217190
rect 604000 217126 604052 217132
rect 604012 210202 604040 217126
rect 604472 210202 604500 217654
rect 605024 210202 605052 222022
rect 606116 221604 606168 221610
rect 606116 221546 606168 221552
rect 605932 221468 605984 221474
rect 605932 221410 605984 221416
rect 605944 214470 605972 221410
rect 605932 214464 605984 214470
rect 605932 214406 605984 214412
rect 606128 210202 606156 221546
rect 609428 220856 609480 220862
rect 609428 220798 609480 220804
rect 608600 220516 608652 220522
rect 608600 220458 608652 220464
rect 607496 219632 607548 219638
rect 607496 219574 607548 219580
rect 607312 219496 607364 219502
rect 607312 219438 607364 219444
rect 606760 217592 606812 217598
rect 606760 217534 606812 217540
rect 606300 214464 606352 214470
rect 606300 214406 606352 214412
rect 593984 210174 594412 210202
rect 594812 210174 594964 210202
rect 595180 210174 595516 210202
rect 595732 210174 596068 210202
rect 596376 210174 596620 210202
rect 596836 210174 597172 210202
rect 597572 210174 597724 210202
rect 597940 210174 598276 210202
rect 598492 210174 598828 210202
rect 599044 210174 599380 210202
rect 599504 210174 599932 210202
rect 600332 210174 600484 210202
rect 600700 210174 601036 210202
rect 601252 210174 601588 210202
rect 601712 210174 602140 210202
rect 602356 210174 602692 210202
rect 603184 210174 603244 210202
rect 603460 210174 603796 210202
rect 604012 210174 604348 210202
rect 604472 210174 604900 210202
rect 605024 210174 605452 210202
rect 606004 210174 606156 210202
rect 606312 210202 606340 214406
rect 606772 210202 606800 217534
rect 607324 214470 607352 219438
rect 607312 214464 607364 214470
rect 607312 214406 607364 214412
rect 607508 210202 607536 219574
rect 607864 214464 607916 214470
rect 607864 214406 607916 214412
rect 607876 210202 607904 214406
rect 608612 210202 608640 220458
rect 608968 217048 609020 217054
rect 608968 216990 609020 216996
rect 608980 210202 609008 216990
rect 609440 210202 609468 220798
rect 610532 220652 610584 220658
rect 610532 220594 610584 220600
rect 610072 220380 610124 220386
rect 610072 220322 610124 220328
rect 609888 218476 609940 218482
rect 609888 218418 609940 218424
rect 609900 217054 609928 218418
rect 609888 217048 609940 217054
rect 609888 216990 609940 216996
rect 610084 210202 610112 220322
rect 610544 210202 610572 220594
rect 611636 220244 611688 220250
rect 611636 220186 611688 220192
rect 611450 219736 611506 219745
rect 611450 219671 611506 219680
rect 611464 214470 611492 219671
rect 611452 214464 611504 214470
rect 611452 214406 611504 214412
rect 611648 210202 611676 220186
rect 614488 218340 614540 218346
rect 614488 218282 614540 218288
rect 613384 217864 613436 217870
rect 613384 217806 613436 217812
rect 612280 216912 612332 216918
rect 612280 216854 612332 216860
rect 611820 214464 611872 214470
rect 611820 214406 611872 214412
rect 606312 210174 606556 210202
rect 606772 210174 607108 210202
rect 607508 210174 607660 210202
rect 607876 210174 608212 210202
rect 608612 210174 608764 210202
rect 608980 210174 609316 210202
rect 609440 210174 609868 210202
rect 610084 210174 610420 210202
rect 610544 210174 610972 210202
rect 611524 210174 611676 210202
rect 611832 210202 611860 214406
rect 612292 210202 612320 216854
rect 612832 213376 612884 213382
rect 612832 213318 612884 213324
rect 612844 210202 612872 213318
rect 613396 210202 613424 217806
rect 614120 217048 614172 217054
rect 614120 216990 614172 216996
rect 614132 210202 614160 216990
rect 614500 210202 614528 218282
rect 614960 210202 614988 223586
rect 615684 218204 615736 218210
rect 615684 218146 615736 218152
rect 615696 210202 615724 218146
rect 616880 217728 616932 217734
rect 616880 217670 616932 217676
rect 616696 214736 616748 214742
rect 616696 214678 616748 214684
rect 616708 214470 616736 214678
rect 616696 214464 616748 214470
rect 616696 214406 616748 214412
rect 616144 213240 616196 213246
rect 616144 213182 616196 213188
rect 616156 210202 616184 213182
rect 616892 210202 616920 217670
rect 617076 214742 617104 224130
rect 619640 224052 619692 224058
rect 619640 223994 619692 224000
rect 618258 221504 618314 221513
rect 618258 221439 618314 221448
rect 617246 219464 617302 219473
rect 617246 219399 617302 219408
rect 617064 214736 617116 214742
rect 617064 214678 617116 214684
rect 617260 210202 617288 219399
rect 617800 214736 617852 214742
rect 617800 214678 617852 214684
rect 617812 210202 617840 214678
rect 618272 210202 618300 221439
rect 618902 215384 618958 215393
rect 618902 215319 618958 215328
rect 618916 210202 618944 215319
rect 619652 210202 619680 223994
rect 619824 219904 619876 219910
rect 619824 219846 619876 219852
rect 619836 214742 619864 219846
rect 620008 219768 620060 219774
rect 620008 219710 620060 219716
rect 619824 214736 619876 214742
rect 619824 214678 619876 214684
rect 620020 210202 620048 219710
rect 621032 214742 621060 224878
rect 626540 224664 626592 224670
rect 626540 224606 626592 224612
rect 625252 224528 625304 224534
rect 625252 224470 625304 224476
rect 622492 223916 622544 223922
rect 622492 223858 622544 223864
rect 621204 222488 621256 222494
rect 621204 222430 621256 222436
rect 620560 214736 620612 214742
rect 620560 214678 620612 214684
rect 621020 214736 621072 214742
rect 621020 214678 621072 214684
rect 620572 210202 620600 214678
rect 621216 210202 621244 222430
rect 622308 214872 622360 214878
rect 622308 214814 622360 214820
rect 621664 214736 621716 214742
rect 621664 214678 621716 214684
rect 621676 210202 621704 214678
rect 622320 214554 622348 214814
rect 622504 214742 622532 223858
rect 622676 223780 622728 223786
rect 622676 223722 622728 223728
rect 622492 214736 622544 214742
rect 622492 214678 622544 214684
rect 622320 214526 622532 214554
rect 622504 210202 622532 214526
rect 622688 210202 622716 223722
rect 623872 216776 623924 216782
rect 623872 216718 623924 216724
rect 623320 214736 623372 214742
rect 623320 214678 623372 214684
rect 623332 210202 623360 214678
rect 623884 210202 623912 216718
rect 624424 214464 624476 214470
rect 624424 214406 624476 214412
rect 624436 210202 624464 214406
rect 625264 210202 625292 224470
rect 625988 224392 626040 224398
rect 625988 224334 626040 224340
rect 625528 214600 625580 214606
rect 625528 214542 625580 214548
rect 625540 210202 625568 214542
rect 626000 210202 626028 224334
rect 626356 218884 626408 218890
rect 626356 218826 626408 218832
rect 626368 214334 626396 218826
rect 626356 214328 626408 214334
rect 626356 214270 626408 214276
rect 626552 210202 626580 224606
rect 629852 222352 629904 222358
rect 629852 222294 629904 222300
rect 627092 222216 627144 222222
rect 627092 222158 627144 222164
rect 627104 210202 627132 222158
rect 627458 218104 627514 218113
rect 627458 218039 627514 218048
rect 627472 213994 627500 218039
rect 628288 217456 628340 217462
rect 628288 217398 628340 217404
rect 627918 216200 627974 216209
rect 627918 216135 627974 216144
rect 627460 213988 627512 213994
rect 627460 213930 627512 213936
rect 627932 210202 627960 216135
rect 628300 210202 628328 217398
rect 628840 214328 628892 214334
rect 628840 214270 628892 214276
rect 628852 210202 628880 214270
rect 629392 213988 629444 213994
rect 629392 213930 629444 213936
rect 629404 210202 629432 213930
rect 629864 210202 629892 222294
rect 630048 214742 630076 229066
rect 632704 222896 632756 222902
rect 632704 222838 632756 222844
rect 630680 222624 630732 222630
rect 630680 222566 630732 222572
rect 630036 214736 630088 214742
rect 630036 214678 630088 214684
rect 630692 212430 630720 222566
rect 631322 220960 631378 220969
rect 631322 220895 631378 220904
rect 631138 218376 631194 218385
rect 631138 218311 631194 218320
rect 630680 212424 630732 212430
rect 630680 212366 630732 212372
rect 631152 210202 631180 218311
rect 611832 210174 612076 210202
rect 612292 210174 612628 210202
rect 612844 210174 613180 210202
rect 613396 210174 613732 210202
rect 614132 210174 614284 210202
rect 614500 210174 614836 210202
rect 614960 210174 615388 210202
rect 615696 210174 615940 210202
rect 616156 210174 616492 210202
rect 616892 210174 617044 210202
rect 617260 210174 617596 210202
rect 617812 210174 618148 210202
rect 618272 210174 618700 210202
rect 618916 210174 619252 210202
rect 619652 210174 619804 210202
rect 620020 210174 620356 210202
rect 620572 210174 620908 210202
rect 621216 210174 621460 210202
rect 621676 210174 622012 210202
rect 622504 210174 622564 210202
rect 622688 210174 623116 210202
rect 623332 210174 623668 210202
rect 623884 210174 624220 210202
rect 624436 210174 624772 210202
rect 625264 210174 625324 210202
rect 625540 210174 625876 210202
rect 626000 210174 626428 210202
rect 626552 210174 626980 210202
rect 627104 210174 627532 210202
rect 627932 210174 628084 210202
rect 628300 210174 628636 210202
rect 628852 210174 629188 210202
rect 629404 210174 629740 210202
rect 629864 210174 630292 210202
rect 630844 210174 631180 210202
rect 631336 210202 631364 220895
rect 632716 212566 632744 222838
rect 633440 220108 633492 220114
rect 633440 220050 633492 220056
rect 633452 219434 633480 220050
rect 633452 219406 633572 219434
rect 632888 214736 632940 214742
rect 632888 214678 632940 214684
rect 632704 212560 632756 212566
rect 632704 212502 632756 212508
rect 631600 212424 631652 212430
rect 631600 212366 631652 212372
rect 631612 210202 631640 212366
rect 632900 210202 632928 214678
rect 633544 212534 633572 219406
rect 633452 212506 633572 212534
rect 633452 211070 633480 212506
rect 633440 211064 633492 211070
rect 633440 211006 633492 211012
rect 633636 210746 633664 231474
rect 652036 227050 652064 287127
rect 652220 232558 652248 291479
rect 652404 233918 652432 292703
rect 663064 289876 663116 289882
rect 663064 289818 663116 289824
rect 652574 280392 652630 280401
rect 652574 280327 652630 280336
rect 652392 233912 652444 233918
rect 652392 233854 652444 233860
rect 652208 232552 652260 232558
rect 652208 232494 652260 232500
rect 652588 228585 652616 280327
rect 663076 232694 663104 289818
rect 664456 248305 664484 293966
rect 665836 268569 665864 296686
rect 667216 278186 667244 570522
rect 667400 535838 667428 597518
rect 667676 570586 667704 639775
rect 667664 570580 667716 570586
rect 667664 570522 667716 570528
rect 667676 570246 667704 570522
rect 667664 570240 667716 570246
rect 667664 570182 667716 570188
rect 667570 553888 667626 553897
rect 667570 553823 667626 553832
rect 667388 535832 667440 535838
rect 667388 535774 667440 535780
rect 667584 481846 667612 553823
rect 667572 481840 667624 481846
rect 667572 481782 667624 481788
rect 667860 456618 667888 703802
rect 668044 671158 668072 733382
rect 668412 705566 668440 774959
rect 669228 741124 669280 741130
rect 669228 741066 669280 741072
rect 668676 733916 668728 733922
rect 668676 733858 668728 733864
rect 668400 705560 668452 705566
rect 668400 705502 668452 705508
rect 668398 696960 668454 696969
rect 668398 696895 668454 696904
rect 668216 685976 668268 685982
rect 668216 685918 668268 685924
rect 668032 671152 668084 671158
rect 668032 671094 668084 671100
rect 668228 619750 668256 685918
rect 668216 619744 668268 619750
rect 668216 619686 668268 619692
rect 668412 618322 668440 696895
rect 668688 662794 668716 733858
rect 668950 730144 669006 730153
rect 668950 730079 669006 730088
rect 668676 662788 668728 662794
rect 668676 662730 668728 662736
rect 668964 660142 668992 730079
rect 669240 663814 669268 741066
rect 669594 735720 669650 735729
rect 669594 735655 669650 735664
rect 669410 688392 669466 688401
rect 669410 688327 669466 688336
rect 669228 663808 669280 663814
rect 669228 663750 669280 663756
rect 669228 661156 669280 661162
rect 669228 661098 669280 661104
rect 668952 660136 669004 660142
rect 668952 660078 669004 660084
rect 668584 640348 668636 640354
rect 668584 640290 668636 640296
rect 668400 618316 668452 618322
rect 668400 618258 668452 618264
rect 668596 580310 668624 640290
rect 668950 600944 669006 600953
rect 668950 600879 669006 600888
rect 668766 594824 668822 594833
rect 668766 594759 668822 594768
rect 668584 580304 668636 580310
rect 668584 580246 668636 580252
rect 668398 554704 668454 554713
rect 668398 554639 668454 554648
rect 668412 481982 668440 554639
rect 668780 524414 668808 594759
rect 668964 529990 668992 600879
rect 668952 529984 669004 529990
rect 668952 529926 669004 529932
rect 668768 524408 668820 524414
rect 668768 524350 668820 524356
rect 668780 520946 668808 524350
rect 668768 520940 668820 520946
rect 668768 520882 668820 520888
rect 668400 481976 668452 481982
rect 668400 481918 668452 481924
rect 667848 456612 667900 456618
rect 667848 456554 667900 456560
rect 669240 455666 669268 661098
rect 669424 616758 669452 688327
rect 669608 665242 669636 735655
rect 669792 711686 669820 775775
rect 669964 775600 670016 775606
rect 669964 775542 670016 775548
rect 669976 715766 670004 775542
rect 670330 728784 670386 728793
rect 670330 728719 670386 728728
rect 669964 715760 670016 715766
rect 669964 715702 670016 715708
rect 670148 714876 670200 714882
rect 670148 714818 670200 714824
rect 669780 711680 669832 711686
rect 669780 711622 669832 711628
rect 669964 687268 670016 687274
rect 669964 687210 670016 687216
rect 669780 668704 669832 668710
rect 669780 668646 669832 668652
rect 669596 665236 669648 665242
rect 669596 665178 669648 665184
rect 669792 624646 669820 668646
rect 669976 625258 670004 687210
rect 670160 670206 670188 714818
rect 670148 670200 670200 670206
rect 670148 670142 670200 670148
rect 670148 669724 670200 669730
rect 670148 669666 670200 669672
rect 670160 649994 670188 669666
rect 670344 664358 670372 728719
rect 670620 709646 670648 789346
rect 670792 775600 670844 775606
rect 670792 775542 670844 775548
rect 670804 710054 670832 775542
rect 670988 713726 671016 892842
rect 671804 885692 671856 885698
rect 671804 885634 671856 885640
rect 671344 744048 671396 744054
rect 671344 743990 671396 743996
rect 671160 743232 671212 743238
rect 671160 743174 671212 743180
rect 670976 713720 671028 713726
rect 670976 713662 671028 713668
rect 670792 710048 670844 710054
rect 670792 709990 670844 709996
rect 670608 709640 670660 709646
rect 670608 709582 670660 709588
rect 670606 696144 670662 696153
rect 670606 696079 670662 696088
rect 670332 664352 670384 664358
rect 670332 664294 670384 664300
rect 670160 649966 670280 649994
rect 669964 625252 670016 625258
rect 669964 625194 670016 625200
rect 670252 625122 670280 649966
rect 670422 638752 670478 638761
rect 670422 638687 670478 638696
rect 670240 625116 670292 625122
rect 670240 625058 670292 625064
rect 669780 624640 669832 624646
rect 669780 624582 669832 624588
rect 669872 624300 669924 624306
rect 669872 624242 669924 624248
rect 669412 616752 669464 616758
rect 669412 616694 669464 616700
rect 669884 579902 669912 624242
rect 670240 623892 670292 623898
rect 670240 623834 670292 623840
rect 670056 623076 670108 623082
rect 670056 623018 670108 623024
rect 669872 579896 669924 579902
rect 669872 579838 669924 579844
rect 669596 579420 669648 579426
rect 669596 579362 669648 579368
rect 669412 577788 669464 577794
rect 669412 577730 669464 577736
rect 669424 533390 669452 577730
rect 669608 535022 669636 579362
rect 670068 578202 670096 623018
rect 670252 579086 670280 623834
rect 670240 579080 670292 579086
rect 670240 579022 670292 579028
rect 670240 578604 670292 578610
rect 670240 578546 670292 578552
rect 670056 578196 670108 578202
rect 670056 578138 670108 578144
rect 669780 569628 669832 569634
rect 669780 569570 669832 569576
rect 669596 535016 669648 535022
rect 669596 534958 669648 534964
rect 669412 533384 669464 533390
rect 669412 533326 669464 533332
rect 669228 455660 669280 455666
rect 669228 455602 669280 455608
rect 669792 455433 669820 569570
rect 669964 550656 670016 550662
rect 669964 550598 670016 550604
rect 669976 491502 670004 550598
rect 670252 534342 670280 578546
rect 670436 574598 670464 638687
rect 670620 620838 670648 696079
rect 670974 689208 671030 689217
rect 670974 689143 671030 689152
rect 670608 620832 670660 620838
rect 670608 620774 670660 620780
rect 670988 618118 671016 689143
rect 671172 665718 671200 743174
rect 671356 731338 671384 743990
rect 671618 733816 671674 733825
rect 671618 733751 671674 733760
rect 671344 731332 671396 731338
rect 671344 731274 671396 731280
rect 671344 713244 671396 713250
rect 671344 713186 671396 713192
rect 671356 668302 671384 713186
rect 671344 668296 671396 668302
rect 671344 668238 671396 668244
rect 671436 667956 671488 667962
rect 671436 667898 671488 667904
rect 671160 665712 671212 665718
rect 671160 665654 671212 665660
rect 671252 665372 671304 665378
rect 671252 665314 671304 665320
rect 671264 663794 671292 665314
rect 671264 663766 671384 663794
rect 671356 630674 671384 663766
rect 671264 630646 671384 630674
rect 671264 622878 671292 630646
rect 671448 623694 671476 667898
rect 671632 661570 671660 733751
rect 671816 728346 671844 885634
rect 671804 728340 671856 728346
rect 671804 728282 671856 728288
rect 671804 714060 671856 714066
rect 671804 714002 671856 714008
rect 671816 669390 671844 714002
rect 672000 712910 672028 892978
rect 672184 716174 672212 894406
rect 672736 866658 672764 895630
rect 675850 895520 675906 895529
rect 675850 895455 675906 895464
rect 675864 894470 675892 895455
rect 676034 894704 676090 894713
rect 676034 894639 676090 894648
rect 675852 894464 675904 894470
rect 675852 894406 675904 894412
rect 676048 894334 676076 894639
rect 673368 894328 673420 894334
rect 673368 894270 673420 894276
rect 676036 894328 676088 894334
rect 676036 894270 676088 894276
rect 673184 886916 673236 886922
rect 673184 886858 673236 886864
rect 672724 866652 672776 866658
rect 672724 866594 672776 866600
rect 672998 778832 673054 778841
rect 672998 778767 673054 778776
rect 672356 742824 672408 742830
rect 672356 742766 672408 742772
rect 672172 716168 672224 716174
rect 672172 716110 672224 716116
rect 671988 712904 672040 712910
rect 671988 712846 672040 712852
rect 671988 712428 672040 712434
rect 671988 712370 672040 712376
rect 671804 669384 671856 669390
rect 671804 669326 671856 669332
rect 672000 666942 672028 712370
rect 672172 670200 672224 670206
rect 672170 670168 672172 670177
rect 672224 670168 672226 670177
rect 672170 670103 672226 670112
rect 672170 669760 672226 669769
rect 672170 669695 672172 669704
rect 672224 669695 672226 669704
rect 672172 669666 672224 669672
rect 671988 666936 672040 666942
rect 671988 666878 672040 666884
rect 671804 666732 671856 666738
rect 671804 666674 671856 666680
rect 671816 665378 671844 666674
rect 671804 665372 671856 665378
rect 671804 665314 671856 665320
rect 672368 664193 672396 742766
rect 672538 739936 672594 739945
rect 672538 739871 672594 739880
rect 672552 665553 672580 739871
rect 672816 715760 672868 715766
rect 672814 715728 672816 715737
rect 672868 715728 672870 715737
rect 672814 715663 672870 715672
rect 673012 706761 673040 778767
rect 673196 728142 673224 886858
rect 673184 728136 673236 728142
rect 673184 728078 673236 728084
rect 673380 721754 673408 894270
rect 675850 893888 675906 893897
rect 675850 893823 675906 893832
rect 675864 892906 675892 893823
rect 676034 893072 676090 893081
rect 676034 893007 676036 893016
rect 676088 893007 676090 893016
rect 676036 892978 676088 892984
rect 675852 892900 675904 892906
rect 675852 892842 675904 892848
rect 676034 892664 676090 892673
rect 676090 892622 676260 892650
rect 676034 892599 676090 892608
rect 676232 891546 676260 892622
rect 679622 891848 679678 891857
rect 679622 891783 679678 891792
rect 676220 891540 676272 891546
rect 676220 891482 676272 891488
rect 676864 891540 676916 891546
rect 676864 891482 676916 891488
rect 676034 891440 676090 891449
rect 676034 891375 676090 891384
rect 675850 891032 675906 891041
rect 675850 890967 675906 890976
rect 674840 890792 674892 890798
rect 674840 890734 674892 890740
rect 674656 888956 674708 888962
rect 674656 888898 674708 888904
rect 674288 888548 674340 888554
rect 674288 888490 674340 888496
rect 674300 870330 674328 888490
rect 674470 888040 674526 888049
rect 674470 887975 674526 887984
rect 674484 876246 674512 887975
rect 674472 876240 674524 876246
rect 674472 876182 674524 876188
rect 674668 872174 674696 888898
rect 674852 879238 674880 890734
rect 675864 888826 675892 890967
rect 676048 890798 676076 891375
rect 676036 890792 676088 890798
rect 676036 890734 676088 890740
rect 676034 890624 676090 890633
rect 676090 890582 676260 890610
rect 676034 890559 676090 890568
rect 676034 890216 676090 890225
rect 676034 890151 676090 890160
rect 676048 890050 676076 890151
rect 676036 890044 676088 890050
rect 676036 889986 676088 889992
rect 676034 888992 676090 889001
rect 676034 888927 676036 888936
rect 676088 888927 676090 888936
rect 676036 888898 676088 888904
rect 675024 888820 675076 888826
rect 675024 888762 675076 888768
rect 675852 888820 675904 888826
rect 675852 888762 675904 888768
rect 674840 879232 674892 879238
rect 674840 879174 674892 879180
rect 674840 879096 674892 879102
rect 674840 879038 674892 879044
rect 674852 876625 674880 879038
rect 675036 877010 675064 888762
rect 676034 888584 676090 888593
rect 676034 888519 676036 888528
rect 676088 888519 676090 888528
rect 676036 888490 676088 888496
rect 676034 887496 676090 887505
rect 676232 887482 676260 890582
rect 676494 887768 676550 887777
rect 676494 887703 676550 887712
rect 676090 887454 676260 887482
rect 676034 887431 676090 887440
rect 676310 887360 676366 887369
rect 676310 887295 676366 887304
rect 676034 886952 676090 886961
rect 676034 886887 676036 886896
rect 676088 886887 676090 886896
rect 676036 886858 676088 886864
rect 676034 885728 676090 885737
rect 676034 885663 676036 885672
rect 676088 885663 676090 885672
rect 676036 885634 676088 885640
rect 676324 883289 676352 887295
rect 676508 883425 676536 887703
rect 676494 883416 676550 883425
rect 676494 883351 676550 883360
rect 676310 883280 676366 883289
rect 676310 883215 676366 883224
rect 675208 881068 675260 881074
rect 675208 881010 675260 881016
rect 675220 879322 675248 881010
rect 675576 880592 675628 880598
rect 675576 880534 675628 880540
rect 674944 876982 675064 877010
rect 675128 879294 675248 879322
rect 675392 879368 675444 879374
rect 675444 879316 675524 879322
rect 675392 879310 675524 879316
rect 675404 879294 675524 879310
rect 675128 877010 675156 879294
rect 675300 879232 675352 879238
rect 675220 879180 675300 879186
rect 675220 879174 675352 879180
rect 675220 879158 675340 879174
rect 675220 877282 675248 879158
rect 675496 878370 675524 879294
rect 675312 878342 675524 878370
rect 675312 877418 675340 878342
rect 675588 878084 675616 880534
rect 675760 880456 675812 880462
rect 675760 880398 675812 880404
rect 675772 878529 675800 880398
rect 676876 878558 676904 891482
rect 677048 890044 677100 890050
rect 677048 889986 677100 889992
rect 677060 879374 677088 889986
rect 678242 889808 678298 889817
rect 678242 889743 678298 889752
rect 677048 879368 677100 879374
rect 677048 879310 677100 879316
rect 678256 879102 678284 889743
rect 679636 880462 679664 891783
rect 683302 889400 683358 889409
rect 683302 889335 683358 889344
rect 683026 886136 683082 886145
rect 683026 886071 683082 886080
rect 683040 881929 683068 886071
rect 683026 881920 683082 881929
rect 683026 881855 683082 881864
rect 683316 881074 683344 889335
rect 683304 881068 683356 881074
rect 683304 881010 683356 881016
rect 679624 880456 679676 880462
rect 679624 880398 679676 880404
rect 678244 879096 678296 879102
rect 678244 879038 678296 879044
rect 676864 878552 676916 878558
rect 675758 878520 675814 878529
rect 676864 878494 676916 878500
rect 675758 878455 675814 878464
rect 675666 877840 675722 877849
rect 675666 877775 675722 877784
rect 675680 877540 675708 877775
rect 675312 877390 675432 877418
rect 675220 877254 675340 877282
rect 675128 876982 675248 877010
rect 674944 876738 674972 876982
rect 675220 876738 675248 876982
rect 674944 876710 675064 876738
rect 674838 876616 674894 876625
rect 674838 876551 674894 876560
rect 674840 876240 674892 876246
rect 674840 876182 674892 876188
rect 674852 872914 674880 876182
rect 674840 872908 674892 872914
rect 674840 872850 674892 872856
rect 675036 872794 675064 876710
rect 675128 876710 675248 876738
rect 675128 873610 675156 876710
rect 675312 874290 675340 877254
rect 675404 876860 675432 877390
rect 675484 876580 675536 876586
rect 675484 876522 675536 876528
rect 675496 876248 675524 876522
rect 675404 874290 675432 874412
rect 675312 874262 675432 874290
rect 675482 874168 675538 874177
rect 675482 874103 675538 874112
rect 675496 873868 675524 874103
rect 675128 873582 675432 873610
rect 675404 873188 675432 873582
rect 675392 872908 675444 872914
rect 675392 872850 675444 872856
rect 674576 872146 674696 872174
rect 674852 872766 675064 872794
rect 675404 872794 675432 872850
rect 675404 872766 675524 872794
rect 674288 870324 674340 870330
rect 674288 870266 674340 870272
rect 674576 869666 674604 872146
rect 674852 870505 674880 872766
rect 675496 872576 675524 872766
rect 675206 872400 675262 872409
rect 675206 872335 675262 872344
rect 674838 870496 674894 870505
rect 674838 870431 674894 870440
rect 674932 870324 674984 870330
rect 674932 870266 674984 870272
rect 674576 869638 674880 869666
rect 674852 868889 674880 869638
rect 674944 869414 674972 870266
rect 674944 869386 675064 869414
rect 675036 869281 675064 869386
rect 675220 869378 675248 872335
rect 675482 870496 675538 870505
rect 675482 870431 675538 870440
rect 675496 870060 675524 870431
rect 675574 869816 675630 869825
rect 675574 869751 675630 869760
rect 675588 869516 675616 869751
rect 675208 869372 675260 869378
rect 675208 869314 675260 869320
rect 675022 869272 675078 869281
rect 675022 869207 675078 869216
rect 675390 869272 675446 869281
rect 675390 869207 675446 869216
rect 675208 869168 675260 869174
rect 675208 869110 675260 869116
rect 675024 869032 675076 869038
rect 675024 868974 675076 868980
rect 674852 868861 674972 868889
rect 674944 868442 674972 868861
rect 675036 868850 675064 868974
rect 675036 868822 675156 868850
rect 674944 868414 675064 868442
rect 674840 868080 674892 868086
rect 674840 868022 674892 868028
rect 674852 866289 674880 868022
rect 675036 867354 675064 868414
rect 675128 867694 675156 868822
rect 675220 868238 675248 869110
rect 675404 868875 675432 869207
rect 675220 868210 675418 868238
rect 675128 867666 675418 867694
rect 675036 867326 675432 867354
rect 675114 867232 675170 867241
rect 675114 867167 675170 867176
rect 674838 866280 674894 866289
rect 674838 866215 674894 866224
rect 675128 866130 675156 867167
rect 675404 867035 675432 867326
rect 675390 866280 675446 866289
rect 675390 866215 675446 866224
rect 675128 866102 675340 866130
rect 675114 865736 675170 865745
rect 675114 865671 675170 865680
rect 675128 863342 675156 865671
rect 675312 864566 675340 866102
rect 675404 865844 675432 866215
rect 675758 865464 675814 865473
rect 675758 865399 675814 865408
rect 675772 865195 675800 865399
rect 675312 864538 675418 864566
rect 675312 863382 675432 863410
rect 675312 863342 675340 863382
rect 675128 863314 675340 863342
rect 675404 863328 675432 863382
rect 675392 790832 675444 790838
rect 675392 790774 675444 790780
rect 675116 789404 675168 789410
rect 675116 789346 675168 789352
rect 675128 787693 675156 789346
rect 675404 788868 675432 790774
rect 675772 788089 675800 788324
rect 675758 788080 675814 788089
rect 675758 788015 675814 788024
rect 675128 787665 675418 787693
rect 675128 787018 675418 787046
rect 675128 786729 675156 787018
rect 675114 786720 675170 786729
rect 675114 786655 675170 786664
rect 674944 785182 675418 785210
rect 674472 783896 674524 783902
rect 674472 783838 674524 783844
rect 673734 780056 673790 780065
rect 673734 779991 673790 780000
rect 673550 738712 673606 738721
rect 673550 738647 673606 738656
rect 673196 721726 673408 721754
rect 673196 714513 673224 721726
rect 673368 716168 673420 716174
rect 673368 716110 673420 716116
rect 673380 715329 673408 716110
rect 673366 715320 673422 715329
rect 673366 715255 673422 715264
rect 673366 714912 673422 714921
rect 673366 714847 673368 714856
rect 673420 714847 673422 714856
rect 673368 714818 673420 714824
rect 673182 714504 673238 714513
rect 673182 714439 673238 714448
rect 672998 706752 673054 706761
rect 672998 706687 673054 706696
rect 673368 705560 673420 705566
rect 673366 705528 673368 705537
rect 673420 705528 673422 705537
rect 673366 705463 673422 705472
rect 673366 705256 673422 705265
rect 673366 705191 673422 705200
rect 673182 703896 673238 703905
rect 673182 703831 673184 703840
rect 673236 703831 673238 703840
rect 673184 703802 673236 703808
rect 673184 701208 673236 701214
rect 673182 701176 673184 701185
rect 673236 701176 673238 701185
rect 673182 701111 673238 701120
rect 673000 701072 673052 701078
rect 673000 701014 673052 701020
rect 673012 700913 673040 701014
rect 672998 700904 673054 700913
rect 672998 700839 673054 700848
rect 673380 695534 673408 705191
rect 673288 695506 673408 695534
rect 672998 695328 673054 695337
rect 672998 695263 673054 695272
rect 672814 695056 672870 695065
rect 672814 694991 672870 695000
rect 672828 692774 672856 694991
rect 672828 692746 672948 692774
rect 672722 684992 672778 685001
rect 672722 684927 672778 684936
rect 672538 665544 672594 665553
rect 672538 665479 672594 665488
rect 672354 664184 672410 664193
rect 672354 664119 672410 664128
rect 672736 663794 672764 684927
rect 672920 678974 672948 692746
rect 673012 688634 673040 695263
rect 673288 690690 673316 695506
rect 673564 693297 673592 738647
rect 673748 724418 673776 779991
rect 674288 777028 674340 777034
rect 674288 776970 674340 776976
rect 674102 734904 674158 734913
rect 674102 734839 674158 734848
rect 673918 734224 673974 734233
rect 673918 734159 673974 734168
rect 673932 727274 673960 734159
rect 673840 727246 673960 727274
rect 673840 724514 673868 727246
rect 673840 724486 674052 724514
rect 673748 724390 673960 724418
rect 673932 723058 673960 724390
rect 673840 723030 673960 723058
rect 673840 722401 673868 723030
rect 673826 722392 673882 722401
rect 673826 722327 673882 722336
rect 674024 722242 674052 724486
rect 673932 722226 674052 722242
rect 673736 722220 673788 722226
rect 673736 722162 673788 722168
rect 673920 722220 674052 722226
rect 673972 722214 674052 722220
rect 673920 722162 673972 722168
rect 673748 721754 673776 722162
rect 674116 721857 674144 734839
rect 674300 726578 674328 776970
rect 674484 727938 674512 783838
rect 674748 782672 674800 782678
rect 674748 782614 674800 782620
rect 674760 782474 674788 782614
rect 674760 782446 674880 782474
rect 674654 779240 674710 779249
rect 674654 779175 674710 779184
rect 674472 727932 674524 727938
rect 674472 727874 674524 727880
rect 674668 726714 674696 779175
rect 674852 776257 674880 782446
rect 674944 776506 674972 785182
rect 675114 784680 675170 784689
rect 675170 784638 675418 784666
rect 675114 784615 675170 784624
rect 675312 784094 675432 784122
rect 675312 783986 675340 784094
rect 675128 783958 675340 783986
rect 675404 783972 675432 784094
rect 675128 783902 675156 783958
rect 675116 783896 675168 783902
rect 675116 783838 675168 783844
rect 675220 783346 675418 783374
rect 675220 782678 675248 783346
rect 675208 782672 675260 782678
rect 675208 782614 675260 782620
rect 675208 781108 675260 781114
rect 675208 781050 675260 781056
rect 675220 778478 675248 781050
rect 675496 780609 675524 780844
rect 675482 780600 675538 780609
rect 675482 780535 675538 780544
rect 675496 780065 675524 780300
rect 675482 780056 675538 780065
rect 675482 779991 675538 780000
rect 675404 779249 675432 779688
rect 675390 779240 675446 779249
rect 675390 779175 675446 779184
rect 675496 778841 675524 779008
rect 675482 778832 675538 778841
rect 675482 778767 675538 778776
rect 675220 778450 675418 778478
rect 675208 778388 675260 778394
rect 675208 778330 675260 778336
rect 675220 778274 675248 778330
rect 675128 778246 675248 778274
rect 675128 776914 675156 778246
rect 675404 777322 675432 777852
rect 675312 777294 675432 777322
rect 675312 777034 675340 777294
rect 675300 777028 675352 777034
rect 675300 776970 675352 776976
rect 675128 776886 675248 776914
rect 675220 776642 675248 776886
rect 675220 776614 675418 776642
rect 674944 776478 675340 776506
rect 674838 776248 674894 776257
rect 674838 776183 674894 776192
rect 674840 775600 674892 775606
rect 674840 775542 674892 775548
rect 675114 775568 675170 775577
rect 674852 774625 674880 775542
rect 675114 775503 675170 775512
rect 674838 774616 674894 774625
rect 674838 774551 674894 774560
rect 675128 772814 675156 775503
rect 675128 772786 675248 772814
rect 675220 760394 675248 772786
rect 675036 760366 675248 760394
rect 674840 741124 674892 741130
rect 674840 741066 674892 741072
rect 674852 740654 674880 741066
rect 674840 740648 674892 740654
rect 674840 740590 674892 740596
rect 675036 739786 675064 760366
rect 675312 750734 675340 776478
rect 675496 775849 675524 776016
rect 675482 775840 675538 775849
rect 675482 775775 675538 775784
rect 675496 775033 675524 775336
rect 675482 775024 675538 775033
rect 675482 774959 675538 774968
rect 675482 774616 675538 774625
rect 675482 774551 675538 774560
rect 675496 774180 675524 774551
rect 674852 739758 675064 739786
rect 675128 750706 675340 750734
rect 674852 727530 674880 739758
rect 675128 738970 675156 750706
rect 675392 744048 675444 744054
rect 675392 743990 675444 743996
rect 675404 743852 675432 743990
rect 675312 743294 675418 743322
rect 675312 743238 675340 743294
rect 675300 743232 675352 743238
rect 675300 743174 675352 743180
rect 675484 742824 675536 742830
rect 675484 742766 675536 742772
rect 675496 742696 675524 742766
rect 675390 742248 675446 742257
rect 675390 742183 675446 742192
rect 675404 742016 675432 742183
rect 675392 740648 675444 740654
rect 675312 740596 675392 740602
rect 675312 740590 675444 740596
rect 675312 740574 675432 740590
rect 675312 739786 675340 740574
rect 675496 739945 675524 740180
rect 675482 739936 675538 739945
rect 675482 739871 675538 739880
rect 675312 739758 675432 739786
rect 675404 739636 675432 739758
rect 674944 738942 675156 738970
rect 674944 728226 674972 738942
rect 675496 738721 675524 739024
rect 675482 738712 675538 738721
rect 675482 738647 675538 738656
rect 675496 738177 675524 738344
rect 675482 738168 675538 738177
rect 675482 738103 675538 738112
rect 675208 735752 675260 735758
rect 675404 735729 675432 735896
rect 675208 735694 675260 735700
rect 675390 735720 675446 735729
rect 675220 735570 675248 735694
rect 675390 735655 675446 735664
rect 675220 735542 675340 735570
rect 675116 734256 675168 734262
rect 675116 734198 675168 734204
rect 675128 731626 675156 734198
rect 675312 733493 675340 735542
rect 675496 734913 675524 735319
rect 675482 734904 675538 734913
rect 675482 734839 675538 734848
rect 675496 734233 675524 734672
rect 675482 734224 675538 734233
rect 675482 734159 675538 734168
rect 675588 733825 675616 734031
rect 675574 733816 675630 733825
rect 675574 733751 675630 733760
rect 675312 733465 675418 733493
rect 675300 733372 675352 733378
rect 675300 733314 675352 733320
rect 675312 732850 675340 733314
rect 675312 732822 675418 732850
rect 675312 731734 675432 731762
rect 675312 731626 675340 731734
rect 675128 731598 675340 731626
rect 675404 731612 675432 731734
rect 675312 730986 675418 731014
rect 675312 728328 675340 730986
rect 675496 730153 675524 730351
rect 675482 730144 675538 730153
rect 675482 730079 675538 730088
rect 675496 728793 675524 729164
rect 675482 728784 675538 728793
rect 675482 728719 675538 728728
rect 675312 728300 675524 728328
rect 674944 728198 675340 728226
rect 674840 727524 674892 727530
rect 674840 727466 674892 727472
rect 675116 727524 675168 727530
rect 675116 727466 675168 727472
rect 674930 727288 674986 727297
rect 674930 727223 674986 727232
rect 674656 726708 674708 726714
rect 674656 726650 674708 726656
rect 674288 726572 674340 726578
rect 674288 726514 674340 726520
rect 674102 721848 674158 721857
rect 674102 721783 674158 721792
rect 673656 721726 673776 721754
rect 673656 695534 673684 721726
rect 674944 721721 674972 727223
rect 675128 721750 675156 727466
rect 675312 721750 675340 728198
rect 675496 727530 675524 728300
rect 683488 727932 683540 727938
rect 683488 727874 683540 727880
rect 675484 727524 675536 727530
rect 675484 727466 675536 727472
rect 678244 727252 678296 727258
rect 678244 727194 678296 727200
rect 675116 721744 675168 721750
rect 674930 721712 674986 721721
rect 675116 721686 675168 721692
rect 675300 721744 675352 721750
rect 675300 721686 675352 721692
rect 674930 721647 674986 721656
rect 675116 721268 675168 721274
rect 675116 721210 675168 721216
rect 675300 721268 675352 721274
rect 675300 721210 675352 721216
rect 675128 720866 675156 721210
rect 675312 720866 675340 721210
rect 675116 720860 675168 720866
rect 675116 720802 675168 720808
rect 675300 720860 675352 720866
rect 675300 720802 675352 720808
rect 675116 720520 675168 720526
rect 675116 720462 675168 720468
rect 675300 720520 675352 720526
rect 675300 720462 675352 720468
rect 674194 720080 674250 720089
rect 674194 720015 674250 720024
rect 674010 717088 674066 717097
rect 674010 717023 674066 717032
rect 673826 716544 673882 716553
rect 673826 716479 673882 716488
rect 673840 716310 673868 716479
rect 673828 716304 673880 716310
rect 673828 716246 673880 716252
rect 673826 716136 673882 716145
rect 673826 716071 673882 716080
rect 673840 715018 673868 716071
rect 673828 715012 673880 715018
rect 673828 714954 673880 714960
rect 673826 714096 673882 714105
rect 673826 714031 673828 714040
rect 673880 714031 673882 714040
rect 673828 714002 673880 714008
rect 673828 713720 673880 713726
rect 673826 713688 673828 713697
rect 673880 713688 673882 713697
rect 673826 713623 673882 713632
rect 673826 713280 673882 713289
rect 673826 713215 673828 713224
rect 673880 713215 673882 713224
rect 673828 713186 673880 713192
rect 673828 712904 673880 712910
rect 673826 712872 673828 712881
rect 673880 712872 673882 712881
rect 673826 712807 673882 712816
rect 673826 712464 673882 712473
rect 673826 712399 673828 712408
rect 673880 712399 673882 712408
rect 673828 712370 673880 712376
rect 673828 711680 673880 711686
rect 673826 711648 673828 711657
rect 673880 711648 673882 711657
rect 673826 711583 673882 711592
rect 673828 710048 673880 710054
rect 673826 710016 673828 710025
rect 673880 710016 673882 710025
rect 673826 709951 673882 709960
rect 673828 709640 673880 709646
rect 673826 709608 673828 709617
rect 673880 709608 673882 709617
rect 673826 709543 673882 709552
rect 674024 702434 674052 717023
rect 674208 713474 674236 720015
rect 674116 713446 674236 713474
rect 674116 707954 674144 713446
rect 674288 708008 674340 708014
rect 674288 707954 674340 707956
rect 674116 707950 674340 707954
rect 674116 707926 674328 707950
rect 674472 705628 674524 705634
rect 674472 705570 674524 705576
rect 674286 705528 674342 705537
rect 674286 705463 674342 705472
rect 674300 705362 674328 705463
rect 674288 705356 674340 705362
rect 674288 705298 674340 705304
rect 674484 705265 674512 705570
rect 674470 705256 674526 705265
rect 674470 705191 674526 705200
rect 674288 703928 674340 703934
rect 674286 703896 674288 703905
rect 674340 703896 674342 703905
rect 674286 703831 674342 703840
rect 674024 702406 674144 702434
rect 673656 695506 673960 695534
rect 673550 693288 673606 693297
rect 673550 693223 673606 693232
rect 673550 693016 673606 693025
rect 673550 692951 673606 692960
rect 673564 692774 673592 692951
rect 673932 692866 673960 695506
rect 673472 692746 673592 692774
rect 673840 692838 673960 692866
rect 673288 690662 673408 690690
rect 673184 690056 673236 690062
rect 673182 690024 673184 690033
rect 673236 690024 673238 690033
rect 673182 689959 673238 689968
rect 673184 688832 673236 688838
rect 673182 688800 673184 688809
rect 673236 688800 673238 688809
rect 673182 688735 673238 688744
rect 673012 688606 673224 688634
rect 672920 678946 673040 678974
rect 672644 663766 672764 663794
rect 671620 661564 671672 661570
rect 671620 661506 671672 661512
rect 672644 659002 672672 663766
rect 672814 659696 672870 659705
rect 672814 659631 672870 659640
rect 672644 658974 672764 659002
rect 671986 652488 672042 652497
rect 671986 652423 672042 652432
rect 671802 649768 671858 649777
rect 671802 649703 671858 649712
rect 671618 647864 671674 647873
rect 671618 647799 671674 647808
rect 671436 623688 671488 623694
rect 671436 623630 671488 623636
rect 671252 622872 671304 622878
rect 671252 622814 671304 622820
rect 671436 622260 671488 622266
rect 671436 622202 671488 622208
rect 670976 618112 671028 618118
rect 670976 618054 671028 618060
rect 670608 614916 670660 614922
rect 670608 614858 670660 614864
rect 670424 574592 670476 574598
rect 670424 574534 670476 574540
rect 670422 549808 670478 549817
rect 670422 549743 670478 549752
rect 670240 534336 670292 534342
rect 670240 534278 670292 534284
rect 669964 491496 670016 491502
rect 669964 491438 670016 491444
rect 670436 480962 670464 549743
rect 670424 480956 670476 480962
rect 670424 480898 670476 480904
rect 669778 455424 669834 455433
rect 669778 455359 669834 455368
rect 670620 455025 670648 614858
rect 671158 607336 671214 607345
rect 671158 607271 671214 607280
rect 670882 600400 670938 600409
rect 670882 600335 670884 600344
rect 670936 600335 670938 600344
rect 670884 600306 670936 600312
rect 670790 599176 670846 599185
rect 670790 599111 670792 599120
rect 670844 599111 670846 599120
rect 670792 599082 670844 599088
rect 670974 593600 671030 593609
rect 670974 593535 671030 593544
rect 670790 533896 670846 533905
rect 670790 533831 670846 533840
rect 670804 490958 670832 533831
rect 670988 529514 671016 593535
rect 670976 529508 671028 529514
rect 670976 529450 671028 529456
rect 671172 529242 671200 607271
rect 671448 577454 671476 622202
rect 671436 577448 671488 577454
rect 671436 577390 671488 577396
rect 671344 576972 671396 576978
rect 671344 576914 671396 576920
rect 671356 532273 671384 576914
rect 671632 572150 671660 647799
rect 671816 575414 671844 649703
rect 671804 575408 671856 575414
rect 671804 575350 671856 575356
rect 672000 574326 672028 652423
rect 672538 649224 672594 649233
rect 672538 649159 672594 649168
rect 672356 637424 672408 637430
rect 672356 637366 672408 637372
rect 672368 632738 672396 637366
rect 672356 632732 672408 632738
rect 672356 632674 672408 632680
rect 672354 604344 672410 604353
rect 672354 604279 672410 604288
rect 672368 596290 672396 604279
rect 672356 596284 672408 596290
rect 672356 596226 672408 596232
rect 671988 574320 672040 574326
rect 671988 574262 672040 574268
rect 672552 573782 672580 649159
rect 672736 637514 672764 658974
rect 672644 637486 672764 637514
rect 672644 632890 672672 637486
rect 672828 637430 672856 659631
rect 672816 637424 672868 637430
rect 672816 637366 672868 637372
rect 672644 632862 672948 632890
rect 672724 632732 672776 632738
rect 672724 632674 672776 632680
rect 672736 627914 672764 632674
rect 672736 627886 672856 627914
rect 672828 625954 672856 627886
rect 672644 625926 672856 625954
rect 672644 600930 672672 625926
rect 672920 621014 672948 632862
rect 672828 620986 672948 621014
rect 672828 615670 672856 620986
rect 673012 618633 673040 678946
rect 673196 619342 673224 688606
rect 673184 619336 673236 619342
rect 673184 619278 673236 619284
rect 672998 618624 673054 618633
rect 672998 618559 673054 618568
rect 672816 615664 672868 615670
rect 672816 615606 672868 615612
rect 673182 608152 673238 608161
rect 673182 608087 673238 608096
rect 672998 604072 673054 604081
rect 672998 604007 673054 604016
rect 672644 600902 672948 600930
rect 672724 596284 672776 596290
rect 672724 596226 672776 596232
rect 672540 573776 672592 573782
rect 672540 573718 672592 573724
rect 671620 572144 671672 572150
rect 671620 572086 671672 572092
rect 671988 570852 672040 570858
rect 671988 570794 672040 570800
rect 671802 562456 671858 562465
rect 671802 562391 671858 562400
rect 671526 533080 671582 533089
rect 671526 533015 671582 533024
rect 671342 532264 671398 532273
rect 671342 532199 671398 532208
rect 671342 531584 671398 531593
rect 671342 531519 671398 531528
rect 671160 529236 671212 529242
rect 671160 529178 671212 529184
rect 670792 490952 670844 490958
rect 670792 490894 670844 490900
rect 671356 488510 671384 531519
rect 671540 489326 671568 533015
rect 671528 489320 671580 489326
rect 671528 489262 671580 489268
rect 671344 488504 671396 488510
rect 671344 488446 671396 488452
rect 671816 486878 671844 562391
rect 671804 486872 671856 486878
rect 671804 486814 671856 486820
rect 672000 455138 672028 570794
rect 672262 555248 672318 555257
rect 672262 555183 672318 555192
rect 672276 486062 672304 555183
rect 672736 549254 672764 596226
rect 672920 596174 672948 600902
rect 672644 549226 672764 549254
rect 672828 596146 672948 596174
rect 672828 549254 672856 596146
rect 672828 549226 672948 549254
rect 672644 544610 672672 549226
rect 672632 544604 672684 544610
rect 672632 544546 672684 544552
rect 672920 544490 672948 549226
rect 672644 544462 672948 544490
rect 672644 536058 672672 544462
rect 672816 544400 672868 544406
rect 672868 544348 672948 544354
rect 672816 544342 672948 544348
rect 672828 544326 672948 544342
rect 672644 536030 672856 536058
rect 672632 535016 672684 535022
rect 672630 534984 672632 534993
rect 672684 534984 672686 534993
rect 672630 534919 672686 534928
rect 672632 534336 672684 534342
rect 672632 534278 672684 534284
rect 672644 534177 672672 534278
rect 672630 534168 672686 534177
rect 672630 534103 672686 534112
rect 672632 533384 672684 533390
rect 672630 533352 672632 533361
rect 672684 533352 672686 533361
rect 672630 533287 672686 533296
rect 672538 532808 672594 532817
rect 672538 532743 672594 532752
rect 672552 499574 672580 532743
rect 672552 499546 672672 499574
rect 672644 490142 672672 499546
rect 672632 490136 672684 490142
rect 672632 490078 672684 490084
rect 672632 489932 672684 489938
rect 672632 489874 672684 489880
rect 672448 489660 672500 489666
rect 672448 489602 672500 489608
rect 672264 486056 672316 486062
rect 672264 485998 672316 486004
rect 672000 455122 672120 455138
rect 672000 455116 672132 455122
rect 672000 455110 672080 455116
rect 672080 455058 672132 455064
rect 670606 455016 670662 455025
rect 670606 454951 670662 454960
rect 672264 453960 672316 453966
rect 672262 453928 672264 453937
rect 672316 453928 672318 453937
rect 672262 453863 672318 453872
rect 672460 401713 672488 489602
rect 672644 402121 672672 489874
rect 672828 455802 672856 536030
rect 672920 529802 672948 544326
rect 673012 529972 673040 604007
rect 673196 543734 673224 608087
rect 673104 543706 673224 543734
rect 673104 534018 673132 543706
rect 673104 533990 673224 534018
rect 673196 530126 673224 533990
rect 673184 530120 673236 530126
rect 673184 530062 673236 530068
rect 673012 529944 673316 529972
rect 672920 529774 673040 529802
rect 673012 528902 673040 529774
rect 673000 528896 673052 528902
rect 673000 528838 673052 528844
rect 673288 528554 673316 529944
rect 673196 528526 673316 528554
rect 673196 527241 673224 528526
rect 673182 527232 673238 527241
rect 673182 527167 673238 527176
rect 673184 493332 673236 493338
rect 673184 493274 673236 493280
rect 673196 492153 673224 493274
rect 673182 492144 673238 492153
rect 673182 492079 673238 492088
rect 673182 490512 673238 490521
rect 673182 490447 673238 490456
rect 673196 489938 673224 490447
rect 673184 489932 673236 489938
rect 673184 489874 673236 489880
rect 673380 475522 673408 690662
rect 673472 678974 673500 692746
rect 673644 685976 673696 685982
rect 673644 685918 673696 685924
rect 673656 685817 673684 685918
rect 673642 685808 673698 685817
rect 673642 685743 673698 685752
rect 673472 678946 673592 678974
rect 673564 670834 673592 678946
rect 673840 676214 673868 692838
rect 674116 692774 674144 702406
rect 675128 701457 675156 720462
rect 675312 710841 675340 720462
rect 675298 710832 675354 710841
rect 675298 710767 675354 710776
rect 678256 710433 678284 727194
rect 683304 726708 683356 726714
rect 683304 726650 683356 726656
rect 682382 726608 682438 726617
rect 682382 726543 682438 726552
rect 682396 711249 682424 726543
rect 682382 711240 682438 711249
rect 682382 711175 682438 711184
rect 678242 710424 678298 710433
rect 678242 710359 678298 710368
rect 676036 708008 676088 708014
rect 683316 707985 683344 726650
rect 683500 708801 683528 727874
rect 684132 726572 684184 726578
rect 684132 726514 684184 726520
rect 683486 708792 683542 708801
rect 683486 708727 683542 708736
rect 684144 708393 684172 726514
rect 703694 717196 703722 717264
rect 704154 717196 704182 717264
rect 704614 717196 704642 717264
rect 705074 717196 705102 717264
rect 705534 717196 705562 717264
rect 705994 717196 706022 717264
rect 706454 717196 706482 717264
rect 706914 717196 706942 717264
rect 707374 717196 707402 717264
rect 707834 717196 707862 717264
rect 708294 717196 708322 717264
rect 708754 717196 708782 717264
rect 709214 717196 709242 717264
rect 684130 708384 684186 708393
rect 684130 708319 684186 708328
rect 676036 707950 676088 707956
rect 683302 707976 683358 707985
rect 676048 707169 676076 707950
rect 683302 707911 683358 707920
rect 676034 707160 676090 707169
rect 676034 707095 676090 707104
rect 676034 706344 676090 706353
rect 676034 706279 676090 706288
rect 676048 705634 676076 706279
rect 676036 705628 676088 705634
rect 676036 705570 676088 705576
rect 683118 705528 683174 705537
rect 683118 705463 683174 705472
rect 683132 705362 683160 705463
rect 683120 705356 683172 705362
rect 683120 705298 683172 705304
rect 676034 705120 676090 705129
rect 676034 705055 676090 705064
rect 676048 703934 676076 705055
rect 676036 703928 676088 703934
rect 676036 703870 676088 703876
rect 675114 701448 675170 701457
rect 675114 701383 675170 701392
rect 675114 701176 675170 701185
rect 675114 701111 675170 701120
rect 674930 700904 674986 700913
rect 674930 700839 674986 700848
rect 674944 698337 674972 700839
rect 675128 698889 675156 701111
rect 675128 698861 675418 698889
rect 674944 698309 675418 698337
rect 675128 697666 675418 697694
rect 675128 696969 675156 697666
rect 675114 696960 675170 696969
rect 675114 696895 675170 696904
rect 675496 696833 675524 697035
rect 675482 696824 675538 696833
rect 675482 696759 675538 696768
rect 675114 696144 675170 696153
rect 675114 696079 675170 696088
rect 675128 695209 675156 696079
rect 675128 695181 675418 695209
rect 675114 695056 675170 695065
rect 675114 694991 675170 695000
rect 675298 695056 675354 695065
rect 675298 694991 675354 695000
rect 675128 694022 675156 694991
rect 675312 694906 675340 694991
rect 675312 694878 675432 694906
rect 675404 694620 675432 694878
rect 675128 693994 675418 694022
rect 675496 693025 675524 693328
rect 675482 693016 675538 693025
rect 675482 692951 675538 692960
rect 673932 692746 674144 692774
rect 673932 688634 673960 692746
rect 674300 690866 675418 690894
rect 674102 690432 674158 690441
rect 674102 690367 674158 690376
rect 674116 688634 674144 690367
rect 674300 688634 674328 690866
rect 675298 690432 675354 690441
rect 675298 690367 675354 690376
rect 675312 690282 675340 690367
rect 675404 690282 675432 690336
rect 675312 690254 675432 690282
rect 674930 690024 674986 690033
rect 674930 689959 674986 689968
rect 674654 688800 674710 688809
rect 674710 688758 674880 688786
rect 674654 688735 674710 688744
rect 673932 688606 674052 688634
rect 674116 688606 674236 688634
rect 674300 688606 674420 688634
rect 674024 678974 674052 688606
rect 674208 678974 674236 688606
rect 674392 687290 674420 688606
rect 674654 688120 674710 688129
rect 674654 688055 674710 688064
rect 673748 676186 673868 676214
rect 673932 678946 674052 678974
rect 674116 678946 674236 678974
rect 674300 687262 674420 687290
rect 673748 674393 673776 676186
rect 673734 674384 673790 674393
rect 673734 674319 673790 674328
rect 673734 671392 673790 671401
rect 673734 671327 673736 671336
rect 673788 671327 673790 671336
rect 673736 671298 673788 671304
rect 673736 671152 673788 671158
rect 673736 671094 673788 671100
rect 673748 670993 673776 671094
rect 673734 670984 673790 670993
rect 673734 670919 673790 670928
rect 673564 670806 673776 670834
rect 673550 670576 673606 670585
rect 673550 670511 673606 670520
rect 673564 669594 673592 670511
rect 673552 669588 673604 669594
rect 673552 669530 673604 669536
rect 673552 669248 673604 669254
rect 673550 669216 673552 669225
rect 673604 669216 673606 669225
rect 673550 669151 673606 669160
rect 673550 668944 673606 668953
rect 673550 668879 673606 668888
rect 673564 668710 673592 668879
rect 673552 668704 673604 668710
rect 673552 668646 673604 668652
rect 673550 668536 673606 668545
rect 673550 668471 673606 668480
rect 673564 668302 673592 668471
rect 673552 668296 673604 668302
rect 673552 668238 673604 668244
rect 673550 668128 673606 668137
rect 673550 668063 673606 668072
rect 673564 667962 673592 668063
rect 673552 667956 673604 667962
rect 673552 667898 673604 667904
rect 673550 667720 673606 667729
rect 673550 667655 673606 667664
rect 673564 666942 673592 667655
rect 673552 666936 673604 666942
rect 673552 666878 673604 666884
rect 673550 666768 673606 666777
rect 673550 666703 673552 666712
rect 673604 666703 673606 666712
rect 673552 666674 673604 666680
rect 673748 666618 673776 670806
rect 673656 666590 673776 666618
rect 673656 666346 673684 666590
rect 673656 666318 673776 666346
rect 673550 666088 673606 666097
rect 673550 666023 673606 666032
rect 673564 665718 673592 666023
rect 673552 665712 673604 665718
rect 673552 665654 673604 665660
rect 673550 665272 673606 665281
rect 673550 665207 673552 665216
rect 673604 665207 673606 665216
rect 673552 665178 673604 665184
rect 673550 664864 673606 664873
rect 673550 664799 673606 664808
rect 673564 664358 673592 664799
rect 673552 664352 673604 664358
rect 673552 664294 673604 664300
rect 673552 663808 673604 663814
rect 673552 663750 673604 663756
rect 673564 663649 673592 663750
rect 673550 663640 673606 663649
rect 673550 663575 673606 663584
rect 673552 663400 673604 663406
rect 673552 663342 673604 663348
rect 673564 662017 673592 663342
rect 673550 662008 673606 662017
rect 673550 661943 673606 661952
rect 673550 644872 673606 644881
rect 673550 644807 673606 644816
rect 673564 630578 673592 644807
rect 673748 635497 673776 666318
rect 673932 663406 673960 678946
rect 673920 663400 673972 663406
rect 673920 663342 673972 663348
rect 673918 663096 673974 663105
rect 673918 663031 673974 663040
rect 673932 662794 673960 663031
rect 673920 662788 673972 662794
rect 673920 662730 673972 662736
rect 673918 661600 673974 661609
rect 673918 661535 673920 661544
rect 673972 661535 673974 661544
rect 673920 661506 673972 661512
rect 673918 661192 673974 661201
rect 673918 661127 673920 661136
rect 673972 661127 673974 661136
rect 673920 661098 673972 661104
rect 673920 660136 673972 660142
rect 673918 660104 673920 660113
rect 673972 660104 673974 660113
rect 673918 660039 673974 660048
rect 673918 655616 673974 655625
rect 673918 655551 673920 655560
rect 673972 655551 673974 655560
rect 673920 655522 673972 655528
rect 674116 654134 674144 678946
rect 674116 654106 674236 654134
rect 674012 647352 674064 647358
rect 674010 647320 674012 647329
rect 674064 647320 674066 647329
rect 674010 647255 674066 647264
rect 674012 645924 674064 645930
rect 674012 645866 674064 645872
rect 674024 645561 674052 645866
rect 674010 645552 674066 645561
rect 674010 645487 674066 645496
rect 674012 643136 674064 643142
rect 674010 643104 674012 643113
rect 674064 643104 674066 643113
rect 674010 643039 674066 643048
rect 673918 641744 673974 641753
rect 673918 641679 673974 641688
rect 673734 635488 673790 635497
rect 673734 635423 673790 635432
rect 673564 630550 673776 630578
rect 673552 627700 673604 627706
rect 673552 627642 673604 627648
rect 673564 626534 673592 627642
rect 673472 626506 673592 626534
rect 673472 616026 673500 626506
rect 673472 615998 673592 616026
rect 673564 613562 673592 615998
rect 673552 613556 673604 613562
rect 673552 613498 673604 613504
rect 673748 613442 673776 630550
rect 673932 627706 673960 641679
rect 674208 640334 674236 654106
rect 674300 649994 674328 687262
rect 674472 687132 674524 687138
rect 674472 687074 674524 687080
rect 674484 649994 674512 687074
rect 674668 682446 674696 688055
rect 674852 686678 674880 688758
rect 674944 688242 674972 689959
rect 675312 689710 675432 689738
rect 675312 689670 675340 689710
rect 675128 689642 675340 689670
rect 675404 689656 675432 689710
rect 675128 689217 675156 689642
rect 675114 689208 675170 689217
rect 675114 689143 675170 689152
rect 675128 689030 675418 689058
rect 675128 688401 675156 689030
rect 675114 688392 675170 688401
rect 675114 688327 675170 688336
rect 675404 688242 675432 688500
rect 674944 688214 675432 688242
rect 675128 687806 675418 687834
rect 675128 687274 675156 687806
rect 675116 687268 675168 687274
rect 675116 687210 675168 687216
rect 674852 686650 675340 686678
rect 675312 686610 675340 686650
rect 675404 686610 675432 686664
rect 675312 686582 675432 686610
rect 675036 686038 675340 686066
rect 675036 685998 675064 686038
rect 674852 685970 675064 685998
rect 675312 685998 675340 686038
rect 675312 685970 675418 685998
rect 674656 682440 674708 682446
rect 674656 682382 674708 682388
rect 674852 676433 674880 685970
rect 675298 685808 675354 685817
rect 675298 685743 675354 685752
rect 675312 684570 675340 685743
rect 675496 685001 675524 685372
rect 675482 684992 675538 685001
rect 675482 684927 675538 684936
rect 675312 684542 675432 684570
rect 675404 684148 675432 684542
rect 683212 682440 683264 682446
rect 683212 682382 683264 682388
rect 683394 682408 683450 682417
rect 675758 681456 675814 681465
rect 675758 681391 675814 681400
rect 675390 681048 675446 681057
rect 675390 680983 675446 680992
rect 674838 676424 674894 676433
rect 674838 676359 674894 676368
rect 675404 676214 675432 680983
rect 675772 676433 675800 681391
rect 675758 676424 675814 676433
rect 675758 676359 675814 676368
rect 675312 676186 675432 676214
rect 674654 674384 674710 674393
rect 674654 674319 674710 674328
rect 674668 662998 674696 674319
rect 675312 669314 675340 676186
rect 675220 669286 675340 669314
rect 675220 667894 675248 669286
rect 675208 667888 675260 667894
rect 675208 667830 675260 667836
rect 676036 667888 676088 667894
rect 676036 667830 676088 667836
rect 676048 666777 676076 667830
rect 676034 666768 676090 666777
rect 676034 666703 676090 666712
rect 674840 663944 674892 663950
rect 674840 663886 674892 663892
rect 676220 663944 676272 663950
rect 676220 663886 676272 663892
rect 674852 663649 674880 663886
rect 676232 663785 676260 663886
rect 683224 663785 683252 682382
rect 683394 682343 683450 682352
rect 676218 663776 676274 663785
rect 676218 663711 676274 663720
rect 683210 663776 683266 663785
rect 683210 663711 683266 663720
rect 674838 663640 674894 663649
rect 674838 663575 674894 663584
rect 674656 662992 674708 662998
rect 676220 662992 676272 662998
rect 674656 662934 674708 662940
rect 676218 662960 676220 662969
rect 676272 662960 676274 662969
rect 676218 662895 676274 662904
rect 683408 662561 683436 682343
rect 703694 671908 703722 672044
rect 704154 671908 704182 672044
rect 704614 671908 704642 672044
rect 705074 671908 705102 672044
rect 705534 671908 705562 672044
rect 705994 671908 706022 672044
rect 706454 671908 706482 672044
rect 706914 671908 706942 672044
rect 707374 671908 707402 672044
rect 707834 671908 707862 672044
rect 708294 671908 708322 672044
rect 708754 671908 708782 672044
rect 709214 671908 709242 672044
rect 683394 662552 683450 662561
rect 683394 662487 683450 662496
rect 674654 660104 674710 660113
rect 674654 660039 674710 660048
rect 683118 660104 683174 660113
rect 683118 660039 683174 660048
rect 674668 659870 674696 660039
rect 683132 659870 683160 660039
rect 674656 659864 674708 659870
rect 674656 659806 674708 659812
rect 683120 659864 683172 659870
rect 683120 659806 683172 659812
rect 675114 655616 675170 655625
rect 675114 655551 675170 655560
rect 675128 653698 675156 655551
rect 675128 653670 675418 653698
rect 675404 652905 675432 653140
rect 675390 652896 675446 652905
rect 675390 652831 675446 652840
rect 675312 652582 675432 652610
rect 675114 652488 675170 652497
rect 675312 652474 675340 652582
rect 675170 652446 675340 652474
rect 675404 652460 675432 652582
rect 675114 652423 675170 652432
rect 675036 651834 675418 651862
rect 675036 649994 675064 651834
rect 675206 650176 675262 650185
rect 675206 650111 675262 650120
rect 674300 649966 674420 649994
rect 674484 649966 674604 649994
rect 674116 640306 674236 640334
rect 674116 636698 674144 640306
rect 674392 636886 674420 649966
rect 674380 636880 674432 636886
rect 674380 636822 674432 636828
rect 674288 636744 674340 636750
rect 674116 636692 674288 636698
rect 674116 636686 674340 636692
rect 674116 636670 674328 636686
rect 674286 635488 674342 635497
rect 674286 635423 674342 635432
rect 673920 627700 673972 627706
rect 673920 627642 673972 627648
rect 674300 626278 674328 635423
rect 674288 626272 674340 626278
rect 674288 626214 674340 626220
rect 674288 626068 674340 626074
rect 674288 626010 674340 626016
rect 674300 625954 674328 626010
rect 674024 625926 674328 625954
rect 674024 625666 674052 625926
rect 674012 625660 674064 625666
rect 674012 625602 674064 625608
rect 674288 625660 674340 625666
rect 674288 625602 674340 625608
rect 674300 625546 674328 625602
rect 674024 625518 674328 625546
rect 674024 625394 674052 625518
rect 674012 625388 674064 625394
rect 674012 625330 674064 625336
rect 674024 625258 674328 625274
rect 674012 625252 674340 625258
rect 674064 625246 674288 625252
rect 674012 625194 674064 625200
rect 674288 625194 674340 625200
rect 674024 625122 674328 625138
rect 674012 625116 674340 625122
rect 674064 625110 674288 625116
rect 674012 625058 674064 625064
rect 674288 625058 674340 625064
rect 674012 624640 674064 624646
rect 674064 624588 674328 624594
rect 674012 624582 674328 624588
rect 674024 624566 674328 624582
rect 674300 624510 674328 624566
rect 674288 624504 674340 624510
rect 674288 624446 674340 624452
rect 674288 624368 674340 624374
rect 674024 624316 674288 624322
rect 674024 624310 674340 624316
rect 674024 624306 674328 624310
rect 674012 624300 674328 624306
rect 674064 624294 674328 624300
rect 674012 624242 674064 624248
rect 674010 623928 674066 623937
rect 674010 623863 674012 623872
rect 674064 623863 674066 623872
rect 674012 623834 674064 623840
rect 674012 623688 674064 623694
rect 674064 623636 674328 623642
rect 674012 623630 674328 623636
rect 674024 623626 674328 623630
rect 674024 623620 674340 623626
rect 674024 623614 674288 623620
rect 674288 623562 674340 623568
rect 674010 623112 674066 623121
rect 674010 623047 674012 623056
rect 674064 623047 674066 623056
rect 674012 623018 674064 623024
rect 674012 622872 674064 622878
rect 674288 622872 674340 622878
rect 674064 622820 674288 622826
rect 674012 622814 674340 622820
rect 674024 622798 674328 622814
rect 674010 622296 674066 622305
rect 674010 622231 674012 622240
rect 674064 622231 674066 622240
rect 674012 622202 674064 622208
rect 674288 621240 674340 621246
rect 674024 621188 674288 621194
rect 674024 621182 674340 621188
rect 674024 621178 674328 621182
rect 674012 621172 674328 621178
rect 674064 621166 674328 621172
rect 674012 621114 674064 621120
rect 674576 621014 674604 649966
rect 674944 649966 675064 649994
rect 674746 643648 674802 643657
rect 674746 643583 674802 643592
rect 674760 640334 674788 643583
rect 674484 620986 674604 621014
rect 674668 640306 674788 640334
rect 674012 620832 674064 620838
rect 674288 620832 674340 620838
rect 674064 620780 674288 620786
rect 674012 620774 674340 620780
rect 674024 620758 674328 620774
rect 674288 619812 674340 619818
rect 674288 619754 674340 619760
rect 674012 619744 674064 619750
rect 674300 619698 674328 619754
rect 674064 619692 674328 619698
rect 674012 619686 674328 619692
rect 674024 619670 674328 619686
rect 674012 619336 674064 619342
rect 674064 619284 674328 619290
rect 674012 619278 674328 619284
rect 674024 619262 674328 619278
rect 674300 619206 674328 619262
rect 674288 619200 674340 619206
rect 674288 619142 674340 619148
rect 674288 618384 674340 618390
rect 674024 618332 674288 618338
rect 674024 618326 674340 618332
rect 674024 618322 674328 618326
rect 674012 618316 674328 618322
rect 674064 618310 674328 618316
rect 674012 618258 674064 618264
rect 674484 618254 674512 620986
rect 674472 618248 674524 618254
rect 674472 618190 674524 618196
rect 674012 618112 674064 618118
rect 674064 618060 674328 618066
rect 674012 618054 674328 618060
rect 674024 618038 674328 618054
rect 674300 617982 674328 618038
rect 674288 617976 674340 617982
rect 674288 617918 674340 617924
rect 674012 616752 674064 616758
rect 674064 616700 674328 616706
rect 674012 616694 674328 616700
rect 674024 616690 674328 616694
rect 674024 616684 674340 616690
rect 674024 616678 674288 616684
rect 674288 616626 674340 616632
rect 674012 615664 674064 615670
rect 674064 615612 674328 615618
rect 674012 615606 674328 615612
rect 674024 615590 674328 615606
rect 674300 615534 674328 615590
rect 674288 615528 674340 615534
rect 674288 615470 674340 615476
rect 674010 614952 674066 614961
rect 674010 614887 674012 614896
rect 674064 614887 674066 614896
rect 674012 614858 674064 614864
rect 673564 613414 673776 613442
rect 673564 588577 673592 613414
rect 673736 613352 673788 613358
rect 673736 613294 673788 613300
rect 673748 603809 673776 613294
rect 674012 611380 674064 611386
rect 674012 611322 674064 611328
rect 674288 611380 674340 611386
rect 674288 611322 674340 611328
rect 674024 611266 674052 611322
rect 674300 611266 674328 611322
rect 674024 611238 674328 611266
rect 673734 603800 673790 603809
rect 673734 603735 673790 603744
rect 674470 603800 674526 603809
rect 674470 603735 674526 603744
rect 673734 599856 673790 599865
rect 673734 599791 673790 599800
rect 673550 588568 673606 588577
rect 673550 588503 673606 588512
rect 673550 580680 673606 580689
rect 673550 580615 673606 580624
rect 673564 579698 673592 580615
rect 673552 579692 673604 579698
rect 673552 579634 673604 579640
rect 673552 574592 673604 574598
rect 673550 574560 673552 574569
rect 673604 574560 673606 574569
rect 673550 574495 673606 574504
rect 673552 574320 673604 574326
rect 673552 574262 673604 574268
rect 673564 574161 673592 574262
rect 673550 574152 673606 574161
rect 673550 574087 673606 574096
rect 673550 569664 673606 569673
rect 673550 569599 673552 569608
rect 673604 569599 673606 569608
rect 673552 569570 673604 569576
rect 673552 565888 673604 565894
rect 673550 565856 673552 565865
rect 673604 565856 673606 565865
rect 673550 565791 673606 565800
rect 673550 559056 673606 559065
rect 673550 558991 673606 559000
rect 673564 484809 673592 558991
rect 673748 536353 673776 599791
rect 674102 599176 674158 599185
rect 674102 599111 674158 599120
rect 674286 599176 674342 599185
rect 674286 599111 674342 599120
rect 674116 598934 674144 599111
rect 674024 598906 674144 598934
rect 674024 598097 674052 598906
rect 674010 598088 674066 598097
rect 674010 598023 674066 598032
rect 674102 597408 674158 597417
rect 674102 597343 674158 597352
rect 673918 581088 673974 581097
rect 673918 581023 673920 581032
rect 673972 581023 673974 581032
rect 673920 580994 673972 581000
rect 673920 580304 673972 580310
rect 673918 580272 673920 580281
rect 673972 580272 673974 580281
rect 673918 580207 673974 580216
rect 673920 579896 673972 579902
rect 673918 579864 673920 579873
rect 673972 579864 673974 579873
rect 673918 579799 673974 579808
rect 673918 579456 673974 579465
rect 673918 579391 673920 579400
rect 673972 579391 673974 579400
rect 673920 579362 673972 579368
rect 673920 579080 673972 579086
rect 673918 579048 673920 579057
rect 673972 579048 673974 579057
rect 673918 578983 673974 578992
rect 673918 578640 673974 578649
rect 673918 578575 673920 578584
rect 673972 578575 673974 578584
rect 673920 578546 673972 578552
rect 673918 578232 673974 578241
rect 673918 578167 673920 578176
rect 673972 578167 673974 578176
rect 673920 578138 673972 578144
rect 673918 577824 673974 577833
rect 673918 577759 673920 577768
rect 673972 577759 673974 577768
rect 673920 577730 673972 577736
rect 673920 577448 673972 577454
rect 673918 577416 673920 577425
rect 673972 577416 673974 577425
rect 673918 577351 673974 577360
rect 673918 577008 673974 577017
rect 673918 576943 673920 576952
rect 673972 576943 673974 576952
rect 673920 576914 673972 576920
rect 673920 575408 673972 575414
rect 673918 575376 673920 575385
rect 673972 575376 673974 575385
rect 673918 575311 673974 575320
rect 673918 574968 673974 574977
rect 673918 574903 673974 574912
rect 673932 574122 673960 574903
rect 673920 574116 673972 574122
rect 673920 574058 673972 574064
rect 673920 573776 673972 573782
rect 673918 573744 673920 573753
rect 673972 573744 673974 573753
rect 673918 573679 673974 573688
rect 673920 572144 673972 572150
rect 673918 572112 673920 572121
rect 673972 572112 673974 572121
rect 673918 572047 673974 572056
rect 673918 570888 673974 570897
rect 673918 570823 673920 570832
rect 673972 570823 673974 570832
rect 673920 570794 673972 570800
rect 673920 570240 673972 570246
rect 673918 570208 673920 570217
rect 673972 570208 673974 570217
rect 673918 570143 673974 570152
rect 674116 569954 674144 597343
rect 674300 582374 674328 599111
rect 674484 598822 674512 603735
rect 674668 598942 674696 640306
rect 674944 631417 674972 649966
rect 675220 647442 675248 650111
rect 675404 649777 675432 650012
rect 675390 649768 675446 649777
rect 675390 649703 675446 649712
rect 675404 649233 675432 649468
rect 675390 649224 675446 649233
rect 675390 649159 675446 649168
rect 675772 648689 675800 648788
rect 675758 648680 675814 648689
rect 675758 648615 675814 648624
rect 675404 647873 675432 648176
rect 675390 647864 675446 647873
rect 675390 647799 675446 647808
rect 675036 647414 675248 647442
rect 675036 637574 675064 647414
rect 675206 647320 675262 647329
rect 675206 647255 675262 647264
rect 675220 645674 675248 647255
rect 675220 645646 675418 645674
rect 675206 645552 675262 645561
rect 675206 645487 675262 645496
rect 675220 643294 675248 645487
rect 675404 644881 675432 645116
rect 675390 644872 675446 644881
rect 675390 644807 675446 644816
rect 675758 644736 675814 644745
rect 675758 644671 675814 644680
rect 675772 644475 675800 644671
rect 675404 643657 675432 643824
rect 675390 643648 675446 643657
rect 675390 643583 675446 643592
rect 675220 643266 675418 643294
rect 675298 643104 675354 643113
rect 675128 643062 675298 643090
rect 675128 641458 675156 643062
rect 675298 643039 675354 643048
rect 675312 642621 675418 642649
rect 675312 641753 675340 642621
rect 675298 641744 675354 641753
rect 675298 641679 675354 641688
rect 675128 641430 675418 641458
rect 675220 640781 675418 640809
rect 675220 637574 675248 640781
rect 675496 639849 675524 640152
rect 675482 639840 675538 639849
rect 675482 639775 675538 639784
rect 675496 638761 675524 638928
rect 675482 638752 675538 638761
rect 675482 638687 675538 638696
rect 675036 637546 675156 637574
rect 675220 637546 675340 637574
rect 675128 635526 675156 637546
rect 675116 635520 675168 635526
rect 675116 635462 675168 635468
rect 674930 631408 674986 631417
rect 675312 631394 675340 637546
rect 675484 637016 675536 637022
rect 675484 636958 675536 636964
rect 683304 637016 683356 637022
rect 683304 636958 683356 636964
rect 675496 636750 675524 636958
rect 675484 636744 675536 636750
rect 675484 636686 675536 636692
rect 682382 636168 682438 636177
rect 682382 636103 682438 636112
rect 675484 635520 675536 635526
rect 675484 635462 675536 635468
rect 674930 631343 674986 631352
rect 675128 631366 675340 631394
rect 674840 626272 674892 626278
rect 674760 626220 674840 626226
rect 674760 626214 674892 626220
rect 674760 626198 674880 626214
rect 674760 620242 674788 626198
rect 675128 621014 675156 631366
rect 675496 627914 675524 635462
rect 675312 627886 675524 627914
rect 675312 621489 675340 627886
rect 676218 626104 676274 626113
rect 676218 626039 676220 626048
rect 676272 626039 676274 626048
rect 676220 626010 676272 626016
rect 676218 625696 676274 625705
rect 676218 625631 676220 625640
rect 676272 625631 676274 625640
rect 676220 625602 676272 625608
rect 676218 625288 676274 625297
rect 676218 625223 676220 625232
rect 676272 625223 676274 625232
rect 676494 625288 676550 625297
rect 676494 625223 676550 625232
rect 676220 625194 676272 625200
rect 676508 625122 676536 625223
rect 676496 625116 676548 625122
rect 676496 625058 676548 625064
rect 676034 624744 676090 624753
rect 676034 624679 676090 624688
rect 676048 624374 676076 624679
rect 676220 624504 676272 624510
rect 676218 624472 676220 624481
rect 676272 624472 676274 624481
rect 676218 624407 676274 624416
rect 676036 624368 676088 624374
rect 676036 624310 676088 624316
rect 676218 623656 676274 623665
rect 676218 623591 676220 623600
rect 676272 623591 676274 623600
rect 676220 623562 676272 623568
rect 676220 622872 676272 622878
rect 676218 622840 676220 622849
rect 676272 622840 676274 622849
rect 676218 622775 676274 622784
rect 682396 622033 682424 636103
rect 682382 622024 682438 622033
rect 682382 621959 682438 621968
rect 675298 621480 675354 621489
rect 675298 621415 675354 621424
rect 676220 621240 676272 621246
rect 676218 621208 676220 621217
rect 676272 621208 676274 621217
rect 676218 621143 676274 621152
rect 675036 620986 675156 621014
rect 674760 620226 674880 620242
rect 674760 620220 674892 620226
rect 674760 620214 674840 620220
rect 674840 620162 674892 620168
rect 675036 611354 675064 620986
rect 676220 620832 676272 620838
rect 676218 620800 676220 620809
rect 676272 620800 676274 620809
rect 676218 620735 676274 620744
rect 683120 620220 683172 620226
rect 683120 620162 683172 620168
rect 676034 619848 676090 619857
rect 676034 619783 676036 619792
rect 676088 619783 676090 619792
rect 676036 619754 676088 619760
rect 676496 619200 676548 619206
rect 676218 619168 676274 619177
rect 676218 619103 676274 619112
rect 676494 619168 676496 619177
rect 676548 619168 676550 619177
rect 676494 619103 676550 619112
rect 676232 618390 676260 619103
rect 676220 618384 676272 618390
rect 676220 618326 676272 618332
rect 676036 618248 676088 618254
rect 676034 618216 676036 618225
rect 676088 618216 676090 618225
rect 676034 618151 676090 618160
rect 676220 617976 676272 617982
rect 676218 617944 676220 617953
rect 676272 617944 676274 617953
rect 676218 617879 676274 617888
rect 683132 617545 683160 620162
rect 683118 617536 683174 617545
rect 683118 617471 683174 617480
rect 683316 617137 683344 636958
rect 683948 636880 684000 636886
rect 683948 636822 684000 636828
rect 683960 620401 683988 636822
rect 703694 626892 703722 627028
rect 704154 626892 704182 627028
rect 704614 626892 704642 627028
rect 705074 626892 705102 627028
rect 705534 626892 705562 627028
rect 705994 626892 706022 627028
rect 706454 626892 706482 627028
rect 706914 626892 706942 627028
rect 707374 626892 707402 627028
rect 707834 626892 707862 627028
rect 708294 626892 708322 627028
rect 708754 626892 708782 627028
rect 709214 626892 709242 627028
rect 683946 620392 684002 620401
rect 683946 620327 684002 620336
rect 683302 617128 683358 617137
rect 683302 617063 683358 617072
rect 676218 616720 676274 616729
rect 676218 616655 676220 616664
rect 676272 616655 676274 616664
rect 676220 616626 676272 616632
rect 683120 615528 683172 615534
rect 683118 615496 683120 615505
rect 683172 615496 683174 615505
rect 683118 615431 683174 615440
rect 674852 611326 675064 611354
rect 675392 611380 675444 611386
rect 674852 607073 674880 611326
rect 675392 611322 675444 611328
rect 675404 608668 675432 611322
rect 675114 608152 675170 608161
rect 675170 608110 675418 608138
rect 675114 608087 675170 608096
rect 675128 607465 675418 607493
rect 675128 607345 675156 607465
rect 675114 607336 675170 607345
rect 675114 607271 675170 607280
rect 674838 607064 674894 607073
rect 674838 606999 674894 607008
rect 674944 606818 675418 606846
rect 674944 599502 674972 606818
rect 675220 604982 675418 605010
rect 675220 603378 675248 604982
rect 675404 604353 675432 604452
rect 675390 604344 675446 604353
rect 675390 604279 675446 604288
rect 675482 604072 675538 604081
rect 675482 604007 675538 604016
rect 675496 603772 675524 604007
rect 675128 603350 675248 603378
rect 674944 599474 675064 599502
rect 674656 598936 674708 598942
rect 674656 598878 674708 598884
rect 674484 598794 674880 598822
rect 674656 598664 674708 598670
rect 674470 598632 674526 598641
rect 674656 598606 674708 598612
rect 674470 598567 674526 598576
rect 674484 582374 674512 598567
rect 674208 582346 674328 582374
rect 674392 582346 674512 582374
rect 674208 572714 674236 582346
rect 674392 572714 674420 582346
rect 674208 572686 674328 572714
rect 674392 572686 674512 572714
rect 674116 569926 674236 569954
rect 674208 565298 674236 569926
rect 674116 565270 674236 565298
rect 673918 565176 673974 565185
rect 673918 565111 673974 565120
rect 673932 560294 673960 565111
rect 673932 560266 674052 560294
rect 674024 554933 674052 560266
rect 674116 558914 674144 565270
rect 674300 565185 674328 572686
rect 674286 565176 674342 565185
rect 674286 565111 674342 565120
rect 674116 558886 674328 558914
rect 674024 554905 674236 554933
rect 674012 554804 674064 554810
rect 674012 554746 674064 554752
rect 674024 554441 674052 554746
rect 674010 554432 674066 554441
rect 674010 554367 674066 554376
rect 674010 553480 674066 553489
rect 674010 553415 674012 553424
rect 674064 553415 674066 553424
rect 674012 553386 674064 553392
rect 674208 553330 674236 554905
rect 674116 553302 674236 553330
rect 673918 551848 673974 551857
rect 673918 551783 673974 551792
rect 673932 540974 673960 551783
rect 674116 549254 674144 553302
rect 674300 549254 674328 558886
rect 674484 550066 674512 572686
rect 674668 571606 674696 598606
rect 674852 592550 674880 598794
rect 674840 592544 674892 592550
rect 674840 592486 674892 592492
rect 675036 592034 675064 599474
rect 675128 596578 675156 603350
rect 675404 602857 675432 603160
rect 675390 602848 675446 602857
rect 675390 602783 675446 602792
rect 675482 600944 675538 600953
rect 675482 600879 675538 600888
rect 675496 600644 675524 600879
rect 675390 600400 675446 600409
rect 675220 600358 675390 600386
rect 675220 598346 675248 600358
rect 675390 600335 675446 600344
rect 675496 599865 675524 600100
rect 675482 599856 675538 599865
rect 675482 599791 675538 599800
rect 675404 599185 675432 599488
rect 675390 599176 675446 599185
rect 675390 599111 675446 599120
rect 675496 598641 675524 598808
rect 675482 598632 675538 598641
rect 675482 598567 675538 598576
rect 675220 598318 675432 598346
rect 675404 598264 675432 598318
rect 675298 598088 675354 598097
rect 675298 598023 675354 598032
rect 675312 596850 675340 598023
rect 675496 597417 675524 597652
rect 675482 597408 675538 597417
rect 675482 597343 675538 597352
rect 675312 596822 675432 596850
rect 675128 596550 675248 596578
rect 675220 596306 675248 596550
rect 675404 596428 675432 596822
rect 674944 592006 675064 592034
rect 675128 596278 675248 596306
rect 674944 586537 674972 592006
rect 674930 586528 674986 586537
rect 674930 586463 674986 586472
rect 675128 586265 675156 596278
rect 675220 595802 675340 595830
rect 675220 593042 675248 595802
rect 675312 595762 675340 595802
rect 675404 595762 675432 595816
rect 675312 595734 675432 595762
rect 675496 594833 675524 595136
rect 675482 594824 675538 594833
rect 675482 594759 675538 594768
rect 675496 593609 675524 593980
rect 675482 593600 675538 593609
rect 675482 593535 675538 593544
rect 675220 593014 675432 593042
rect 675114 586256 675170 586265
rect 675114 586191 675170 586200
rect 675404 582374 675432 593014
rect 677506 592920 677562 592929
rect 677506 592855 677562 592864
rect 675576 588600 675628 588606
rect 675574 588568 675576 588577
rect 675628 588568 675630 588577
rect 675574 588503 675630 588512
rect 675036 582346 675432 582374
rect 674656 571600 674708 571606
rect 674656 571542 674708 571548
rect 674654 570208 674710 570217
rect 674654 570143 674710 570152
rect 674668 569974 674696 570143
rect 674656 569968 674708 569974
rect 675036 569954 675064 582346
rect 677520 573617 677548 592855
rect 678242 592648 678298 592657
rect 678242 592583 678298 592592
rect 678256 576881 678284 592583
rect 683396 592544 683448 592550
rect 683396 592486 683448 592492
rect 678242 576872 678298 576881
rect 678242 576807 678298 576816
rect 677506 573608 677562 573617
rect 677506 573543 677562 573552
rect 683408 573209 683436 592486
rect 684222 591288 684278 591297
rect 684222 591223 684278 591232
rect 684040 588600 684092 588606
rect 684040 588542 684092 588548
rect 683394 573200 683450 573209
rect 683394 573135 683450 573144
rect 684052 571985 684080 588542
rect 684236 576065 684264 591223
rect 703694 581740 703722 581876
rect 704154 581740 704182 581876
rect 704614 581740 704642 581876
rect 705074 581740 705102 581876
rect 705534 581740 705562 581876
rect 705994 581740 706022 581876
rect 706454 581740 706482 581876
rect 706914 581740 706942 581876
rect 707374 581740 707402 581876
rect 707834 581740 707862 581876
rect 708294 581740 708322 581876
rect 708754 581740 708782 581876
rect 709214 581740 709242 581876
rect 684222 576056 684278 576065
rect 684222 575991 684278 576000
rect 684038 571976 684094 571985
rect 684038 571911 684094 571920
rect 676220 571600 676272 571606
rect 676218 571568 676220 571577
rect 676272 571568 676274 571577
rect 676218 571503 676274 571512
rect 683118 570344 683174 570353
rect 683118 570279 683174 570288
rect 683132 569974 683160 570279
rect 674656 569910 674708 569916
rect 674944 569926 675064 569954
rect 683120 569968 683172 569974
rect 674656 558068 674708 558074
rect 674656 558010 674708 558016
rect 674668 553093 674696 558010
rect 674944 555529 674972 569926
rect 683120 569910 683172 569916
rect 675390 565856 675446 565865
rect 675390 565791 675446 565800
rect 675404 563448 675432 565791
rect 675312 562958 675432 562986
rect 675312 562918 675340 562958
rect 675128 562890 675340 562918
rect 675404 562904 675432 562958
rect 675128 562465 675156 562890
rect 675114 562456 675170 562465
rect 675114 562391 675170 562400
rect 675404 562193 675432 562292
rect 675390 562184 675446 562193
rect 675390 562119 675446 562128
rect 675390 561912 675446 561921
rect 675390 561847 675446 561856
rect 675404 561612 675432 561847
rect 675496 559473 675524 559776
rect 675482 559464 675538 559473
rect 675482 559399 675538 559408
rect 675220 559218 675418 559246
rect 675220 559065 675248 559218
rect 675206 559056 675262 559065
rect 675206 558991 675262 559000
rect 675404 558260 675432 558620
rect 675312 558232 675432 558260
rect 675312 558074 675340 558232
rect 675300 558068 675352 558074
rect 675300 558010 675352 558016
rect 675220 557926 675418 557954
rect 674930 555520 674986 555529
rect 674930 555455 674986 555464
rect 675220 555234 675248 557926
rect 675404 555257 675432 555492
rect 674944 555206 675248 555234
rect 675390 555248 675446 555257
rect 674944 554418 674972 555206
rect 675390 555183 675446 555192
rect 675128 554905 675418 554933
rect 675128 554713 675156 554905
rect 675114 554704 675170 554713
rect 675114 554639 675170 554648
rect 674576 553065 674696 553093
rect 674760 554390 674972 554418
rect 675298 554432 675354 554441
rect 674576 551698 674604 553065
rect 674760 551857 674788 554390
rect 675298 554367 675354 554376
rect 675114 553480 675170 553489
rect 675114 553415 675170 553424
rect 674746 551848 674802 551857
rect 674746 551783 674802 551792
rect 674576 551670 674788 551698
rect 674484 550038 674604 550066
rect 674576 549254 674604 550038
rect 674760 549982 674788 551670
rect 675128 551253 675156 553415
rect 675312 553093 675340 554367
rect 675772 554033 675800 554268
rect 675758 554024 675814 554033
rect 675758 553959 675814 553968
rect 675482 553888 675538 553897
rect 675482 553823 675538 553832
rect 675496 553656 675524 553823
rect 675312 553065 675418 553093
rect 675772 552129 675800 552432
rect 675758 552120 675814 552129
rect 675758 552055 675814 552064
rect 675128 551225 675418 551253
rect 675036 550582 675418 550610
rect 674748 549976 674800 549982
rect 674748 549918 674800 549924
rect 674840 549840 674892 549846
rect 674806 549788 674840 549794
rect 674806 549782 674892 549788
rect 674806 549766 674880 549782
rect 674806 549522 674834 549766
rect 674806 549494 674972 549522
rect 674748 549296 674800 549302
rect 674116 549226 674236 549254
rect 674300 549226 674420 549254
rect 674208 548978 674236 549226
rect 674024 548950 674236 548978
rect 674024 543734 674052 548950
rect 674392 547330 674420 549226
rect 674484 549226 674604 549254
rect 674668 549244 674748 549254
rect 674668 549238 674800 549244
rect 674944 549254 674972 549494
rect 675036 549386 675064 550582
rect 675390 550488 675446 550497
rect 675390 550423 675446 550432
rect 675404 550202 675432 550423
rect 675312 550174 675432 550202
rect 675312 550118 675340 550174
rect 675300 550112 675352 550118
rect 675300 550054 675352 550060
rect 675312 549937 675418 549965
rect 675312 549817 675340 549937
rect 675298 549808 675354 549817
rect 675298 549743 675354 549752
rect 675298 549536 675354 549545
rect 675298 549471 675354 549480
rect 675036 549358 675156 549386
rect 674668 549226 674788 549238
rect 674944 549226 675064 549254
rect 674484 548706 674512 549226
rect 674484 548678 674604 548706
rect 674380 547324 674432 547330
rect 674380 547266 674432 547272
rect 674024 543706 674144 543734
rect 674116 540974 674144 543706
rect 673932 540946 674052 540974
rect 674116 540946 674328 540974
rect 674024 536466 674052 540946
rect 674300 537198 674328 540946
rect 674288 537192 674340 537198
rect 674288 537134 674340 537140
rect 673932 536450 674052 536466
rect 673920 536444 674052 536450
rect 673972 536438 674052 536444
rect 673920 536386 673972 536392
rect 673734 536344 673790 536353
rect 673734 536279 673790 536288
rect 674286 536344 674342 536353
rect 674286 536279 674342 536288
rect 673920 536172 673972 536178
rect 673920 536114 673972 536120
rect 673734 536072 673790 536081
rect 673734 536007 673736 536016
rect 673788 536007 673790 536016
rect 673736 535978 673788 535984
rect 673736 535832 673788 535838
rect 673734 535800 673736 535809
rect 673788 535800 673790 535809
rect 673734 535735 673790 535744
rect 673734 535256 673790 535265
rect 673734 535191 673790 535200
rect 673748 534138 673776 535191
rect 673736 534132 673788 534138
rect 673736 534074 673788 534080
rect 673734 530768 673790 530777
rect 673734 530703 673790 530712
rect 673748 530126 673776 530703
rect 673736 530120 673788 530126
rect 673736 530062 673788 530068
rect 673736 529984 673788 529990
rect 673734 529952 673736 529961
rect 673788 529952 673790 529961
rect 673734 529887 673790 529896
rect 673734 529544 673790 529553
rect 673734 529479 673736 529488
rect 673788 529479 673790 529488
rect 673736 529450 673788 529456
rect 673734 529272 673790 529281
rect 673734 529207 673736 529216
rect 673788 529207 673790 529216
rect 673736 529178 673788 529184
rect 673734 528864 673790 528873
rect 673734 528799 673736 528808
rect 673788 528799 673790 528808
rect 673736 528770 673788 528776
rect 673932 524702 673960 536114
rect 674300 535922 674328 536279
rect 674024 535894 674328 535922
rect 674024 528554 674052 535894
rect 674288 534268 674340 534274
rect 674288 534210 674340 534216
rect 674300 533905 674328 534210
rect 674286 533896 674342 533905
rect 674286 533831 674342 533840
rect 674288 532840 674340 532846
rect 674286 532808 674288 532817
rect 674340 532808 674342 532817
rect 674286 532743 674342 532752
rect 674024 528526 674236 528554
rect 674208 527082 674236 528526
rect 674380 527604 674432 527610
rect 674380 527546 674432 527552
rect 674392 527241 674420 527546
rect 674378 527232 674434 527241
rect 674378 527167 674434 527176
rect 674576 527082 674604 548678
rect 674208 527054 674328 527082
rect 674300 526794 674328 527054
rect 674484 527054 674604 527082
rect 674288 526788 674340 526794
rect 674288 526730 674340 526736
rect 674484 526386 674512 527054
rect 674472 526380 674524 526386
rect 674472 526322 674524 526328
rect 673840 524674 673960 524702
rect 673840 518894 673868 524674
rect 674288 524612 674340 524618
rect 674024 524572 674288 524600
rect 674024 524482 674052 524572
rect 674288 524554 674340 524560
rect 674012 524476 674064 524482
rect 674012 524418 674064 524424
rect 673840 518866 673960 518894
rect 673932 499574 673960 518866
rect 673932 499546 674512 499574
rect 673828 491496 673880 491502
rect 674288 491496 674340 491502
rect 673828 491438 673880 491444
rect 674024 491444 674288 491450
rect 674024 491438 674340 491444
rect 673840 491337 673868 491438
rect 674024 491422 674328 491438
rect 674024 491366 674052 491422
rect 674012 491360 674064 491366
rect 673826 491328 673882 491337
rect 674012 491302 674064 491308
rect 673826 491263 673882 491272
rect 674012 490952 674064 490958
rect 674010 490920 674012 490929
rect 674064 490920 674066 490929
rect 674010 490855 674066 490864
rect 674012 490136 674064 490142
rect 674010 490104 674012 490113
rect 674064 490104 674066 490113
rect 674010 490039 674066 490048
rect 674010 489696 674066 489705
rect 674010 489631 674012 489640
rect 674064 489631 674066 489640
rect 674012 489602 674064 489608
rect 674012 489320 674064 489326
rect 674010 489288 674012 489297
rect 674064 489288 674066 489297
rect 674010 489223 674066 489232
rect 674012 488504 674064 488510
rect 674010 488472 674012 488481
rect 674064 488472 674066 488481
rect 674010 488407 674066 488416
rect 674012 486872 674064 486878
rect 674010 486840 674012 486849
rect 674064 486840 674066 486849
rect 674010 486775 674066 486784
rect 674012 486056 674064 486062
rect 674010 486024 674012 486033
rect 674064 486024 674066 486033
rect 674010 485959 674066 485968
rect 674288 485172 674340 485178
rect 674288 485114 674340 485120
rect 674300 485058 674328 485114
rect 674024 485030 674328 485058
rect 673550 484800 673606 484809
rect 673550 484735 673606 484744
rect 674024 484430 674052 485030
rect 674484 484430 674512 499546
rect 674012 484424 674064 484430
rect 674012 484366 674064 484372
rect 674472 484424 674524 484430
rect 674668 484401 674696 549226
rect 674838 548448 674894 548457
rect 674838 548383 674894 548392
rect 674852 543734 674880 548383
rect 675036 544610 675064 549226
rect 675128 546394 675156 549358
rect 675312 546922 675340 549471
rect 675772 548321 675800 548760
rect 675758 548312 675814 548321
rect 675758 548247 675814 548256
rect 677414 547632 677470 547641
rect 677414 547567 677470 547576
rect 675300 546916 675352 546922
rect 675300 546858 675352 546864
rect 675128 546366 675248 546394
rect 675024 544604 675076 544610
rect 675024 544546 675076 544552
rect 674852 543706 674972 543734
rect 674944 503878 674972 543706
rect 675220 541249 675248 546366
rect 675392 544604 675444 544610
rect 675392 544546 675444 544552
rect 675206 541240 675262 541249
rect 675206 541175 675262 541184
rect 675114 539608 675170 539617
rect 675404 539594 675432 544546
rect 675114 539543 675170 539552
rect 675312 539566 675432 539594
rect 674932 503872 674984 503878
rect 674932 503814 674984 503820
rect 675128 503674 675156 539543
rect 675116 503668 675168 503674
rect 675116 503610 675168 503616
rect 675312 503538 675340 539566
rect 675484 537192 675536 537198
rect 675484 537134 675536 537140
rect 675496 533390 675524 537134
rect 676218 534304 676274 534313
rect 676218 534239 676220 534248
rect 676272 534239 676274 534248
rect 676220 534210 676272 534216
rect 676034 533692 676090 533701
rect 676034 533627 676090 533636
rect 675484 533384 675536 533390
rect 675484 533326 675536 533332
rect 676048 532846 676076 533627
rect 676036 532840 676088 532846
rect 676036 532782 676088 532788
rect 676218 528184 676274 528193
rect 676218 528119 676274 528128
rect 676232 527610 676260 528119
rect 676220 527604 676272 527610
rect 676220 527546 676272 527552
rect 676036 526788 676088 526794
rect 676034 526756 676036 526765
rect 676088 526756 676090 526765
rect 676034 526691 676090 526700
rect 676036 526380 676088 526386
rect 676034 526348 676036 526357
rect 676088 526348 676090 526357
rect 676034 526283 676090 526292
rect 675668 520260 675720 520266
rect 675668 520202 675720 520208
rect 675484 520124 675536 520130
rect 675484 520066 675536 520072
rect 675300 503532 675352 503538
rect 675300 503474 675352 503480
rect 674472 484366 674524 484372
rect 674654 484392 674710 484401
rect 674654 484327 674710 484336
rect 674288 482520 674340 482526
rect 674288 482462 674340 482468
rect 674300 482202 674328 482462
rect 674024 482186 674328 482202
rect 674012 482180 674328 482186
rect 674064 482174 674328 482180
rect 674012 482122 674064 482128
rect 674288 482112 674340 482118
rect 674024 482060 674288 482066
rect 674024 482054 674340 482060
rect 674024 482038 674328 482054
rect 674024 481846 674052 482038
rect 674012 481840 674064 481846
rect 674012 481782 674064 481788
rect 674012 480956 674064 480962
rect 674012 480898 674064 480904
rect 674024 480842 674052 480898
rect 674024 480814 674328 480842
rect 674300 480418 674328 480814
rect 674288 480412 674340 480418
rect 674288 480354 674340 480360
rect 673368 475516 673420 475522
rect 673368 475458 673420 475464
rect 674012 475516 674064 475522
rect 674288 475516 674340 475522
rect 674064 475476 674288 475504
rect 674012 475458 674064 475464
rect 674288 475458 674340 475464
rect 674288 456136 674340 456142
rect 673840 456084 674288 456090
rect 673840 456078 674340 456084
rect 673840 456074 674328 456078
rect 673828 456068 674328 456074
rect 673880 456062 674328 456068
rect 673828 456010 673880 456016
rect 672816 455796 672868 455802
rect 672816 455738 672868 455744
rect 673274 455424 673330 455433
rect 673274 455359 673276 455368
rect 673328 455359 673330 455368
rect 673276 455330 673328 455336
rect 673386 455288 673442 455297
rect 673386 455223 673388 455232
rect 673440 455223 673442 455232
rect 673506 455252 673558 455258
rect 673388 455194 673440 455200
rect 673506 455194 673558 455200
rect 673518 455025 673546 455194
rect 673504 455016 673560 455025
rect 673504 454951 673560 454960
rect 673046 454776 673098 454782
rect 673044 454744 673046 454753
rect 674288 454776 674340 454782
rect 673098 454744 673100 454753
rect 673044 454679 673100 454688
rect 674286 454744 674288 454753
rect 674340 454744 674342 454753
rect 674286 454679 674342 454688
rect 675496 454510 675524 520066
rect 675680 454782 675708 520202
rect 676034 491736 676090 491745
rect 676034 491671 676090 491680
rect 676048 491502 676076 491671
rect 676036 491496 676088 491502
rect 676036 491438 676088 491444
rect 676034 488880 676090 488889
rect 676034 488815 676090 488824
rect 676048 485382 676076 488815
rect 676036 485376 676088 485382
rect 676036 485318 676088 485324
rect 677140 485376 677192 485382
rect 677140 485318 677192 485324
rect 676034 485208 676090 485217
rect 676034 485143 676036 485152
rect 676088 485143 676090 485152
rect 676036 485114 676088 485120
rect 675852 484424 675904 484430
rect 675852 484366 675904 484372
rect 675864 483177 675892 484366
rect 676220 484356 676272 484362
rect 676220 484298 676272 484304
rect 676034 483576 676090 483585
rect 676232 483562 676260 484298
rect 676090 483534 676260 483562
rect 676034 483511 676090 483520
rect 675850 483168 675906 483177
rect 675850 483103 675906 483112
rect 676034 482760 676090 482769
rect 676034 482695 676090 482704
rect 676048 482526 676076 482695
rect 677152 482531 677180 485318
rect 677428 484362 677456 547567
rect 683394 547360 683450 547369
rect 683212 547324 683264 547330
rect 683394 547295 683450 547304
rect 683212 547266 683264 547272
rect 681002 547088 681058 547097
rect 681002 547023 681058 547032
rect 679622 546816 679678 546825
rect 679622 546751 679678 546760
rect 679636 530641 679664 546751
rect 681016 531865 681044 547023
rect 682384 546916 682436 546922
rect 682384 546858 682436 546864
rect 681002 531856 681058 531865
rect 681002 531791 681058 531800
rect 682396 531457 682424 546858
rect 682382 531448 682438 531457
rect 682382 531383 682438 531392
rect 679622 530632 679678 530641
rect 679622 530567 679678 530576
rect 683224 528193 683252 547266
rect 683210 528184 683266 528193
rect 683210 528119 683266 528128
rect 683408 527377 683436 547295
rect 703694 536724 703722 536860
rect 704154 536724 704182 536860
rect 704614 536724 704642 536860
rect 705074 536724 705102 536860
rect 705534 536724 705562 536860
rect 705994 536724 706022 536860
rect 706454 536724 706482 536860
rect 706914 536724 706942 536860
rect 707374 536724 707402 536860
rect 707834 536724 707862 536860
rect 708294 536724 708322 536860
rect 708754 536724 708782 536860
rect 709214 536724 709242 536860
rect 683580 533384 683632 533390
rect 683580 533326 683632 533332
rect 683592 527785 683620 533326
rect 683578 527776 683634 527785
rect 683578 527711 683634 527720
rect 683394 527368 683450 527377
rect 683394 527303 683450 527312
rect 678978 525736 679034 525745
rect 678978 525671 679034 525680
rect 678992 520130 679020 525671
rect 683118 524920 683174 524929
rect 683118 524855 683174 524864
rect 683132 524618 683160 524855
rect 683120 524612 683172 524618
rect 683120 524554 683172 524560
rect 680358 524512 680414 524521
rect 680358 524447 680414 524456
rect 680372 520266 680400 524447
rect 680360 520260 680412 520266
rect 680360 520202 680412 520208
rect 678980 520124 679032 520130
rect 678980 520066 679032 520072
rect 678244 503872 678296 503878
rect 678244 503814 678296 503820
rect 678256 487665 678284 503814
rect 683210 503704 683266 503713
rect 679624 503668 679676 503674
rect 683210 503639 683266 503648
rect 679624 503610 679676 503616
rect 678242 487656 678298 487665
rect 678242 487591 678298 487600
rect 679636 487257 679664 503610
rect 681004 503532 681056 503538
rect 681004 503474 681056 503480
rect 679622 487248 679678 487257
rect 679622 487183 679678 487192
rect 681016 486441 681044 503474
rect 681002 486432 681058 486441
rect 681002 486367 681058 486376
rect 683224 485625 683252 503639
rect 703694 492796 703722 492864
rect 704154 492796 704182 492864
rect 704614 492796 704642 492864
rect 705074 492796 705102 492864
rect 705534 492796 705562 492864
rect 705994 492796 706022 492864
rect 706454 492796 706482 492864
rect 706914 492796 706942 492864
rect 707374 492796 707402 492864
rect 707834 492796 707862 492864
rect 708294 492796 708322 492864
rect 708754 492796 708782 492864
rect 709214 492796 709242 492864
rect 683210 485616 683266 485625
rect 683210 485551 683266 485560
rect 677416 484356 677468 484362
rect 677416 484298 677468 484304
rect 676036 482520 676088 482526
rect 676036 482462 676088 482468
rect 677138 482522 677194 482531
rect 677138 482457 677194 482466
rect 676034 482352 676090 482361
rect 676034 482287 676090 482296
rect 676048 482118 676076 482287
rect 676036 482112 676088 482118
rect 676036 482054 676088 482060
rect 680358 481944 680414 481953
rect 680358 481879 680414 481888
rect 675850 480720 675906 480729
rect 675850 480655 675906 480664
rect 675668 454776 675720 454782
rect 675668 454718 675720 454724
rect 674288 454504 674340 454510
rect 672952 454472 673008 454481
rect 672952 454407 672954 454416
rect 673006 454407 673008 454416
rect 674286 454472 674288 454481
rect 675484 454504 675536 454510
rect 674340 454472 674342 454481
rect 675484 454446 675536 454452
rect 674286 454407 674342 454416
rect 672954 454378 673006 454384
rect 675864 454238 675892 480655
rect 676220 475516 676272 475522
rect 676220 475458 676272 475464
rect 676036 475176 676088 475182
rect 676036 475118 676088 475124
rect 672816 454232 672868 454238
rect 672814 454200 672816 454209
rect 674288 454232 674340 454238
rect 672868 454200 672870 454209
rect 672814 454135 672870 454144
rect 674286 454200 674288 454209
rect 675852 454232 675904 454238
rect 674340 454200 674342 454209
rect 675852 454174 675904 454180
rect 674286 454135 674342 454144
rect 676048 453966 676076 475118
rect 676232 456142 676260 475458
rect 680372 475182 680400 481879
rect 683118 481128 683174 481137
rect 683118 481063 683174 481072
rect 683132 480418 683160 481063
rect 683120 480412 683172 480418
rect 683120 480354 683172 480360
rect 680360 475176 680412 475182
rect 680360 475118 680412 475124
rect 676220 456136 676272 456142
rect 676220 456078 676272 456084
rect 674288 453960 674340 453966
rect 674286 453928 674288 453937
rect 676036 453960 676088 453966
rect 674340 453928 674342 453937
rect 676036 453902 676088 453908
rect 674286 453863 674342 453872
rect 703694 404532 703722 404668
rect 704154 404532 704182 404668
rect 704614 404532 704642 404668
rect 705074 404532 705102 404668
rect 705534 404532 705562 404668
rect 705994 404532 706022 404668
rect 706454 404532 706482 404668
rect 706914 404532 706942 404668
rect 707374 404532 707402 404668
rect 707834 404532 707862 404668
rect 708294 404532 708322 404668
rect 708754 404532 708782 404668
rect 709214 404532 709242 404668
rect 676218 403336 676274 403345
rect 674564 403300 674616 403306
rect 676218 403271 676220 403280
rect 674564 403242 674616 403248
rect 676272 403271 676274 403280
rect 676220 403242 676272 403248
rect 673182 402384 673238 402393
rect 673182 402319 673238 402328
rect 672630 402112 672686 402121
rect 672630 402047 672686 402056
rect 672446 401704 672502 401713
rect 672446 401639 672502 401648
rect 672814 399664 672870 399673
rect 672814 399599 672870 399608
rect 672630 393952 672686 393961
rect 672630 393887 672686 393896
rect 671342 392592 671398 392601
rect 671342 392527 671398 392536
rect 668582 391232 668638 391241
rect 668582 391167 668638 391176
rect 667386 358728 667442 358737
rect 667386 358663 667442 358672
rect 667400 328438 667428 358663
rect 667388 328432 667440 328438
rect 667388 328374 667440 328380
rect 667386 313712 667442 313721
rect 667386 313647 667442 313656
rect 667400 302190 667428 313647
rect 667388 302184 667440 302190
rect 667388 302126 667440 302132
rect 667388 282940 667440 282946
rect 667388 282882 667440 282888
rect 667204 278180 667256 278186
rect 667204 278122 667256 278128
rect 665822 268560 665878 268569
rect 665822 268495 665878 268504
rect 664442 248296 664498 248305
rect 664442 248231 664498 248240
rect 663064 232688 663116 232694
rect 663064 232630 663116 232636
rect 662328 231668 662380 231674
rect 662328 231610 662380 231616
rect 659566 230480 659622 230489
rect 659566 230415 659622 230424
rect 652574 228576 652630 228585
rect 652574 228511 652630 228520
rect 652024 227044 652076 227050
rect 652024 226986 652076 226992
rect 656162 226400 656218 226409
rect 656162 226335 656218 226344
rect 653402 225312 653458 225321
rect 653402 225247 653458 225256
rect 651470 225040 651526 225049
rect 651470 224975 651526 224984
rect 651288 222896 651340 222902
rect 651288 222838 651340 222844
rect 647240 220516 647292 220522
rect 647240 220458 647292 220464
rect 646042 219872 646098 219881
rect 646042 219807 646098 219816
rect 644940 218748 644992 218754
rect 644940 218690 644992 218696
rect 643836 213240 643888 213246
rect 643836 213182 643888 213188
rect 634360 212560 634412 212566
rect 634360 212502 634412 212508
rect 633808 211064 633860 211070
rect 633808 211006 633860 211012
rect 633636 210718 633756 210746
rect 633728 210202 633756 210718
rect 631336 210174 631396 210202
rect 631612 210174 631948 210202
rect 632900 210174 633052 210202
rect 633604 210174 633756 210202
rect 633820 210202 633848 211006
rect 634372 210202 634400 212502
rect 643848 210202 643876 213182
rect 644952 210202 644980 218690
rect 646056 213586 646084 219807
rect 646320 214260 646372 214266
rect 646320 214202 646372 214208
rect 646044 213580 646096 213586
rect 646044 213522 646096 213528
rect 645492 212900 645544 212906
rect 645492 212842 645544 212848
rect 645504 210202 645532 212842
rect 646332 210202 646360 214202
rect 646504 213580 646556 213586
rect 646504 213522 646556 213528
rect 633820 210174 634156 210202
rect 634372 210174 634708 210202
rect 643540 210174 643876 210202
rect 644644 210174 644980 210202
rect 645196 210174 645532 210202
rect 646300 210174 646360 210202
rect 646516 210202 646544 213522
rect 647252 210338 647280 220458
rect 648618 218648 648674 218657
rect 648618 218583 648674 218592
rect 648632 212650 648660 218583
rect 651102 217832 651158 217841
rect 651102 217767 651158 217776
rect 649908 215960 649960 215966
rect 649908 215902 649960 215908
rect 648448 212622 648660 212650
rect 647252 210310 647556 210338
rect 647528 210202 647556 210310
rect 648448 210202 648476 212622
rect 649920 210202 649948 215902
rect 650460 212764 650512 212770
rect 650460 212706 650512 212712
rect 650472 210202 650500 212706
rect 646516 210174 646852 210202
rect 647528 210174 647956 210202
rect 648448 210174 648508 210202
rect 649612 210174 649948 210202
rect 650164 210174 650500 210202
rect 651116 210202 651144 217767
rect 651300 212770 651328 222838
rect 651484 220522 651512 224975
rect 651930 221640 651986 221649
rect 651930 221575 651986 221584
rect 651472 220516 651524 220522
rect 651472 220458 651524 220464
rect 651944 212906 651972 221575
rect 653220 214464 653272 214470
rect 653220 214406 653272 214412
rect 652116 213580 652168 213586
rect 652116 213522 652168 213528
rect 651932 212900 651984 212906
rect 651932 212842 651984 212848
rect 651288 212764 651340 212770
rect 651288 212706 651340 212712
rect 652128 210202 652156 213522
rect 653232 210202 653260 214406
rect 653416 214266 653444 225247
rect 654322 221096 654378 221105
rect 654322 221031 654378 221040
rect 654138 220416 654194 220425
rect 654138 220351 654194 220360
rect 653770 217560 653826 217569
rect 653770 217495 653826 217504
rect 653404 214260 653456 214266
rect 653404 214202 653456 214208
rect 653784 210202 653812 217495
rect 654152 213042 654180 220351
rect 654336 213586 654364 221031
rect 656176 218754 656204 226335
rect 657542 223680 657598 223689
rect 657542 223615 657598 223624
rect 656806 218920 656862 218929
rect 656806 218855 656862 218864
rect 656164 218748 656216 218754
rect 656164 218690 656216 218696
rect 656530 215928 656586 215937
rect 656530 215863 656586 215872
rect 654324 213580 654376 213586
rect 654324 213522 654376 213528
rect 654600 213172 654652 213178
rect 654600 213114 654652 213120
rect 654140 213036 654192 213042
rect 654140 212978 654192 212984
rect 654612 210202 654640 213114
rect 654784 213036 654836 213042
rect 654784 212978 654836 212984
rect 651116 210174 651268 210202
rect 651820 210174 652156 210202
rect 652924 210174 653260 210202
rect 653476 210174 653812 210202
rect 654580 210174 654640 210202
rect 654796 210202 654824 212978
rect 656544 210202 656572 215863
rect 656820 210202 656848 218855
rect 657556 213178 657584 223615
rect 658186 222320 658242 222329
rect 658186 222255 658242 222264
rect 657544 213172 657596 213178
rect 657544 213114 657596 213120
rect 658200 210202 658228 222255
rect 659382 213752 659438 213761
rect 659382 213687 659438 213696
rect 658740 212764 658792 212770
rect 658740 212706 658792 212712
rect 658752 210202 658780 212706
rect 654796 210174 655132 210202
rect 656236 210174 656572 210202
rect 656788 210174 656848 210202
rect 657892 210174 658228 210202
rect 658444 210174 658780 210202
rect 659396 210202 659424 213687
rect 659580 212770 659608 230415
rect 660948 229764 661000 229770
rect 660948 229706 661000 229712
rect 660210 224088 660266 224097
rect 660210 224023 660266 224032
rect 660224 214470 660252 224023
rect 660394 215112 660450 215121
rect 660394 215047 660450 215056
rect 660212 214464 660264 214470
rect 660212 214406 660264 214412
rect 659568 212764 659620 212770
rect 659568 212706 659620 212712
rect 660408 210202 660436 215047
rect 660960 210202 660988 229706
rect 661498 213480 661554 213489
rect 661498 213415 661554 213424
rect 661512 210202 661540 213415
rect 662052 213036 662104 213042
rect 662052 212978 662104 212984
rect 662064 210202 662092 212978
rect 662340 210202 662368 231610
rect 664996 231532 665048 231538
rect 664996 231474 665048 231480
rect 663706 229392 663762 229401
rect 663706 229327 663762 229336
rect 663062 225720 663118 225729
rect 663062 225655 663118 225664
rect 663076 215966 663104 225655
rect 663064 215960 663116 215966
rect 663064 215902 663116 215908
rect 663720 215294 663748 229327
rect 665008 229094 665036 231474
rect 667204 231260 667256 231266
rect 667204 231202 667256 231208
rect 665824 230648 665876 230654
rect 665824 230590 665876 230596
rect 665178 230208 665234 230217
rect 665178 230143 665234 230152
rect 665192 229094 665220 230143
rect 665008 229066 665128 229094
rect 665192 229066 665312 229094
rect 664904 227792 664956 227798
rect 664904 227734 664956 227740
rect 664258 217832 664314 217841
rect 664258 217767 664314 217776
rect 664272 217297 664300 217767
rect 664258 217288 664314 217297
rect 664258 217223 664314 217232
rect 664718 216472 664774 216481
rect 664718 216407 664774 216416
rect 663628 215266 663748 215294
rect 663432 214464 663484 214470
rect 663432 214406 663484 214412
rect 663156 213920 663208 213926
rect 663156 213862 663208 213868
rect 663168 210202 663196 213862
rect 663444 210202 663472 214406
rect 663628 213926 663656 215266
rect 663616 213920 663668 213926
rect 663616 213862 663668 213868
rect 664732 213042 664760 216407
rect 664720 213036 664772 213042
rect 664720 212978 664772 212984
rect 664260 212764 664312 212770
rect 664260 212706 664312 212712
rect 664272 210202 664300 212706
rect 664916 210202 664944 227734
rect 665100 212770 665128 229066
rect 665284 227798 665312 229066
rect 665272 227792 665324 227798
rect 665272 227734 665324 227740
rect 665836 214470 665864 230590
rect 666468 225072 666520 225078
rect 666468 225014 666520 225020
rect 666480 222902 666508 225014
rect 667020 224392 667072 224398
rect 666834 224360 666890 224369
rect 667020 224334 667072 224340
rect 666834 224295 666890 224304
rect 666848 224058 666876 224295
rect 667032 224097 667060 224334
rect 667018 224088 667074 224097
rect 666836 224052 666888 224058
rect 667018 224023 667074 224032
rect 666836 223994 666888 224000
rect 667020 223780 667072 223786
rect 667020 223722 667072 223728
rect 666468 222896 666520 222902
rect 666468 222838 666520 222844
rect 666006 222728 666062 222737
rect 666006 222663 666062 222672
rect 665824 214464 665876 214470
rect 665824 214406 665876 214412
rect 666020 213382 666048 222663
rect 667032 220425 667060 223722
rect 667018 220416 667074 220425
rect 667018 220351 667074 220360
rect 667018 219464 667074 219473
rect 667018 219399 667074 219408
rect 666834 216744 666890 216753
rect 666834 216679 666890 216688
rect 666650 215656 666706 215665
rect 666650 215591 666706 215600
rect 666008 213376 666060 213382
rect 666008 213318 666060 213324
rect 665088 212764 665140 212770
rect 665088 212706 665140 212712
rect 659396 210174 659548 210202
rect 660100 210174 660436 210202
rect 660652 210174 660988 210202
rect 661204 210174 661540 210202
rect 661756 210174 662092 210202
rect 662308 210174 662368 210202
rect 662860 210174 663196 210202
rect 663412 210174 663472 210202
rect 663964 210174 664300 210202
rect 664516 210174 664944 210202
rect 582288 209840 582340 209846
rect 582288 209782 582340 209788
rect 581644 208616 581696 208622
rect 581644 208558 581696 208564
rect 580908 206916 580960 206922
rect 580908 206858 580960 206864
rect 581000 205828 581052 205834
rect 581000 205770 581052 205776
rect 579712 204264 579764 204270
rect 579712 204206 579764 204212
rect 578330 203280 578386 203289
rect 578330 203215 578386 203224
rect 578344 202910 578372 203215
rect 578332 202904 578384 202910
rect 578332 202846 578384 202852
rect 580264 202904 580316 202910
rect 580264 202846 580316 202852
rect 578790 200832 578846 200841
rect 578790 200767 578846 200776
rect 578804 200190 578832 200767
rect 578792 200184 578844 200190
rect 578792 200126 578844 200132
rect 580276 200054 580304 202846
rect 581012 202842 581040 205770
rect 581000 202836 581052 202842
rect 581000 202778 581052 202784
rect 580264 200048 580316 200054
rect 580264 199990 580316 199996
rect 579526 198928 579582 198937
rect 579526 198863 579582 198872
rect 579540 198762 579568 198863
rect 579528 198756 579580 198762
rect 579528 198698 579580 198704
rect 578514 196480 578570 196489
rect 578514 196415 578570 196424
rect 578528 196042 578556 196415
rect 578516 196036 578568 196042
rect 578516 195978 578568 195984
rect 579526 194984 579582 194993
rect 579526 194919 579582 194928
rect 579540 194614 579568 194919
rect 579528 194608 579580 194614
rect 579528 194550 579580 194556
rect 579526 192264 579582 192273
rect 579526 192199 579582 192208
rect 579540 191894 579568 192199
rect 579528 191888 579580 191894
rect 579528 191830 579580 191836
rect 579526 190768 579582 190777
rect 579526 190703 579582 190712
rect 579540 190534 579568 190703
rect 579528 190528 579580 190534
rect 579528 190470 579580 190476
rect 579526 188048 579582 188057
rect 579526 187983 579582 187992
rect 579540 187746 579568 187983
rect 579528 187740 579580 187746
rect 579528 187682 579580 187688
rect 579528 186312 579580 186318
rect 579526 186280 579528 186289
rect 579580 186280 579582 186289
rect 579526 186215 579582 186224
rect 579528 184884 579580 184890
rect 579528 184826 579580 184832
rect 579540 184385 579568 184826
rect 579526 184376 579582 184385
rect 579526 184311 579582 184320
rect 579528 182164 579580 182170
rect 579528 182106 579580 182112
rect 579540 181937 579568 182106
rect 579526 181928 579582 181937
rect 579526 181863 579582 181872
rect 578792 180804 578844 180810
rect 578792 180746 578844 180752
rect 578804 180169 578832 180746
rect 578790 180160 578846 180169
rect 578790 180095 578846 180104
rect 578792 178084 578844 178090
rect 578792 178026 578844 178032
rect 578804 175137 578832 178026
rect 579528 177948 579580 177954
rect 579528 177890 579580 177896
rect 579540 177721 579568 177890
rect 579526 177712 579582 177721
rect 579526 177647 579582 177656
rect 579988 175296 580040 175302
rect 579988 175238 580040 175244
rect 578790 175128 578846 175137
rect 578790 175063 578846 175072
rect 578424 174548 578476 174554
rect 578424 174490 578476 174496
rect 578436 173505 578464 174490
rect 578422 173496 578478 173505
rect 578422 173431 578478 173440
rect 580000 172922 580028 175238
rect 578240 172916 578292 172922
rect 578240 172858 578292 172864
rect 579988 172916 580040 172922
rect 579988 172858 580040 172864
rect 578252 171057 578280 172858
rect 580908 172576 580960 172582
rect 580908 172518 580960 172524
rect 580264 171148 580316 171154
rect 580264 171090 580316 171096
rect 578238 171048 578294 171057
rect 578238 170983 578294 170992
rect 578700 169788 578752 169794
rect 578700 169730 578752 169736
rect 578712 169289 578740 169730
rect 578698 169280 578754 169289
rect 578698 169215 578754 169224
rect 580276 167346 580304 171090
rect 580920 169794 580948 172518
rect 580908 169788 580960 169794
rect 580908 169730 580960 169736
rect 578240 167340 578292 167346
rect 578240 167282 578292 167288
rect 580264 167340 580316 167346
rect 580264 167282 580316 167288
rect 578252 166977 578280 167282
rect 579988 167068 580040 167074
rect 579988 167010 580040 167016
rect 578238 166968 578294 166977
rect 578238 166903 578294 166912
rect 579528 166320 579580 166326
rect 579528 166262 579580 166268
rect 579344 165232 579396 165238
rect 579344 165174 579396 165180
rect 578240 163668 578292 163674
rect 578240 163610 578292 163616
rect 578252 159905 578280 163610
rect 579356 162761 579384 165174
rect 579540 164529 579568 166262
rect 579526 164520 579582 164529
rect 579526 164455 579582 164464
rect 580000 163674 580028 167010
rect 579988 163668 580040 163674
rect 579988 163610 580040 163616
rect 580908 162920 580960 162926
rect 580908 162862 580960 162868
rect 579342 162752 579398 162761
rect 578424 162716 578476 162722
rect 579342 162687 579398 162696
rect 578424 162658 578476 162664
rect 578238 159896 578294 159905
rect 578238 159831 578294 159840
rect 578436 158409 578464 162658
rect 580540 161492 580592 161498
rect 580540 161434 580592 161440
rect 578884 158772 578936 158778
rect 578884 158714 578936 158720
rect 578422 158400 578478 158409
rect 578422 158335 578478 158344
rect 578896 155961 578924 158714
rect 578882 155952 578938 155961
rect 578882 155887 578938 155896
rect 580552 154834 580580 161434
rect 580724 160132 580776 160138
rect 580724 160074 580776 160080
rect 578332 154828 578384 154834
rect 578332 154770 578384 154776
rect 580540 154828 580592 154834
rect 580540 154770 580592 154776
rect 578344 153649 578372 154770
rect 578330 153640 578386 153649
rect 578330 153575 578386 153584
rect 580736 152794 580764 160074
rect 580920 158778 580948 162862
rect 580908 158772 580960 158778
rect 580908 158714 580960 158720
rect 578240 152788 578292 152794
rect 578240 152730 578292 152736
rect 580724 152788 580776 152794
rect 580724 152730 580776 152736
rect 578252 151745 578280 152730
rect 580264 151836 580316 151842
rect 580264 151778 580316 151784
rect 578238 151736 578294 151745
rect 578238 151671 578294 151680
rect 578884 150612 578936 150618
rect 578884 150554 578936 150560
rect 578896 149705 578924 150554
rect 578882 149696 578938 149705
rect 578882 149631 578938 149640
rect 579528 148368 579580 148374
rect 579528 148310 579580 148316
rect 579540 147529 579568 148310
rect 579526 147520 579582 147529
rect 579526 147455 579582 147464
rect 578884 146328 578936 146334
rect 578884 146270 578936 146276
rect 578608 140752 578660 140758
rect 578608 140694 578660 140700
rect 578620 140593 578648 140694
rect 578606 140584 578662 140593
rect 578606 140519 578662 140528
rect 578608 139324 578660 139330
rect 578608 139266 578660 139272
rect 578620 138825 578648 139266
rect 578606 138816 578662 138825
rect 578606 138751 578662 138760
rect 578896 136649 578924 146270
rect 579252 144696 579304 144702
rect 579250 144664 579252 144673
rect 579304 144664 579306 144673
rect 579250 144599 579306 144608
rect 579528 143472 579580 143478
rect 579528 143414 579580 143420
rect 579540 143041 579568 143414
rect 579526 143032 579582 143041
rect 579526 142967 579582 142976
rect 580276 140758 580304 151778
rect 580448 140820 580500 140826
rect 580448 140762 580500 140768
rect 580264 140752 580316 140758
rect 580264 140694 580316 140700
rect 579528 138712 579580 138718
rect 579528 138654 579580 138660
rect 579068 137352 579120 137358
rect 579068 137294 579120 137300
rect 578882 136640 578938 136649
rect 578882 136575 578938 136584
rect 579080 132297 579108 137294
rect 579540 134473 579568 138654
rect 580264 134564 580316 134570
rect 580264 134506 580316 134512
rect 579526 134464 579582 134473
rect 579526 134399 579582 134408
rect 579066 132288 579122 132297
rect 579066 132223 579122 132232
rect 578884 131164 578936 131170
rect 578884 131106 578936 131112
rect 578896 129713 578924 131106
rect 578882 129704 578938 129713
rect 578882 129639 578938 129648
rect 579528 129056 579580 129062
rect 579528 128998 579580 129004
rect 579540 127945 579568 128998
rect 579526 127936 579582 127945
rect 579526 127871 579582 127880
rect 578332 125656 578384 125662
rect 578332 125598 578384 125604
rect 578344 125361 578372 125598
rect 578330 125352 578386 125361
rect 578330 125287 578386 125296
rect 579068 124908 579120 124914
rect 579068 124850 579120 124856
rect 578700 124160 578752 124166
rect 578700 124102 578752 124108
rect 578712 123593 578740 124102
rect 578698 123584 578754 123593
rect 578698 123519 578754 123528
rect 578884 122188 578936 122194
rect 578884 122130 578936 122136
rect 578896 121417 578924 122130
rect 578882 121408 578938 121417
rect 578882 121343 578938 121352
rect 578516 118584 578568 118590
rect 578516 118526 578568 118532
rect 578528 118425 578556 118526
rect 578514 118416 578570 118425
rect 578514 118351 578570 118360
rect 578332 108996 578384 109002
rect 578332 108938 578384 108944
rect 578344 108361 578372 108938
rect 578330 108352 578386 108361
rect 578330 108287 578386 108296
rect 579080 105913 579108 124850
rect 580276 118590 580304 134506
rect 580460 125662 580488 140762
rect 580448 125656 580500 125662
rect 580448 125598 580500 125604
rect 580632 122052 580684 122058
rect 580632 121994 580684 122000
rect 580264 118584 580316 118590
rect 580264 118526 580316 118532
rect 579528 116952 579580 116958
rect 579526 116920 579528 116929
rect 579580 116920 579582 116929
rect 579526 116855 579582 116864
rect 579252 114504 579304 114510
rect 579250 114472 579252 114481
rect 579304 114472 579306 114481
rect 579250 114407 579306 114416
rect 579528 112872 579580 112878
rect 579528 112814 579580 112820
rect 579540 112577 579568 112814
rect 579526 112568 579582 112577
rect 579526 112503 579582 112512
rect 579344 110288 579396 110294
rect 579344 110230 579396 110236
rect 579356 110129 579384 110230
rect 579342 110120 579398 110129
rect 579342 110055 579398 110064
rect 580448 109132 580500 109138
rect 580448 109074 580500 109080
rect 580264 106344 580316 106350
rect 580264 106286 580316 106292
rect 579066 105904 579122 105913
rect 579066 105839 579122 105848
rect 579344 105664 579396 105670
rect 579344 105606 579396 105612
rect 578516 103420 578568 103426
rect 578516 103362 578568 103368
rect 578528 103193 578556 103362
rect 578514 103184 578570 103193
rect 578514 103119 578570 103128
rect 579160 102128 579212 102134
rect 579160 102070 579212 102076
rect 579172 101697 579200 102070
rect 579158 101688 579214 101697
rect 579158 101623 579214 101632
rect 578608 100020 578660 100026
rect 578608 99962 578660 99968
rect 577504 99136 577556 99142
rect 577504 99078 577556 99084
rect 578620 97481 578648 99962
rect 578606 97472 578662 97481
rect 578606 97407 578662 97416
rect 578332 95192 578384 95198
rect 578332 95134 578384 95140
rect 578344 95033 578372 95134
rect 578330 95024 578386 95033
rect 578330 94959 578386 94968
rect 579356 93854 579384 105606
rect 579528 99272 579580 99278
rect 579526 99240 579528 99249
rect 579580 99240 579582 99249
rect 579526 99175 579582 99184
rect 579356 93826 579476 93854
rect 579252 93424 579304 93430
rect 579252 93366 579304 93372
rect 579264 93129 579292 93366
rect 579250 93120 579306 93129
rect 579250 93055 579306 93064
rect 578608 91180 578660 91186
rect 578608 91122 578660 91128
rect 578620 90953 578648 91122
rect 578606 90944 578662 90953
rect 578606 90879 578662 90888
rect 579252 88324 579304 88330
rect 579252 88266 579304 88272
rect 579264 88097 579292 88266
rect 579250 88088 579306 88097
rect 579250 88023 579306 88032
rect 578332 86964 578384 86970
rect 578332 86906 578384 86912
rect 578344 86465 578372 86906
rect 578330 86456 578386 86465
rect 578330 86391 578386 86400
rect 579252 84040 579304 84046
rect 579250 84008 579252 84017
rect 579304 84008 579306 84017
rect 579250 83943 579306 83952
rect 578884 82816 578936 82822
rect 578884 82758 578936 82764
rect 578896 82249 578924 82758
rect 578882 82240 578938 82249
rect 578882 82175 578938 82184
rect 579252 82136 579304 82142
rect 579252 82078 579304 82084
rect 578240 78124 578292 78130
rect 578240 78066 578292 78072
rect 578252 77897 578280 78066
rect 578238 77888 578294 77897
rect 578238 77823 578294 77832
rect 579264 75721 579292 82078
rect 579448 80073 579476 93826
rect 579434 80064 579490 80073
rect 579434 79999 579490 80008
rect 580276 78130 580304 106286
rect 580460 86970 580488 109074
rect 580644 109002 580672 121994
rect 581656 114510 581684 208558
rect 582300 205562 582328 209782
rect 632152 209568 632204 209574
rect 632204 209516 632500 209522
rect 632152 209510 632500 209516
rect 632164 209494 632500 209510
rect 589464 208344 589516 208350
rect 589464 208286 589516 208292
rect 589476 208049 589504 208286
rect 589462 208040 589518 208049
rect 589462 207975 589518 207984
rect 589464 206916 589516 206922
rect 589464 206858 589516 206864
rect 589476 206417 589504 206858
rect 589462 206408 589518 206417
rect 589462 206343 589518 206352
rect 582288 205556 582340 205562
rect 582288 205498 582340 205504
rect 589464 205556 589516 205562
rect 589464 205498 589516 205504
rect 589476 204785 589504 205498
rect 589462 204776 589518 204785
rect 589462 204711 589518 204720
rect 589464 204264 589516 204270
rect 589464 204206 589516 204212
rect 589476 203153 589504 204206
rect 589462 203144 589518 203153
rect 589462 203079 589518 203088
rect 589464 202836 589516 202842
rect 589464 202778 589516 202784
rect 589476 201521 589504 202778
rect 589462 201512 589518 201521
rect 589462 201447 589518 201456
rect 590384 200184 590436 200190
rect 590384 200126 590436 200132
rect 589464 200048 589516 200054
rect 589464 199990 589516 199996
rect 589476 199889 589504 199990
rect 589462 199880 589518 199889
rect 589462 199815 589518 199824
rect 589464 198756 589516 198762
rect 589464 198698 589516 198704
rect 589476 196625 589504 198698
rect 590396 198257 590424 200126
rect 666664 198665 666692 215591
rect 666650 198656 666706 198665
rect 666650 198591 666706 198600
rect 666848 198393 666876 216679
rect 666834 198384 666890 198393
rect 666834 198319 666890 198328
rect 590382 198248 590438 198257
rect 590382 198183 590438 198192
rect 589462 196616 589518 196625
rect 589462 196551 589518 196560
rect 589280 196036 589332 196042
rect 589280 195978 589332 195984
rect 589292 194993 589320 195978
rect 589278 194984 589334 194993
rect 589278 194919 589334 194928
rect 589464 194608 589516 194614
rect 589464 194550 589516 194556
rect 589476 193361 589504 194550
rect 589462 193352 589518 193361
rect 589462 193287 589518 193296
rect 589464 191888 589516 191894
rect 589464 191830 589516 191836
rect 589476 191729 589504 191830
rect 589462 191720 589518 191729
rect 589462 191655 589518 191664
rect 590568 190528 590620 190534
rect 590568 190470 590620 190476
rect 590580 190097 590608 190470
rect 590566 190088 590622 190097
rect 590566 190023 590622 190032
rect 589646 188456 589702 188465
rect 589646 188391 589702 188400
rect 589464 187740 589516 187746
rect 589464 187682 589516 187688
rect 589476 186833 589504 187682
rect 589462 186824 589518 186833
rect 589462 186759 589518 186768
rect 589660 186318 589688 188391
rect 589648 186312 589700 186318
rect 589648 186254 589700 186260
rect 589462 185192 589518 185201
rect 589462 185127 589518 185136
rect 589476 184890 589504 185127
rect 589464 184884 589516 184890
rect 589464 184826 589516 184832
rect 589462 183560 589518 183569
rect 589462 183495 589518 183504
rect 589476 182170 589504 183495
rect 589464 182164 589516 182170
rect 589464 182106 589516 182112
rect 590566 181928 590622 181937
rect 590566 181863 590622 181872
rect 590580 180810 590608 181863
rect 590568 180804 590620 180810
rect 590568 180746 590620 180752
rect 589646 180296 589702 180305
rect 589646 180231 589702 180240
rect 589462 178664 589518 178673
rect 589462 178599 589518 178608
rect 589476 178090 589504 178599
rect 589464 178084 589516 178090
rect 589464 178026 589516 178032
rect 589660 177954 589688 180231
rect 589648 177948 589700 177954
rect 589648 177890 589700 177896
rect 589646 177032 589702 177041
rect 589646 176967 589702 176976
rect 589462 175400 589518 175409
rect 589462 175335 589464 175344
rect 589516 175335 589518 175344
rect 589464 175306 589516 175312
rect 589660 174554 589688 176967
rect 667032 175001 667060 219399
rect 667018 174992 667074 175001
rect 667018 174927 667074 174936
rect 589648 174548 589700 174554
rect 589648 174490 589700 174496
rect 589462 173768 589518 173777
rect 589462 173703 589518 173712
rect 589476 172582 589504 173703
rect 589464 172576 589516 172582
rect 589464 172518 589516 172524
rect 589462 172136 589518 172145
rect 589462 172071 589518 172080
rect 589476 171154 589504 172071
rect 589464 171148 589516 171154
rect 589464 171090 589516 171096
rect 589646 170504 589702 170513
rect 589646 170439 589702 170448
rect 589462 168872 589518 168881
rect 589462 168807 589518 168816
rect 589476 168434 589504 168807
rect 582380 168428 582432 168434
rect 582380 168370 582432 168376
rect 589464 168428 589516 168434
rect 589464 168370 589516 168376
rect 582392 165238 582420 168370
rect 589462 167240 589518 167249
rect 589462 167175 589518 167184
rect 589476 167074 589504 167175
rect 589464 167068 589516 167074
rect 589464 167010 589516 167016
rect 589660 166326 589688 170439
rect 589648 166320 589700 166326
rect 589648 166262 589700 166268
rect 589462 165608 589518 165617
rect 589462 165543 589518 165552
rect 582380 165232 582432 165238
rect 582380 165174 582432 165180
rect 589476 164286 589504 165543
rect 582472 164280 582524 164286
rect 582472 164222 582524 164228
rect 589464 164280 589516 164286
rect 589464 164222 589516 164228
rect 582484 162722 582512 164222
rect 589462 163976 589518 163985
rect 589462 163911 589518 163920
rect 589476 162926 589504 163911
rect 589464 162920 589516 162926
rect 589464 162862 589516 162868
rect 582472 162716 582524 162722
rect 582472 162658 582524 162664
rect 589462 162344 589518 162353
rect 589462 162279 589518 162288
rect 589476 161498 589504 162279
rect 589464 161492 589516 161498
rect 589464 161434 589516 161440
rect 589462 160712 589518 160721
rect 589462 160647 589518 160656
rect 589476 160138 589504 160647
rect 589464 160132 589516 160138
rect 589464 160074 589516 160080
rect 589462 159080 589518 159089
rect 589462 159015 589518 159024
rect 589476 158778 589504 159015
rect 585784 158772 585836 158778
rect 585784 158714 585836 158720
rect 589464 158772 589516 158778
rect 589464 158714 589516 158720
rect 584404 154624 584456 154630
rect 584404 154566 584456 154572
rect 583024 153264 583076 153270
rect 583024 153206 583076 153212
rect 583036 143478 583064 153206
rect 584416 144702 584444 154566
rect 585796 150618 585824 158714
rect 589278 157448 589334 157457
rect 587164 157412 587216 157418
rect 589278 157383 589280 157392
rect 587164 157354 587216 157360
rect 589332 157383 589334 157392
rect 589280 157354 589332 157360
rect 585784 150612 585836 150618
rect 585784 150554 585836 150560
rect 585140 149116 585192 149122
rect 585140 149058 585192 149064
rect 585152 146334 585180 149058
rect 587176 148374 587204 157354
rect 589462 155816 589518 155825
rect 589462 155751 589518 155760
rect 589476 154630 589504 155751
rect 589464 154624 589516 154630
rect 589464 154566 589516 154572
rect 589462 154184 589518 154193
rect 589462 154119 589518 154128
rect 589476 153270 589504 154119
rect 589464 153264 589516 153270
rect 589464 153206 589516 153212
rect 589462 152552 589518 152561
rect 589462 152487 589518 152496
rect 589476 151842 589504 152487
rect 589464 151836 589516 151842
rect 589464 151778 589516 151784
rect 590014 150920 590070 150929
rect 590014 150855 590070 150864
rect 589462 149288 589518 149297
rect 589462 149223 589518 149232
rect 589476 149122 589504 149223
rect 589464 149116 589516 149122
rect 589464 149058 589516 149064
rect 587164 148368 587216 148374
rect 587164 148310 587216 148316
rect 588542 147656 588598 147665
rect 588542 147591 588598 147600
rect 585140 146328 585192 146334
rect 585140 146270 585192 146276
rect 584772 144968 584824 144974
rect 584772 144910 584824 144916
rect 584404 144696 584456 144702
rect 584404 144638 584456 144644
rect 583024 143472 583076 143478
rect 583024 143414 583076 143420
rect 583024 139460 583076 139466
rect 583024 139402 583076 139408
rect 581828 131300 581880 131306
rect 581828 131242 581880 131248
rect 581644 114504 581696 114510
rect 581644 114446 581696 114452
rect 581644 110492 581696 110498
rect 581644 110434 581696 110440
rect 580632 108996 580684 109002
rect 580632 108938 580684 108944
rect 580448 86964 580500 86970
rect 580448 86906 580500 86912
rect 581656 84046 581684 110434
rect 581840 110294 581868 131242
rect 583036 124166 583064 139402
rect 584784 137358 584812 144910
rect 585784 143608 585836 143614
rect 585784 143550 585836 143556
rect 584772 137352 584824 137358
rect 584772 137294 584824 137300
rect 584588 136672 584640 136678
rect 584588 136614 584640 136620
rect 583392 129192 583444 129198
rect 583392 129134 583444 129140
rect 583024 124160 583076 124166
rect 583024 124102 583076 124108
rect 583208 120760 583260 120766
rect 583208 120702 583260 120708
rect 583024 113212 583076 113218
rect 583024 113154 583076 113160
rect 581828 110288 581880 110294
rect 581828 110230 581880 110236
rect 582288 107704 582340 107710
rect 582288 107646 582340 107652
rect 582300 105670 582328 107646
rect 582288 105664 582340 105670
rect 582288 105606 582340 105612
rect 581644 84040 581696 84046
rect 581644 83982 581696 83988
rect 583036 82822 583064 113154
rect 583220 99278 583248 120702
rect 583404 116958 583432 129134
rect 584404 122868 584456 122874
rect 584404 122810 584456 122816
rect 583392 116952 583444 116958
rect 583392 116894 583444 116900
rect 584416 102134 584444 122810
rect 584600 122194 584628 136614
rect 585796 131170 585824 143550
rect 587164 142452 587216 142458
rect 587164 142394 587216 142400
rect 585968 132524 586020 132530
rect 585968 132466 586020 132472
rect 585784 131164 585836 131170
rect 585784 131106 585836 131112
rect 584588 122188 584640 122194
rect 584588 122130 584640 122136
rect 585784 116000 585836 116006
rect 585784 115942 585836 115948
rect 584588 115252 584640 115258
rect 584588 115194 584640 115200
rect 584404 102128 584456 102134
rect 584404 102070 584456 102076
rect 584404 100156 584456 100162
rect 584404 100098 584456 100104
rect 583208 99272 583260 99278
rect 583208 99214 583260 99220
rect 583024 82816 583076 82822
rect 583024 82758 583076 82764
rect 583024 79348 583076 79354
rect 583024 79290 583076 79296
rect 580264 78124 580316 78130
rect 580264 78066 580316 78072
rect 580446 77888 580502 77897
rect 580446 77823 580502 77832
rect 579250 75712 579306 75721
rect 579250 75647 579306 75656
rect 578884 75200 578936 75206
rect 578884 75142 578936 75148
rect 578516 71596 578568 71602
rect 578516 71538 578568 71544
rect 578528 71233 578556 71538
rect 578514 71224 578570 71233
rect 578514 71159 578570 71168
rect 578896 60489 578924 75142
rect 579528 73160 579580 73166
rect 579526 73128 579528 73137
rect 579580 73128 579582 73137
rect 579526 73063 579582 73072
rect 579528 66904 579580 66910
rect 579526 66872 579528 66881
rect 579580 66872 579582 66881
rect 579526 66807 579582 66816
rect 579528 64864 579580 64870
rect 579528 64806 579580 64812
rect 579540 64569 579568 64806
rect 579526 64560 579582 64569
rect 579526 64495 579582 64504
rect 579528 62076 579580 62082
rect 579528 62018 579580 62024
rect 579540 61849 579568 62018
rect 579526 61840 579582 61849
rect 579526 61775 579582 61784
rect 578882 60480 578938 60489
rect 578882 60415 578938 60424
rect 578332 60036 578384 60042
rect 578332 59978 578384 59984
rect 576124 58812 576176 58818
rect 576124 58754 576176 58760
rect 574928 57248 574980 57254
rect 574928 57190 574980 57196
rect 574744 56024 574796 56030
rect 574744 55966 574796 55972
rect 574468 55888 574520 55894
rect 574468 55830 574520 55836
rect 574480 54777 574508 55830
rect 574466 54768 574522 54777
rect 574466 54703 574522 54712
rect 574756 53990 574784 55966
rect 574744 53984 574796 53990
rect 574744 53926 574796 53932
rect 574940 53854 574968 57190
rect 576136 54233 576164 58754
rect 577504 58676 577556 58682
rect 577504 58618 577556 58624
rect 577516 55049 577544 58618
rect 578344 56137 578372 59978
rect 579528 57928 579580 57934
rect 579526 57896 579528 57905
rect 579580 57896 579582 57905
rect 579526 57831 579582 57840
rect 578330 56128 578386 56137
rect 578330 56063 578386 56072
rect 577502 55040 577558 55049
rect 577502 54975 577558 54984
rect 576122 54224 576178 54233
rect 576122 54159 576178 54168
rect 580460 54126 580488 77823
rect 583036 54262 583064 79290
rect 584416 71602 584444 100098
rect 584600 95198 584628 115194
rect 584588 95192 584640 95198
rect 584588 95134 584640 95140
rect 585796 91186 585824 115942
rect 585980 112878 586008 132466
rect 587176 129062 587204 142394
rect 588556 138718 588584 147591
rect 589462 146024 589518 146033
rect 589462 145959 589518 145968
rect 589476 144974 589504 145959
rect 589464 144968 589516 144974
rect 589464 144910 589516 144916
rect 589462 144392 589518 144401
rect 589462 144327 589518 144336
rect 589476 143614 589504 144327
rect 589464 143608 589516 143614
rect 589464 143550 589516 143556
rect 589830 142760 589886 142769
rect 589830 142695 589886 142704
rect 589844 142458 589872 142695
rect 589832 142452 589884 142458
rect 589832 142394 589884 142400
rect 590028 142154 590056 150855
rect 589936 142126 590056 142154
rect 589462 141128 589518 141137
rect 589462 141063 589518 141072
rect 589476 140826 589504 141063
rect 589464 140820 589516 140826
rect 589464 140762 589516 140768
rect 589462 139496 589518 139505
rect 589462 139431 589464 139440
rect 589516 139431 589518 139440
rect 589464 139402 589516 139408
rect 589936 139330 589964 142126
rect 589924 139324 589976 139330
rect 589924 139266 589976 139272
rect 588544 138712 588596 138718
rect 588544 138654 588596 138660
rect 589462 137864 589518 137873
rect 589462 137799 589518 137808
rect 589476 136678 589504 137799
rect 589464 136672 589516 136678
rect 589464 136614 589516 136620
rect 589462 136232 589518 136241
rect 589462 136167 589518 136176
rect 589476 134570 589504 136167
rect 590382 134600 590438 134609
rect 589464 134564 589516 134570
rect 590382 134535 590438 134544
rect 589464 134506 589516 134512
rect 589462 132968 589518 132977
rect 589462 132903 589518 132912
rect 589476 132530 589504 132903
rect 589464 132524 589516 132530
rect 589464 132466 589516 132472
rect 589462 131336 589518 131345
rect 589462 131271 589464 131280
rect 589516 131271 589518 131280
rect 589464 131242 589516 131248
rect 588726 129704 588782 129713
rect 588726 129639 588782 129648
rect 587164 129056 587216 129062
rect 587164 128998 587216 129004
rect 587808 127016 587860 127022
rect 587808 126958 587860 126964
rect 587820 124914 587848 126958
rect 587808 124908 587860 124914
rect 587808 124850 587860 124856
rect 587348 121508 587400 121514
rect 587348 121450 587400 121456
rect 585968 112872 586020 112878
rect 585968 112814 586020 112820
rect 586152 112464 586204 112470
rect 586152 112406 586204 112412
rect 586164 93430 586192 112406
rect 587164 104916 587216 104922
rect 587164 104858 587216 104864
rect 586152 93424 586204 93430
rect 586152 93366 586204 93372
rect 585784 91180 585836 91186
rect 585784 91122 585836 91128
rect 587176 82142 587204 104858
rect 587360 100026 587388 121450
rect 588542 103592 588598 103601
rect 588542 103527 588598 103536
rect 587348 100020 587400 100026
rect 587348 99962 587400 99968
rect 587164 82136 587216 82142
rect 587164 82078 587216 82084
rect 587164 76560 587216 76566
rect 587164 76502 587216 76508
rect 584404 71596 584456 71602
rect 584404 71538 584456 71544
rect 587176 62082 587204 76502
rect 588556 73166 588584 103527
rect 588740 103426 588768 129639
rect 590396 129198 590424 134535
rect 590384 129192 590436 129198
rect 590384 129134 590436 129140
rect 589462 128072 589518 128081
rect 589462 128007 589518 128016
rect 589476 127022 589504 128007
rect 589464 127016 589516 127022
rect 589464 126958 589516 126964
rect 590106 126440 590162 126449
rect 590106 126375 590162 126384
rect 589462 123176 589518 123185
rect 589462 123111 589518 123120
rect 589476 122874 589504 123111
rect 589464 122868 589516 122874
rect 589464 122810 589516 122816
rect 590120 122058 590148 126375
rect 590566 124808 590622 124817
rect 590566 124743 590622 124752
rect 590108 122052 590160 122058
rect 590108 121994 590160 122000
rect 589278 121544 589334 121553
rect 589278 121479 589280 121488
rect 589332 121479 589334 121488
rect 589280 121450 589332 121456
rect 590580 120766 590608 124743
rect 667216 122097 667244 231202
rect 667400 132705 667428 282882
rect 667756 281580 667808 281586
rect 667756 281522 667808 281528
rect 667572 280220 667624 280226
rect 667572 280162 667624 280168
rect 667584 133113 667612 280162
rect 667768 134609 667796 281522
rect 668216 234592 668268 234598
rect 668216 234534 668268 234540
rect 668032 234456 668084 234462
rect 668032 234398 668084 234404
rect 668044 177993 668072 234398
rect 668030 177984 668086 177993
rect 668030 177919 668086 177928
rect 668032 174752 668084 174758
rect 668030 174720 668032 174729
rect 668084 174720 668086 174729
rect 668030 174655 668086 174664
rect 667940 173120 667992 173126
rect 667938 173088 667940 173097
rect 667992 173088 667994 173097
rect 667938 173023 667994 173032
rect 668228 169697 668256 234534
rect 668400 231668 668452 231674
rect 668400 231610 668452 231616
rect 668412 230994 668440 231610
rect 668400 230988 668452 230994
rect 668400 230930 668452 230936
rect 668400 230852 668452 230858
rect 668400 230794 668452 230800
rect 668214 169688 668270 169697
rect 668214 169623 668270 169632
rect 668216 168224 668268 168230
rect 668214 168192 668216 168201
rect 668268 168192 668270 168201
rect 668214 168127 668270 168136
rect 667940 164960 667992 164966
rect 667938 164928 667940 164937
rect 667992 164928 667994 164937
rect 667938 164863 667994 164872
rect 668412 163305 668440 230794
rect 668398 163296 668454 163305
rect 668398 163231 668454 163240
rect 668398 160440 668454 160449
rect 668398 160375 668454 160384
rect 668412 158409 668440 160375
rect 668398 158400 668454 158409
rect 668398 158335 668454 158344
rect 668400 149116 668452 149122
rect 668400 149058 668452 149064
rect 668216 140684 668268 140690
rect 668216 140626 668268 140632
rect 668228 140457 668256 140626
rect 668214 140448 668270 140457
rect 668214 140383 668270 140392
rect 668412 138825 668440 149058
rect 668596 143721 668624 391167
rect 670606 347304 670662 347313
rect 670606 347239 670662 347248
rect 669318 344992 669374 345001
rect 669318 344927 669374 344936
rect 669332 338774 669360 344927
rect 669320 338768 669372 338774
rect 669320 338710 669372 338716
rect 669962 302152 670018 302161
rect 669962 302087 670018 302096
rect 668766 300792 668822 300801
rect 668766 300727 668822 300736
rect 668780 229094 668808 300727
rect 669320 235612 669372 235618
rect 669320 235554 669372 235560
rect 668950 234560 669006 234569
rect 668950 234495 669006 234504
rect 668964 230858 668992 234495
rect 669136 231668 669188 231674
rect 669136 231610 669188 231616
rect 669148 231402 669176 231610
rect 669136 231396 669188 231402
rect 669136 231338 669188 231344
rect 668952 230852 669004 230858
rect 668952 230794 669004 230800
rect 668688 229066 668808 229094
rect 668688 224954 668716 229066
rect 669136 227792 669188 227798
rect 669136 227734 669188 227740
rect 668952 227044 669004 227050
rect 668952 226986 669004 226992
rect 668688 224926 668808 224954
rect 668582 143712 668638 143721
rect 668582 143647 668638 143656
rect 668398 138816 668454 138825
rect 668398 138751 668454 138760
rect 668584 138032 668636 138038
rect 668584 137974 668636 137980
rect 667754 134600 667810 134609
rect 667754 134535 667810 134544
rect 667570 133104 667626 133113
rect 667570 133039 667626 133048
rect 667386 132696 667442 132705
rect 667386 132631 667442 132640
rect 667940 130688 667992 130694
rect 667938 130656 667940 130665
rect 667992 130656 667994 130665
rect 667938 130591 667994 130600
rect 668596 129033 668624 137974
rect 668780 133793 668808 224926
rect 668964 220250 668992 226986
rect 668952 220244 669004 220250
rect 668952 220186 669004 220192
rect 669148 220130 669176 227734
rect 668964 220102 669176 220130
rect 668964 148617 668992 220102
rect 669136 220040 669188 220046
rect 669136 219982 669188 219988
rect 669148 150249 669176 219982
rect 669332 160041 669360 235554
rect 669780 235136 669832 235142
rect 669780 235078 669832 235084
rect 669596 233232 669648 233238
rect 669596 233174 669648 233180
rect 669608 173126 669636 233174
rect 669596 173120 669648 173126
rect 669596 173062 669648 173068
rect 669594 172408 669650 172417
rect 669594 172343 669650 172352
rect 669318 160032 669374 160041
rect 669318 159967 669374 159976
rect 669608 150385 669636 172343
rect 669792 164966 669820 235078
rect 669780 164960 669832 164966
rect 669780 164902 669832 164908
rect 669594 150376 669650 150385
rect 669594 150311 669650 150320
rect 669134 150240 669190 150249
rect 669134 150175 669190 150184
rect 668950 148608 669006 148617
rect 668950 148543 669006 148552
rect 668766 133784 668822 133793
rect 668766 133719 668822 133728
rect 669976 130694 670004 302087
rect 670422 260536 670478 260545
rect 670422 260471 670478 260480
rect 670146 258496 670202 258505
rect 670146 258431 670202 258440
rect 670160 138038 670188 258431
rect 670436 240281 670464 260471
rect 670422 240272 670478 240281
rect 670422 240207 670478 240216
rect 670332 234184 670384 234190
rect 670332 234126 670384 234132
rect 670344 174758 670372 234126
rect 670620 224954 670648 347239
rect 671356 263594 671384 392527
rect 672644 376281 672672 393887
rect 672630 376272 672686 376281
rect 672630 376207 672686 376216
rect 672538 357096 672594 357105
rect 672538 357031 672594 357040
rect 672170 352608 672226 352617
rect 672170 352543 672226 352552
rect 671526 348528 671582 348537
rect 671526 348463 671582 348472
rect 671356 263566 671476 263594
rect 671158 259720 671214 259729
rect 671158 259655 671214 259664
rect 670974 250744 671030 250753
rect 670974 250679 671030 250688
rect 670988 248305 671016 250679
rect 670974 248296 671030 248305
rect 670974 248231 671030 248240
rect 671172 245585 671200 259655
rect 671158 245576 671214 245585
rect 671158 245511 671214 245520
rect 671068 235952 671120 235958
rect 671068 235894 671120 235900
rect 670884 235476 670936 235482
rect 670884 235418 670936 235424
rect 670436 224926 670648 224954
rect 670896 224954 670924 235418
rect 670896 224926 671016 224954
rect 670436 215294 670464 224926
rect 670700 224868 670752 224874
rect 670700 224810 670752 224816
rect 670712 224720 670740 224810
rect 670620 224692 670740 224720
rect 670620 217569 670648 224692
rect 670792 224188 670844 224194
rect 670792 224130 670844 224136
rect 670804 223961 670832 224130
rect 670790 223952 670846 223961
rect 670790 223887 670846 223896
rect 670790 223680 670846 223689
rect 670790 223615 670792 223624
rect 670844 223615 670846 223624
rect 670792 223586 670844 223592
rect 670792 223168 670844 223174
rect 670792 223110 670844 223116
rect 670804 222329 670832 223110
rect 670790 222320 670846 222329
rect 670790 222255 670846 222264
rect 670792 222148 670844 222154
rect 670792 222090 670844 222096
rect 670804 218929 670832 222090
rect 670790 218920 670846 218929
rect 670790 218855 670846 218864
rect 670606 217560 670662 217569
rect 670606 217495 670662 217504
rect 670436 215266 670648 215294
rect 670332 174752 670384 174758
rect 670332 174694 670384 174700
rect 670620 171057 670648 215266
rect 670790 214160 670846 214169
rect 670790 214095 670846 214104
rect 670804 197577 670832 214095
rect 670790 197568 670846 197577
rect 670790 197503 670846 197512
rect 670988 180794 671016 224926
rect 671080 215294 671108 235894
rect 671252 235816 671304 235822
rect 671252 235758 671304 235764
rect 671264 234569 671292 235758
rect 671250 234560 671306 234569
rect 671250 234495 671306 234504
rect 671252 226092 671304 226098
rect 671252 226034 671304 226040
rect 671264 225321 671292 226034
rect 671250 225312 671306 225321
rect 671250 225247 671306 225256
rect 671448 224954 671476 263566
rect 671172 224926 671476 224954
rect 671172 220130 671200 224926
rect 671540 224754 671568 348463
rect 672184 333441 672212 352543
rect 672354 349344 672410 349353
rect 672354 349279 672410 349288
rect 672170 333432 672226 333441
rect 672170 333367 672226 333376
rect 672368 332761 672396 349279
rect 672354 332752 672410 332761
rect 672354 332687 672410 332696
rect 672552 312497 672580 357031
rect 672828 355065 672856 399599
rect 672998 394768 673054 394777
rect 672998 394703 673054 394712
rect 673012 381041 673040 394703
rect 672998 381032 673054 381041
rect 672998 380967 673054 380976
rect 673196 357513 673224 402319
rect 673918 401432 673974 401441
rect 673918 401367 673974 401376
rect 673366 400480 673422 400489
rect 673366 400415 673422 400424
rect 673182 357504 673238 357513
rect 673182 357439 673238 357448
rect 673380 355881 673408 400415
rect 673932 364334 673960 401367
rect 674576 396681 674604 403242
rect 676586 402928 676642 402937
rect 676586 402863 676642 402872
rect 674838 402656 674894 402665
rect 674838 402591 674894 402600
rect 674852 402121 674880 402591
rect 674838 402112 674894 402121
rect 674838 402047 674894 402056
rect 676600 400897 676628 402863
rect 676586 400888 676642 400897
rect 676586 400823 676642 400832
rect 676034 399392 676090 399401
rect 676034 399327 676090 399336
rect 676048 398886 676076 399327
rect 674932 398880 674984 398886
rect 674932 398822 674984 398828
rect 676036 398880 676088 398886
rect 676036 398822 676088 398828
rect 674746 397352 674802 397361
rect 674746 397287 674802 397296
rect 674562 396672 674618 396681
rect 674562 396607 674618 396616
rect 674380 396092 674432 396098
rect 674380 396034 674432 396040
rect 674102 395856 674158 395865
rect 674102 395791 674158 395800
rect 674116 379386 674144 395791
rect 674392 395706 674420 396034
rect 674208 395678 674420 395706
rect 674208 393314 674236 395678
rect 674472 394324 674524 394330
rect 674472 394266 674524 394272
rect 674208 393286 674328 393314
rect 674300 383654 674328 393286
rect 674484 383654 674512 394266
rect 674760 393314 674788 397287
rect 674944 395842 674972 398822
rect 679622 398440 679678 398449
rect 679622 398375 679678 398384
rect 676218 398032 676274 398041
rect 676218 397967 676274 397976
rect 676034 396128 676090 396137
rect 676034 396063 676036 396072
rect 676088 396063 676090 396072
rect 676036 396034 676088 396040
rect 674668 393286 674788 393314
rect 674852 395814 674972 395842
rect 674668 383654 674696 393286
rect 674852 386170 674880 395814
rect 676232 395758 676260 397967
rect 678242 397624 678298 397633
rect 678242 397559 678298 397568
rect 675024 395752 675076 395758
rect 675024 395694 675076 395700
rect 676220 395752 676272 395758
rect 676220 395694 676272 395700
rect 674840 386164 674892 386170
rect 674840 386106 674892 386112
rect 674300 383626 674420 383654
rect 674484 383626 674604 383654
rect 674668 383626 674788 383654
rect 674392 382226 674420 383626
rect 674380 382220 674432 382226
rect 674380 382162 674432 382168
rect 674116 379358 674420 379386
rect 674392 375358 674420 379358
rect 674576 378146 674604 383626
rect 674564 378140 674616 378146
rect 674564 378082 674616 378088
rect 674380 375352 674432 375358
rect 674380 375294 674432 375300
rect 674760 372570 674788 383626
rect 675036 382582 675064 395694
rect 676218 394360 676274 394369
rect 676218 394295 676220 394304
rect 676272 394295 676274 394304
rect 676220 394266 676272 394272
rect 676678 393544 676734 393553
rect 676678 393479 676734 393488
rect 676692 391241 676720 393479
rect 676678 391232 676734 391241
rect 676678 391167 676734 391176
rect 678256 387705 678284 397559
rect 678242 387696 678298 387705
rect 678242 387631 678298 387640
rect 679636 386782 679664 398375
rect 679624 386776 679676 386782
rect 679624 386718 679676 386724
rect 675128 386261 675418 386289
rect 675128 383654 675156 386261
rect 675300 386164 675352 386170
rect 675300 386106 675352 386112
rect 675312 384449 675340 386106
rect 675484 386028 675536 386034
rect 675484 385970 675536 385976
rect 675496 385696 675524 385970
rect 675772 384985 675800 385084
rect 675758 384976 675814 384985
rect 675758 384911 675814 384920
rect 675312 384421 675418 384449
rect 675128 383626 675248 383654
rect 675220 382945 675248 383626
rect 675206 382936 675262 382945
rect 675206 382871 675262 382880
rect 675312 382622 675432 382650
rect 675312 382582 675340 382622
rect 675036 382554 675340 382582
rect 675404 382568 675432 382622
rect 675758 382256 675814 382265
rect 675116 382220 675168 382226
rect 675758 382191 675814 382200
rect 675116 382162 675168 382168
rect 675128 381426 675156 382162
rect 675772 382024 675800 382191
rect 675128 381398 675418 381426
rect 675390 381032 675446 381041
rect 675390 380967 675446 380976
rect 675404 380732 675432 380967
rect 675758 378720 675814 378729
rect 675758 378655 675814 378664
rect 675772 378284 675800 378655
rect 675116 378140 675168 378146
rect 675116 378082 675168 378088
rect 675128 377754 675156 378082
rect 675128 377726 675340 377754
rect 675312 377618 675340 377726
rect 675404 377618 675432 377740
rect 675312 377590 675432 377618
rect 675758 377360 675814 377369
rect 675758 377295 675814 377304
rect 675772 377060 675800 377295
rect 675404 376281 675432 376448
rect 675390 376272 675446 376281
rect 675390 376207 675446 376216
rect 675116 375352 675168 375358
rect 675116 375294 675168 375300
rect 675128 375238 675156 375294
rect 675128 375210 675418 375238
rect 675758 373688 675814 373697
rect 675758 373623 675814 373632
rect 675772 373388 675800 373623
rect 675666 373008 675722 373017
rect 675666 372943 675722 372952
rect 675680 372790 675708 372943
rect 675036 372762 675340 372790
rect 675418 372776 675708 372790
rect 674748 372564 674800 372570
rect 674748 372506 674800 372512
rect 675036 364334 675064 372762
rect 675312 372722 675340 372762
rect 675404 372762 675694 372776
rect 675404 372722 675432 372762
rect 675312 372694 675432 372722
rect 675300 372564 675352 372570
rect 675300 372506 675352 372512
rect 675312 371566 675340 372506
rect 675312 371538 675418 371566
rect 673932 364306 674420 364334
rect 675036 364306 675248 364334
rect 673918 358320 673974 358329
rect 673918 358255 673974 358264
rect 673366 355872 673422 355881
rect 673366 355807 673422 355816
rect 673366 355464 673422 355473
rect 673366 355399 673422 355408
rect 672814 355056 672870 355065
rect 672814 354991 672870 355000
rect 673182 354648 673238 354657
rect 673182 354583 673238 354592
rect 672722 353424 672778 353433
rect 672722 353359 672778 353368
rect 672736 340785 672764 353359
rect 672906 348936 672962 348945
rect 672906 348871 672962 348880
rect 672722 340776 672778 340785
rect 672722 340711 672778 340720
rect 672920 331265 672948 348871
rect 672906 331256 672962 331265
rect 672906 331191 672962 331200
rect 672906 325000 672962 325009
rect 672906 324935 672962 324944
rect 672538 312488 672594 312497
rect 672538 312423 672594 312432
rect 672538 304328 672594 304337
rect 672538 304263 672594 304272
rect 672080 288448 672132 288454
rect 672080 288390 672132 288396
rect 671894 262168 671950 262177
rect 671894 262103 671950 262112
rect 671710 257272 671766 257281
rect 671710 257207 671766 257216
rect 671724 234614 671752 257207
rect 671908 245313 671936 262103
rect 672092 246265 672120 288390
rect 672552 287881 672580 304263
rect 672538 287872 672594 287881
rect 672538 287807 672594 287816
rect 672448 287700 672500 287706
rect 672448 287642 672500 287648
rect 672264 285728 672316 285734
rect 672262 285696 672264 285705
rect 672316 285696 672318 285705
rect 672262 285631 672318 285640
rect 672264 284368 672316 284374
rect 672264 284310 672316 284316
rect 672078 246256 672134 246265
rect 672078 246191 672134 246200
rect 671894 245304 671950 245313
rect 671894 245239 671950 245248
rect 672080 237040 672132 237046
rect 672080 236982 672132 236988
rect 671896 236904 671948 236910
rect 671896 236846 671948 236852
rect 671632 234586 671752 234614
rect 671632 224954 671660 234586
rect 671632 224926 671752 224954
rect 671540 224726 671660 224754
rect 671482 224664 671534 224670
rect 671356 224624 671482 224652
rect 671356 221105 671384 224624
rect 671482 224606 671534 224612
rect 671632 222194 671660 224726
rect 671540 222166 671660 222194
rect 671342 221096 671398 221105
rect 671342 221031 671398 221040
rect 671172 220102 671384 220130
rect 671080 215266 671200 215294
rect 670804 180766 671016 180794
rect 670606 171048 670662 171057
rect 670606 170983 670662 170992
rect 670330 170776 670386 170785
rect 670330 170711 670386 170720
rect 670344 170082 670372 170711
rect 670252 170054 670372 170082
rect 670252 157334 670280 170054
rect 670422 169960 670478 169969
rect 670422 169895 670478 169904
rect 670436 166994 670464 169895
rect 670804 168230 670832 180766
rect 670974 171184 671030 171193
rect 670974 171119 671030 171128
rect 670792 168224 670844 168230
rect 670792 168166 670844 168172
rect 670436 166966 670648 166994
rect 670252 157306 670464 157334
rect 670436 155145 670464 157306
rect 670422 155136 670478 155145
rect 670422 155071 670478 155080
rect 670620 151745 670648 166966
rect 670988 157334 671016 171119
rect 670804 157306 671016 157334
rect 670804 154465 670832 157306
rect 671172 155417 671200 215266
rect 671158 155408 671214 155417
rect 671158 155343 671214 155352
rect 670790 154456 670846 154465
rect 670790 154391 670846 154400
rect 670606 151736 670662 151745
rect 670606 151671 670662 151680
rect 670790 149152 670846 149161
rect 670790 149087 670792 149096
rect 670844 149087 670846 149096
rect 670792 149058 670844 149064
rect 671356 142154 671384 220102
rect 671540 149161 671568 222166
rect 671526 149152 671582 149161
rect 671526 149087 671582 149096
rect 670804 142126 671384 142154
rect 670804 140690 670832 142126
rect 670792 140684 670844 140690
rect 670792 140626 670844 140632
rect 670148 138032 670200 138038
rect 671724 138014 671752 224926
rect 671908 145353 671936 236846
rect 672092 236337 672120 236982
rect 672078 236328 672134 236337
rect 672078 236263 672134 236272
rect 672080 234864 672132 234870
rect 672080 234806 672132 234812
rect 672092 233238 672120 234806
rect 672080 233232 672132 233238
rect 672080 233174 672132 233180
rect 672080 230852 672132 230858
rect 672080 230794 672132 230800
rect 672092 229770 672120 230794
rect 672080 229764 672132 229770
rect 672080 229706 672132 229712
rect 672276 227089 672304 284310
rect 672262 227080 672318 227089
rect 672262 227015 672318 227024
rect 672264 225888 672316 225894
rect 672262 225856 672264 225865
rect 672316 225856 672318 225865
rect 672262 225791 672318 225800
rect 672264 225548 672316 225554
rect 672264 225490 672316 225496
rect 672032 225448 672088 225457
rect 672032 225383 672088 225392
rect 672046 225282 672074 225383
rect 672156 225344 672208 225350
rect 672154 225312 672156 225321
rect 672208 225312 672210 225321
rect 672034 225276 672086 225282
rect 672154 225247 672210 225256
rect 672034 225218 672086 225224
rect 672276 225049 672304 225490
rect 672262 225040 672318 225049
rect 672262 224975 672318 224984
rect 672078 223952 672134 223961
rect 672078 223887 672134 223896
rect 672092 217841 672120 223887
rect 672262 223680 672318 223689
rect 672262 223615 672318 223624
rect 672078 217832 672134 217841
rect 672078 217767 672134 217776
rect 672078 217560 672134 217569
rect 672078 217495 672134 217504
rect 672092 213761 672120 217495
rect 672276 215937 672304 223615
rect 672262 215928 672318 215937
rect 672262 215863 672318 215872
rect 672078 213752 672134 213761
rect 672078 213687 672134 213696
rect 672078 213344 672134 213353
rect 672078 213279 672134 213288
rect 671894 145344 671950 145353
rect 671894 145279 671950 145288
rect 670148 137974 670200 137980
rect 670804 137986 671752 138014
rect 670146 130928 670202 130937
rect 670146 130863 670202 130872
rect 669964 130688 670016 130694
rect 669964 130630 670016 130636
rect 668582 129024 668638 129033
rect 668582 128959 668638 128968
rect 668768 128648 668820 128654
rect 668768 128590 668820 128596
rect 668582 127800 668638 127809
rect 668582 127735 668638 127744
rect 667202 122088 667258 122097
rect 667202 122023 667258 122032
rect 590568 120760 590620 120766
rect 590568 120702 590620 120708
rect 589646 119912 589702 119921
rect 589646 119847 589702 119856
rect 589462 116648 589518 116657
rect 589462 116583 589518 116592
rect 589476 116006 589504 116583
rect 589464 116000 589516 116006
rect 589464 115942 589516 115948
rect 589660 115258 589688 119847
rect 590106 118280 590162 118289
rect 590106 118215 590162 118224
rect 589648 115252 589700 115258
rect 589648 115194 589700 115200
rect 589462 113384 589518 113393
rect 589462 113319 589518 113328
rect 589476 113218 589504 113319
rect 589464 113212 589516 113218
rect 589464 113154 589516 113160
rect 590120 112470 590148 118215
rect 590290 115016 590346 115025
rect 590290 114951 590346 114960
rect 590108 112464 590160 112470
rect 590108 112406 590160 112412
rect 589462 111752 589518 111761
rect 589462 111687 589518 111696
rect 589476 110498 589504 111687
rect 589464 110492 589516 110498
rect 589464 110434 589516 110440
rect 589462 110120 589518 110129
rect 589462 110055 589518 110064
rect 589476 109138 589504 110055
rect 589464 109132 589516 109138
rect 589464 109074 589516 109080
rect 589462 108488 589518 108497
rect 589462 108423 589518 108432
rect 589476 107710 589504 108423
rect 589464 107704 589516 107710
rect 589464 107646 589516 107652
rect 589462 106856 589518 106865
rect 589462 106791 589518 106800
rect 589476 106350 589504 106791
rect 589464 106344 589516 106350
rect 589464 106286 589516 106292
rect 589830 105224 589886 105233
rect 589830 105159 589886 105168
rect 589844 104922 589872 105159
rect 589832 104916 589884 104922
rect 589832 104858 589884 104864
rect 590304 103514 590332 114951
rect 666650 109372 666706 109381
rect 666650 109307 666706 109316
rect 666664 103514 666692 109307
rect 667940 108044 667992 108050
rect 667940 107986 667992 107992
rect 667952 107817 667980 107986
rect 667938 107808 667994 107817
rect 667938 107743 667994 107752
rect 668400 106208 668452 106214
rect 668122 106176 668178 106185
rect 668122 106111 668178 106120
rect 668398 106176 668400 106185
rect 668452 106176 668454 106185
rect 668398 106111 668454 106120
rect 589936 103486 590332 103514
rect 666572 103486 666692 103514
rect 588728 103420 588780 103426
rect 588728 103362 588780 103368
rect 589462 101960 589518 101969
rect 589462 101895 589518 101904
rect 589476 100162 589504 101895
rect 589464 100156 589516 100162
rect 589464 100098 589516 100104
rect 589936 88330 589964 103486
rect 592684 100020 592736 100026
rect 592684 99962 592736 99968
rect 595272 100014 595608 100042
rect 596192 100014 596344 100042
rect 596468 100014 597080 100042
rect 591304 96076 591356 96082
rect 591304 96018 591356 96024
rect 589924 88324 589976 88330
rect 589924 88266 589976 88272
rect 588544 73160 588596 73166
rect 588544 73102 588596 73108
rect 587164 62076 587216 62082
rect 587164 62018 587216 62024
rect 591316 54505 591344 96018
rect 592696 64870 592724 99962
rect 595272 99142 595300 100014
rect 595260 99136 595312 99142
rect 595260 99078 595312 99084
rect 594064 95940 594116 95946
rect 594064 95882 594116 95888
rect 592684 64864 592736 64870
rect 592684 64806 592736 64812
rect 594076 57934 594104 95882
rect 595272 93854 595300 99078
rect 595272 93826 595484 93854
rect 595456 80714 595484 93826
rect 595444 80708 595496 80714
rect 595444 80650 595496 80656
rect 594064 57928 594116 57934
rect 594064 57870 594116 57876
rect 591302 54496 591358 54505
rect 591302 54431 591358 54440
rect 596192 54398 596220 100014
rect 596468 55214 596496 100014
rect 597802 99770 597830 100028
rect 598216 100014 598552 100042
rect 599136 100014 599288 100042
rect 599688 100014 600024 100042
rect 600516 100014 600760 100042
rect 601160 100014 601496 100042
rect 601896 100014 602232 100042
rect 602632 100014 602968 100042
rect 603092 100014 603704 100042
rect 597802 99742 597876 99770
rect 597652 96960 597704 96966
rect 597652 96902 597704 96908
rect 596456 55208 596508 55214
rect 596456 55150 596508 55156
rect 597664 54942 597692 96902
rect 597848 55078 597876 99742
rect 598216 96966 598244 100014
rect 598204 96960 598256 96966
rect 598204 96902 598256 96908
rect 598940 95804 598992 95810
rect 598940 95746 598992 95752
rect 598952 56030 598980 95746
rect 598940 56024 598992 56030
rect 598940 55966 598992 55972
rect 597836 55072 597888 55078
rect 597836 55014 597888 55020
rect 597652 54936 597704 54942
rect 597652 54878 597704 54884
rect 599136 54806 599164 100014
rect 599688 95810 599716 100014
rect 600320 96960 600372 96966
rect 600320 96902 600372 96908
rect 599676 95804 599728 95810
rect 599676 95746 599728 95752
rect 600332 79354 600360 96902
rect 600320 79348 600372 79354
rect 600320 79290 600372 79296
rect 600516 57254 600544 100014
rect 601160 96966 601188 100014
rect 601148 96960 601200 96966
rect 601148 96902 601200 96908
rect 600504 57248 600556 57254
rect 600504 57190 600556 57196
rect 601896 55894 601924 100014
rect 602632 96082 602660 100014
rect 602620 96076 602672 96082
rect 602620 96018 602672 96024
rect 603092 58818 603120 100014
rect 604426 99770 604454 100028
rect 605176 100014 605512 100042
rect 605912 100014 606248 100042
rect 606648 100014 606984 100042
rect 607384 100014 607720 100042
rect 608120 100014 608548 100042
rect 608856 100014 609192 100042
rect 609592 100014 609928 100042
rect 610328 100014 610664 100042
rect 611064 100014 611308 100042
rect 611800 100014 612136 100042
rect 612536 100014 612688 100042
rect 613272 100014 613884 100042
rect 604426 99742 604500 99770
rect 603080 58812 603132 58818
rect 603080 58754 603132 58760
rect 604472 58682 604500 99742
rect 605484 97442 605512 100014
rect 605472 97436 605524 97442
rect 605472 97378 605524 97384
rect 606220 96966 606248 100014
rect 606208 96960 606260 96966
rect 606208 96902 606260 96908
rect 606956 91798 606984 100014
rect 607128 96960 607180 96966
rect 607128 96902 607180 96908
rect 606944 91792 606996 91798
rect 606944 91734 606996 91740
rect 607140 75342 607168 96902
rect 607692 94518 607720 100014
rect 607680 94512 607732 94518
rect 607680 94454 607732 94460
rect 608520 84182 608548 100014
rect 609164 96762 609192 100014
rect 609152 96756 609204 96762
rect 609152 96698 609204 96704
rect 609704 96756 609756 96762
rect 609704 96698 609756 96704
rect 609716 93158 609744 96698
rect 609704 93152 609756 93158
rect 609704 93094 609756 93100
rect 609900 85542 609928 100014
rect 610636 96082 610664 100014
rect 610624 96076 610676 96082
rect 610624 96018 610676 96024
rect 611280 91050 611308 100014
rect 611912 97436 611964 97442
rect 611912 97378 611964 97384
rect 611924 93854 611952 97378
rect 612108 96898 612136 100014
rect 612660 97442 612688 100014
rect 612648 97436 612700 97442
rect 612648 97378 612700 97384
rect 612096 96892 612148 96898
rect 612096 96834 612148 96840
rect 612648 96892 612700 96898
rect 612648 96834 612700 96840
rect 611924 93826 612044 93854
rect 611268 91044 611320 91050
rect 611268 90986 611320 90992
rect 609888 85536 609940 85542
rect 609888 85478 609940 85484
rect 608508 84176 608560 84182
rect 608508 84118 608560 84124
rect 612016 76702 612044 93826
rect 612660 79354 612688 96834
rect 613856 80850 613884 100014
rect 613994 99770 614022 100028
rect 614744 100014 615264 100042
rect 615480 100014 615816 100042
rect 616216 100014 616552 100042
rect 616952 100014 617288 100042
rect 617688 100014 618024 100042
rect 618424 100014 618760 100042
rect 619160 100014 619588 100042
rect 619896 100014 620140 100042
rect 620632 100014 620968 100042
rect 621368 100014 621704 100042
rect 622104 100014 622348 100042
rect 622840 100014 623176 100042
rect 623576 100014 623728 100042
rect 624312 100014 624648 100042
rect 613994 99742 614068 99770
rect 613844 80844 613896 80850
rect 613844 80786 613896 80792
rect 614040 79490 614068 99742
rect 615236 93854 615264 100014
rect 615788 96966 615816 100014
rect 615776 96960 615828 96966
rect 615776 96902 615828 96908
rect 616524 94994 616552 100014
rect 616788 96960 616840 96966
rect 616788 96902 616840 96908
rect 616512 94988 616564 94994
rect 616512 94930 616564 94936
rect 615236 93826 615448 93854
rect 615420 80986 615448 93826
rect 615408 80980 615460 80986
rect 615408 80922 615460 80928
rect 614028 79484 614080 79490
rect 614028 79426 614080 79432
rect 612648 79348 612700 79354
rect 612648 79290 612700 79296
rect 612004 76696 612056 76702
rect 612004 76638 612056 76644
rect 616800 75478 616828 96902
rect 617260 96898 617288 100014
rect 617248 96892 617300 96898
rect 617248 96834 617300 96840
rect 617996 92478 618024 100014
rect 618732 97986 618760 100014
rect 618720 97980 618772 97986
rect 618720 97922 618772 97928
rect 618168 96892 618220 96898
rect 618168 96834 618220 96840
rect 617984 92472 618036 92478
rect 617984 92414 618036 92420
rect 618180 91186 618208 96834
rect 619560 93838 619588 100014
rect 620112 97170 620140 100014
rect 620284 97436 620336 97442
rect 620284 97378 620336 97384
rect 620100 97164 620152 97170
rect 620100 97106 620152 97112
rect 619548 93832 619600 93838
rect 619548 93774 619600 93780
rect 618628 93152 618680 93158
rect 618628 93094 618680 93100
rect 618168 91180 618220 91186
rect 618168 91122 618220 91128
rect 618168 91044 618220 91050
rect 618168 90986 618220 90992
rect 618180 88194 618208 90986
rect 618168 88188 618220 88194
rect 618168 88130 618220 88136
rect 618640 85406 618668 93094
rect 618628 85400 618680 85406
rect 618628 85342 618680 85348
rect 620296 76838 620324 97378
rect 620940 95198 620968 100014
rect 621676 97442 621704 100014
rect 622320 99346 622348 100014
rect 622308 99340 622360 99346
rect 622308 99282 622360 99288
rect 621664 97436 621716 97442
rect 621664 97378 621716 97384
rect 623148 97306 623176 100014
rect 623700 99210 623728 100014
rect 623688 99204 623740 99210
rect 623688 99146 623740 99152
rect 624620 99074 624648 100014
rect 625034 99770 625062 100028
rect 625784 100014 626120 100042
rect 626520 100014 626856 100042
rect 627256 100014 627592 100042
rect 627992 100014 628328 100042
rect 628728 100014 629064 100042
rect 629464 100014 629800 100042
rect 630200 100014 630536 100042
rect 630936 100014 631272 100042
rect 631672 100014 632008 100042
rect 632408 100014 632744 100042
rect 633144 100014 633296 100042
rect 633880 100014 634216 100042
rect 634616 100014 634768 100042
rect 635352 100014 635596 100042
rect 625034 99742 625108 99770
rect 624608 99068 624660 99074
rect 624608 99010 624660 99016
rect 625080 98938 625108 99742
rect 625068 98932 625120 98938
rect 625068 98874 625120 98880
rect 625804 97980 625856 97986
rect 625804 97922 625856 97928
rect 623136 97300 623188 97306
rect 623136 97242 623188 97248
rect 621664 96076 621716 96082
rect 621664 96018 621716 96024
rect 620928 95192 620980 95198
rect 620928 95134 620980 95140
rect 620652 94512 620704 94518
rect 620652 94454 620704 94460
rect 620664 89690 620692 94454
rect 620652 89684 620704 89690
rect 620652 89626 620704 89632
rect 621676 86358 621704 96018
rect 625436 95192 625488 95198
rect 625436 95134 625488 95140
rect 624976 94988 625028 94994
rect 624976 94930 625028 94936
rect 622400 91792 622452 91798
rect 622400 91734 622452 91740
rect 622412 88330 622440 91734
rect 624988 88641 625016 94930
rect 625448 94489 625476 95134
rect 625434 94480 625490 94489
rect 625434 94415 625490 94424
rect 625816 92041 625844 97922
rect 626092 97034 626120 100014
rect 626448 97164 626500 97170
rect 626448 97106 626500 97112
rect 626080 97028 626132 97034
rect 626080 96970 626132 96976
rect 626264 93832 626316 93838
rect 626264 93774 626316 93780
rect 626276 92857 626304 93774
rect 626460 93673 626488 97106
rect 626828 96898 626856 100014
rect 627564 97578 627592 100014
rect 628300 97850 628328 100014
rect 629036 98802 629064 100014
rect 629024 98796 629076 98802
rect 629024 98738 629076 98744
rect 629772 97986 629800 100014
rect 630508 98666 630536 100014
rect 630772 99340 630824 99346
rect 630772 99282 630824 99288
rect 630496 98660 630548 98666
rect 630496 98602 630548 98608
rect 629760 97980 629812 97986
rect 629760 97922 629812 97928
rect 628288 97844 628340 97850
rect 628288 97786 628340 97792
rect 627552 97572 627604 97578
rect 627552 97514 627604 97520
rect 629300 97436 629352 97442
rect 629300 97378 629352 97384
rect 626816 96892 626868 96898
rect 626816 96834 626868 96840
rect 629312 95826 629340 97378
rect 630784 95826 630812 99282
rect 631244 97714 631272 100014
rect 631416 98320 631468 98326
rect 631416 98262 631468 98268
rect 631428 97850 631456 98262
rect 631416 97844 631468 97850
rect 631416 97786 631468 97792
rect 631232 97708 631284 97714
rect 631232 97650 631284 97656
rect 631980 97442 632008 100014
rect 632716 97850 632744 100014
rect 632704 97844 632756 97850
rect 632704 97786 632756 97792
rect 631968 97436 632020 97442
rect 631968 97378 632020 97384
rect 633268 97306 633296 100014
rect 633440 99204 633492 99210
rect 633440 99146 633492 99152
rect 632060 97300 632112 97306
rect 632060 97242 632112 97248
rect 633256 97300 633308 97306
rect 633256 97242 633308 97248
rect 629280 95798 629340 95826
rect 630752 95798 630812 95826
rect 632072 95826 632100 97242
rect 633452 95826 633480 99146
rect 633624 98184 633676 98190
rect 633624 98126 633676 98132
rect 633636 97578 633664 98126
rect 633624 97572 633676 97578
rect 633624 97514 633676 97520
rect 633808 97572 633860 97578
rect 633808 97514 633860 97520
rect 633820 97034 633848 97514
rect 634188 97170 634216 100014
rect 634176 97164 634228 97170
rect 634176 97106 634228 97112
rect 634740 97034 634768 100014
rect 635004 99068 635056 99074
rect 635004 99010 635056 99016
rect 633808 97028 633860 97034
rect 633808 96970 633860 96976
rect 634728 97028 634780 97034
rect 634728 96970 634780 96976
rect 635016 95826 635044 99010
rect 635568 96937 635596 100014
rect 635752 100014 636088 100042
rect 636824 100014 637068 100042
rect 635554 96928 635610 96937
rect 635554 96863 635610 96872
rect 635752 95985 635780 100014
rect 636292 98932 636344 98938
rect 636292 98874 636344 98880
rect 635738 95976 635794 95985
rect 635738 95911 635794 95920
rect 636304 95826 636332 98874
rect 637040 96937 637068 100014
rect 637546 99770 637574 100028
rect 638296 100014 638632 100042
rect 637546 99742 637620 99770
rect 637026 96928 637082 96937
rect 637026 96863 637082 96872
rect 637592 96354 637620 99742
rect 637764 97572 637816 97578
rect 637764 97514 637816 97520
rect 637580 96348 637632 96354
rect 637580 96290 637632 96296
rect 637776 95826 637804 97514
rect 638604 96490 638632 100014
rect 639018 99770 639046 100028
rect 639768 100014 640104 100042
rect 639018 99742 639092 99770
rect 638592 96484 638644 96490
rect 638592 96426 638644 96432
rect 632072 95798 632224 95826
rect 633452 95798 633696 95826
rect 635016 95798 635168 95826
rect 636304 95798 636640 95826
rect 637776 95798 638112 95826
rect 639064 95810 639092 99742
rect 639236 96892 639288 96898
rect 639236 96834 639288 96840
rect 639248 95826 639276 96834
rect 640076 96626 640104 100014
rect 640490 99770 640518 100028
rect 641240 100014 641576 100042
rect 640490 99742 640564 99770
rect 640064 96620 640116 96626
rect 640064 96562 640116 96568
rect 640536 96150 640564 99742
rect 640708 98184 640760 98190
rect 640708 98126 640760 98132
rect 640524 96144 640576 96150
rect 640524 96086 640576 96092
rect 640720 95826 640748 98126
rect 641548 96490 641576 100014
rect 641962 99770 641990 100028
rect 642712 100014 643048 100042
rect 641962 99742 642036 99770
rect 642008 96529 642036 99742
rect 642180 98320 642232 98326
rect 642180 98262 642232 98268
rect 641994 96520 642050 96529
rect 641352 96484 641404 96490
rect 641352 96426 641404 96432
rect 641536 96484 641588 96490
rect 641994 96455 642050 96464
rect 641536 96426 641588 96432
rect 639052 95804 639104 95810
rect 639248 95798 639584 95826
rect 640720 95798 641056 95826
rect 639052 95746 639104 95752
rect 641364 95470 641392 96426
rect 642192 95826 642220 98262
rect 643020 97578 643048 100014
rect 643434 99770 643462 100028
rect 644184 100014 644336 100042
rect 644920 100014 645532 100042
rect 645656 100014 645808 100042
rect 643434 99742 643508 99770
rect 643008 97572 643060 97578
rect 643008 97514 643060 97520
rect 642192 95798 642528 95826
rect 643480 95470 643508 99742
rect 643652 98796 643704 98802
rect 643652 98738 643704 98744
rect 643664 95826 643692 98738
rect 644308 96898 644336 100014
rect 645308 98048 645360 98054
rect 645308 97990 645360 97996
rect 644296 96892 644348 96898
rect 644296 96834 644348 96840
rect 645124 96620 645176 96626
rect 645124 96562 645176 96568
rect 644940 96144 644992 96150
rect 644938 96112 644940 96121
rect 644992 96112 644994 96121
rect 644938 96047 644994 96056
rect 643664 95798 644000 95826
rect 645136 95674 645164 96562
rect 645320 95826 645348 97990
rect 645504 96218 645532 100014
rect 645492 96212 645544 96218
rect 645492 96154 645544 96160
rect 645780 96082 645808 100014
rect 646378 99770 646406 100028
rect 647114 99770 647142 100028
rect 647864 100014 648476 100042
rect 648600 100014 648936 100042
rect 649336 100014 649764 100042
rect 650072 100014 650408 100042
rect 650808 100014 651328 100042
rect 651544 100014 651880 100042
rect 652280 100014 652616 100042
rect 653016 100014 653352 100042
rect 653752 100014 653996 100042
rect 654488 100014 654824 100042
rect 655224 100014 655468 100042
rect 646378 99742 646452 99770
rect 647114 99742 647188 99770
rect 646424 96626 646452 99742
rect 647160 98802 647188 99742
rect 647148 98796 647200 98802
rect 647148 98738 647200 98744
rect 646596 98660 646648 98666
rect 646596 98602 646648 98608
rect 646412 96620 646464 96626
rect 646412 96562 646464 96568
rect 645768 96076 645820 96082
rect 645768 96018 645820 96024
rect 646608 95826 646636 98602
rect 647516 97844 647568 97850
rect 647516 97786 647568 97792
rect 647332 97708 647384 97714
rect 647332 97650 647384 97656
rect 647056 97028 647108 97034
rect 647056 96970 647108 96976
rect 645320 95798 645472 95826
rect 646608 95798 646944 95826
rect 645124 95668 645176 95674
rect 645124 95610 645176 95616
rect 641352 95464 641404 95470
rect 641352 95406 641404 95412
rect 643468 95464 643520 95470
rect 643468 95406 643520 95412
rect 647068 95198 647096 96970
rect 647056 95192 647108 95198
rect 647056 95134 647108 95140
rect 647344 95033 647372 97650
rect 647330 95024 647386 95033
rect 647330 94959 647386 94968
rect 647528 93770 647556 97786
rect 648066 96520 648122 96529
rect 648066 96455 648068 96464
rect 648120 96455 648122 96464
rect 648068 96426 648120 96432
rect 647884 96212 647936 96218
rect 647884 96154 647936 96160
rect 647896 95849 647924 96154
rect 648068 96076 648120 96082
rect 648068 96018 648120 96024
rect 647882 95840 647938 95849
rect 647882 95775 647938 95784
rect 647884 95464 647936 95470
rect 647884 95406 647936 95412
rect 647700 95328 647752 95334
rect 647700 95270 647752 95276
rect 647516 93764 647568 93770
rect 647516 93706 647568 93712
rect 626446 93664 626502 93673
rect 626446 93599 626502 93608
rect 626262 92848 626318 92857
rect 626262 92783 626318 92792
rect 647712 92478 647740 95270
rect 626448 92472 626500 92478
rect 626448 92414 626500 92420
rect 647700 92472 647752 92478
rect 647700 92414 647752 92420
rect 625802 92032 625858 92041
rect 625802 91967 625858 91976
rect 626460 91225 626488 92414
rect 626446 91216 626502 91225
rect 626446 91151 626502 91160
rect 626448 91044 626500 91050
rect 626448 90986 626500 90992
rect 626460 90409 626488 90986
rect 626446 90400 626502 90409
rect 626446 90335 626502 90344
rect 625436 89684 625488 89690
rect 625436 89626 625488 89632
rect 625250 89584 625306 89593
rect 625250 89519 625306 89528
rect 625264 88641 625292 89519
rect 625448 88777 625476 89626
rect 625434 88768 625490 88777
rect 625434 88703 625490 88712
rect 624974 88632 625030 88641
rect 624974 88567 625030 88576
rect 625250 88632 625306 88641
rect 625250 88567 625306 88576
rect 622400 88324 622452 88330
rect 622400 88266 622452 88272
rect 626448 88324 626500 88330
rect 626448 88266 626500 88272
rect 626264 88188 626316 88194
rect 626264 88130 626316 88136
rect 626276 87145 626304 88130
rect 626460 87961 626488 88266
rect 626446 87952 626502 87961
rect 626446 87887 626502 87896
rect 626262 87136 626318 87145
rect 626262 87071 626318 87080
rect 647896 86630 647924 95406
rect 648080 95402 648108 96018
rect 648068 95396 648120 95402
rect 648068 95338 648120 95344
rect 648252 93764 648304 93770
rect 648252 93706 648304 93712
rect 648264 89593 648292 93706
rect 648250 89584 648306 89593
rect 648250 89519 648306 89528
rect 648448 87038 648476 100014
rect 648620 97436 648672 97442
rect 648620 97378 648672 97384
rect 648632 96370 648660 97378
rect 648908 96490 648936 100014
rect 649080 97164 649132 97170
rect 649080 97106 649132 97112
rect 648896 96484 648948 96490
rect 648896 96426 648948 96432
rect 648632 96342 648844 96370
rect 648618 96112 648674 96121
rect 648618 96047 648620 96056
rect 648672 96047 648674 96056
rect 648620 96018 648672 96024
rect 648620 95804 648672 95810
rect 648620 95746 648672 95752
rect 648632 90846 648660 95746
rect 648816 92041 648844 96342
rect 648802 92032 648858 92041
rect 648802 91967 648858 91976
rect 648620 90840 648672 90846
rect 648620 90782 648672 90788
rect 649092 89714 649120 97106
rect 649262 96520 649318 96529
rect 649262 96455 649318 96464
rect 649276 96218 649304 96455
rect 649264 96212 649316 96218
rect 649264 96154 649316 96160
rect 648632 89686 649120 89714
rect 648436 87032 648488 87038
rect 648436 86974 648488 86980
rect 647884 86624 647936 86630
rect 647884 86566 647936 86572
rect 621664 86352 621716 86358
rect 626448 86352 626500 86358
rect 621664 86294 621716 86300
rect 626446 86320 626448 86329
rect 626500 86320 626502 86329
rect 626446 86255 626502 86264
rect 626448 85536 626500 85542
rect 626446 85504 626448 85513
rect 626500 85504 626502 85513
rect 626446 85439 626502 85448
rect 625252 85400 625304 85406
rect 625252 85342 625304 85348
rect 625264 84697 625292 85342
rect 648632 84697 648660 89686
rect 649736 88806 649764 100014
rect 650380 97306 650408 100014
rect 650368 97300 650420 97306
rect 650368 97242 650420 97248
rect 650552 97164 650604 97170
rect 650552 97106 650604 97112
rect 650276 95192 650328 95198
rect 650276 95134 650328 95140
rect 649724 88800 649776 88806
rect 649724 88742 649776 88748
rect 625250 84688 625306 84697
rect 625250 84623 625306 84632
rect 648618 84688 648674 84697
rect 648618 84623 648674 84632
rect 626448 84176 626500 84182
rect 626448 84118 626500 84124
rect 626460 83881 626488 84118
rect 626446 83872 626502 83881
rect 626446 83807 626502 83816
rect 628746 83328 628802 83337
rect 628746 83263 628802 83272
rect 628760 81122 628788 83263
rect 650288 82249 650316 95134
rect 650564 87145 650592 97106
rect 651300 93634 651328 100014
rect 651852 97714 651880 100014
rect 651840 97708 651892 97714
rect 651840 97650 651892 97656
rect 652588 96626 652616 100014
rect 652208 96620 652260 96626
rect 652208 96562 652260 96568
rect 652576 96620 652628 96626
rect 652576 96562 652628 96568
rect 652024 95668 652076 95674
rect 652024 95610 652076 95616
rect 651288 93628 651340 93634
rect 651288 93570 651340 93576
rect 650550 87136 650606 87145
rect 650550 87071 650606 87080
rect 652036 86766 652064 95610
rect 652024 86760 652076 86766
rect 652024 86702 652076 86708
rect 652220 86494 652248 96562
rect 653324 95810 653352 100014
rect 653968 97442 653996 100014
rect 653956 97436 654008 97442
rect 653956 97378 654008 97384
rect 654796 96762 654824 100014
rect 655244 97844 655296 97850
rect 655244 97786 655296 97792
rect 655256 97578 655284 97786
rect 655440 97578 655468 100014
rect 655808 100014 655960 100042
rect 656696 100014 656848 100042
rect 657432 100014 657768 100042
rect 655244 97572 655296 97578
rect 655244 97514 655296 97520
rect 655428 97572 655480 97578
rect 655428 97514 655480 97520
rect 655244 97436 655296 97442
rect 655244 97378 655296 97384
rect 654784 96756 654836 96762
rect 654784 96698 654836 96704
rect 653312 95804 653364 95810
rect 653312 95746 653364 95752
rect 655256 94217 655284 97378
rect 655428 96756 655480 96762
rect 655428 96698 655480 96704
rect 655242 94208 655298 94217
rect 655242 94143 655298 94152
rect 655440 93854 655468 96698
rect 655256 93826 655468 93854
rect 654692 93628 654744 93634
rect 654692 93570 654744 93576
rect 654704 93401 654732 93570
rect 654690 93392 654746 93401
rect 654690 93327 654746 93336
rect 655256 88330 655284 93826
rect 655428 92472 655480 92478
rect 655428 92414 655480 92420
rect 655440 91497 655468 92414
rect 655426 91488 655482 91497
rect 655426 91423 655482 91432
rect 655428 90840 655480 90846
rect 655428 90782 655480 90788
rect 655440 90681 655468 90782
rect 655426 90672 655482 90681
rect 655426 90607 655482 90616
rect 655808 89865 655836 100014
rect 656820 97170 656848 100014
rect 656808 97164 656860 97170
rect 656808 97106 656860 97112
rect 656716 96960 656768 96966
rect 656716 96902 656768 96908
rect 656346 95840 656402 95849
rect 656346 95775 656402 95784
rect 656164 95532 656216 95538
rect 656164 95474 656216 95480
rect 655794 89856 655850 89865
rect 655794 89791 655850 89800
rect 656176 88670 656204 95474
rect 656164 88664 656216 88670
rect 656164 88606 656216 88612
rect 655244 88324 655296 88330
rect 655244 88266 655296 88272
rect 652208 86488 652260 86494
rect 652208 86430 652260 86436
rect 656360 86358 656388 95775
rect 656728 86902 656756 96902
rect 657740 95132 657768 100014
rect 658154 99770 658182 100028
rect 658904 100014 659240 100042
rect 659640 100014 659976 100042
rect 658154 99742 658228 99770
rect 658200 97442 658228 99742
rect 659212 97986 659240 100014
rect 659200 97980 659252 97986
rect 659200 97922 659252 97928
rect 659948 97850 659976 100014
rect 660132 100014 660376 100042
rect 659752 97844 659804 97850
rect 659752 97786 659804 97792
rect 659936 97844 659988 97850
rect 659936 97786 659988 97792
rect 659568 97708 659620 97714
rect 659568 97650 659620 97656
rect 658188 97436 658240 97442
rect 658188 97378 658240 97384
rect 658280 97300 658332 97306
rect 658280 97242 658332 97248
rect 658292 95132 658320 97242
rect 658832 96824 658884 96830
rect 658832 96766 658884 96772
rect 658844 95132 658872 96766
rect 659580 95132 659608 97650
rect 659764 95146 659792 97786
rect 660132 96966 660160 100014
rect 661960 98796 662012 98802
rect 661960 98738 662012 98744
rect 661408 97164 661460 97170
rect 661408 97106 661460 97112
rect 660120 96960 660172 96966
rect 660120 96902 660172 96908
rect 660672 96348 660724 96354
rect 660672 96290 660724 96296
rect 659764 95118 660146 95146
rect 660684 95132 660712 96290
rect 661420 95132 661448 97106
rect 661972 95132 662000 98738
rect 664168 97980 664220 97986
rect 664168 97922 664220 97928
rect 662512 97572 662564 97578
rect 662512 97514 662564 97520
rect 662524 95132 662552 97514
rect 663064 97436 663116 97442
rect 663064 97378 663116 97384
rect 663076 95132 663104 97378
rect 663800 96212 663852 96218
rect 663800 96154 663852 96160
rect 663812 93129 663840 96154
rect 663984 96076 664036 96082
rect 663984 96018 664036 96024
rect 663798 93120 663854 93129
rect 663798 93055 663854 93064
rect 663996 91769 664024 96018
rect 663982 91760 664038 91769
rect 663982 91695 664038 91704
rect 664180 88806 664208 97922
rect 665364 97844 665416 97850
rect 665364 97786 665416 97792
rect 664352 96620 664404 96626
rect 664352 96562 664404 96568
rect 664364 90681 664392 96562
rect 664536 96484 664588 96490
rect 664536 96426 664588 96432
rect 664350 90672 664406 90681
rect 664350 90607 664406 90616
rect 664548 89865 664576 96426
rect 665180 95804 665232 95810
rect 665180 95746 665232 95752
rect 664534 89856 664590 89865
rect 664534 89791 664590 89800
rect 665192 89049 665220 95746
rect 665376 93401 665404 97786
rect 665362 93392 665418 93401
rect 665362 93327 665418 93336
rect 665178 89040 665234 89049
rect 665178 88975 665234 88984
rect 658556 88800 658608 88806
rect 662328 88800 662380 88806
rect 658608 88748 658858 88754
rect 658556 88742 658858 88748
rect 658568 88726 658858 88742
rect 661986 88748 662328 88754
rect 661986 88742 662380 88748
rect 664168 88800 664220 88806
rect 664168 88742 664220 88748
rect 661986 88726 662368 88742
rect 657452 88664 657504 88670
rect 657504 88612 657754 88618
rect 657452 88606 657754 88612
rect 657464 88590 657754 88606
rect 658306 88330 658504 88346
rect 658306 88324 658516 88330
rect 658306 88318 658464 88324
rect 658464 88266 658516 88272
rect 656716 86896 656768 86902
rect 656716 86838 656768 86844
rect 657188 86494 657216 88196
rect 659580 86902 659608 88196
rect 659568 86896 659620 86902
rect 659568 86838 659620 86844
rect 660132 86766 660160 88196
rect 660120 86760 660172 86766
rect 660120 86702 660172 86708
rect 657176 86488 657228 86494
rect 657176 86430 657228 86436
rect 660684 86358 660712 88196
rect 661420 86630 661448 88196
rect 662524 87038 662552 88196
rect 662512 87032 662564 87038
rect 662512 86974 662564 86980
rect 661408 86624 661460 86630
rect 661408 86566 661460 86572
rect 656348 86352 656400 86358
rect 656348 86294 656400 86300
rect 660672 86352 660724 86358
rect 660672 86294 660724 86300
rect 650274 82240 650330 82249
rect 650274 82175 650330 82184
rect 629206 81696 629262 81705
rect 629206 81631 629262 81640
rect 628748 81116 628800 81122
rect 628748 81058 628800 81064
rect 629220 80034 629248 81631
rect 642456 81116 642508 81122
rect 642456 81058 642508 81064
rect 632808 80974 633144 81002
rect 629208 80028 629260 80034
rect 629208 79970 629260 79976
rect 631048 77988 631100 77994
rect 631048 77930 631100 77936
rect 628472 77648 628524 77654
rect 628472 77590 628524 77596
rect 628484 77450 628512 77590
rect 628472 77444 628524 77450
rect 628472 77386 628524 77392
rect 623042 77344 623098 77353
rect 623042 77279 623098 77288
rect 624424 77308 624476 77314
rect 620284 76832 620336 76838
rect 620284 76774 620336 76780
rect 616788 75472 616840 75478
rect 616788 75414 616840 75420
rect 607128 75336 607180 75342
rect 607128 75278 607180 75284
rect 604460 58676 604512 58682
rect 604460 58618 604512 58624
rect 601884 55888 601936 55894
rect 601884 55830 601936 55836
rect 599124 54800 599176 54806
rect 599124 54742 599176 54748
rect 623056 54670 623084 77279
rect 624424 77250 624476 77256
rect 625804 77308 625856 77314
rect 625804 77250 625856 77256
rect 624436 60042 624464 77250
rect 624424 60036 624476 60042
rect 624424 59978 624476 59984
rect 623044 54664 623096 54670
rect 623044 54606 623096 54612
rect 625816 54534 625844 77250
rect 628484 75290 628512 77386
rect 631060 77314 631088 77930
rect 632808 77654 632836 80974
rect 636752 80708 636804 80714
rect 636752 80650 636804 80656
rect 633440 80028 633492 80034
rect 633440 79970 633492 79976
rect 633452 78130 633480 79970
rect 633898 78568 633954 78577
rect 633898 78503 633954 78512
rect 633440 78124 633492 78130
rect 633440 78066 633492 78072
rect 632796 77648 632848 77654
rect 632796 77590 632848 77596
rect 633912 77353 633940 78503
rect 633898 77344 633954 77353
rect 631048 77308 631100 77314
rect 633898 77279 633954 77288
rect 631048 77250 631100 77256
rect 631060 75290 631088 77250
rect 633912 75290 633940 77279
rect 636764 75290 636792 80650
rect 639602 77616 639658 77625
rect 639602 77551 639658 77560
rect 639616 75290 639644 77551
rect 642468 75290 642496 81058
rect 643080 80974 643140 81002
rect 643112 77994 643140 80974
rect 646320 80980 646372 80986
rect 646320 80922 646372 80928
rect 646044 79484 646096 79490
rect 646044 79426 646096 79432
rect 645308 78124 645360 78130
rect 645308 78066 645360 78072
rect 643100 77988 643152 77994
rect 643100 77930 643152 77936
rect 645320 75290 645348 78066
rect 628176 75262 628512 75290
rect 631028 75262 631088 75290
rect 633880 75262 633940 75290
rect 636732 75262 636792 75290
rect 639584 75262 639644 75290
rect 642436 75262 642496 75290
rect 645288 75262 645348 75290
rect 646056 74534 646084 79426
rect 646056 74506 646176 74534
rect 646148 67153 646176 74506
rect 646332 69193 646360 80922
rect 647332 80844 647384 80850
rect 647332 80786 647384 80792
rect 646688 75472 646740 75478
rect 646688 75414 646740 75420
rect 646504 75336 646556 75342
rect 646504 75278 646556 75284
rect 646516 74225 646544 75278
rect 646502 74216 646558 74225
rect 646502 74151 646558 74160
rect 646700 71777 646728 75414
rect 646686 71768 646742 71777
rect 646686 71703 646742 71712
rect 646318 69184 646374 69193
rect 646318 69119 646374 69128
rect 646134 67144 646190 67153
rect 646134 67079 646190 67088
rect 625988 66904 626040 66910
rect 625988 66846 626040 66852
rect 625804 54528 625856 54534
rect 625804 54470 625856 54476
rect 596180 54392 596232 54398
rect 596180 54334 596232 54340
rect 583024 54256 583076 54262
rect 583024 54198 583076 54204
rect 580448 54120 580500 54126
rect 580448 54062 580500 54068
rect 574928 53848 574980 53854
rect 574928 53790 574980 53796
rect 459834 53680 459890 53689
rect 459834 53615 459890 53624
rect 460754 53680 460810 53689
rect 460754 53615 460810 53624
rect 461674 53680 461730 53689
rect 461674 53615 461730 53624
rect 462594 53680 462650 53689
rect 462594 53615 462650 53624
rect 463884 53644 463936 53650
rect 129004 53236 129056 53242
rect 129004 53178 129056 53184
rect 51724 52012 51776 52018
rect 51724 51954 51776 51960
rect 50528 51876 50580 51882
rect 50528 51818 50580 51824
rect 128360 44872 128412 44878
rect 128360 44814 128412 44820
rect 128372 44470 128400 44814
rect 129016 44674 129044 53178
rect 312360 53168 312412 53174
rect 312018 53116 312360 53122
rect 312018 53110 312412 53116
rect 313740 53168 313792 53174
rect 316316 53168 316368 53174
rect 313792 53116 314042 53122
rect 313740 53110 314042 53116
rect 130384 53100 130436 53106
rect 130384 53042 130436 53048
rect 129372 52012 129424 52018
rect 129372 51954 129424 51960
rect 129188 51740 129240 51746
rect 129188 51682 129240 51688
rect 129200 47870 129228 51682
rect 129188 47864 129240 47870
rect 129188 47806 129240 47812
rect 129384 45354 129412 51954
rect 129648 50380 129700 50386
rect 129648 50322 129700 50328
rect 129660 46102 129688 50322
rect 129648 46096 129700 46102
rect 129648 46038 129700 46044
rect 130396 45558 130424 53042
rect 130568 51876 130620 51882
rect 130568 51818 130620 51824
rect 130384 45552 130436 45558
rect 130384 45494 130436 45500
rect 129372 45348 129424 45354
rect 129372 45290 129424 45296
rect 129372 45008 129424 45014
rect 129372 44950 129424 44956
rect 129004 44668 129056 44674
rect 129004 44610 129056 44616
rect 50344 44464 50396 44470
rect 50344 44406 50396 44412
rect 128360 44464 128412 44470
rect 128360 44406 128412 44412
rect 43628 44328 43680 44334
rect 43628 44270 43680 44276
rect 43444 44192 43496 44198
rect 43444 44134 43496 44140
rect 129384 44062 129412 44950
rect 130580 44441 130608 51818
rect 306024 51746 306052 53108
rect 145380 51740 145432 51746
rect 145380 51682 145432 51688
rect 306012 51740 306064 51746
rect 306012 51682 306064 51688
rect 145392 50810 145420 51682
rect 145084 50782 145420 50810
rect 308048 50289 308076 53108
rect 312018 53094 312400 53110
rect 313752 53108 314042 53110
rect 316020 53116 316316 53122
rect 316020 53110 316368 53116
rect 317696 53168 317748 53174
rect 317748 53116 318380 53122
rect 317696 53110 318380 53116
rect 313752 53094 314056 53108
rect 316020 53094 316356 53110
rect 317708 53094 318380 53110
rect 314028 50386 314056 53094
rect 318352 50522 318380 53094
rect 459146 52828 459198 52834
rect 459146 52770 459198 52776
rect 459158 52564 459186 52770
rect 459848 52578 459876 53615
rect 460388 52964 460440 52970
rect 460388 52906 460440 52912
rect 460400 52578 460428 52906
rect 460768 52578 460796 53615
rect 461308 53100 461360 53106
rect 461308 53042 461360 53048
rect 461320 52578 461348 53042
rect 461688 52578 461716 53615
rect 462228 53372 462280 53378
rect 462228 53314 462280 53320
rect 462240 52578 462268 53314
rect 462608 52578 462636 53615
rect 463884 53586 463936 53592
rect 464528 53644 464580 53650
rect 464528 53586 464580 53592
rect 464804 53644 464856 53650
rect 464804 53586 464856 53592
rect 474280 53644 474332 53650
rect 474280 53586 474332 53592
rect 474464 53644 474516 53650
rect 474464 53586 474516 53592
rect 475200 53644 475252 53650
rect 475200 53586 475252 53592
rect 475384 53644 475436 53650
rect 475384 53586 475436 53592
rect 480076 53644 480128 53650
rect 480076 53586 480128 53592
rect 463608 53508 463660 53514
rect 463608 53450 463660 53456
rect 463148 53236 463200 53242
rect 463148 53178 463200 53184
rect 463160 52578 463188 53178
rect 463620 52578 463648 53450
rect 463896 52578 463924 53586
rect 459632 52550 459876 52578
rect 460092 52550 460428 52578
rect 460552 52550 460796 52578
rect 461012 52550 461348 52578
rect 461472 52550 461716 52578
rect 461932 52550 462268 52578
rect 462392 52550 462636 52578
rect 462852 52550 463188 52578
rect 463312 52550 463648 52578
rect 463772 52550 463924 52578
rect 464540 52442 464568 53586
rect 464816 52834 464844 53586
rect 464988 53508 465040 53514
rect 464988 53450 465040 53456
rect 464804 52828 464856 52834
rect 464804 52770 464856 52776
rect 465000 52578 465028 53450
rect 468298 53272 468354 53281
rect 468298 53207 468300 53216
rect 468352 53207 468354 53216
rect 468300 53178 468352 53184
rect 465126 52828 465178 52834
rect 465126 52770 465178 52776
rect 464692 52550 465028 52578
rect 465138 52564 465166 52770
rect 474292 52698 474320 53586
rect 474476 52970 474504 53586
rect 475212 53281 475240 53586
rect 475198 53272 475254 53281
rect 475198 53207 475254 53216
rect 474464 52964 474516 52970
rect 474464 52906 474516 52912
rect 475396 52834 475424 53586
rect 480088 53106 480116 53586
rect 480076 53100 480128 53106
rect 480076 53042 480128 53048
rect 475384 52828 475436 52834
rect 475384 52770 475436 52776
rect 465908 52692 465960 52698
rect 465908 52634 465960 52640
rect 474280 52692 474332 52698
rect 474280 52634 474332 52640
rect 465920 52578 465948 52634
rect 465612 52550 465948 52578
rect 464232 52414 464568 52442
rect 318340 50516 318392 50522
rect 318340 50458 318392 50464
rect 458364 50516 458416 50522
rect 458364 50458 458416 50464
rect 314016 50380 314068 50386
rect 314016 50322 314068 50328
rect 458180 50380 458232 50386
rect 458180 50322 458232 50328
rect 308034 50280 308090 50289
rect 308034 50215 308090 50224
rect 131028 49020 131080 49026
rect 131028 48962 131080 48968
rect 131040 45506 131068 48962
rect 131580 47864 131632 47870
rect 131580 47806 131632 47812
rect 131040 45478 131344 45506
rect 131316 45422 131344 45478
rect 131304 45416 131356 45422
rect 131304 45358 131356 45364
rect 130936 45348 130988 45354
rect 130936 45290 130988 45296
rect 130948 45122 130976 45290
rect 130936 45116 130988 45122
rect 130936 45058 130988 45064
rect 131396 44736 131448 44742
rect 131396 44678 131448 44684
rect 130566 44432 130622 44441
rect 130566 44367 130622 44376
rect 131408 44198 131436 44678
rect 131592 44334 131620 47806
rect 458192 47025 458220 50322
rect 458178 47016 458234 47025
rect 458178 46951 458234 46960
rect 458376 46753 458404 50458
rect 544028 50386 544056 53108
rect 545684 53094 546020 53122
rect 547892 53094 548044 53122
rect 522948 50380 523000 50386
rect 522948 50322 523000 50328
rect 544016 50380 544068 50386
rect 544016 50322 544068 50328
rect 522960 47841 522988 50322
rect 522946 47832 523002 47841
rect 522946 47767 523002 47776
rect 459172 47654 459232 47682
rect 459632 47654 459968 47682
rect 460092 47654 460152 47682
rect 460552 47654 460888 47682
rect 461012 47654 461164 47682
rect 461472 47654 461808 47682
rect 461932 47654 461992 47682
rect 458362 46744 458418 46753
rect 142370 46702 142660 46730
rect 132040 46096 132092 46102
rect 132040 46038 132092 46044
rect 131580 44328 131632 44334
rect 131580 44270 131632 44276
rect 132052 44266 132080 46038
rect 132224 45552 132276 45558
rect 132224 45494 132276 45500
rect 132236 44266 132264 45494
rect 132960 45416 133012 45422
rect 132960 45358 133012 45364
rect 132590 44432 132646 44441
rect 132590 44367 132592 44376
rect 132644 44367 132646 44376
rect 132592 44358 132644 44364
rect 132972 44310 133000 45358
rect 132960 44304 133012 44310
rect 142632 44305 142660 46702
rect 458362 46679 458418 46688
rect 459204 44441 459232 47654
rect 459190 44432 459246 44441
rect 459190 44367 459246 44376
rect 132040 44260 132092 44266
rect 132040 44202 132092 44208
rect 132224 44260 132276 44266
rect 132960 44246 133012 44252
rect 142618 44296 142674 44305
rect 142618 44231 142674 44240
rect 132224 44202 132276 44208
rect 131396 44192 131448 44198
rect 131396 44134 131448 44140
rect 255870 44160 255926 44169
rect 255870 44095 255926 44104
rect 129372 44056 129424 44062
rect 129372 43998 129424 44004
rect 255884 42838 255912 44095
rect 307298 43888 307354 43897
rect 307298 43823 307354 43832
rect 440238 43888 440294 43897
rect 440238 43823 440240 43832
rect 187332 42832 187384 42838
rect 187332 42774 187384 42780
rect 255872 42832 255924 42838
rect 255872 42774 255924 42780
rect 187344 42092 187372 42774
rect 194322 42120 194378 42129
rect 194074 42078 194322 42106
rect 307312 42106 307340 43823
rect 440292 43823 440294 43832
rect 441066 43888 441122 43897
rect 441066 43823 441068 43832
rect 440240 43794 440292 43800
rect 441120 43823 441122 43832
rect 441068 43794 441120 43800
rect 410892 42900 410944 42906
rect 410892 42842 410944 42848
rect 415584 42900 415636 42906
rect 415584 42842 415636 42848
rect 310428 42764 310480 42770
rect 310428 42706 310480 42712
rect 364524 42764 364576 42770
rect 364524 42706 364576 42712
rect 310440 42106 310468 42706
rect 361764 42492 361816 42498
rect 361764 42434 361816 42440
rect 307004 42078 307340 42106
rect 310132 42078 310468 42106
rect 361776 42092 361804 42434
rect 364536 42362 364564 42706
rect 364892 42628 364944 42634
rect 364892 42570 364944 42576
rect 364524 42356 364576 42362
rect 364524 42298 364576 42304
rect 364904 42092 364932 42570
rect 410904 42498 410932 42842
rect 410892 42492 410944 42498
rect 410892 42434 410944 42440
rect 415596 42362 415624 42842
rect 431224 42764 431276 42770
rect 431224 42706 431276 42712
rect 441068 42764 441120 42770
rect 441068 42706 441120 42712
rect 449164 42764 449216 42770
rect 449164 42706 449216 42712
rect 453580 42764 453632 42770
rect 453580 42706 453632 42712
rect 427084 42628 427136 42634
rect 427084 42570 427136 42576
rect 416594 42392 416650 42401
rect 415584 42356 415636 42362
rect 416594 42327 416650 42336
rect 415584 42298 415636 42304
rect 415766 42120 415822 42129
rect 415426 42078 415766 42106
rect 194322 42055 194378 42064
rect 416608 42092 416636 42327
rect 415766 42055 415822 42064
rect 427096 42022 427124 42570
rect 429108 42492 429160 42498
rect 429108 42434 429160 42440
rect 427084 42016 427136 42022
rect 427084 41958 427136 41964
rect 405646 41848 405702 41857
rect 405582 41806 405646 41834
rect 419906 41848 419962 41857
rect 419750 41806 419906 41834
rect 405646 41783 405702 41792
rect 419906 41783 419962 41792
rect 429120 41750 429148 42434
rect 431236 42022 431264 42706
rect 441080 42022 441108 42706
rect 441252 42628 441304 42634
rect 441252 42570 441304 42576
rect 446404 42628 446456 42634
rect 446404 42570 446456 42576
rect 431224 42016 431276 42022
rect 431224 41958 431276 41964
rect 441068 42016 441120 42022
rect 441068 41958 441120 41964
rect 441264 41886 441292 42570
rect 446218 42256 446274 42265
rect 446218 42191 446274 42200
rect 441252 41880 441304 41886
rect 441252 41822 441304 41828
rect 429108 41744 429160 41750
rect 429108 41686 429160 41692
rect 446232 41585 446260 42191
rect 446416 42022 446444 42570
rect 446404 42016 446456 42022
rect 446404 41958 446456 41964
rect 449176 41750 449204 42706
rect 453592 41750 453620 42706
rect 454684 42628 454736 42634
rect 454684 42570 454736 42576
rect 454500 42492 454552 42498
rect 454500 42434 454552 42440
rect 454512 42022 454540 42434
rect 454500 42016 454552 42022
rect 454500 41958 454552 41964
rect 454696 41886 454724 42570
rect 459940 42106 459968 47654
rect 460124 44169 460152 47654
rect 460110 44160 460166 44169
rect 460110 44095 460166 44104
rect 460860 43489 460888 47654
rect 460846 43480 460902 43489
rect 460846 43415 460902 43424
rect 461136 42265 461164 47654
rect 461780 42945 461808 47654
rect 461964 44441 461992 47654
rect 462378 47410 462406 47668
rect 462332 47382 462406 47410
rect 462516 47654 462852 47682
rect 462976 47654 463312 47682
rect 461950 44432 462006 44441
rect 461950 44367 462006 44376
rect 462332 43217 462360 47382
rect 462516 44441 462544 47654
rect 462502 44432 462558 44441
rect 462502 44367 462558 44376
rect 462318 43208 462374 43217
rect 462318 43143 462374 43152
rect 461766 42936 461822 42945
rect 461766 42871 461822 42880
rect 462976 42634 463004 47654
rect 463758 47410 463786 47668
rect 463712 47382 463786 47410
rect 463896 47654 464232 47682
rect 464356 47654 464692 47682
rect 462964 42628 463016 42634
rect 462964 42570 463016 42576
rect 463712 42498 463740 47382
rect 463896 44169 463924 47654
rect 463882 44160 463938 44169
rect 463882 44095 463938 44104
rect 463974 42936 464030 42945
rect 463974 42871 464030 42880
rect 463988 42514 464016 42871
rect 464356 42770 464384 47654
rect 465138 47410 465166 47668
rect 465092 47382 465166 47410
rect 465276 47654 465612 47682
rect 465092 46753 465120 47382
rect 465276 47025 465304 47654
rect 545684 47297 545712 53094
rect 547892 47569 547920 53094
rect 550008 48929 550036 53108
rect 549994 48920 550050 48929
rect 549994 48855 550050 48864
rect 552032 47841 552060 53108
rect 553688 53094 554024 53122
rect 553688 48113 553716 53094
rect 553674 48104 553730 48113
rect 553674 48039 553730 48048
rect 552018 47832 552074 47841
rect 552018 47767 552074 47776
rect 547878 47560 547934 47569
rect 547878 47495 547934 47504
rect 545670 47288 545726 47297
rect 545670 47223 545726 47232
rect 465262 47016 465318 47025
rect 465262 46951 465318 46960
rect 465078 46744 465134 46753
rect 465078 46679 465134 46688
rect 626000 46510 626028 66846
rect 647344 64433 647372 80786
rect 648620 79348 648672 79354
rect 648620 79290 648672 79296
rect 647514 78160 647570 78169
rect 647514 78095 647570 78104
rect 647330 64424 647386 64433
rect 647330 64359 647386 64368
rect 647528 57361 647556 78095
rect 648632 59265 648660 79290
rect 648988 76832 649040 76838
rect 648988 76774 649040 76780
rect 649000 62121 649028 76774
rect 662420 76696 662472 76702
rect 662420 76638 662472 76644
rect 648986 62112 649042 62121
rect 648986 62047 649042 62056
rect 648618 59256 648674 59265
rect 648618 59191 648674 59200
rect 647514 57352 647570 57361
rect 647514 57287 647570 57296
rect 661590 48510 661646 48519
rect 661590 48445 661646 48454
rect 625988 46504 626040 46510
rect 625988 46446 626040 46452
rect 661604 45554 661632 48445
rect 661774 47789 661830 47798
rect 661774 47724 661830 47733
rect 661788 46510 661816 47724
rect 662432 47433 662460 76638
rect 666572 75206 666600 103486
rect 667938 102776 667994 102785
rect 667938 102711 667994 102720
rect 667952 100026 667980 102711
rect 667940 100020 667992 100026
rect 667940 99962 667992 99968
rect 668136 95946 668164 106111
rect 668308 104848 668360 104854
rect 668308 104790 668360 104796
rect 668320 104417 668348 104790
rect 668306 104408 668362 104417
rect 668306 104343 668362 104352
rect 668124 95940 668176 95946
rect 668124 95882 668176 95888
rect 668320 84194 668348 104343
rect 668596 102785 668624 127735
rect 668780 125769 668808 128590
rect 668950 126984 669006 126993
rect 668950 126919 669006 126928
rect 668766 125760 668822 125769
rect 668766 125695 668822 125704
rect 668964 120873 668992 126919
rect 668950 120864 669006 120873
rect 668950 120799 669006 120808
rect 668766 120592 668822 120601
rect 668766 120527 668822 120536
rect 668780 111081 668808 120527
rect 669042 116512 669098 116521
rect 669042 116447 669098 116456
rect 669056 114345 669084 116447
rect 669226 115832 669282 115841
rect 669226 115767 669282 115776
rect 669240 114617 669268 115767
rect 669226 114608 669282 114617
rect 669226 114543 669282 114552
rect 669042 114336 669098 114345
rect 669042 114271 669098 114280
rect 669226 114336 669282 114345
rect 669226 114271 669282 114280
rect 669240 112713 669268 114271
rect 669226 112704 669282 112713
rect 669226 112639 669282 112648
rect 668766 111072 668822 111081
rect 668766 111007 668822 111016
rect 670160 108050 670188 130863
rect 670804 128654 670832 137986
rect 671342 131744 671398 131753
rect 671342 131679 671398 131688
rect 670792 128648 670844 128654
rect 670792 128590 670844 128596
rect 671356 109034 671384 131679
rect 671526 129296 671582 129305
rect 671526 129231 671582 129240
rect 671540 109034 671568 129231
rect 672092 124137 672120 213279
rect 672262 212120 672318 212129
rect 672262 212055 672318 212064
rect 672276 126993 672304 212055
rect 672460 206961 672488 287642
rect 672920 287054 672948 324935
rect 673196 310049 673224 354583
rect 673380 310865 673408 355399
rect 673734 351384 673790 351393
rect 673734 351319 673790 351328
rect 673748 338065 673776 351319
rect 673932 351121 673960 358255
rect 674392 356561 674420 364306
rect 674378 356552 674434 356561
rect 674378 356487 674434 356496
rect 674102 356280 674158 356289
rect 674102 356215 674158 356224
rect 673918 351112 673974 351121
rect 673918 351047 673974 351056
rect 674116 350962 674144 356215
rect 674654 352200 674710 352209
rect 674654 352135 674710 352144
rect 673932 350934 674144 350962
rect 674470 350976 674526 350985
rect 673734 338056 673790 338065
rect 673734 337991 673790 338000
rect 673932 325694 673960 350934
rect 674470 350911 674526 350920
rect 674484 350690 674512 350911
rect 674116 350662 674512 350690
rect 674116 336546 674144 350662
rect 674470 350568 674526 350577
rect 674470 350503 674526 350512
rect 674286 349752 674342 349761
rect 674286 349687 674342 349696
rect 674300 340874 674328 349687
rect 674300 340846 674420 340874
rect 674392 336734 674420 340846
rect 674484 338114 674512 350503
rect 674668 338114 674696 352135
rect 675220 345001 675248 364306
rect 703694 359380 703722 359516
rect 704154 359380 704182 359516
rect 704614 359380 704642 359516
rect 705074 359380 705102 359516
rect 705534 359380 705562 359516
rect 705994 359380 706022 359516
rect 706454 359380 706482 359516
rect 706914 359380 706942 359516
rect 707374 359380 707402 359516
rect 707834 359380 707862 359516
rect 708294 359380 708322 359516
rect 708754 359380 708782 359516
rect 709214 359380 709242 359516
rect 675942 357912 675998 357921
rect 675942 357847 675998 357856
rect 675956 356833 675984 357847
rect 675942 356824 675998 356833
rect 675942 356759 675998 356768
rect 676034 350160 676090 350169
rect 676034 350095 676090 350104
rect 676048 346633 676076 350095
rect 676034 346624 676090 346633
rect 676034 346559 676090 346568
rect 675206 344992 675262 345001
rect 675206 344927 675262 344936
rect 674944 341074 675418 341102
rect 674944 338745 674972 341074
rect 675114 340776 675170 340785
rect 675114 340711 675170 340720
rect 675128 340558 675156 340711
rect 675128 340530 675340 340558
rect 675312 340490 675340 340530
rect 675404 340490 675432 340544
rect 675312 340462 675432 340490
rect 675758 340368 675814 340377
rect 675758 340303 675814 340312
rect 675772 339864 675800 340303
rect 675482 339416 675538 339425
rect 675482 339351 675538 339360
rect 675496 339252 675524 339351
rect 674930 338736 674986 338745
rect 674930 338671 674986 338680
rect 674484 338086 674604 338114
rect 674668 338086 674788 338114
rect 674380 336728 674432 336734
rect 674380 336670 674432 336676
rect 674116 336530 674420 336546
rect 674116 336524 674432 336530
rect 674116 336518 674380 336524
rect 674380 336466 674432 336472
rect 674576 331889 674604 338086
rect 674484 331861 674604 331889
rect 674484 331158 674512 331861
rect 674472 331152 674524 331158
rect 674472 331094 674524 331100
rect 674760 328454 674788 338086
rect 675114 338056 675170 338065
rect 675114 337991 675170 338000
rect 675128 336857 675156 337991
rect 675758 337920 675814 337929
rect 675758 337855 675814 337864
rect 675772 337416 675800 337855
rect 675128 336829 675418 336857
rect 675116 336728 675168 336734
rect 675116 336670 675168 336676
rect 675128 335594 675156 336670
rect 675300 336524 675352 336530
rect 675300 336466 675352 336472
rect 675312 336206 675340 336466
rect 675312 336178 675418 336206
rect 675128 335566 675340 335594
rect 675312 335458 675340 335566
rect 675404 335458 675432 335580
rect 675312 335430 675432 335458
rect 675298 335336 675354 335345
rect 675298 335271 675354 335280
rect 675312 331889 675340 335271
rect 675482 333432 675538 333441
rect 675482 333367 675538 333376
rect 675496 333064 675524 333367
rect 675482 332752 675538 332761
rect 675482 332687 675538 332696
rect 675496 332520 675524 332687
rect 675312 331861 675418 331889
rect 675114 331256 675170 331265
rect 675170 331214 675418 331242
rect 675114 331191 675170 331200
rect 675300 331152 675352 331158
rect 675300 331094 675352 331100
rect 675312 330049 675340 331094
rect 675312 330021 675418 330049
rect 674668 328426 674788 328454
rect 674668 326913 674696 328426
rect 675312 328222 675432 328250
rect 675312 328182 675340 328222
rect 675220 328154 675340 328182
rect 675404 328168 675432 328222
rect 675022 327992 675078 328001
rect 675022 327927 675078 327936
rect 674654 326904 674710 326913
rect 674654 326839 674710 326848
rect 673932 325666 674420 325694
rect 674392 311681 674420 325666
rect 675036 325009 675064 327927
rect 675220 325689 675248 328154
rect 675390 327992 675446 328001
rect 675390 327927 675446 327936
rect 675404 327556 675432 327927
rect 675390 326904 675446 326913
rect 675390 326839 675446 326848
rect 675404 326332 675432 326839
rect 675206 325680 675262 325689
rect 675206 325615 675262 325624
rect 675022 325000 675078 325009
rect 675022 324935 675078 324944
rect 703694 314364 703722 314500
rect 704154 314364 704182 314500
rect 704614 314364 704642 314500
rect 705074 314364 705102 314500
rect 705534 314364 705562 314500
rect 705994 314364 706022 314500
rect 706454 314364 706482 314500
rect 706914 314364 706942 314500
rect 707374 314364 707402 314500
rect 707834 314364 707862 314500
rect 708294 314364 708322 314500
rect 708754 314364 708782 314500
rect 709214 314364 709242 314500
rect 676034 313304 676090 313313
rect 676090 313262 676260 313290
rect 676034 313239 676090 313248
rect 674838 312896 674894 312905
rect 674838 312831 674894 312840
rect 674564 312044 674616 312050
rect 674564 311986 674616 311992
rect 674378 311672 674434 311681
rect 674378 311607 674434 311616
rect 673366 310856 673422 310865
rect 673366 310791 673422 310800
rect 673918 310448 673974 310457
rect 673918 310383 673974 310392
rect 673182 310040 673238 310049
rect 673182 309975 673238 309984
rect 673366 309632 673422 309641
rect 673366 309567 673422 309576
rect 673182 303920 673238 303929
rect 673182 303855 673238 303864
rect 672644 287026 672948 287054
rect 672644 278594 672672 287026
rect 673196 286521 673224 303855
rect 673182 286512 673238 286521
rect 673182 286447 673238 286456
rect 672814 285696 672870 285705
rect 672814 285631 672870 285640
rect 672632 278588 672684 278594
rect 672632 278530 672684 278536
rect 672828 277394 672856 285631
rect 672736 277366 672856 277394
rect 672736 229786 672764 277366
rect 672998 266112 673054 266121
rect 672998 266047 673054 266056
rect 673012 244274 673040 266047
rect 673380 265033 673408 309567
rect 673734 305960 673790 305969
rect 673734 305895 673790 305904
rect 673748 291553 673776 305895
rect 673734 291544 673790 291553
rect 673734 291479 673790 291488
rect 673550 290456 673606 290465
rect 673550 290391 673606 290400
rect 673564 287054 673592 290391
rect 673564 287026 673684 287054
rect 673656 268161 673684 287026
rect 673642 268152 673698 268161
rect 673642 268087 673698 268096
rect 673932 265849 673960 310383
rect 674576 307034 674604 311986
rect 674852 311953 674880 312831
rect 675482 312080 675538 312089
rect 675482 312015 675484 312024
rect 675536 312015 675538 312024
rect 675484 311986 675536 311992
rect 674838 311944 674894 311953
rect 674838 311879 674894 311888
rect 674746 311400 674802 311409
rect 674746 311335 674802 311344
rect 674208 307006 674604 307034
rect 674208 287054 674236 307006
rect 674760 306490 674788 311335
rect 675942 311128 675998 311137
rect 676232 311114 676260 313262
rect 675998 311086 676260 311114
rect 675942 311063 675998 311072
rect 675022 309224 675078 309233
rect 675022 309159 675078 309168
rect 674668 306462 674788 306490
rect 674378 305552 674434 305561
rect 674378 305487 674434 305496
rect 674392 303634 674420 305487
rect 674300 303606 674420 303634
rect 674300 292574 674328 303606
rect 674470 303512 674526 303521
rect 674470 303447 674526 303456
rect 674484 300801 674512 303447
rect 674470 300792 674526 300801
rect 674470 300727 674526 300736
rect 674472 295724 674524 295730
rect 674472 295666 674524 295672
rect 674484 293865 674512 295666
rect 674470 293856 674526 293865
rect 674470 293791 674526 293800
rect 674300 292546 674512 292574
rect 674208 287026 674420 287054
rect 674392 267481 674420 287026
rect 674484 285070 674512 292546
rect 674668 285190 674696 306462
rect 674840 306400 674892 306406
rect 674840 306342 674892 306348
rect 674852 302234 674880 306342
rect 674852 302206 674972 302234
rect 674944 299418 674972 302206
rect 674852 299390 674972 299418
rect 674852 297401 674880 299390
rect 674838 297392 674894 297401
rect 675036 297362 675064 309159
rect 676678 308408 676734 308417
rect 676678 308343 676734 308352
rect 675482 308000 675538 308009
rect 675482 307935 675538 307944
rect 675496 306406 675524 307935
rect 676034 307592 676090 307601
rect 676090 307550 676444 307578
rect 676034 307527 676090 307536
rect 676034 307184 676090 307193
rect 676090 307142 676260 307170
rect 676034 307119 676090 307128
rect 676232 306406 676260 307142
rect 675484 306400 675536 306406
rect 675484 306342 675536 306348
rect 676220 306400 676272 306406
rect 676220 306342 676272 306348
rect 676416 304910 676444 307550
rect 675852 304904 675904 304910
rect 675852 304846 675904 304852
rect 676404 304904 676456 304910
rect 676404 304846 676456 304852
rect 675864 302234 675892 304846
rect 676402 304736 676458 304745
rect 676402 304671 676458 304680
rect 675128 302206 675892 302234
rect 675128 297514 675156 302206
rect 676416 301617 676444 304671
rect 676402 301608 676458 301617
rect 676402 301543 676458 301552
rect 676692 301481 676720 308343
rect 678242 306776 678298 306785
rect 678242 306711 678298 306720
rect 676864 306400 676916 306406
rect 676864 306342 676916 306348
rect 676678 301472 676734 301481
rect 676678 301407 676734 301416
rect 676128 298104 676180 298110
rect 676128 298046 676180 298052
rect 675944 297968 675996 297974
rect 675944 297910 675996 297916
rect 675128 297486 675248 297514
rect 674838 297327 674894 297336
rect 675024 297356 675076 297362
rect 675024 297298 675076 297304
rect 675220 297158 675248 297486
rect 675208 297152 675260 297158
rect 675208 297094 675260 297100
rect 675024 297016 675076 297022
rect 675024 296958 675076 296964
rect 675206 296984 675262 296993
rect 674840 296880 674892 296886
rect 674840 296822 674892 296828
rect 674852 288062 674880 296822
rect 675036 295202 675064 296958
rect 675206 296919 675262 296928
rect 675220 295338 675248 296919
rect 675956 296585 675984 297910
rect 676140 296993 676168 298046
rect 676876 297401 676904 306342
rect 678256 298110 678284 306711
rect 678978 306368 679034 306377
rect 678978 306303 679034 306312
rect 678992 298110 679020 306303
rect 678244 298104 678296 298110
rect 678244 298046 678296 298052
rect 678980 298104 679032 298110
rect 678980 298046 679032 298052
rect 676862 297392 676918 297401
rect 676862 297327 676918 297336
rect 676126 296984 676182 296993
rect 676126 296919 676182 296928
rect 675942 296576 675998 296585
rect 675942 296511 675998 296520
rect 675496 295730 675524 296072
rect 675758 295760 675814 295769
rect 675484 295724 675536 295730
rect 675758 295695 675814 295704
rect 675484 295666 675536 295672
rect 675772 295528 675800 295695
rect 675220 295310 675432 295338
rect 675036 295174 675340 295202
rect 675312 294250 675340 295174
rect 675404 294879 675432 295310
rect 675312 294222 675418 294250
rect 675390 292904 675446 292913
rect 675390 292839 675446 292848
rect 675404 292400 675432 292839
rect 675574 292224 675630 292233
rect 675574 292159 675630 292168
rect 675588 291856 675616 292159
rect 675482 291544 675538 291553
rect 675482 291479 675538 291488
rect 675496 291176 675524 291479
rect 675758 291000 675814 291009
rect 675758 290935 675814 290944
rect 675772 290564 675800 290935
rect 675312 288102 675432 288130
rect 675312 288062 675340 288102
rect 674852 288034 675340 288062
rect 675404 288048 675432 288102
rect 675114 287872 675170 287881
rect 675114 287807 675170 287816
rect 675128 287518 675156 287807
rect 675128 287490 675418 287518
rect 675758 287056 675814 287065
rect 675758 286991 675814 287000
rect 675772 286892 675800 286991
rect 675390 286512 675446 286521
rect 675390 286447 675446 286456
rect 675404 286212 675432 286447
rect 674656 285184 674708 285190
rect 674656 285126 674708 285132
rect 674484 285042 675340 285070
rect 675312 285002 675340 285042
rect 675404 285002 675432 285056
rect 674656 284980 674708 284986
rect 675312 284974 675432 285002
rect 674656 284922 674708 284928
rect 674378 267472 674434 267481
rect 674378 267407 674434 267416
rect 674470 267064 674526 267073
rect 674470 266999 674526 267008
rect 673918 265840 673974 265849
rect 673918 265775 673974 265784
rect 673918 265432 673974 265441
rect 673918 265367 673974 265376
rect 673366 265024 673422 265033
rect 673366 264959 673422 264968
rect 673550 261624 673606 261633
rect 673550 261559 673606 261568
rect 673182 259312 673238 259321
rect 673182 259247 673238 259256
rect 672828 244246 673040 244274
rect 672828 234614 672856 244246
rect 673196 242729 673224 259247
rect 673564 247081 673592 261559
rect 673734 258904 673790 258913
rect 673734 258839 673790 258848
rect 673550 247072 673606 247081
rect 673550 247007 673606 247016
rect 673182 242720 673238 242729
rect 673182 242655 673238 242664
rect 673748 241505 673776 258839
rect 673734 241496 673790 241505
rect 673734 241431 673790 241440
rect 672954 236768 673006 236774
rect 673182 236736 673238 236745
rect 673006 236716 673182 236722
rect 672954 236710 673182 236716
rect 672966 236694 673182 236710
rect 673182 236671 673238 236680
rect 673184 236496 673236 236502
rect 673236 236444 673868 236450
rect 673184 236438 673868 236444
rect 673196 236422 673868 236438
rect 673642 236328 673698 236337
rect 673642 236263 673698 236272
rect 673092 236224 673144 236230
rect 673144 236172 673500 236178
rect 673092 236166 673500 236172
rect 673104 236150 673500 236166
rect 673472 235226 673500 236150
rect 673472 235198 673568 235226
rect 673540 234954 673568 235198
rect 673472 234926 673568 234954
rect 672828 234586 673040 234614
rect 672736 229758 672948 229786
rect 672724 226432 672776 226438
rect 672722 226400 672724 226409
rect 672776 226400 672778 226409
rect 672722 226335 672778 226344
rect 672604 226160 672656 226166
rect 672602 226128 672604 226137
rect 672656 226128 672658 226137
rect 672602 226063 672658 226072
rect 672920 215294 672948 229758
rect 673012 224954 673040 234586
rect 673472 230602 673500 234926
rect 673288 230574 673500 230602
rect 673288 230058 673316 230574
rect 673460 230444 673512 230450
rect 673460 230386 673512 230392
rect 673472 230217 673500 230386
rect 673458 230208 673514 230217
rect 673458 230143 673514 230152
rect 673288 230030 673500 230058
rect 673472 227050 673500 230030
rect 673656 229242 673684 236263
rect 673840 229786 673868 236422
rect 673932 229922 673960 265367
rect 674102 264616 674158 264625
rect 674102 264551 674158 264560
rect 674116 235249 674144 264551
rect 674484 263594 674512 266999
rect 674668 266665 674696 284922
rect 675758 283656 675814 283665
rect 675758 283591 675814 283600
rect 675772 283220 675800 283591
rect 675666 282704 675722 282713
rect 675666 282639 675722 282648
rect 675680 282554 675708 282639
rect 675128 282540 675708 282554
rect 675128 282526 675694 282540
rect 675128 278361 675156 282526
rect 675666 281616 675722 281625
rect 675666 281551 675722 281560
rect 675680 281355 675708 281551
rect 676862 279440 676918 279449
rect 676862 279375 676918 279384
rect 675114 278352 675170 278361
rect 675114 278287 675170 278296
rect 676876 268569 676904 279375
rect 703694 269348 703722 269484
rect 704154 269348 704182 269484
rect 704614 269348 704642 269484
rect 705074 269348 705102 269484
rect 705534 269348 705562 269484
rect 705994 269348 706022 269484
rect 706454 269348 706482 269484
rect 706914 269348 706942 269484
rect 707374 269348 707402 269484
rect 707834 269348 707862 269484
rect 708294 269348 708322 269484
rect 708754 269348 708782 269484
rect 709214 269348 709242 269484
rect 676862 268560 676918 268569
rect 676862 268495 676918 268504
rect 676218 268152 676274 268161
rect 676218 268087 676274 268096
rect 676232 267753 676260 268087
rect 676218 267744 676274 267753
rect 676218 267679 676274 267688
rect 674654 266656 674710 266665
rect 674654 266591 674710 266600
rect 675482 264072 675538 264081
rect 675482 264007 675538 264016
rect 675496 263594 675524 264007
rect 676218 263664 676274 263673
rect 676218 263599 676274 263608
rect 674484 263566 674696 263594
rect 674470 262576 674526 262585
rect 674470 262511 674526 262520
rect 674286 260128 674342 260137
rect 674286 260063 674342 260072
rect 674300 243522 674328 260063
rect 674484 243710 674512 262511
rect 674472 243704 674524 243710
rect 674472 243646 674524 243652
rect 674300 243494 674420 243522
rect 674392 242894 674420 243494
rect 674380 242888 674432 242894
rect 674380 242830 674432 242836
rect 674102 235240 674158 235249
rect 674102 235175 674158 235184
rect 674102 230480 674158 230489
rect 674102 230415 674158 230424
rect 674286 230480 674342 230489
rect 674286 230415 674342 230424
rect 674116 230042 674144 230415
rect 674300 230246 674328 230415
rect 674288 230240 674340 230246
rect 674288 230182 674340 230188
rect 674470 230208 674526 230217
rect 674470 230143 674526 230152
rect 674484 230058 674512 230143
rect 674104 230036 674156 230042
rect 674104 229978 674156 229984
rect 674346 230030 674512 230058
rect 673932 229894 674052 229922
rect 673840 229758 673960 229786
rect 673564 229214 673684 229242
rect 673564 227882 673592 229214
rect 673736 229152 673788 229158
rect 673736 229094 673788 229100
rect 673748 228585 673776 229094
rect 673734 228576 673790 228585
rect 673734 228511 673790 228520
rect 673564 227854 673684 227882
rect 673656 227798 673684 227854
rect 673644 227792 673696 227798
rect 673644 227734 673696 227740
rect 673460 227044 673512 227050
rect 673460 226986 673512 226992
rect 673552 226840 673604 226846
rect 673552 226782 673604 226788
rect 673012 224926 673132 224954
rect 673104 221513 673132 224926
rect 673090 221504 673146 221513
rect 673090 221439 673146 221448
rect 673564 220153 673592 226782
rect 673736 226568 673788 226574
rect 673734 226536 673736 226545
rect 673788 226536 673790 226545
rect 673734 226471 673790 226480
rect 673734 221912 673790 221921
rect 673734 221847 673790 221856
rect 673550 220144 673606 220153
rect 673550 220079 673606 220088
rect 673182 217560 673238 217569
rect 673182 217495 673238 217504
rect 672736 215266 672948 215294
rect 672446 206952 672502 206961
rect 672446 206887 672502 206896
rect 672538 203008 672594 203017
rect 672538 202943 672594 202952
rect 672552 182073 672580 202943
rect 672538 182064 672594 182073
rect 672538 181999 672594 182008
rect 672736 177721 672764 215266
rect 672998 214568 673054 214577
rect 672998 214503 673054 214512
rect 673012 200569 673040 214503
rect 672998 200560 673054 200569
rect 672998 200495 673054 200504
rect 673196 195265 673224 217495
rect 673366 217016 673422 217025
rect 673366 216951 673422 216960
rect 673182 195256 673238 195265
rect 673182 195191 673238 195200
rect 673380 191185 673408 216951
rect 673550 214976 673606 214985
rect 673550 214911 673606 214920
rect 673564 197169 673592 214911
rect 673550 197160 673606 197169
rect 673550 197095 673606 197104
rect 673366 191176 673422 191185
rect 673366 191111 673422 191120
rect 673748 180794 673776 221847
rect 673932 215294 673960 229758
rect 674024 224954 674052 229894
rect 674346 229838 674374 230030
rect 674452 229968 674504 229974
rect 674452 229910 674504 229916
rect 674334 229832 674386 229838
rect 674334 229774 674386 229780
rect 674464 229650 674492 229910
rect 674464 229622 674512 229650
rect 674242 229560 674294 229566
rect 674242 229502 674294 229508
rect 674254 229242 674282 229502
rect 674484 229401 674512 229622
rect 674470 229392 674526 229401
rect 674470 229327 674526 229336
rect 674254 229214 674328 229242
rect 674300 224954 674328 229214
rect 674024 224926 674144 224954
rect 674300 224926 674512 224954
rect 674116 220697 674144 224926
rect 674102 220688 674158 220697
rect 674102 220623 674158 220632
rect 674102 220144 674158 220153
rect 674102 220079 674158 220088
rect 673656 180766 673776 180794
rect 673840 215266 673960 215294
rect 672722 177712 672778 177721
rect 672722 177647 672778 177656
rect 673656 177313 673684 180766
rect 673642 177304 673698 177313
rect 673642 177239 673698 177248
rect 673642 176896 673698 176905
rect 673642 176831 673698 176840
rect 672538 175264 672594 175273
rect 672538 175199 672594 175208
rect 672552 130529 672580 175199
rect 673366 174448 673422 174457
rect 673366 174383 673422 174392
rect 672998 169552 673054 169561
rect 672998 169487 673054 169496
rect 672722 168328 672778 168337
rect 672722 168263 672778 168272
rect 672538 130520 672594 130529
rect 672538 130455 672594 130464
rect 672262 126984 672318 126993
rect 672262 126919 672318 126928
rect 672078 124128 672134 124137
rect 672078 124063 672134 124072
rect 672538 122904 672594 122913
rect 672538 122839 672594 122848
rect 672078 121680 672134 121689
rect 672078 121615 672134 121624
rect 672092 114345 672120 121615
rect 672552 116521 672580 122839
rect 672736 119241 672764 168263
rect 673012 155553 673040 169487
rect 673182 168736 673238 168745
rect 673182 168671 673238 168680
rect 672998 155544 673054 155553
rect 672998 155479 673054 155488
rect 673196 151065 673224 168671
rect 673182 151056 673238 151065
rect 673182 150991 673238 151000
rect 673380 129713 673408 174383
rect 673656 132161 673684 176831
rect 673840 160449 673868 215266
rect 674116 178537 674144 220079
rect 674286 213752 674342 213761
rect 674286 213687 674342 213696
rect 674300 196081 674328 213687
rect 674484 213081 674512 224926
rect 674668 222329 674696 263566
rect 674852 263566 675524 263594
rect 674852 250646 674880 263566
rect 676232 261225 676260 263599
rect 679622 263256 679678 263265
rect 679622 263191 679678 263200
rect 676402 262848 676458 262857
rect 676402 262783 676458 262792
rect 676218 261216 676274 261225
rect 676218 261151 676274 261160
rect 676416 259486 676444 262783
rect 675852 259480 675904 259486
rect 675852 259422 675904 259428
rect 676404 259480 676456 259486
rect 676404 259422 676456 259428
rect 675864 255377 675892 259422
rect 675022 255368 675078 255377
rect 675022 255303 675078 255312
rect 675850 255368 675906 255377
rect 675850 255303 675906 255312
rect 674840 250640 674892 250646
rect 674840 250582 674892 250588
rect 674838 249928 674894 249937
rect 674838 249863 674894 249872
rect 674852 238649 674880 249863
rect 675036 249234 675064 255303
rect 679636 252550 679664 263191
rect 675852 252544 675904 252550
rect 675852 252486 675904 252492
rect 679624 252544 679676 252550
rect 679624 252486 679676 252492
rect 675864 251546 675892 252486
rect 675496 251518 675892 251546
rect 675496 251394 675524 251518
rect 675484 251388 675536 251394
rect 675484 251330 675536 251336
rect 675484 250776 675536 250782
rect 675680 250753 675708 251056
rect 675484 250718 675536 250724
rect 675666 250744 675722 250753
rect 675300 250640 675352 250646
rect 675300 250582 675352 250588
rect 675312 249642 675340 250582
rect 675496 250512 675524 250718
rect 675666 250679 675722 250688
rect 675758 250200 675814 250209
rect 675758 250135 675814 250144
rect 675772 249900 675800 250135
rect 675312 249614 675432 249642
rect 675036 249206 675340 249234
rect 675404 249220 675432 249614
rect 675114 248976 675170 248985
rect 675114 248911 675170 248920
rect 675128 247194 675156 248911
rect 675312 247398 675340 249206
rect 675312 247370 675418 247398
rect 674944 247166 675156 247194
rect 674944 239578 674972 247166
rect 675114 247072 675170 247081
rect 675114 247007 675170 247016
rect 675128 246854 675156 247007
rect 675128 246826 675418 246854
rect 675758 246664 675814 246673
rect 675758 246599 675814 246608
rect 675772 246199 675800 246599
rect 675114 245576 675170 245585
rect 675170 245534 675418 245562
rect 675114 245511 675170 245520
rect 675114 245304 675170 245313
rect 675114 245239 675170 245248
rect 675128 244274 675156 245239
rect 675036 244246 675156 244274
rect 675036 239850 675064 244246
rect 675208 243704 675260 243710
rect 675208 243646 675260 243652
rect 675220 243085 675248 243646
rect 675220 243057 675418 243085
rect 675208 242888 675260 242894
rect 675208 242830 675260 242836
rect 675220 241890 675248 242830
rect 675390 242720 675446 242729
rect 675390 242655 675446 242664
rect 675404 242519 675432 242655
rect 675220 241862 675418 241890
rect 675206 241496 675262 241505
rect 675206 241431 675262 241440
rect 675220 241245 675248 241431
rect 675220 241217 675418 241245
rect 675206 240272 675262 240281
rect 675206 240207 675262 240216
rect 675220 240054 675248 240207
rect 675220 240026 675418 240054
rect 675036 239822 675248 239850
rect 674944 239550 675064 239578
rect 674838 238640 674894 238649
rect 674838 238575 674894 238584
rect 675036 238105 675064 239550
rect 675022 238096 675078 238105
rect 675022 238031 675078 238040
rect 675220 236382 675248 239822
rect 675390 238640 675446 238649
rect 675390 238575 675446 238584
rect 675404 238204 675432 238575
rect 675390 238096 675446 238105
rect 675390 238031 675446 238040
rect 675404 237524 675432 238031
rect 675220 236354 675418 236382
rect 675850 235240 675906 235249
rect 675850 235175 675906 235184
rect 675864 233986 675892 235175
rect 683304 234048 683356 234054
rect 683304 233990 683356 233996
rect 675852 233980 675904 233986
rect 675852 233922 675904 233928
rect 675484 233912 675536 233918
rect 675536 233860 675892 233866
rect 675484 233854 675892 233860
rect 675496 233838 675892 233854
rect 675864 233782 675892 233838
rect 675852 233776 675904 233782
rect 675852 233718 675904 233724
rect 678244 233776 678296 233782
rect 678244 233718 678296 233724
rect 675496 232762 675892 232778
rect 675484 232756 675892 232762
rect 675536 232750 675892 232756
rect 675484 232698 675536 232704
rect 675864 232694 675892 232750
rect 675852 232688 675904 232694
rect 675852 232630 675904 232636
rect 675484 232416 675536 232422
rect 675852 232416 675904 232422
rect 675536 232364 675852 232370
rect 675484 232358 675904 232364
rect 675496 232342 675892 232358
rect 675392 231668 675444 231674
rect 675392 231610 675444 231616
rect 674932 231124 674984 231130
rect 674932 231066 674984 231072
rect 674944 228993 674972 231066
rect 674930 228984 674986 228993
rect 674930 228919 674986 228928
rect 675206 226536 675262 226545
rect 675206 226471 675262 226480
rect 674838 226128 674894 226137
rect 674838 226063 674894 226072
rect 674654 222320 674710 222329
rect 674654 222255 674710 222264
rect 674852 221241 674880 226063
rect 675022 225856 675078 225865
rect 675022 225791 675078 225800
rect 674838 221232 674894 221241
rect 674838 221167 674894 221176
rect 674654 220280 674710 220289
rect 674654 220215 674710 220224
rect 674668 219450 674696 220215
rect 675036 219881 675064 225791
rect 675220 222737 675248 226471
rect 675206 222728 675262 222737
rect 675206 222663 675262 222672
rect 675022 219872 675078 219881
rect 675022 219807 675078 219816
rect 675404 219722 675432 231610
rect 676954 230480 677010 230489
rect 676954 230415 677010 230424
rect 676218 230208 676274 230217
rect 676218 230143 676274 230152
rect 676036 226840 676088 226846
rect 676036 226782 676088 226788
rect 675666 225312 675722 225321
rect 675666 225247 675722 225256
rect 675680 224954 675708 225247
rect 674576 219422 674696 219450
rect 675128 219694 675432 219722
rect 675588 224926 675708 224954
rect 674576 215294 674604 219422
rect 674930 219056 674986 219065
rect 674930 218991 674986 219000
rect 674746 216200 674802 216209
rect 674746 216135 674802 216144
rect 674576 215266 674696 215294
rect 674470 213072 674526 213081
rect 674470 213007 674526 213016
rect 674668 212534 674696 215266
rect 674392 212506 674696 212534
rect 674392 211154 674420 212506
rect 674392 211126 674512 211154
rect 674484 201494 674512 211126
rect 674760 201929 674788 216135
rect 674944 215294 674972 218991
rect 675128 218362 675156 219694
rect 675390 218648 675446 218657
rect 675588 218634 675616 224926
rect 676048 223145 676076 226782
rect 676034 223136 676090 223145
rect 676034 223071 676090 223080
rect 676034 221096 676090 221105
rect 676034 221031 676090 221040
rect 675446 218606 675616 218634
rect 675390 218583 675446 218592
rect 675128 218334 675524 218362
rect 675298 218240 675354 218249
rect 675298 218175 675354 218184
rect 674852 215266 674972 215294
rect 674852 204049 674880 215266
rect 675312 205337 675340 218175
rect 675496 211449 675524 218334
rect 675852 218000 675904 218006
rect 675666 217968 675722 217977
rect 675722 217948 675852 217954
rect 675722 217942 675904 217948
rect 675722 217926 675892 217942
rect 675666 217903 675722 217912
rect 676048 217569 676076 221031
rect 676034 217560 676090 217569
rect 676034 217495 676090 217504
rect 675852 216504 675904 216510
rect 675666 216472 675722 216481
rect 675722 216452 675852 216458
rect 675722 216446 675904 216452
rect 675722 216430 675892 216446
rect 675666 216407 675722 216416
rect 676034 215384 676090 215393
rect 676034 215319 676036 215328
rect 676088 215319 676090 215328
rect 676036 215290 676088 215296
rect 675666 215248 675722 215257
rect 676232 215234 676260 230143
rect 676678 228576 676734 228585
rect 676678 228511 676734 228520
rect 676692 218006 676720 228511
rect 676680 218000 676732 218006
rect 676680 217942 676732 217948
rect 676968 216510 676996 230415
rect 678256 226846 678284 233718
rect 679256 232416 679308 232422
rect 679256 232358 679308 232364
rect 678244 226840 678296 226846
rect 678244 226782 678296 226788
rect 679268 223825 679296 232358
rect 679254 223816 679310 223825
rect 679254 223751 679310 223760
rect 683316 219881 683344 233990
rect 683672 232688 683724 232694
rect 683672 232630 683724 232636
rect 683684 222737 683712 232630
rect 703694 224196 703722 224264
rect 704154 224196 704182 224264
rect 704614 224196 704642 224264
rect 705074 224196 705102 224264
rect 705534 224196 705562 224264
rect 705994 224196 706022 224264
rect 706454 224196 706482 224264
rect 706914 224196 706942 224264
rect 707374 224196 707402 224264
rect 707834 224196 707862 224264
rect 708294 224196 708322 224264
rect 708754 224196 708782 224264
rect 709214 224196 709242 224264
rect 683670 222728 683726 222737
rect 683670 222663 683726 222672
rect 683302 219872 683358 219881
rect 683302 219807 683358 219816
rect 676956 216504 677008 216510
rect 676956 216446 677008 216452
rect 676588 215348 676640 215354
rect 676588 215290 676640 215296
rect 675722 215206 676260 215234
rect 675666 215183 675722 215192
rect 675482 211440 675538 211449
rect 675482 211375 675538 211384
rect 676600 211177 676628 215290
rect 683118 212528 683174 212537
rect 683118 212463 683174 212472
rect 683132 211449 683160 212463
rect 683118 211440 683174 211449
rect 683118 211375 683174 211384
rect 676586 211168 676642 211177
rect 676586 211103 676642 211112
rect 675482 206952 675538 206961
rect 675482 206887 675538 206896
rect 675496 205875 675524 206887
rect 675312 205309 675418 205337
rect 675758 205048 675814 205057
rect 675758 204983 675814 204992
rect 675772 204680 675800 204983
rect 674852 204021 675418 204049
rect 675758 202736 675814 202745
rect 675758 202671 675814 202680
rect 675772 202195 675800 202671
rect 674746 201920 674802 201929
rect 674746 201855 674802 201864
rect 675390 201920 675446 201929
rect 675390 201855 675446 201864
rect 675404 201620 675432 201855
rect 674484 201466 674696 201494
rect 674286 196072 674342 196081
rect 674286 196007 674342 196016
rect 674668 180794 674696 201466
rect 675128 200994 675418 201022
rect 675128 198665 675156 200994
rect 675482 200560 675538 200569
rect 675482 200495 675538 200504
rect 675496 200328 675524 200495
rect 675114 198656 675170 198665
rect 675114 198591 675170 198600
rect 675390 198384 675446 198393
rect 675390 198319 675446 198328
rect 675404 197880 675432 198319
rect 675482 197568 675538 197577
rect 675482 197503 675538 197512
rect 675496 197336 675524 197503
rect 675390 197160 675446 197169
rect 675390 197095 675446 197104
rect 675404 196656 675432 197095
rect 675114 196072 675170 196081
rect 675170 196030 675418 196058
rect 675114 196007 675170 196016
rect 675772 194585 675800 194820
rect 675758 194576 675814 194585
rect 675758 194511 675814 194520
rect 675758 193216 675814 193225
rect 675758 193151 675814 193160
rect 675772 192984 675800 193151
rect 675666 192808 675722 192817
rect 675666 192743 675722 192752
rect 675680 192372 675708 192743
rect 675114 191176 675170 191185
rect 675170 191134 675418 191162
rect 675114 191111 675170 191120
rect 676126 189136 676182 189145
rect 676126 189071 676182 189080
rect 674484 180766 674696 180794
rect 674102 178528 674158 178537
rect 674102 178463 674158 178472
rect 674484 175681 674512 180766
rect 675942 180296 675998 180305
rect 675942 180231 675998 180240
rect 675956 178129 675984 180231
rect 675942 178120 675998 178129
rect 675942 178055 675998 178064
rect 676140 176654 676168 189071
rect 703694 179180 703722 179316
rect 704154 179180 704182 179316
rect 704614 179180 704642 179316
rect 705074 179180 705102 179316
rect 705534 179180 705562 179316
rect 705994 179180 706022 179316
rect 706454 179180 706482 179316
rect 706914 179180 706942 179316
rect 707374 179180 707402 179316
rect 707834 179180 707862 179316
rect 708294 179180 708322 179316
rect 708754 179180 708782 179316
rect 709214 179180 709242 179316
rect 675680 176626 676168 176654
rect 674654 176080 674710 176089
rect 674654 176015 674710 176024
rect 674470 175672 674526 175681
rect 674470 175607 674526 175616
rect 674668 172122 674696 176015
rect 674838 174040 674894 174049
rect 674838 173975 674894 173984
rect 674668 172094 674788 172122
rect 674562 172000 674618 172009
rect 674562 171935 674618 171944
rect 674378 169144 674434 169153
rect 674378 169079 674434 169088
rect 674392 166994 674420 169079
rect 674102 166968 674158 166977
rect 674392 166966 674512 166994
rect 674102 166903 674158 166912
rect 674116 162854 674144 166903
rect 674286 165608 674342 165617
rect 674286 165543 674342 165552
rect 674024 162826 674144 162854
rect 673826 160440 673882 160449
rect 673826 160375 673882 160384
rect 674024 157842 674052 162826
rect 673932 157814 674052 157842
rect 673932 153194 673960 157814
rect 674300 157706 674328 165543
rect 674484 162854 674512 166966
rect 674024 157678 674328 157706
rect 674392 162826 674512 162854
rect 674024 154986 674052 157678
rect 674392 157593 674420 162826
rect 674378 157584 674434 157593
rect 674576 157570 674604 171935
rect 674760 162058 674788 172094
rect 674852 162194 674880 173975
rect 675680 167521 675708 176626
rect 678242 173632 678298 173641
rect 678242 173567 678298 173576
rect 676034 173224 676090 173233
rect 676090 173182 676260 173210
rect 676034 173159 676090 173168
rect 676232 168450 676260 173182
rect 675864 168422 676260 168450
rect 675864 167634 675892 168422
rect 676034 167920 676090 167929
rect 676034 167855 676090 167864
rect 675864 167606 675984 167634
rect 675666 167512 675722 167521
rect 675666 167447 675722 167456
rect 675956 166994 675984 167606
rect 675220 166966 675984 166994
rect 674852 162166 675064 162194
rect 674760 162030 674972 162058
rect 674746 157584 674802 157593
rect 674576 157542 674746 157570
rect 674378 157519 674434 157528
rect 674746 157519 674802 157528
rect 674392 157406 674788 157434
rect 674392 155394 674420 157406
rect 674760 157334 674788 157406
rect 674944 157334 674972 162030
rect 675036 159066 675064 162166
rect 675220 161378 675248 166966
rect 676048 165617 676076 167855
rect 676034 165608 676090 165617
rect 676034 165543 676090 165552
rect 678256 162217 678284 173567
rect 679622 171592 679678 171601
rect 679622 171527 679678 171536
rect 678242 162208 678298 162217
rect 678242 162143 678298 162152
rect 679636 161770 679664 171527
rect 675944 161764 675996 161770
rect 675944 161706 675996 161712
rect 679624 161764 679676 161770
rect 679624 161706 679676 161712
rect 675956 161401 675984 161706
rect 675128 161350 675248 161378
rect 675942 161392 675998 161401
rect 675128 160358 675156 161350
rect 675942 161327 675998 161336
rect 675390 161120 675446 161129
rect 675390 161055 675446 161064
rect 675404 160888 675432 161055
rect 675128 160330 675340 160358
rect 675312 160290 675340 160330
rect 675404 160290 675432 160344
rect 675312 160262 675432 160290
rect 675666 160032 675722 160041
rect 675666 159967 675722 159976
rect 675680 159664 675708 159967
rect 675036 159038 675340 159066
rect 675312 158930 675340 159038
rect 675404 158930 675432 159052
rect 675312 158902 675432 158930
rect 674760 157306 674972 157334
rect 674746 157176 674802 157185
rect 674576 157134 674746 157162
rect 674576 156346 674604 157134
rect 674746 157111 674802 157120
rect 675772 157049 675800 157216
rect 675758 157040 675814 157049
rect 675758 156975 675814 156984
rect 674852 156629 675418 156657
rect 674576 156318 674788 156346
rect 674392 155366 674696 155394
rect 674024 154958 674328 154986
rect 673932 153166 674144 153194
rect 673642 132152 673698 132161
rect 673642 132087 673698 132096
rect 673366 129704 673422 129713
rect 673366 129639 673422 129648
rect 673918 128344 673974 128353
rect 673918 128279 673974 128288
rect 673366 126576 673422 126585
rect 673366 126511 673422 126520
rect 673182 124808 673238 124817
rect 673182 124743 673238 124752
rect 672998 123584 673054 123593
rect 672998 123519 673054 123528
rect 672722 119232 672778 119241
rect 672722 119167 672778 119176
rect 672538 116512 672594 116521
rect 672538 116447 672594 116456
rect 672078 114336 672134 114345
rect 672078 114271 672134 114280
rect 670804 109006 671384 109034
rect 671448 109006 671568 109034
rect 670148 108044 670200 108050
rect 670148 107986 670200 107992
rect 670804 106214 670832 109006
rect 670792 106208 670844 106214
rect 670792 106150 670844 106156
rect 671448 104938 671476 109006
rect 673012 106049 673040 123519
rect 673196 107001 673224 124743
rect 673182 106992 673238 107001
rect 673182 106927 673238 106936
rect 672998 106040 673054 106049
rect 672998 105975 673054 105984
rect 670804 104910 671476 104938
rect 670804 104854 670832 104910
rect 670792 104848 670844 104854
rect 670792 104790 670844 104796
rect 668582 102776 668638 102785
rect 668582 102711 668638 102720
rect 673380 101017 673408 126511
rect 673932 102830 673960 128279
rect 674116 114617 674144 153166
rect 674300 117473 674328 154958
rect 674470 154864 674526 154873
rect 674470 154799 674526 154808
rect 674484 152697 674512 154799
rect 674470 152688 674526 152697
rect 674470 152623 674526 152632
rect 674668 131345 674696 155366
rect 674760 149002 674788 156318
rect 674852 154442 674880 156629
rect 674944 155978 675418 156006
rect 674944 155258 674972 155978
rect 675114 155544 675170 155553
rect 675114 155479 675170 155488
rect 675128 155394 675156 155479
rect 675128 155366 675340 155394
rect 675312 155258 675340 155366
rect 675404 155258 675432 155380
rect 674944 155230 675064 155258
rect 675312 155230 675432 155258
rect 675036 155145 675064 155230
rect 675022 155136 675078 155145
rect 675022 155071 675078 155080
rect 675022 154456 675078 154465
rect 674852 154414 675022 154442
rect 675022 154391 675078 154400
rect 674944 152850 675418 152878
rect 674944 150385 674972 152850
rect 675114 152688 675170 152697
rect 675114 152623 675170 152632
rect 675128 152334 675156 152623
rect 675128 152306 675418 152334
rect 675114 151736 675170 151745
rect 675170 151680 675418 151689
rect 675114 151671 675418 151680
rect 675128 151661 675418 151671
rect 675114 151056 675170 151065
rect 675170 151014 675418 151042
rect 675114 150991 675170 151000
rect 674930 150376 674986 150385
rect 674930 150311 674986 150320
rect 675758 150376 675814 150385
rect 675758 150311 675814 150320
rect 675772 149835 675800 150311
rect 674760 148974 674880 149002
rect 674852 146146 674880 148974
rect 675758 148472 675814 148481
rect 675758 148407 675814 148416
rect 675772 147968 675800 148407
rect 675390 147656 675446 147665
rect 675390 147591 675446 147600
rect 675404 147356 675432 147591
rect 675312 146254 675432 146282
rect 675312 146146 675340 146254
rect 674852 146118 675340 146146
rect 675404 146132 675432 146254
rect 674838 134600 674894 134609
rect 674838 134535 674894 134544
rect 674852 133929 674880 134535
rect 674838 133920 674894 133929
rect 703694 133892 703722 134028
rect 704154 133892 704182 134028
rect 704614 133892 704642 134028
rect 705074 133892 705102 134028
rect 705534 133892 705562 134028
rect 705994 133892 706022 134028
rect 706454 133892 706482 134028
rect 706914 133892 706942 134028
rect 707374 133892 707402 134028
rect 707834 133892 707862 134028
rect 708294 133892 708322 134028
rect 708754 133892 708782 134028
rect 709214 133892 709242 134028
rect 674838 133855 674894 133864
rect 676494 133104 676550 133113
rect 676494 133039 676550 133048
rect 676508 132705 676536 133039
rect 676494 132696 676550 132705
rect 676494 132631 676550 132640
rect 674654 131336 674710 131345
rect 674654 131271 674710 131280
rect 676218 130248 676274 130257
rect 676218 130183 676274 130192
rect 675850 128888 675906 128897
rect 675850 128823 675906 128832
rect 675864 125882 675892 128823
rect 676232 127809 676260 130183
rect 676218 127800 676274 127809
rect 676218 127735 676274 127744
rect 676402 127800 676458 127809
rect 676402 127735 676458 127744
rect 674852 125854 675892 125882
rect 674654 125216 674710 125225
rect 674654 125151 674710 125160
rect 674470 123992 674526 124001
rect 674470 123927 674526 123936
rect 674286 117464 674342 117473
rect 674286 117399 674342 117408
rect 674102 114608 674158 114617
rect 674102 114543 674158 114552
rect 674484 107545 674512 123927
rect 674470 107536 674526 107545
rect 674470 107471 674526 107480
rect 674668 104666 674696 125151
rect 674852 113846 674880 125854
rect 676416 125458 676444 127735
rect 678242 126168 678298 126177
rect 678242 126103 678298 126112
rect 676036 125452 676088 125458
rect 676036 125394 676088 125400
rect 676404 125452 676456 125458
rect 676404 125394 676456 125400
rect 675022 122496 675078 122505
rect 675022 122431 675078 122440
rect 675036 121689 675064 122431
rect 675022 121680 675078 121689
rect 675022 121615 675078 121624
rect 675852 116680 675904 116686
rect 675852 116622 675904 116628
rect 675864 116385 675892 116622
rect 675114 116376 675170 116385
rect 675114 116311 675170 116320
rect 675850 116376 675906 116385
rect 675850 116311 675906 116320
rect 675128 116226 675156 116311
rect 674944 116198 675156 116226
rect 674944 115934 674972 116198
rect 676048 116113 676076 125394
rect 678256 116686 678284 126103
rect 682382 125352 682438 125361
rect 682382 125287 682438 125296
rect 682396 117337 682424 125287
rect 682382 117328 682438 117337
rect 682382 117263 682438 117272
rect 678244 116680 678296 116686
rect 678244 116622 678296 116628
rect 675114 116104 675170 116113
rect 675114 116039 675170 116048
rect 676034 116104 676090 116113
rect 676034 116039 676090 116048
rect 674944 115906 675064 115934
rect 675036 114493 675064 115906
rect 675128 115274 675156 116039
rect 675482 115832 675538 115841
rect 675482 115767 675538 115776
rect 675496 115668 675524 115767
rect 675128 115246 675432 115274
rect 675404 115124 675432 115246
rect 675036 114465 675418 114493
rect 674852 113818 675418 113846
rect 675758 112432 675814 112441
rect 675758 112367 675814 112376
rect 675772 111996 675800 112367
rect 675758 111752 675814 111761
rect 675758 111687 675814 111696
rect 675772 111452 675800 111687
rect 675758 111344 675814 111353
rect 675758 111279 675814 111288
rect 675772 110772 675800 111279
rect 675758 110392 675814 110401
rect 675758 110327 675814 110336
rect 675772 110160 675800 110327
rect 675758 108216 675814 108225
rect 675758 108151 675814 108160
rect 675772 107644 675800 108151
rect 675390 107536 675446 107545
rect 675390 107471 675446 107480
rect 675404 107100 675432 107471
rect 675390 106992 675446 107001
rect 675390 106927 675446 106936
rect 675404 106488 675432 106927
rect 675390 106040 675446 106049
rect 675390 105975 675446 105984
rect 675404 105808 675432 105975
rect 674668 104638 675340 104666
rect 675312 104530 675340 104638
rect 675404 104530 675432 104652
rect 675312 104502 675432 104530
rect 673932 102802 675340 102830
rect 675312 102762 675340 102802
rect 675404 102762 675432 102816
rect 675312 102734 675432 102762
rect 675390 102640 675446 102649
rect 675390 102575 675446 102584
rect 675404 102136 675432 102575
rect 673366 101008 673422 101017
rect 673366 100943 673422 100952
rect 675114 101008 675170 101017
rect 675170 100966 675340 100994
rect 675114 100943 675170 100952
rect 675312 100858 675340 100966
rect 675404 100858 675432 100980
rect 675312 100830 675432 100858
rect 668228 84166 668348 84194
rect 668228 76566 668256 84166
rect 668216 76560 668268 76566
rect 668216 76502 668268 76508
rect 666560 75200 666612 75206
rect 666560 75142 666612 75148
rect 662418 47424 662474 47433
rect 662418 47359 662474 47368
rect 661776 46504 661828 46510
rect 661776 46446 661828 46452
rect 661420 45526 661632 45554
rect 471058 43480 471114 43489
rect 471058 43415 471114 43424
rect 465814 43208 465870 43217
rect 465814 43143 465870 43152
rect 464344 42764 464396 42770
rect 464344 42706 464396 42712
rect 463700 42492 463752 42498
rect 463988 42486 464050 42514
rect 463700 42434 463752 42440
rect 461122 42256 461178 42265
rect 464022 42228 464050 42486
rect 465828 42364 465856 43143
rect 461122 42191 461178 42200
rect 471072 42106 471100 43415
rect 518806 42800 518862 42809
rect 518806 42735 518862 42744
rect 518820 42228 518848 42735
rect 661420 42187 661448 45526
rect 661408 42181 661460 42187
rect 515402 42120 515458 42129
rect 459940 42078 460368 42106
rect 471072 42078 471408 42106
rect 515154 42078 515402 42106
rect 520922 42120 520978 42129
rect 520674 42078 520922 42106
rect 515402 42055 515458 42064
rect 522026 42120 522082 42129
rect 521870 42078 522026 42106
rect 520922 42055 520978 42064
rect 526442 42120 526498 42129
rect 526194 42078 526442 42106
rect 522026 42055 522082 42064
rect 529570 42120 529626 42129
rect 661408 42123 661460 42129
rect 529322 42078 529570 42106
rect 526442 42055 526498 42064
rect 529570 42055 529626 42064
rect 454684 41880 454736 41886
rect 454684 41822 454736 41828
rect 449164 41744 449216 41750
rect 449164 41686 449216 41692
rect 453580 41744 453632 41750
rect 453580 41686 453632 41692
rect 446218 41576 446274 41585
rect 446218 41511 446274 41520
rect 141698 40352 141754 40361
rect 141698 40287 141754 40296
rect 141712 39984 141740 40287
<< via2 >>
rect 676034 897116 676090 897152
rect 676034 897096 676036 897116
rect 676036 897096 676088 897116
rect 676088 897096 676090 897116
rect 651470 868536 651526 868592
rect 675850 896688 675906 896744
rect 676034 896280 676090 896336
rect 652022 867584 652078 867640
rect 651470 866224 651526 866280
rect 651378 865172 651380 865192
rect 651380 865172 651432 865192
rect 651432 865172 651434 865192
rect 651378 865136 651434 865172
rect 651470 863812 651472 863832
rect 651472 863812 651524 863832
rect 651524 863812 651526 863832
rect 651470 863776 651526 863812
rect 651470 862280 651526 862336
rect 35622 817944 35678 818000
rect 35806 817264 35862 817320
rect 35622 816856 35678 816912
rect 35806 816040 35862 816096
rect 35622 815224 35678 815280
rect 35806 814428 35862 814464
rect 35806 814408 35808 814428
rect 35808 814408 35860 814428
rect 35860 814408 35862 814428
rect 41326 813592 41382 813648
rect 31666 812776 31722 812832
rect 31022 809920 31078 809976
rect 30286 809104 30342 809160
rect 41326 812368 41382 812424
rect 35162 811960 35218 812016
rect 32218 811144 32274 811200
rect 33782 809342 33838 809398
rect 39302 811552 39358 811608
rect 35162 802440 35218 802496
rect 41786 811280 41842 811336
rect 41786 810736 41842 810792
rect 41326 808716 41382 808752
rect 41326 808696 41328 808716
rect 41328 808696 41380 808716
rect 41380 808696 41382 808716
rect 41142 808288 41198 808344
rect 41326 807492 41382 807528
rect 41326 807472 41328 807492
rect 41328 807472 41380 807492
rect 41380 807472 41382 807492
rect 41142 806656 41198 806712
rect 41326 806248 41382 806304
rect 42154 810328 42210 810384
rect 41970 807880 42026 807936
rect 41786 805568 41842 805624
rect 41970 804752 42026 804808
rect 41970 804480 42026 804536
rect 40498 800672 40554 800728
rect 39302 800536 39358 800592
rect 41786 800264 41842 800320
rect 41786 799856 41842 799912
rect 42154 797272 42210 797328
rect 42154 795368 42210 795424
rect 41786 794824 41842 794880
rect 42062 793464 42118 793520
rect 42706 793464 42762 793520
rect 41786 793056 41842 793112
rect 42430 792648 42486 792704
rect 42246 791288 42302 791344
rect 42062 790608 42118 790664
rect 42614 791560 42670 791616
rect 42246 788160 42302 788216
rect 41786 786800 41842 786856
rect 41786 786120 41842 786176
rect 35806 774696 35862 774752
rect 35254 773880 35310 773936
rect 35622 773472 35678 773528
rect 35438 773064 35494 773120
rect 35806 773100 35808 773120
rect 35808 773100 35860 773120
rect 35860 773100 35862 773120
rect 35806 773064 35862 773100
rect 41510 773064 41566 773120
rect 35622 772248 35678 772304
rect 35806 771860 35862 771896
rect 35806 771840 35808 771860
rect 35808 771840 35860 771860
rect 35860 771840 35862 771860
rect 35806 771452 35862 771488
rect 35806 771432 35808 771452
rect 35808 771432 35860 771452
rect 35860 771432 35862 771452
rect 35622 771024 35678 771080
rect 35806 770616 35862 770672
rect 39118 770616 39174 770672
rect 43074 790608 43130 790664
rect 35806 770228 35862 770264
rect 35806 770208 35808 770228
rect 35808 770208 35860 770228
rect 35860 770208 35862 770228
rect 39486 770208 39542 770264
rect 35806 769392 35862 769448
rect 39854 769392 39910 769448
rect 35622 768984 35678 769040
rect 35806 768576 35862 768632
rect 35162 768168 35218 768224
rect 32402 767760 32458 767816
rect 33782 766944 33838 767000
rect 35806 767372 35862 767408
rect 35806 767352 35808 767372
rect 35808 767352 35860 767372
rect 35860 767352 35862 767372
rect 35806 766148 35862 766184
rect 35806 766128 35808 766148
rect 35808 766128 35860 766148
rect 35860 766128 35862 766148
rect 35806 765720 35862 765776
rect 35806 764532 35808 764552
rect 35808 764532 35860 764552
rect 35860 764532 35862 764552
rect 35806 764496 35862 764532
rect 35622 764088 35678 764144
rect 35806 763680 35862 763736
rect 35806 762864 35862 762920
rect 39578 764496 39634 764552
rect 40038 766944 40094 767000
rect 39762 764088 39818 764144
rect 40498 763308 40500 763328
rect 40500 763308 40552 763328
rect 40552 763308 40554 763328
rect 40498 763272 40554 763308
rect 40130 761776 40186 761832
rect 39946 758512 40002 758568
rect 36542 757696 36598 757752
rect 39854 757288 39910 757344
rect 41970 757152 42026 757208
rect 41786 757016 41842 757072
rect 41878 756608 41934 756664
rect 42430 764088 42486 764144
rect 43626 797272 43682 797328
rect 43258 770616 43314 770672
rect 43074 770208 43130 770264
rect 42614 761776 42670 761832
rect 42246 754024 42302 754080
rect 43258 758512 43314 758568
rect 42154 753344 42210 753400
rect 42062 752936 42118 752992
rect 41878 751576 41934 751632
rect 42062 751576 42118 751632
rect 42614 753616 42670 753672
rect 41970 750488 42026 750544
rect 41970 749672 42026 749728
rect 42246 749400 42302 749456
rect 41786 746816 41842 746872
rect 41970 745592 42026 745648
rect 42798 745592 42854 745648
rect 42246 745320 42302 745376
rect 41786 743688 41842 743744
rect 42522 744368 42578 744424
rect 41142 730904 41198 730960
rect 40774 728626 40830 728682
rect 41326 728626 41382 728682
rect 41050 727456 41106 727458
rect 41050 727404 41052 727456
rect 41052 727404 41104 727456
rect 41104 727404 41106 727456
rect 41050 727402 41106 727404
rect 41142 726824 41198 726880
rect 40958 726178 41014 726234
rect 35162 724784 35218 724840
rect 33046 724376 33102 724432
rect 33782 723730 33838 723786
rect 33046 716760 33102 716816
rect 39302 723152 39358 723208
rect 41326 726232 41382 726234
rect 41326 726180 41328 726232
rect 41328 726180 41380 726232
rect 41380 726180 41382 726232
rect 41326 726178 41382 726180
rect 41786 725736 41842 725792
rect 41326 725600 41382 725656
rect 41142 725192 41198 725248
rect 40958 717576 41014 717632
rect 40774 715264 40830 715320
rect 41786 722336 41842 722392
rect 41326 718800 41382 718856
rect 42062 720296 42118 720352
rect 42062 718800 42118 718856
rect 41786 718528 41842 718584
rect 41142 714856 41198 714912
rect 42430 715264 42486 715320
rect 42522 714856 42578 714912
rect 42062 714584 42118 714640
rect 39302 714176 39358 714232
rect 42154 710776 42210 710832
rect 41786 709824 41842 709880
rect 41878 708464 41934 708520
rect 42062 708464 42118 708520
rect 42062 707784 42118 707840
rect 41786 707376 41842 707432
rect 42522 706424 42578 706480
rect 41786 704248 41842 704304
rect 42246 703568 42302 703624
rect 42062 703024 42118 703080
rect 41970 702208 42026 702264
rect 42706 703024 42762 703080
rect 42522 702208 42578 702264
rect 42522 701800 42578 701856
rect 42522 701528 42578 701584
rect 42706 688064 42762 688120
rect 40866 686840 40922 686896
rect 41142 686432 41198 686488
rect 41050 685854 41106 685910
rect 41326 683460 41382 683462
rect 41326 683408 41328 683460
rect 41328 683408 41380 683460
rect 41380 683408 41382 683460
rect 41326 683406 41382 683408
rect 35162 681944 35218 682000
rect 31666 681536 31722 681592
rect 32402 680958 32458 681014
rect 33782 680958 33838 681014
rect 32402 672696 32458 672752
rect 41694 680992 41750 681048
rect 42706 682352 42762 682408
rect 41142 677048 41198 677104
rect 42338 671608 42394 671664
rect 42062 668480 42118 668536
rect 42062 666576 42118 666632
rect 41786 665080 41842 665136
rect 41786 663992 41842 664048
rect 42246 662768 42302 662824
rect 41786 658280 41842 658336
rect 41786 657192 41842 657248
rect 42522 658552 42578 658608
rect 35806 644680 35862 644736
rect 39486 644680 39542 644736
rect 38566 644272 38622 644328
rect 35346 643864 35402 643920
rect 35530 643456 35586 643512
rect 35806 643492 35808 643512
rect 35808 643492 35860 643512
rect 35860 643492 35862 643512
rect 35806 643456 35862 643492
rect 35622 642640 35678 642696
rect 35806 642232 35862 642288
rect 40498 643492 40500 643512
rect 40500 643492 40552 643512
rect 40552 643492 40554 643512
rect 40498 643456 40554 643492
rect 35622 641416 35678 641472
rect 35806 641008 35862 641064
rect 39578 641008 39634 641064
rect 35806 640600 35862 640656
rect 39946 640192 40002 640248
rect 35346 639784 35402 639840
rect 35530 639376 35586 639432
rect 35806 639376 35862 639432
rect 35622 638560 35678 638616
rect 32402 637744 32458 637800
rect 35162 637336 35218 637392
rect 32402 629856 32458 629912
rect 35806 638152 35862 638208
rect 35622 636928 35678 636984
rect 35806 636520 35862 636576
rect 35806 635704 35862 635760
rect 35806 634480 35862 634536
rect 35622 633664 35678 633720
rect 35806 633256 35862 633312
rect 39026 636148 39028 636168
rect 39028 636148 39080 636168
rect 39080 636148 39082 636168
rect 39026 636112 39082 636148
rect 39854 635704 39910 635760
rect 39486 634480 39542 634536
rect 40130 633664 40186 633720
rect 39762 632848 39818 632904
rect 41602 633256 41658 633312
rect 40406 632576 40462 632632
rect 42062 633256 42118 633312
rect 42706 632576 42762 632632
rect 37922 629176 37978 629232
rect 40498 628668 40500 628688
rect 40500 628668 40552 628688
rect 40552 628668 40554 628688
rect 40498 628632 40554 628668
rect 42338 628632 42394 628688
rect 41786 627408 41842 627464
rect 41786 627136 41842 627192
rect 42062 624416 42118 624472
rect 41786 623328 41842 623384
rect 41786 621968 41842 622024
rect 42154 621968 42210 622024
rect 41786 620744 41842 620800
rect 41878 615984 41934 616040
rect 42062 615848 42118 615904
rect 42706 615848 42762 615904
rect 42614 615440 42670 615496
rect 41878 613400 41934 613456
rect 43074 729272 43130 729328
rect 43074 686024 43130 686080
rect 43074 680312 43130 680368
rect 43074 635704 43130 635760
rect 43442 731312 43498 731368
rect 43626 730496 43682 730552
rect 43442 723560 43498 723616
rect 43626 710776 43682 710832
rect 43626 707784 43682 707840
rect 43442 687248 43498 687304
rect 43626 679496 43682 679552
rect 43442 676640 43498 676696
rect 43626 633664 43682 633720
rect 45006 795368 45062 795424
rect 62210 790472 62266 790528
rect 62118 789148 62120 789168
rect 62120 789148 62172 789168
rect 62172 789148 62174 789168
rect 62118 789112 62174 789148
rect 62118 787344 62174 787400
rect 62762 787072 62818 787128
rect 61382 786120 61438 786176
rect 62118 784896 62174 784952
rect 44914 773064 44970 773120
rect 44546 769392 44602 769448
rect 44362 764496 44418 764552
rect 44362 752936 44418 752992
rect 44178 751848 44234 751904
rect 44270 728048 44326 728104
rect 45098 751576 45154 751632
rect 44914 730088 44970 730144
rect 45190 729680 45246 729736
rect 44546 727640 44602 727696
rect 44454 722744 44510 722800
rect 44638 721520 44694 721576
rect 44638 708736 44694 708792
rect 44454 708464 44510 708520
rect 44822 687656 44878 687712
rect 44270 685208 44326 685264
rect 44638 684800 44694 684856
rect 44454 683984 44510 684040
rect 44270 680992 44326 681048
rect 43994 677864 44050 677920
rect 44270 644680 44326 644736
rect 45558 763272 45614 763328
rect 45006 684392 45062 684448
rect 45006 679904 45062 679960
rect 45006 666576 45062 666632
rect 45006 643456 45062 643512
rect 44454 641008 44510 641064
rect 44638 636112 44694 636168
rect 44270 634480 44326 634536
rect 44454 624416 44510 624472
rect 44822 632848 44878 632904
rect 44730 621968 44786 622024
rect 43258 612176 43314 612232
rect 43764 612196 43820 612232
rect 43764 612176 43766 612196
rect 43766 612176 43818 612196
rect 43818 612176 43820 612196
rect 43873 612040 43929 612096
rect 33782 601704 33838 601760
rect 32402 595176 32458 595232
rect 31022 594360 31078 594416
rect 38566 601296 38622 601352
rect 35438 595754 35494 595810
rect 33782 589328 33838 589384
rect 39946 600888 40002 600944
rect 45190 640192 45246 640248
rect 45006 600480 45062 600536
rect 44638 600072 44694 600128
rect 42890 597624 42946 597680
rect 42154 596808 42210 596864
rect 41694 595756 41696 595776
rect 41696 595756 41748 595776
rect 41748 595756 41750 595776
rect 41694 595720 41750 595756
rect 39302 594768 39358 594824
rect 36542 593544 36598 593600
rect 41694 594124 41696 594144
rect 41696 594124 41748 594144
rect 41748 594124 41750 594144
rect 41694 594088 41750 594124
rect 41970 592728 42026 592784
rect 41786 592320 41842 592376
rect 41786 590280 41842 590336
rect 41970 589600 42026 589656
rect 41510 589056 41566 589112
rect 41694 589056 41750 589112
rect 41510 586880 41566 586936
rect 39670 586100 39672 586120
rect 39672 586100 39724 586120
rect 39724 586100 39726 586120
rect 39670 586064 39726 586100
rect 42706 595992 42762 596048
rect 43074 596944 43130 597000
rect 42798 586880 42854 586936
rect 39302 585112 39358 585168
rect 39762 584568 39818 584624
rect 42614 584568 42670 584624
rect 42338 581168 42394 581224
rect 42062 580624 42118 580680
rect 41786 580216 41842 580272
rect 42246 578856 42302 578912
rect 42246 578040 42302 578096
rect 41786 577768 41842 577824
rect 41970 577088 42026 577144
rect 41786 574640 41842 574696
rect 41786 573824 41842 573880
rect 42798 577360 42854 577416
rect 42246 572192 42302 572248
rect 41786 570832 41842 570888
rect 42614 571920 42670 571976
rect 42430 571376 42486 571432
rect 41142 558048 41198 558104
rect 40038 553376 40094 553408
rect 40038 553352 40040 553376
rect 40040 553352 40092 553376
rect 40092 553352 40094 553376
rect 37922 552336 37978 552392
rect 29642 551928 29698 551984
rect 44362 593136 44418 593192
rect 44178 591912 44234 591968
rect 43350 591504 43406 591560
rect 43626 589056 43682 589112
rect 43074 556416 43130 556472
rect 42798 554784 42854 554840
rect 41326 552744 41382 552800
rect 41694 551792 41750 551848
rect 41970 550296 42026 550352
rect 41786 549888 41842 549944
rect 42154 550160 42210 550216
rect 41970 545672 42026 545728
rect 41786 545400 41842 545456
rect 37922 542272 37978 542328
rect 42798 551112 42854 551168
rect 42430 539552 42486 539608
rect 42522 537512 42578 537568
rect 42338 537240 42394 537296
rect 41786 536968 41842 537024
rect 42062 535744 42118 535800
rect 42154 535472 42210 535528
rect 42430 533840 42486 533896
rect 41786 533704 41842 533760
rect 42614 532888 42670 532944
rect 42062 530168 42118 530224
rect 42982 549480 43038 549536
rect 42706 530168 42762 530224
rect 42338 529896 42394 529952
rect 41878 529352 41934 529408
rect 42430 528944 42486 529000
rect 42706 527176 42762 527232
rect 35806 430072 35862 430128
rect 41142 425992 41198 426048
rect 35162 425346 35218 425402
rect 39302 425346 39358 425402
rect 33046 424768 33102 424824
rect 33782 423952 33838 424008
rect 40958 424360 41014 424416
rect 41786 423952 41842 424008
rect 41786 421912 41842 421968
rect 41510 418648 41566 418704
rect 40590 415948 40646 415984
rect 40590 415928 40592 415948
rect 40592 415928 40644 415948
rect 40644 415928 40646 415948
rect 42154 423952 42210 424008
rect 42798 423544 42854 423600
rect 42154 422864 42210 422920
rect 39302 415248 39358 415304
rect 35162 414840 35218 414896
rect 33782 414568 33838 414624
rect 42614 415928 42670 415984
rect 42246 409808 42302 409864
rect 42062 408040 42118 408096
rect 41786 406952 41842 407008
rect 42062 406680 42118 406736
rect 42430 407224 42486 407280
rect 42246 404504 42302 404560
rect 41786 403824 41842 403880
rect 43258 420688 43314 420744
rect 43074 419464 43130 419520
rect 42338 402872 42394 402928
rect 41786 401920 41842 401976
rect 42430 399744 42486 399800
rect 41786 399336 41842 399392
rect 41786 398792 41842 398848
rect 42154 395664 42210 395720
rect 41142 387096 41198 387152
rect 40958 385872 41014 385928
rect 40222 382200 40278 382256
rect 40958 382200 41014 382256
rect 40038 381792 40094 381848
rect 32402 381384 32458 381440
rect 37922 380976 37978 381032
rect 35806 376488 35862 376544
rect 35806 376080 35862 376136
rect 41326 386688 41382 386744
rect 41326 385872 41382 385928
rect 41326 382608 41382 382664
rect 41142 381792 41198 381848
rect 42798 379888 42854 379944
rect 40222 378936 40278 378992
rect 40038 376896 40094 376952
rect 39026 376488 39082 376544
rect 39026 376080 39082 376136
rect 41786 365608 41842 365664
rect 41786 364248 41842 364304
rect 42154 364248 42210 364304
rect 41786 363704 41842 363760
rect 42430 363024 42486 363080
rect 42246 362888 42302 362944
rect 42062 359216 42118 359272
rect 41878 358672 41934 358728
rect 42430 358672 42486 358728
rect 41786 356904 41842 356960
rect 41878 355544 41934 355600
rect 42154 353232 42210 353288
rect 43074 353912 43130 353968
rect 44178 581168 44234 581224
rect 44362 578040 44418 578096
rect 44914 598440 44970 598496
rect 44638 558728 44694 558784
rect 44546 556824 44602 556880
rect 44362 551520 44418 551576
rect 44178 549072 44234 549128
rect 43810 548256 43866 548312
rect 43994 547032 44050 547088
rect 44178 537512 44234 537568
rect 44362 528944 44418 529000
rect 44730 556008 44786 556064
rect 47214 721112 47270 721168
rect 47030 719888 47086 719944
rect 45558 612040 45614 612096
rect 45374 598848 45430 598904
rect 45190 598032 45246 598088
rect 45098 580624 45154 580680
rect 45558 578856 45614 578912
rect 54482 558456 54538 558512
rect 44914 555600 44970 555656
rect 45834 555192 45890 555248
rect 45650 554376 45706 554432
rect 44730 535744 44786 535800
rect 44546 429664 44602 429720
rect 44270 429256 44326 429312
rect 45098 550704 45154 550760
rect 45282 548664 45338 548720
rect 45282 535472 45338 535528
rect 45098 533840 45154 533896
rect 45098 527176 45154 527232
rect 44914 428848 44970 428904
rect 44638 428440 44694 428496
rect 44454 421504 44510 421560
rect 44454 406680 44510 406736
rect 44270 386416 44326 386472
rect 47582 547440 47638 547496
rect 45834 428032 45890 428088
rect 45558 427624 45614 427680
rect 44914 423136 44970 423192
rect 45098 422592 45154 422648
rect 45282 421096 45338 421152
rect 45098 409808 45154 409864
rect 45282 408040 45338 408096
rect 45098 407224 45154 407280
rect 44914 402872 44970 402928
rect 44638 385600 44694 385656
rect 45098 385192 45154 385248
rect 44914 382200 44970 382256
rect 44454 380296 44510 380352
rect 44178 377440 44234 377496
rect 44638 379344 44694 379400
rect 44638 364248 44694 364304
rect 45742 427216 45798 427272
rect 45926 426808 45982 426864
rect 45742 426400 45798 426456
rect 45742 399744 45798 399800
rect 45558 384784 45614 384840
rect 45558 384376 45614 384432
rect 45374 363024 45430 363080
rect 44454 359216 44510 359272
rect 43902 354864 43958 354920
rect 45190 354864 45246 354920
rect 43258 353640 43314 353696
rect 42430 352960 42486 353016
rect 35530 344256 35586 344312
rect 35806 344256 35862 344312
rect 39670 344256 39726 344312
rect 35806 343440 35862 343496
rect 39486 341808 39542 341864
rect 35622 341400 35678 341456
rect 35806 340992 35862 341048
rect 44914 343304 44970 343360
rect 45282 353932 45338 353968
rect 45282 353912 45284 353932
rect 45284 353912 45336 353932
rect 45336 353912 45338 353932
rect 45282 353676 45303 353696
rect 45303 353676 45338 353696
rect 45282 353640 45338 353676
rect 46110 404504 46166 404560
rect 53102 539552 53158 539608
rect 47950 430888 48006 430944
rect 47766 419872 47822 419928
rect 45926 383968 45982 384024
rect 46202 383560 46258 383616
rect 46018 380704 46074 380760
rect 45834 376216 45890 376272
rect 46478 378664 46534 378720
rect 45926 352960 45982 353016
rect 45558 344256 45614 344312
rect 45098 342488 45154 342544
rect 40222 342236 40278 342272
rect 40222 342216 40224 342236
rect 40224 342216 40276 342236
rect 40276 342216 40278 342236
rect 45466 342236 45522 342272
rect 45466 342216 45468 342236
rect 45468 342216 45520 342236
rect 45520 342216 45522 342236
rect 40038 341808 40094 341864
rect 39854 341400 39910 341456
rect 40222 340992 40278 341048
rect 47582 376624 47638 376680
rect 46754 362616 46810 362672
rect 46478 358672 46534 358728
rect 46110 340720 46166 340776
rect 39486 340176 39542 340232
rect 35530 339768 35586 339824
rect 35806 339768 35862 339824
rect 35162 338544 35218 338600
rect 35530 335688 35586 335744
rect 35806 335688 35862 335744
rect 35806 334464 35862 334520
rect 35806 332832 35862 332888
rect 35806 331744 35862 331800
rect 45650 339224 45706 339280
rect 45466 338000 45522 338056
rect 38566 335688 38622 335744
rect 40038 334464 40094 334520
rect 39762 332832 39818 332888
rect 44178 334600 44234 334656
rect 42798 334328 42854 334384
rect 40222 332424 40278 332480
rect 36542 331200 36598 331256
rect 35162 330384 35218 330440
rect 42430 326984 42486 327040
rect 41786 324808 41842 324864
rect 41786 322768 41842 322824
rect 42062 321136 42118 321192
rect 42430 320728 42486 320784
rect 42154 320456 42210 320512
rect 42338 320048 42394 320104
rect 42430 319640 42486 319696
rect 42982 332832 43038 332888
rect 43166 332424 43222 332480
rect 42982 321136 43038 321192
rect 43166 320456 43222 320512
rect 45282 326984 45338 327040
rect 46938 338408 46994 338464
rect 41786 316784 41842 316840
rect 41786 315968 41842 316024
rect 41786 315560 41842 315616
rect 41786 313656 41842 313712
rect 42430 312704 42486 312760
rect 46938 319640 46994 319696
rect 42154 312296 42210 312352
rect 45558 312296 45614 312352
rect 42062 310392 42118 310448
rect 35622 300872 35678 300928
rect 46202 300464 46258 300520
rect 44178 299648 44234 299704
rect 35806 298832 35862 298888
rect 41786 298696 41842 298752
rect 41786 297336 41842 297392
rect 42798 297336 42854 297392
rect 35806 297200 35862 297256
rect 41786 296520 41842 296576
rect 35438 296384 35494 296440
rect 31022 294752 31078 294808
rect 35622 295976 35678 296032
rect 35806 295568 35862 295624
rect 35806 295160 35862 295216
rect 35806 293528 35862 293584
rect 35806 292712 35862 292768
rect 35806 290264 35862 290320
rect 40774 292532 40830 292588
rect 41786 292440 41842 292496
rect 41786 292168 41842 292224
rect 41786 291896 41842 291952
rect 42154 291372 42210 291374
rect 42154 291320 42156 291372
rect 42156 291320 42208 291372
rect 42208 291320 42210 291372
rect 42154 291318 42210 291320
rect 41786 291080 41842 291136
rect 39302 284280 39358 284336
rect 41786 279792 41842 279848
rect 42062 278432 42118 278488
rect 42062 277888 42118 277944
rect 41786 277072 41842 277128
rect 42062 276664 42118 276720
rect 42430 278704 42486 278760
rect 42614 276664 42670 276720
rect 42246 275848 42302 275904
rect 41786 274216 41842 274272
rect 42338 273128 42394 273184
rect 42430 272856 42486 272912
rect 41786 272312 41842 272368
rect 41786 270408 41842 270464
rect 42430 270408 42486 270464
rect 42062 269048 42118 269104
rect 40682 267008 40738 267064
rect 35806 257080 35862 257136
rect 42154 266192 42210 266248
rect 43166 296520 43222 296576
rect 42982 292168 43038 292224
rect 42982 277888 43038 277944
rect 35806 255856 35862 255912
rect 39394 255856 39450 255912
rect 42798 255856 42854 255912
rect 35530 254224 35586 254280
rect 35806 254244 35862 254280
rect 35806 254224 35808 254244
rect 35808 254224 35860 254244
rect 35860 254224 35862 254244
rect 43626 291080 43682 291136
rect 43626 273128 43682 273184
rect 39394 253816 39450 253872
rect 42890 253816 42946 253872
rect 35806 253000 35862 253056
rect 35806 252612 35862 252648
rect 35806 252592 35808 252612
rect 35808 252592 35860 252612
rect 35860 252592 35862 252612
rect 35806 250144 35862 250200
rect 35806 248532 35862 248568
rect 35806 248512 35808 248532
rect 35808 248512 35860 248532
rect 35860 248512 35862 248532
rect 35806 247696 35862 247752
rect 35806 246880 35862 246936
rect 39394 244704 39450 244760
rect 40958 247696 41014 247752
rect 40314 245656 40370 245712
rect 42522 244704 42578 244760
rect 39578 244024 39634 244080
rect 42062 240080 42118 240136
rect 42246 238856 42302 238912
rect 43350 247696 43406 247752
rect 43166 245656 43222 245712
rect 43074 244024 43130 244080
rect 41786 236544 41842 236600
rect 42430 235864 42486 235920
rect 42430 233280 42486 233336
rect 42430 231920 42486 231976
rect 41786 229608 41842 229664
rect 42430 228928 42486 228984
rect 42430 227568 42486 227624
rect 41970 226072 42026 226128
rect 42614 226208 42670 226264
rect 42430 224848 42486 224904
rect 42154 223488 42210 223544
rect 35806 217912 35862 217968
rect 35806 214648 35862 214704
rect 35806 214260 35862 214296
rect 35806 214240 35808 214260
rect 35808 214240 35860 214260
rect 35860 214240 35862 214260
rect 39670 214260 39726 214296
rect 39670 214240 39672 214260
rect 39672 214240 39724 214260
rect 39724 214240 39726 214260
rect 35806 212200 35862 212256
rect 35622 211792 35678 211848
rect 44638 298016 44694 298072
rect 44362 294344 44418 294400
rect 44362 270408 44418 270464
rect 44178 256808 44234 256864
rect 44362 256400 44418 256456
rect 44178 254768 44234 254824
rect 43810 237904 43866 237960
rect 43442 230432 43498 230488
rect 40130 211792 40186 211848
rect 42798 211792 42854 211848
rect 35806 211384 35862 211440
rect 35530 210160 35586 210216
rect 35806 210160 35862 210216
rect 35806 209344 35862 209400
rect 33046 208936 33102 208992
rect 35806 207712 35862 207768
rect 40774 209344 40830 209400
rect 40130 207304 40186 207360
rect 41510 208120 41566 208176
rect 40958 206488 41014 206544
rect 40774 205672 40830 205728
rect 42982 209344 43038 209400
rect 42798 205672 42854 205728
rect 35622 205264 35678 205320
rect 35806 204468 35862 204504
rect 35806 204448 35808 204468
rect 35808 204448 35860 204468
rect 35860 204448 35862 204468
rect 41694 204468 41750 204504
rect 41694 204448 41696 204468
rect 41696 204448 41748 204468
rect 41748 204448 41750 204468
rect 41694 204040 41750 204096
rect 35806 203632 35862 203688
rect 33046 202136 33102 202192
rect 41878 202136 41934 202192
rect 35806 200640 35862 200696
rect 42430 197240 42486 197296
rect 41786 195744 41842 195800
rect 41970 195064 42026 195120
rect 42430 193160 42486 193216
rect 42338 191664 42394 191720
rect 41786 191528 41842 191584
rect 42430 190440 42486 190496
rect 42430 189896 42486 189952
rect 42430 187584 42486 187640
rect 41786 187176 41842 187232
rect 41786 186360 41842 186416
rect 41786 185952 41842 186008
rect 43166 206488 43222 206544
rect 42062 179288 42118 179344
rect 43994 230560 44050 230616
rect 43810 214240 43866 214296
rect 44822 293936 44878 293992
rect 45006 291488 45062 291544
rect 45006 278432 45062 278488
rect 44822 272856 44878 272912
rect 46202 258032 46258 258088
rect 54482 430480 54538 430536
rect 47950 387640 48006 387696
rect 50342 331744 50398 331800
rect 48962 289856 49018 289912
rect 47582 257624 47638 257680
rect 44914 255584 44970 255640
rect 44638 255176 44694 255232
rect 44546 251504 44602 251560
rect 44730 248240 44786 248296
rect 44546 240080 44602 240136
rect 44730 235864 44786 235920
rect 45558 253544 45614 253600
rect 44362 213696 44418 213752
rect 47214 252320 47270 252376
rect 45926 251912 45982 251968
rect 45742 249056 45798 249112
rect 47030 251096 47086 251152
rect 46110 249464 46166 249520
rect 46110 233280 46166 233336
rect 45926 231920 45982 231976
rect 45742 228928 45798 228984
rect 45558 227568 45614 227624
rect 47582 246608 47638 246664
rect 47214 226208 47270 226264
rect 47030 224848 47086 224904
rect 44822 212880 44878 212936
rect 44178 212064 44234 212120
rect 46938 208800 46994 208856
rect 44362 206760 44418 206816
rect 44178 205944 44234 206000
rect 43810 204448 43866 204504
rect 43994 204040 44050 204096
rect 43994 190440 44050 190496
rect 44546 205128 44602 205184
rect 44362 193160 44418 193216
rect 44822 204720 44878 204776
rect 44546 191664 44602 191720
rect 44178 187584 44234 187640
rect 46202 203496 46258 203552
rect 47122 208392 47178 208448
rect 47122 197240 47178 197296
rect 46938 189896 46994 189952
rect 47950 214920 48006 214976
rect 47766 213288 47822 213344
rect 47950 210840 48006 210896
rect 48594 202136 48650 202192
rect 48594 196424 48650 196480
rect 48318 194384 48374 194440
rect 47766 190440 47822 190496
rect 49146 247424 49202 247480
rect 49606 208120 49662 208176
rect 49606 192344 49662 192400
rect 50526 290672 50582 290728
rect 51078 395664 51134 395720
rect 51722 353232 51778 353288
rect 51722 334056 51778 334112
rect 50710 179288 50766 179344
rect 53838 320728 53894 320784
rect 53102 320048 53158 320104
rect 53838 310392 53894 310448
rect 53102 275848 53158 275904
rect 54482 266192 54538 266248
rect 55862 264152 55918 264208
rect 62762 747632 62818 747688
rect 62118 746136 62174 746192
rect 62118 744096 62174 744152
rect 62118 743724 62120 743744
rect 62120 743724 62172 743744
rect 62172 743724 62174 743744
rect 62118 743688 62174 743724
rect 62118 742364 62120 742384
rect 62120 742364 62172 742384
rect 62172 742364 62174 742384
rect 62118 742328 62174 742364
rect 63038 741784 63094 741840
rect 62118 704384 62174 704440
rect 62118 703296 62174 703352
rect 62210 701256 62266 701312
rect 62762 700848 62818 700904
rect 61382 699624 61438 699680
rect 62118 698164 62120 698184
rect 62120 698164 62172 698184
rect 62172 698164 62174 698184
rect 62118 698128 62174 698164
rect 62118 660900 62120 660920
rect 62120 660900 62172 660920
rect 62172 660900 62174 660920
rect 62118 660864 62174 660900
rect 62118 659540 62120 659560
rect 62120 659540 62172 659560
rect 62172 659540 62174 659560
rect 62118 659504 62174 659540
rect 62118 658280 62174 658336
rect 62762 657600 62818 657656
rect 61382 656512 61438 656568
rect 62118 655288 62174 655344
rect 62118 616528 62174 616584
rect 62118 614624 62174 614680
rect 61382 613808 61438 613864
rect 62118 612620 62120 612640
rect 62120 612620 62172 612640
rect 62172 612620 62174 612640
rect 62118 612584 62174 612620
rect 63130 618024 63186 618080
rect 62946 612040 63002 612096
rect 62670 595720 62726 595776
rect 62394 574776 62450 574832
rect 62394 573552 62450 573608
rect 63130 594088 63186 594144
rect 62946 590688 63002 590744
rect 62854 590008 62910 590064
rect 62394 571104 62450 571160
rect 62578 569880 62634 569936
rect 62210 556688 62266 556744
rect 62670 550160 62726 550216
rect 62118 531140 62174 531176
rect 62118 531120 62120 531140
rect 62120 531120 62172 531140
rect 62172 531120 62174 531140
rect 62302 530576 62358 530632
rect 62118 528572 62120 528592
rect 62120 528572 62172 528592
rect 62172 528572 62174 528592
rect 62118 528536 62174 528572
rect 62486 527992 62542 528048
rect 62118 527076 62120 527096
rect 62120 527076 62172 527096
rect 62172 527076 62174 527096
rect 62118 527040 62174 527076
rect 62670 525680 62726 525736
rect 62394 422864 62450 422920
rect 62118 404096 62174 404152
rect 62118 402600 62174 402656
rect 62118 400560 62174 400616
rect 62394 400152 62450 400208
rect 62118 399336 62174 399392
rect 62118 398248 62174 398304
rect 62210 385872 62266 385928
rect 62670 381792 62726 381848
rect 62118 360848 62174 360904
rect 62118 359760 62174 359816
rect 62118 357720 62174 357776
rect 62302 357312 62358 357368
rect 62118 355988 62120 356008
rect 62120 355988 62172 356008
rect 62172 355988 62174 356008
rect 62118 355952 62174 355988
rect 62670 354456 62726 354512
rect 62118 317364 62120 317384
rect 62120 317364 62172 317384
rect 62172 317364 62174 317384
rect 62118 317328 62174 317364
rect 62118 315988 62174 316024
rect 62118 315968 62120 315988
rect 62120 315968 62172 315988
rect 62172 315968 62174 315988
rect 62118 314764 62174 314800
rect 62118 314744 62120 314764
rect 62120 314744 62172 314764
rect 62172 314744 62174 314764
rect 62670 341672 62726 341728
rect 62486 341400 62542 341456
rect 62302 314064 62358 314120
rect 62486 312976 62542 313032
rect 62670 311752 62726 311808
rect 60002 300872 60058 300928
rect 62670 298696 62726 298752
rect 61566 295296 61622 295352
rect 61382 280336 61438 280392
rect 60002 223488 60058 223544
rect 62210 294208 62266 294264
rect 62302 292712 62358 292768
rect 62118 292460 62174 292496
rect 62118 292440 62120 292460
rect 62120 292440 62172 292460
rect 62172 292440 62174 292460
rect 62302 290944 62358 291000
rect 62670 289720 62726 289776
rect 62118 288516 62174 288552
rect 62118 288496 62120 288516
rect 62120 288496 62172 288516
rect 62172 288496 62174 288516
rect 62394 287136 62450 287192
rect 62118 285912 62174 285968
rect 62210 282104 62266 282160
rect 62118 280880 62174 280936
rect 61566 278704 61622 278760
rect 63130 568520 63186 568576
rect 63222 332560 63278 332616
rect 62946 284552 63002 284608
rect 62670 283192 62726 283248
rect 62394 267008 62450 267064
rect 62210 237904 62266 237960
rect 61290 217912 61346 217968
rect 63406 278704 63462 278760
rect 651470 778368 651526 778424
rect 652022 777008 652078 777064
rect 651470 776056 651526 776112
rect 651378 775276 651380 775296
rect 651380 775276 651432 775296
rect 651432 775276 651434 775296
rect 651378 775240 651434 775276
rect 651470 774172 651526 774208
rect 651470 774152 651472 774172
rect 651472 774152 651524 774172
rect 651524 774152 651526 774172
rect 651470 773336 651526 773392
rect 651470 734168 651526 734224
rect 651470 732944 651526 733000
rect 651470 731720 651526 731776
rect 651470 731040 651526 731096
rect 651470 729816 651526 729872
rect 651470 728492 651472 728512
rect 651472 728492 651524 728512
rect 651524 728492 651526 728512
rect 651470 728456 651526 728492
rect 651470 689424 651526 689480
rect 651654 688744 651710 688800
rect 651470 687384 651526 687440
rect 651470 686704 651526 686760
rect 651470 685208 651526 685264
rect 652574 684392 652630 684448
rect 651470 643184 651526 643240
rect 652022 641824 652078 641880
rect 651470 640736 651526 640792
rect 651378 640092 651380 640112
rect 651380 640092 651432 640112
rect 651432 640092 651434 640112
rect 651378 640056 651434 640092
rect 651470 638560 651526 638616
rect 651654 638152 651710 638208
rect 651470 597896 651526 597952
rect 651470 596672 651526 596728
rect 651470 595312 651526 595368
rect 651654 595040 651710 595096
rect 651470 594088 651526 594144
rect 651470 592728 651526 592784
rect 669778 775784 669834 775840
rect 668398 774968 668454 775024
rect 651470 553424 651526 553480
rect 652022 552064 652078 552120
rect 651470 551112 651526 551168
rect 651378 550332 651380 550352
rect 651380 550332 651432 550352
rect 651432 550332 651434 550352
rect 651378 550296 651434 550332
rect 651470 549228 651526 549264
rect 651470 549208 651472 549228
rect 651472 549208 651524 549228
rect 651524 549208 651526 549228
rect 651470 548392 651526 548448
rect 667662 639784 667718 639840
rect 667018 562128 667074 562184
rect 657542 403280 657598 403336
rect 652022 400832 652078 400888
rect 651470 373224 651526 373280
rect 652206 396616 652262 396672
rect 654782 382880 654838 382936
rect 652206 373904 652262 373960
rect 652022 372136 652078 372192
rect 651470 370640 651526 370696
rect 652022 356632 652078 356688
rect 651470 328208 651526 328264
rect 652390 351056 652446 351112
rect 653402 338680 653458 338736
rect 652390 329704 652446 329760
rect 652022 326848 652078 326904
rect 651378 325644 651434 325680
rect 651378 325624 651380 325644
rect 651380 325624 651432 325644
rect 651432 325624 651434 325644
rect 651470 301824 651526 301880
rect 651470 300600 651526 300656
rect 651746 297472 651802 297528
rect 651746 296812 651802 296848
rect 651746 296792 651748 296812
rect 651748 296792 651800 296812
rect 651800 296792 651802 296812
rect 651654 295296 651710 295352
rect 651470 294208 651526 294264
rect 651470 290400 651526 290456
rect 651654 290400 651710 290456
rect 651654 289176 651710 289232
rect 651470 288632 651526 288688
rect 651470 285912 651526 285968
rect 651470 284688 651526 284744
rect 651470 283464 651526 283520
rect 651470 282104 651526 282160
rect 651470 280880 651526 280936
rect 660302 311888 660358 311944
rect 652206 311072 652262 311128
rect 652206 303320 652262 303376
rect 652574 298560 652630 298616
rect 652850 293800 652906 293856
rect 652390 292712 652446 292768
rect 652206 291488 652262 291544
rect 652022 287136 652078 287192
rect 651838 279384 651894 279440
rect 461030 272856 461086 272912
rect 460846 272584 460902 272640
rect 461858 272620 461860 272640
rect 461860 272620 461912 272640
rect 461912 272620 461914 272640
rect 461858 272584 461914 272620
rect 464710 272448 464766 272504
rect 466274 272856 466330 272912
rect 470690 272484 470692 272504
rect 470692 272484 470744 272504
rect 470744 272484 470746 272504
rect 470690 272448 470746 272484
rect 470552 271940 470554 271960
rect 470554 271940 470606 271960
rect 470606 271940 470608 271960
rect 470552 271904 470608 271940
rect 478050 271904 478106 271960
rect 479522 271768 479578 271824
rect 480258 272312 480314 272368
rect 483202 271768 483258 271824
rect 484858 272312 484914 272368
rect 489918 272584 489974 272640
rect 499486 273028 499488 273048
rect 499488 273028 499540 273048
rect 499540 273028 499542 273048
rect 499486 272992 499542 273028
rect 499670 272584 499726 272640
rect 503350 273028 503352 273048
rect 503352 273028 503404 273048
rect 503404 273028 503406 273048
rect 503350 272992 503406 273028
rect 509238 269864 509294 269920
rect 509146 269456 509202 269512
rect 509882 269492 509884 269512
rect 509884 269492 509936 269512
rect 509936 269492 509938 269512
rect 509882 269456 509938 269492
rect 516506 269864 516562 269920
rect 532238 270136 532294 270192
rect 534078 270136 534134 270192
rect 536562 272448 536618 272504
rect 539322 273944 539378 274000
rect 538034 269728 538090 269784
rect 541806 269764 541808 269784
rect 541808 269764 541860 269784
rect 541860 269764 541862 269784
rect 541806 269728 541862 269764
rect 545946 273964 546002 274000
rect 545946 273944 545948 273964
rect 545948 273944 546000 273964
rect 546000 273944 546002 273964
rect 547694 272448 547750 272504
rect 547510 271940 547512 271960
rect 547512 271940 547564 271960
rect 547564 271940 547566 271960
rect 547510 271904 547566 271940
rect 547878 271904 547934 271960
rect 554410 262112 554466 262168
rect 554318 259936 554374 259992
rect 553950 257760 554006 257816
rect 553490 255604 553546 255640
rect 553490 255584 553492 255604
rect 553492 255584 553544 255604
rect 553544 255584 553546 255604
rect 554410 253408 554466 253464
rect 554134 251252 554190 251288
rect 554134 251232 554136 251252
rect 554136 251232 554188 251252
rect 554188 251232 554190 251252
rect 554042 249056 554098 249112
rect 553858 246880 553914 246936
rect 553674 242528 553730 242584
rect 140042 229200 140098 229256
rect 139306 228656 139362 228712
rect 141146 226108 141148 226128
rect 141148 226108 141200 226128
rect 141200 226108 141202 226128
rect 141146 226072 141202 226108
rect 142618 230444 142674 230480
rect 142618 230424 142620 230444
rect 142620 230424 142672 230444
rect 142672 230424 142674 230444
rect 140778 219836 140834 219872
rect 140778 219816 140780 219836
rect 140780 219816 140832 219836
rect 140832 219816 140834 219836
rect 141974 220380 142030 220416
rect 141974 220360 141976 220380
rect 141976 220360 142028 220380
rect 142028 220360 142030 220380
rect 142158 219836 142214 219872
rect 142158 219816 142160 219836
rect 142160 219816 142212 219836
rect 142212 219816 142214 219836
rect 142158 219564 142214 219600
rect 142158 219544 142160 219564
rect 142160 219544 142212 219564
rect 142212 219544 142214 219564
rect 144090 230424 144146 230480
rect 145838 229200 145894 229256
rect 145194 226108 145196 226128
rect 145196 226108 145248 226128
rect 145248 226108 145250 226128
rect 145194 226072 145250 226108
rect 145930 222264 145986 222320
rect 144182 220360 144238 220416
rect 147126 229200 147182 229256
rect 146482 228928 146538 228984
rect 147310 228656 147366 228712
rect 149242 228928 149298 228984
rect 147310 222944 147366 223000
rect 147126 222300 147128 222320
rect 147128 222300 147180 222320
rect 147180 222300 147182 222320
rect 147126 222264 147182 222300
rect 146758 220360 146814 220416
rect 147770 219564 147826 219600
rect 147770 219544 147772 219564
rect 147772 219544 147824 219564
rect 147824 219544 147826 219564
rect 150346 229336 150402 229392
rect 149978 229200 150034 229256
rect 151910 223252 151912 223272
rect 151912 223252 151964 223272
rect 151964 223252 151966 223272
rect 151910 223216 151966 223252
rect 151450 222944 151506 223000
rect 151634 222672 151690 222728
rect 152094 222672 152150 222728
rect 151772 220380 151828 220382
rect 151772 220328 151774 220380
rect 151774 220328 151826 220380
rect 151826 220328 151828 220380
rect 151772 220326 151828 220328
rect 151634 219544 151690 219600
rect 153658 219544 153714 219600
rect 154026 220652 154082 220688
rect 154026 220632 154028 220652
rect 154028 220632 154080 220652
rect 154080 220632 154082 220652
rect 156694 229900 156750 229936
rect 156694 229880 156696 229900
rect 156696 229880 156748 229900
rect 156748 229880 156750 229900
rect 156326 229356 156382 229392
rect 156326 229336 156328 229356
rect 156328 229336 156380 229356
rect 156380 229336 156382 229356
rect 156694 227432 156750 227488
rect 157430 229880 157486 229936
rect 157706 229628 157762 229664
rect 157706 229608 157708 229628
rect 157708 229608 157760 229628
rect 157760 229608 157762 229628
rect 158718 229608 158774 229664
rect 156970 220652 157026 220688
rect 156970 220632 156972 220652
rect 156972 220632 157024 220652
rect 157024 220632 157026 220652
rect 158258 221448 158314 221504
rect 160006 228112 160062 228168
rect 159822 223216 159878 223272
rect 161432 221876 161488 221912
rect 161432 221856 161434 221876
rect 161434 221856 161486 221876
rect 161486 221856 161488 221876
rect 161662 221604 161718 221640
rect 161662 221584 161664 221604
rect 161664 221584 161716 221604
rect 161716 221584 161718 221604
rect 166814 228928 166870 228984
rect 166814 228112 166870 228168
rect 166538 227432 166594 227488
rect 164514 221876 164570 221912
rect 164514 221856 164516 221876
rect 164516 221856 164568 221876
rect 164568 221856 164570 221876
rect 164146 220632 164202 220688
rect 167366 228948 167422 228984
rect 167366 228928 167368 228948
rect 167368 228928 167420 228948
rect 167420 228928 167422 228948
rect 169482 227316 169538 227352
rect 169482 227296 169484 227316
rect 169484 227296 169536 227316
rect 169536 227296 169538 227316
rect 167090 220632 167146 220688
rect 166952 220108 167008 220144
rect 166952 220088 166954 220108
rect 166954 220088 167006 220108
rect 167006 220088 167008 220108
rect 171230 227568 171286 227624
rect 172150 227568 172206 227624
rect 171690 227296 171746 227352
rect 170954 218476 171010 218512
rect 170954 218456 170956 218476
rect 170956 218456 171008 218476
rect 171008 218456 171010 218476
rect 173162 228792 173218 228848
rect 174818 228812 174874 228848
rect 174818 228792 174820 228812
rect 174820 228792 174872 228812
rect 174872 228792 174874 228812
rect 172886 218456 172942 218512
rect 176290 224848 176346 224904
rect 176842 224884 176844 224904
rect 176844 224884 176896 224904
rect 176896 224884 176898 224904
rect 176842 224848 176898 224884
rect 175554 220088 175610 220144
rect 176474 221332 176530 221368
rect 176474 221312 176476 221332
rect 176476 221312 176528 221332
rect 176528 221312 176530 221332
rect 177302 221312 177358 221368
rect 176474 220788 176530 220824
rect 176474 220768 176476 220788
rect 176476 220768 176528 220788
rect 176528 220768 176530 220788
rect 179786 220768 179842 220824
rect 180522 220088 180578 220144
rect 180890 219972 180946 220008
rect 180890 219952 180892 219972
rect 180892 219952 180944 219972
rect 180944 219952 180946 219972
rect 181534 220224 181590 220280
rect 184662 221720 184718 221776
rect 185766 221740 185822 221776
rect 185766 221720 185768 221740
rect 185768 221720 185820 221740
rect 185820 221720 185822 221740
rect 185122 219952 185178 220008
rect 202878 229084 202934 229120
rect 202878 229064 202880 229084
rect 202880 229064 202932 229084
rect 202932 229064 202934 229084
rect 203890 225392 203946 225448
rect 205178 229064 205234 229120
rect 205086 225428 205088 225448
rect 205088 225428 205140 225448
rect 205140 225428 205142 225448
rect 205086 225392 205142 225428
rect 219622 228656 219678 228712
rect 220542 228676 220598 228712
rect 220542 228656 220544 228676
rect 220544 228656 220596 228676
rect 220596 228656 220598 228676
rect 486974 219408 487030 219464
rect 487802 218048 487858 218104
rect 490378 218592 490434 218648
rect 492678 218320 492734 218376
rect 488676 217096 488732 217152
rect 493782 218320 493838 218376
rect 493782 217232 493838 217288
rect 494702 218864 494758 218920
rect 495346 217232 495402 217288
rect 497738 220904 497794 220960
rect 496910 218320 496966 218376
rect 498474 217232 498530 217288
rect 505650 217504 505706 217560
rect 508502 217776 508558 217832
rect 510158 217776 510214 217832
rect 513562 221176 513618 221232
rect 515218 219408 515274 219464
rect 519634 221448 519690 221504
rect 520186 221448 520242 221504
rect 522578 217776 522634 217832
rect 542266 222148 542322 222184
rect 542266 222128 542268 222148
rect 542268 222128 542320 222148
rect 542320 222128 542322 222148
rect 543692 222152 543748 222208
rect 543554 220516 543610 220552
rect 543554 220496 543556 220516
rect 543556 220496 543608 220516
rect 543608 220496 543610 220516
rect 544750 220496 544806 220552
rect 547142 221720 547198 221776
rect 550638 221992 550694 222048
rect 550822 221992 550878 222048
rect 554502 244704 554558 244760
rect 554502 240352 554558 240408
rect 554318 238176 554374 238232
rect 554502 236036 554504 236056
rect 554504 236036 554556 236056
rect 554556 236036 554558 236056
rect 554502 236000 554558 236036
rect 554410 233824 554466 233880
rect 553582 220632 553638 220688
rect 555790 224476 555792 224496
rect 555792 224476 555844 224496
rect 555844 224476 555846 224496
rect 555790 224440 555846 224476
rect 557262 224748 557264 224768
rect 557264 224748 557316 224768
rect 557316 224748 557318 224768
rect 557262 224712 557318 224748
rect 555698 217776 555754 217832
rect 558550 224748 558552 224768
rect 558552 224748 558604 224768
rect 558604 224748 558606 224768
rect 558550 224712 558606 224748
rect 558734 221992 558790 222048
rect 558550 221720 558606 221776
rect 558366 220360 558422 220416
rect 561402 224748 561404 224768
rect 561404 224748 561456 224768
rect 561456 224748 561458 224768
rect 561402 224712 561458 224748
rect 561678 224440 561734 224496
rect 562598 224476 562600 224496
rect 562600 224476 562652 224496
rect 562652 224476 562654 224496
rect 562598 224440 562654 224476
rect 563150 224476 563152 224496
rect 563152 224476 563204 224496
rect 563204 224476 563206 224496
rect 563150 224440 563206 224476
rect 560942 221720 560998 221776
rect 561494 220632 561550 220688
rect 562690 224032 562746 224088
rect 563426 224032 563482 224088
rect 563058 220632 563114 220688
rect 563242 220360 563298 220416
rect 563426 220360 563482 220416
rect 562874 219952 562930 220008
rect 563058 219952 563114 220008
rect 562690 217776 562746 217832
rect 562874 217776 562930 217832
rect 563610 217776 563666 217832
rect 565174 224712 565230 224768
rect 564806 220632 564862 220688
rect 565634 220360 565690 220416
rect 564806 219952 564862 220008
rect 567290 219136 567346 219192
rect 568946 221720 569002 221776
rect 569958 220652 570014 220688
rect 569958 220632 569960 220652
rect 569960 220632 570012 220652
rect 570012 220632 570014 220652
rect 571522 219156 571578 219192
rect 571522 219136 571524 219156
rect 571524 219136 571576 219156
rect 571576 219136 571578 219156
rect 570970 217776 571026 217832
rect 571338 217776 571394 217832
rect 573362 220632 573418 220688
rect 576582 220360 576638 220416
rect 572534 219952 572590 220008
rect 576582 219952 576638 220008
rect 572442 217776 572498 217832
rect 574098 217776 574154 217832
rect 574558 217776 574614 217832
rect 574098 216688 574154 216744
rect 574374 216688 574430 216744
rect 574926 216416 574982 216472
rect 582470 220224 582526 220280
rect 581826 219988 581828 220008
rect 581828 219988 581880 220008
rect 581880 219988 581882 220008
rect 581826 219952 581882 219988
rect 582654 219952 582710 220008
rect 591946 219952 592002 220008
rect 578882 213968 578938 214024
rect 578330 211656 578386 211712
rect 579526 209788 579528 209808
rect 579528 209788 579580 209808
rect 579580 209788 579582 209808
rect 579526 209752 579582 209788
rect 579526 207440 579582 207496
rect 579526 205828 579582 205864
rect 579526 205808 579528 205828
rect 579528 205808 579580 205828
rect 579580 205808 579582 205828
rect 599490 221176 599546 221232
rect 594798 218592 594854 218648
rect 595166 217504 595222 217560
rect 596362 217232 596418 217288
rect 595718 216960 595774 217016
rect 598478 215872 598534 215928
rect 600134 220088 600190 220144
rect 601146 220088 601202 220144
rect 603354 218320 603410 218376
rect 611450 219680 611506 219736
rect 618258 221448 618314 221504
rect 617246 219408 617302 219464
rect 618902 215328 618958 215384
rect 627458 218048 627514 218104
rect 627918 216144 627974 216200
rect 631322 220904 631378 220960
rect 631138 218320 631194 218376
rect 652574 280336 652630 280392
rect 667570 553832 667626 553888
rect 668398 696904 668454 696960
rect 668950 730088 669006 730144
rect 669594 735664 669650 735720
rect 669410 688336 669466 688392
rect 668950 600888 669006 600944
rect 668766 594768 668822 594824
rect 668398 554648 668454 554704
rect 670330 728728 670386 728784
rect 670606 696088 670662 696144
rect 670422 638696 670478 638752
rect 670974 689152 671030 689208
rect 671618 733760 671674 733816
rect 675850 895464 675906 895520
rect 676034 894648 676090 894704
rect 672998 778776 673054 778832
rect 672170 670148 672172 670168
rect 672172 670148 672224 670168
rect 672224 670148 672226 670168
rect 672170 670112 672226 670148
rect 672170 669724 672226 669760
rect 672170 669704 672172 669724
rect 672172 669704 672224 669724
rect 672224 669704 672226 669724
rect 672538 739880 672594 739936
rect 672814 715708 672816 715728
rect 672816 715708 672868 715728
rect 672868 715708 672870 715728
rect 672814 715672 672870 715708
rect 675850 893832 675906 893888
rect 676034 893036 676090 893072
rect 676034 893016 676036 893036
rect 676036 893016 676088 893036
rect 676088 893016 676090 893036
rect 676034 892608 676090 892664
rect 679622 891792 679678 891848
rect 676034 891384 676090 891440
rect 675850 890976 675906 891032
rect 674470 887984 674526 888040
rect 676034 890568 676090 890624
rect 676034 890160 676090 890216
rect 676034 888956 676090 888992
rect 676034 888936 676036 888956
rect 676036 888936 676088 888956
rect 676088 888936 676090 888956
rect 676034 888548 676090 888584
rect 676034 888528 676036 888548
rect 676036 888528 676088 888548
rect 676088 888528 676090 888548
rect 676034 887440 676090 887496
rect 676494 887712 676550 887768
rect 676310 887304 676366 887360
rect 676034 886916 676090 886952
rect 676034 886896 676036 886916
rect 676036 886896 676088 886916
rect 676088 886896 676090 886916
rect 676034 885692 676090 885728
rect 676034 885672 676036 885692
rect 676036 885672 676088 885692
rect 676088 885672 676090 885692
rect 676494 883360 676550 883416
rect 676310 883224 676366 883280
rect 678242 889752 678298 889808
rect 683302 889344 683358 889400
rect 683026 886080 683082 886136
rect 683026 881864 683082 881920
rect 675758 878464 675814 878520
rect 675666 877784 675722 877840
rect 674838 876560 674894 876616
rect 675482 874112 675538 874168
rect 675206 872344 675262 872400
rect 674838 870440 674894 870496
rect 675482 870440 675538 870496
rect 675574 869760 675630 869816
rect 675022 869216 675078 869272
rect 675390 869216 675446 869272
rect 675114 867176 675170 867232
rect 674838 866224 674894 866280
rect 675390 866224 675446 866280
rect 675114 865680 675170 865736
rect 675758 865408 675814 865464
rect 675758 788024 675814 788080
rect 675114 786664 675170 786720
rect 673734 780000 673790 780056
rect 673550 738656 673606 738712
rect 673366 715264 673422 715320
rect 673366 714876 673422 714912
rect 673366 714856 673368 714876
rect 673368 714856 673420 714876
rect 673420 714856 673422 714876
rect 673182 714448 673238 714504
rect 672998 706696 673054 706752
rect 673366 705508 673368 705528
rect 673368 705508 673420 705528
rect 673420 705508 673422 705528
rect 673366 705472 673422 705508
rect 673366 705200 673422 705256
rect 673182 703860 673238 703896
rect 673182 703840 673184 703860
rect 673184 703840 673236 703860
rect 673236 703840 673238 703860
rect 673182 701156 673184 701176
rect 673184 701156 673236 701176
rect 673236 701156 673238 701176
rect 673182 701120 673238 701156
rect 672998 700848 673054 700904
rect 672998 695272 673054 695328
rect 672814 695000 672870 695056
rect 672722 684936 672778 684992
rect 672538 665488 672594 665544
rect 672354 664128 672410 664184
rect 674102 734848 674158 734904
rect 673918 734168 673974 734224
rect 673826 722336 673882 722392
rect 674654 779184 674710 779240
rect 675114 784624 675170 784680
rect 675482 780544 675538 780600
rect 675482 780000 675538 780056
rect 675390 779184 675446 779240
rect 675482 778776 675538 778832
rect 674838 776192 674894 776248
rect 675114 775512 675170 775568
rect 674838 774560 674894 774616
rect 675482 775784 675538 775840
rect 675482 774968 675538 775024
rect 675482 774560 675538 774616
rect 675390 742192 675446 742248
rect 675482 739880 675538 739936
rect 675482 738656 675538 738712
rect 675482 738112 675538 738168
rect 675390 735664 675446 735720
rect 675482 734848 675538 734904
rect 675482 734168 675538 734224
rect 675574 733760 675630 733816
rect 675482 730088 675538 730144
rect 675482 728728 675538 728784
rect 674930 727232 674986 727288
rect 674102 721792 674158 721848
rect 674930 721656 674986 721712
rect 674194 720024 674250 720080
rect 674010 717032 674066 717088
rect 673826 716488 673882 716544
rect 673826 716080 673882 716136
rect 673826 714060 673882 714096
rect 673826 714040 673828 714060
rect 673828 714040 673880 714060
rect 673880 714040 673882 714060
rect 673826 713668 673828 713688
rect 673828 713668 673880 713688
rect 673880 713668 673882 713688
rect 673826 713632 673882 713668
rect 673826 713244 673882 713280
rect 673826 713224 673828 713244
rect 673828 713224 673880 713244
rect 673880 713224 673882 713244
rect 673826 712852 673828 712872
rect 673828 712852 673880 712872
rect 673880 712852 673882 712872
rect 673826 712816 673882 712852
rect 673826 712428 673882 712464
rect 673826 712408 673828 712428
rect 673828 712408 673880 712428
rect 673880 712408 673882 712428
rect 673826 711628 673828 711648
rect 673828 711628 673880 711648
rect 673880 711628 673882 711648
rect 673826 711592 673882 711628
rect 673826 709996 673828 710016
rect 673828 709996 673880 710016
rect 673880 709996 673882 710016
rect 673826 709960 673882 709996
rect 673826 709588 673828 709608
rect 673828 709588 673880 709608
rect 673880 709588 673882 709608
rect 673826 709552 673882 709588
rect 674286 705472 674342 705528
rect 674470 705200 674526 705256
rect 674286 703876 674288 703896
rect 674288 703876 674340 703896
rect 674340 703876 674342 703896
rect 674286 703840 674342 703876
rect 673550 693232 673606 693288
rect 673550 692960 673606 693016
rect 673182 690004 673184 690024
rect 673184 690004 673236 690024
rect 673236 690004 673238 690024
rect 673182 689968 673238 690004
rect 673182 688780 673184 688800
rect 673184 688780 673236 688800
rect 673236 688780 673238 688800
rect 673182 688744 673238 688780
rect 672814 659640 672870 659696
rect 671986 652432 672042 652488
rect 671802 649712 671858 649768
rect 671618 647808 671674 647864
rect 670422 549752 670478 549808
rect 669778 455368 669834 455424
rect 671158 607280 671214 607336
rect 670882 600364 670938 600400
rect 670882 600344 670884 600364
rect 670884 600344 670936 600364
rect 670936 600344 670938 600364
rect 670790 599140 670846 599176
rect 670790 599120 670792 599140
rect 670792 599120 670844 599140
rect 670844 599120 670846 599140
rect 670974 593544 671030 593600
rect 670790 533840 670846 533896
rect 672538 649168 672594 649224
rect 672354 604288 672410 604344
rect 672998 618568 673054 618624
rect 673182 608096 673238 608152
rect 672998 604016 673054 604072
rect 671802 562400 671858 562456
rect 671526 533024 671582 533080
rect 671342 532208 671398 532264
rect 671342 531528 671398 531584
rect 672262 555192 672318 555248
rect 672630 534964 672632 534984
rect 672632 534964 672684 534984
rect 672684 534964 672686 534984
rect 672630 534928 672686 534964
rect 672630 534112 672686 534168
rect 672630 533332 672632 533352
rect 672632 533332 672684 533352
rect 672684 533332 672686 533352
rect 672630 533296 672686 533332
rect 672538 532752 672594 532808
rect 670606 454960 670662 455016
rect 672262 453908 672264 453928
rect 672264 453908 672316 453928
rect 672316 453908 672318 453928
rect 672262 453872 672318 453908
rect 673182 527176 673238 527232
rect 673182 492088 673238 492144
rect 673182 490456 673238 490512
rect 673642 685752 673698 685808
rect 675298 710776 675354 710832
rect 682382 726552 682438 726608
rect 682382 711184 682438 711240
rect 678242 710368 678298 710424
rect 683486 708736 683542 708792
rect 684130 708328 684186 708384
rect 683302 707920 683358 707976
rect 676034 707104 676090 707160
rect 676034 706288 676090 706344
rect 683118 705472 683174 705528
rect 676034 705064 676090 705120
rect 675114 701392 675170 701448
rect 675114 701120 675170 701176
rect 674930 700848 674986 700904
rect 675114 696904 675170 696960
rect 675482 696768 675538 696824
rect 675114 696088 675170 696144
rect 675114 695000 675170 695056
rect 675298 695000 675354 695056
rect 675482 692960 675538 693016
rect 674102 690376 674158 690432
rect 675298 690376 675354 690432
rect 674930 689968 674986 690024
rect 674654 688744 674710 688800
rect 674654 688064 674710 688120
rect 673734 674328 673790 674384
rect 673734 671356 673790 671392
rect 673734 671336 673736 671356
rect 673736 671336 673788 671356
rect 673788 671336 673790 671356
rect 673734 670928 673790 670984
rect 673550 670520 673606 670576
rect 673550 669196 673552 669216
rect 673552 669196 673604 669216
rect 673604 669196 673606 669216
rect 673550 669160 673606 669196
rect 673550 668888 673606 668944
rect 673550 668480 673606 668536
rect 673550 668072 673606 668128
rect 673550 667664 673606 667720
rect 673550 666732 673606 666768
rect 673550 666712 673552 666732
rect 673552 666712 673604 666732
rect 673604 666712 673606 666732
rect 673550 666032 673606 666088
rect 673550 665236 673606 665272
rect 673550 665216 673552 665236
rect 673552 665216 673604 665236
rect 673604 665216 673606 665236
rect 673550 664808 673606 664864
rect 673550 663584 673606 663640
rect 673550 661952 673606 662008
rect 673550 644816 673606 644872
rect 673918 663040 673974 663096
rect 673918 661564 673974 661600
rect 673918 661544 673920 661564
rect 673920 661544 673972 661564
rect 673972 661544 673974 661564
rect 673918 661156 673974 661192
rect 673918 661136 673920 661156
rect 673920 661136 673972 661156
rect 673972 661136 673974 661156
rect 673918 660084 673920 660104
rect 673920 660084 673972 660104
rect 673972 660084 673974 660104
rect 673918 660048 673974 660084
rect 673918 655580 673974 655616
rect 673918 655560 673920 655580
rect 673920 655560 673972 655580
rect 673972 655560 673974 655580
rect 674010 647300 674012 647320
rect 674012 647300 674064 647320
rect 674064 647300 674066 647320
rect 674010 647264 674066 647300
rect 674010 645496 674066 645552
rect 674010 643084 674012 643104
rect 674012 643084 674064 643104
rect 674064 643084 674066 643104
rect 674010 643048 674066 643084
rect 673918 641688 673974 641744
rect 673734 635432 673790 635488
rect 675114 689152 675170 689208
rect 675114 688336 675170 688392
rect 675298 685752 675354 685808
rect 675482 684936 675538 684992
rect 675758 681400 675814 681456
rect 675390 680992 675446 681048
rect 674838 676368 674894 676424
rect 675758 676368 675814 676424
rect 674654 674328 674710 674384
rect 676034 666712 676090 666768
rect 683394 682352 683450 682408
rect 676218 663720 676274 663776
rect 683210 663720 683266 663776
rect 674838 663584 674894 663640
rect 676218 662940 676220 662960
rect 676220 662940 676272 662960
rect 676272 662940 676274 662960
rect 676218 662904 676274 662940
rect 683394 662496 683450 662552
rect 674654 660048 674710 660104
rect 683118 660048 683174 660104
rect 675114 655560 675170 655616
rect 675390 652840 675446 652896
rect 675114 652432 675170 652488
rect 675206 650120 675262 650176
rect 674286 635432 674342 635488
rect 674010 623892 674066 623928
rect 674010 623872 674012 623892
rect 674012 623872 674064 623892
rect 674064 623872 674066 623892
rect 674010 623076 674066 623112
rect 674010 623056 674012 623076
rect 674012 623056 674064 623076
rect 674064 623056 674066 623076
rect 674010 622260 674066 622296
rect 674010 622240 674012 622260
rect 674012 622240 674064 622260
rect 674064 622240 674066 622260
rect 674746 643592 674802 643648
rect 674010 614916 674066 614952
rect 674010 614896 674012 614916
rect 674012 614896 674064 614916
rect 674064 614896 674066 614916
rect 673734 603744 673790 603800
rect 674470 603744 674526 603800
rect 673734 599800 673790 599856
rect 673550 588512 673606 588568
rect 673550 580624 673606 580680
rect 673550 574540 673552 574560
rect 673552 574540 673604 574560
rect 673604 574540 673606 574560
rect 673550 574504 673606 574540
rect 673550 574096 673606 574152
rect 673550 569628 673606 569664
rect 673550 569608 673552 569628
rect 673552 569608 673604 569628
rect 673604 569608 673606 569628
rect 673550 565836 673552 565856
rect 673552 565836 673604 565856
rect 673604 565836 673606 565856
rect 673550 565800 673606 565836
rect 673550 559000 673606 559056
rect 674102 599120 674158 599176
rect 674286 599120 674342 599176
rect 674010 598032 674066 598088
rect 674102 597352 674158 597408
rect 673918 581052 673974 581088
rect 673918 581032 673920 581052
rect 673920 581032 673972 581052
rect 673972 581032 673974 581052
rect 673918 580252 673920 580272
rect 673920 580252 673972 580272
rect 673972 580252 673974 580272
rect 673918 580216 673974 580252
rect 673918 579844 673920 579864
rect 673920 579844 673972 579864
rect 673972 579844 673974 579864
rect 673918 579808 673974 579844
rect 673918 579420 673974 579456
rect 673918 579400 673920 579420
rect 673920 579400 673972 579420
rect 673972 579400 673974 579420
rect 673918 579028 673920 579048
rect 673920 579028 673972 579048
rect 673972 579028 673974 579048
rect 673918 578992 673974 579028
rect 673918 578604 673974 578640
rect 673918 578584 673920 578604
rect 673920 578584 673972 578604
rect 673972 578584 673974 578604
rect 673918 578196 673974 578232
rect 673918 578176 673920 578196
rect 673920 578176 673972 578196
rect 673972 578176 673974 578196
rect 673918 577788 673974 577824
rect 673918 577768 673920 577788
rect 673920 577768 673972 577788
rect 673972 577768 673974 577788
rect 673918 577396 673920 577416
rect 673920 577396 673972 577416
rect 673972 577396 673974 577416
rect 673918 577360 673974 577396
rect 673918 576972 673974 577008
rect 673918 576952 673920 576972
rect 673920 576952 673972 576972
rect 673972 576952 673974 576972
rect 673918 575356 673920 575376
rect 673920 575356 673972 575376
rect 673972 575356 673974 575376
rect 673918 575320 673974 575356
rect 673918 574912 673974 574968
rect 673918 573724 673920 573744
rect 673920 573724 673972 573744
rect 673972 573724 673974 573744
rect 673918 573688 673974 573724
rect 673918 572092 673920 572112
rect 673920 572092 673972 572112
rect 673972 572092 673974 572112
rect 673918 572056 673974 572092
rect 673918 570852 673974 570888
rect 673918 570832 673920 570852
rect 673920 570832 673972 570852
rect 673972 570832 673974 570852
rect 673918 570188 673920 570208
rect 673920 570188 673972 570208
rect 673972 570188 673974 570208
rect 673918 570152 673974 570188
rect 675390 649712 675446 649768
rect 675390 649168 675446 649224
rect 675758 648624 675814 648680
rect 675390 647808 675446 647864
rect 675206 647264 675262 647320
rect 675206 645496 675262 645552
rect 675390 644816 675446 644872
rect 675758 644680 675814 644736
rect 675390 643592 675446 643648
rect 675298 643048 675354 643104
rect 675298 641688 675354 641744
rect 675482 639784 675538 639840
rect 675482 638696 675538 638752
rect 674930 631352 674986 631408
rect 682382 636112 682438 636168
rect 676218 626068 676274 626104
rect 676218 626048 676220 626068
rect 676220 626048 676272 626068
rect 676272 626048 676274 626068
rect 676218 625660 676274 625696
rect 676218 625640 676220 625660
rect 676220 625640 676272 625660
rect 676272 625640 676274 625660
rect 676218 625252 676274 625288
rect 676218 625232 676220 625252
rect 676220 625232 676272 625252
rect 676272 625232 676274 625252
rect 676494 625232 676550 625288
rect 676034 624688 676090 624744
rect 676218 624452 676220 624472
rect 676220 624452 676272 624472
rect 676272 624452 676274 624472
rect 676218 624416 676274 624452
rect 676218 623620 676274 623656
rect 676218 623600 676220 623620
rect 676220 623600 676272 623620
rect 676272 623600 676274 623620
rect 676218 622820 676220 622840
rect 676220 622820 676272 622840
rect 676272 622820 676274 622840
rect 676218 622784 676274 622820
rect 682382 621968 682438 622024
rect 675298 621424 675354 621480
rect 676218 621188 676220 621208
rect 676220 621188 676272 621208
rect 676272 621188 676274 621208
rect 676218 621152 676274 621188
rect 676218 620780 676220 620800
rect 676220 620780 676272 620800
rect 676272 620780 676274 620800
rect 676218 620744 676274 620780
rect 676034 619812 676090 619848
rect 676034 619792 676036 619812
rect 676036 619792 676088 619812
rect 676088 619792 676090 619812
rect 676218 619112 676274 619168
rect 676494 619148 676496 619168
rect 676496 619148 676548 619168
rect 676548 619148 676550 619168
rect 676494 619112 676550 619148
rect 676034 618196 676036 618216
rect 676036 618196 676088 618216
rect 676088 618196 676090 618216
rect 676034 618160 676090 618196
rect 676218 617924 676220 617944
rect 676220 617924 676272 617944
rect 676272 617924 676274 617944
rect 676218 617888 676274 617924
rect 683118 617480 683174 617536
rect 683946 620336 684002 620392
rect 683302 617072 683358 617128
rect 676218 616684 676274 616720
rect 676218 616664 676220 616684
rect 676220 616664 676272 616684
rect 676272 616664 676274 616684
rect 683118 615476 683120 615496
rect 683120 615476 683172 615496
rect 683172 615476 683174 615496
rect 683118 615440 683174 615476
rect 675114 608096 675170 608152
rect 675114 607280 675170 607336
rect 674838 607008 674894 607064
rect 675390 604288 675446 604344
rect 675482 604016 675538 604072
rect 674470 598576 674526 598632
rect 673918 565120 673974 565176
rect 674286 565120 674342 565176
rect 674010 554376 674066 554432
rect 674010 553444 674066 553480
rect 674010 553424 674012 553444
rect 674012 553424 674064 553444
rect 674064 553424 674066 553444
rect 673918 551792 673974 551848
rect 675390 602792 675446 602848
rect 675482 600888 675538 600944
rect 675390 600344 675446 600400
rect 675482 599800 675538 599856
rect 675390 599120 675446 599176
rect 675482 598576 675538 598632
rect 675298 598032 675354 598088
rect 675482 597352 675538 597408
rect 674930 586472 674986 586528
rect 675482 594768 675538 594824
rect 675482 593544 675538 593600
rect 675114 586200 675170 586256
rect 677506 592864 677562 592920
rect 675574 588548 675576 588568
rect 675576 588548 675628 588568
rect 675628 588548 675630 588568
rect 675574 588512 675630 588548
rect 674654 570152 674710 570208
rect 678242 592592 678298 592648
rect 678242 576816 678298 576872
rect 677506 573552 677562 573608
rect 684222 591232 684278 591288
rect 683394 573144 683450 573200
rect 684222 576000 684278 576056
rect 684038 571920 684094 571976
rect 676218 571548 676220 571568
rect 676220 571548 676272 571568
rect 676272 571548 676274 571568
rect 676218 571512 676274 571548
rect 683118 570288 683174 570344
rect 675390 565800 675446 565856
rect 675114 562400 675170 562456
rect 675390 562128 675446 562184
rect 675390 561856 675446 561912
rect 675482 559408 675538 559464
rect 675206 559000 675262 559056
rect 674930 555464 674986 555520
rect 675390 555192 675446 555248
rect 675114 554648 675170 554704
rect 675298 554376 675354 554432
rect 675114 553424 675170 553480
rect 674746 551792 674802 551848
rect 675758 553968 675814 554024
rect 675482 553832 675538 553888
rect 675758 552064 675814 552120
rect 675390 550432 675446 550488
rect 675298 549752 675354 549808
rect 675298 549480 675354 549536
rect 673734 536288 673790 536344
rect 674286 536288 674342 536344
rect 673734 536036 673790 536072
rect 673734 536016 673736 536036
rect 673736 536016 673788 536036
rect 673788 536016 673790 536036
rect 673734 535780 673736 535800
rect 673736 535780 673788 535800
rect 673788 535780 673790 535800
rect 673734 535744 673790 535780
rect 673734 535200 673790 535256
rect 673734 530712 673790 530768
rect 673734 529932 673736 529952
rect 673736 529932 673788 529952
rect 673788 529932 673790 529952
rect 673734 529896 673790 529932
rect 673734 529508 673790 529544
rect 673734 529488 673736 529508
rect 673736 529488 673788 529508
rect 673788 529488 673790 529508
rect 673734 529236 673790 529272
rect 673734 529216 673736 529236
rect 673736 529216 673788 529236
rect 673788 529216 673790 529236
rect 673734 528828 673790 528864
rect 673734 528808 673736 528828
rect 673736 528808 673788 528828
rect 673788 528808 673790 528828
rect 674286 533840 674342 533896
rect 674286 532788 674288 532808
rect 674288 532788 674340 532808
rect 674340 532788 674342 532808
rect 674286 532752 674342 532788
rect 674378 527176 674434 527232
rect 673826 491272 673882 491328
rect 674010 490900 674012 490920
rect 674012 490900 674064 490920
rect 674064 490900 674066 490920
rect 674010 490864 674066 490900
rect 674010 490084 674012 490104
rect 674012 490084 674064 490104
rect 674064 490084 674066 490104
rect 674010 490048 674066 490084
rect 674010 489660 674066 489696
rect 674010 489640 674012 489660
rect 674012 489640 674064 489660
rect 674064 489640 674066 489660
rect 674010 489268 674012 489288
rect 674012 489268 674064 489288
rect 674064 489268 674066 489288
rect 674010 489232 674066 489268
rect 674010 488452 674012 488472
rect 674012 488452 674064 488472
rect 674064 488452 674066 488472
rect 674010 488416 674066 488452
rect 674010 486820 674012 486840
rect 674012 486820 674064 486840
rect 674064 486820 674066 486840
rect 674010 486784 674066 486820
rect 674010 486004 674012 486024
rect 674012 486004 674064 486024
rect 674064 486004 674066 486024
rect 674010 485968 674066 486004
rect 673550 484744 673606 484800
rect 674838 548392 674894 548448
rect 675758 548256 675814 548312
rect 677414 547576 677470 547632
rect 675206 541184 675262 541240
rect 675114 539552 675170 539608
rect 676218 534268 676274 534304
rect 676218 534248 676220 534268
rect 676220 534248 676272 534268
rect 676272 534248 676274 534268
rect 676034 533636 676090 533692
rect 676218 528128 676274 528184
rect 676034 526736 676036 526756
rect 676036 526736 676088 526756
rect 676088 526736 676090 526756
rect 676034 526700 676090 526736
rect 676034 526328 676036 526348
rect 676036 526328 676088 526348
rect 676088 526328 676090 526348
rect 676034 526292 676090 526328
rect 674654 484336 674710 484392
rect 673274 455388 673330 455424
rect 673274 455368 673276 455388
rect 673276 455368 673328 455388
rect 673328 455368 673330 455388
rect 673386 455252 673442 455288
rect 673386 455232 673388 455252
rect 673388 455232 673440 455252
rect 673440 455232 673442 455252
rect 673504 454960 673560 455016
rect 673044 454724 673046 454744
rect 673046 454724 673098 454744
rect 673098 454724 673100 454744
rect 673044 454688 673100 454724
rect 674286 454724 674288 454744
rect 674288 454724 674340 454744
rect 674340 454724 674342 454744
rect 674286 454688 674342 454724
rect 676034 491680 676090 491736
rect 676034 488824 676090 488880
rect 676034 485172 676090 485208
rect 676034 485152 676036 485172
rect 676036 485152 676088 485172
rect 676088 485152 676090 485172
rect 676034 483520 676090 483576
rect 675850 483112 675906 483168
rect 676034 482704 676090 482760
rect 683394 547304 683450 547360
rect 681002 547032 681058 547088
rect 679622 546760 679678 546816
rect 681002 531800 681058 531856
rect 682382 531392 682438 531448
rect 679622 530576 679678 530632
rect 683210 528128 683266 528184
rect 683578 527720 683634 527776
rect 683394 527312 683450 527368
rect 678978 525680 679034 525736
rect 683118 524864 683174 524920
rect 680358 524456 680414 524512
rect 683210 503648 683266 503704
rect 678242 487600 678298 487656
rect 679622 487192 679678 487248
rect 681002 486376 681058 486432
rect 683210 485560 683266 485616
rect 677138 482466 677194 482522
rect 676034 482296 676090 482352
rect 680358 481888 680414 481944
rect 675850 480664 675906 480720
rect 672952 454436 673008 454472
rect 672952 454416 672954 454436
rect 672954 454416 673006 454436
rect 673006 454416 673008 454436
rect 674286 454452 674288 454472
rect 674288 454452 674340 454472
rect 674340 454452 674342 454472
rect 674286 454416 674342 454452
rect 672814 454180 672816 454200
rect 672816 454180 672868 454200
rect 672868 454180 672870 454200
rect 672814 454144 672870 454180
rect 674286 454180 674288 454200
rect 674288 454180 674340 454200
rect 674340 454180 674342 454200
rect 674286 454144 674342 454180
rect 683118 481072 683174 481128
rect 674286 453908 674288 453928
rect 674288 453908 674340 453928
rect 674340 453908 674342 453928
rect 674286 453872 674342 453908
rect 676218 403300 676274 403336
rect 676218 403280 676220 403300
rect 676220 403280 676272 403300
rect 676272 403280 676274 403300
rect 673182 402328 673238 402384
rect 672630 402056 672686 402112
rect 672446 401648 672502 401704
rect 672814 399608 672870 399664
rect 672630 393896 672686 393952
rect 671342 392536 671398 392592
rect 668582 391176 668638 391232
rect 667386 358672 667442 358728
rect 667386 313656 667442 313712
rect 665822 268504 665878 268560
rect 664442 248240 664498 248296
rect 659566 230424 659622 230480
rect 652574 228520 652630 228576
rect 656162 226344 656218 226400
rect 653402 225256 653458 225312
rect 651470 224984 651526 225040
rect 646042 219816 646098 219872
rect 648618 218592 648674 218648
rect 651102 217776 651158 217832
rect 651930 221584 651986 221640
rect 654322 221040 654378 221096
rect 654138 220360 654194 220416
rect 653770 217504 653826 217560
rect 657542 223624 657598 223680
rect 656806 218864 656862 218920
rect 656530 215872 656586 215928
rect 658186 222264 658242 222320
rect 659382 213696 659438 213752
rect 660210 224032 660266 224088
rect 660394 215056 660450 215112
rect 661498 213424 661554 213480
rect 663706 229336 663762 229392
rect 663062 225664 663118 225720
rect 665178 230152 665234 230208
rect 664258 217776 664314 217832
rect 664258 217232 664314 217288
rect 664718 216416 664774 216472
rect 666834 224304 666890 224360
rect 667018 224032 667074 224088
rect 666006 222672 666062 222728
rect 667018 220360 667074 220416
rect 667018 219408 667074 219464
rect 666834 216688 666890 216744
rect 666650 215600 666706 215656
rect 578330 203224 578386 203280
rect 578790 200776 578846 200832
rect 579526 198872 579582 198928
rect 578514 196424 578570 196480
rect 579526 194928 579582 194984
rect 579526 192208 579582 192264
rect 579526 190712 579582 190768
rect 579526 187992 579582 188048
rect 579526 186260 579528 186280
rect 579528 186260 579580 186280
rect 579580 186260 579582 186280
rect 579526 186224 579582 186260
rect 579526 184320 579582 184376
rect 579526 181872 579582 181928
rect 578790 180104 578846 180160
rect 579526 177656 579582 177712
rect 578790 175072 578846 175128
rect 578422 173440 578478 173496
rect 578238 170992 578294 171048
rect 578698 169224 578754 169280
rect 578238 166912 578294 166968
rect 579526 164464 579582 164520
rect 579342 162696 579398 162752
rect 578238 159840 578294 159896
rect 578422 158344 578478 158400
rect 578882 155896 578938 155952
rect 578330 153584 578386 153640
rect 578238 151680 578294 151736
rect 578882 149640 578938 149696
rect 579526 147464 579582 147520
rect 578606 140528 578662 140584
rect 578606 138760 578662 138816
rect 579250 144644 579252 144664
rect 579252 144644 579304 144664
rect 579304 144644 579306 144664
rect 579250 144608 579306 144644
rect 579526 142976 579582 143032
rect 578882 136584 578938 136640
rect 579526 134408 579582 134464
rect 579066 132232 579122 132288
rect 578882 129648 578938 129704
rect 579526 127880 579582 127936
rect 578330 125296 578386 125352
rect 578698 123528 578754 123584
rect 578882 121352 578938 121408
rect 578514 118360 578570 118416
rect 578330 108296 578386 108352
rect 579526 116900 579528 116920
rect 579528 116900 579580 116920
rect 579580 116900 579582 116920
rect 579526 116864 579582 116900
rect 579250 114452 579252 114472
rect 579252 114452 579304 114472
rect 579304 114452 579306 114472
rect 579250 114416 579306 114452
rect 579526 112512 579582 112568
rect 579342 110064 579398 110120
rect 579066 105848 579122 105904
rect 578514 103128 578570 103184
rect 579158 101632 579214 101688
rect 578606 97416 578662 97472
rect 578330 94968 578386 95024
rect 579526 99220 579528 99240
rect 579528 99220 579580 99240
rect 579580 99220 579582 99240
rect 579526 99184 579582 99220
rect 579250 93064 579306 93120
rect 578606 90888 578662 90944
rect 579250 88032 579306 88088
rect 578330 86400 578386 86456
rect 579250 83988 579252 84008
rect 579252 83988 579304 84008
rect 579304 83988 579306 84008
rect 579250 83952 579306 83988
rect 578882 82184 578938 82240
rect 578238 77832 578294 77888
rect 579434 80008 579490 80064
rect 589462 207984 589518 208040
rect 589462 206352 589518 206408
rect 589462 204720 589518 204776
rect 589462 203088 589518 203144
rect 589462 201456 589518 201512
rect 589462 199824 589518 199880
rect 666650 198600 666706 198656
rect 666834 198328 666890 198384
rect 590382 198192 590438 198248
rect 589462 196560 589518 196616
rect 589278 194928 589334 194984
rect 589462 193296 589518 193352
rect 589462 191664 589518 191720
rect 590566 190032 590622 190088
rect 589646 188400 589702 188456
rect 589462 186768 589518 186824
rect 589462 185136 589518 185192
rect 589462 183504 589518 183560
rect 590566 181872 590622 181928
rect 589646 180240 589702 180296
rect 589462 178608 589518 178664
rect 589646 176976 589702 177032
rect 589462 175364 589518 175400
rect 589462 175344 589464 175364
rect 589464 175344 589516 175364
rect 589516 175344 589518 175364
rect 667018 174936 667074 174992
rect 589462 173712 589518 173768
rect 589462 172080 589518 172136
rect 589646 170448 589702 170504
rect 589462 168816 589518 168872
rect 589462 167184 589518 167240
rect 589462 165552 589518 165608
rect 589462 163920 589518 163976
rect 589462 162288 589518 162344
rect 589462 160656 589518 160712
rect 589462 159024 589518 159080
rect 589278 157412 589334 157448
rect 589278 157392 589280 157412
rect 589280 157392 589332 157412
rect 589332 157392 589334 157412
rect 589462 155760 589518 155816
rect 589462 154128 589518 154184
rect 589462 152496 589518 152552
rect 590014 150864 590070 150920
rect 589462 149232 589518 149288
rect 588542 147600 588598 147656
rect 580446 77832 580502 77888
rect 579250 75656 579306 75712
rect 578514 71168 578570 71224
rect 579526 73108 579528 73128
rect 579528 73108 579580 73128
rect 579580 73108 579582 73128
rect 579526 73072 579582 73108
rect 579526 66852 579528 66872
rect 579528 66852 579580 66872
rect 579580 66852 579582 66872
rect 579526 66816 579582 66852
rect 579526 64504 579582 64560
rect 579526 61784 579582 61840
rect 578882 60424 578938 60480
rect 574466 54712 574522 54768
rect 579526 57876 579528 57896
rect 579528 57876 579580 57896
rect 579580 57876 579582 57896
rect 579526 57840 579582 57876
rect 578330 56072 578386 56128
rect 577502 54984 577558 55040
rect 576122 54168 576178 54224
rect 589462 145968 589518 146024
rect 589462 144336 589518 144392
rect 589830 142704 589886 142760
rect 589462 141072 589518 141128
rect 589462 139460 589518 139496
rect 589462 139440 589464 139460
rect 589464 139440 589516 139460
rect 589516 139440 589518 139460
rect 589462 137808 589518 137864
rect 589462 136176 589518 136232
rect 590382 134544 590438 134600
rect 589462 132912 589518 132968
rect 589462 131300 589518 131336
rect 589462 131280 589464 131300
rect 589464 131280 589516 131300
rect 589516 131280 589518 131300
rect 588726 129648 588782 129704
rect 588542 103536 588598 103592
rect 589462 128016 589518 128072
rect 590106 126384 590162 126440
rect 589462 123120 589518 123176
rect 590566 124752 590622 124808
rect 589278 121508 589334 121544
rect 589278 121488 589280 121508
rect 589280 121488 589332 121508
rect 589332 121488 589334 121508
rect 668030 177928 668086 177984
rect 668030 174700 668032 174720
rect 668032 174700 668084 174720
rect 668084 174700 668086 174720
rect 668030 174664 668086 174700
rect 667938 173068 667940 173088
rect 667940 173068 667992 173088
rect 667992 173068 667994 173088
rect 667938 173032 667994 173068
rect 668214 169632 668270 169688
rect 668214 168172 668216 168192
rect 668216 168172 668268 168192
rect 668268 168172 668270 168192
rect 668214 168136 668270 168172
rect 667938 164908 667940 164928
rect 667940 164908 667992 164928
rect 667992 164908 667994 164928
rect 667938 164872 667994 164908
rect 668398 163240 668454 163296
rect 668398 160384 668454 160440
rect 668398 158344 668454 158400
rect 668214 140392 668270 140448
rect 670606 347248 670662 347304
rect 669318 344936 669374 344992
rect 669962 302096 670018 302152
rect 668766 300736 668822 300792
rect 668950 234504 669006 234560
rect 668582 143656 668638 143712
rect 668398 138760 668454 138816
rect 667754 134544 667810 134600
rect 667570 133048 667626 133104
rect 667386 132640 667442 132696
rect 667938 130636 667940 130656
rect 667940 130636 667992 130656
rect 667992 130636 667994 130656
rect 667938 130600 667994 130636
rect 669594 172352 669650 172408
rect 669318 159976 669374 160032
rect 669594 150320 669650 150376
rect 669134 150184 669190 150240
rect 668950 148552 669006 148608
rect 668766 133728 668822 133784
rect 670422 260480 670478 260536
rect 670146 258440 670202 258496
rect 670422 240216 670478 240272
rect 672630 376216 672686 376272
rect 672538 357040 672594 357096
rect 672170 352552 672226 352608
rect 671526 348472 671582 348528
rect 671158 259664 671214 259720
rect 670974 250688 671030 250744
rect 670974 248240 671030 248296
rect 671158 245520 671214 245576
rect 670790 223896 670846 223952
rect 670790 223644 670846 223680
rect 670790 223624 670792 223644
rect 670792 223624 670844 223644
rect 670844 223624 670846 223644
rect 670790 222264 670846 222320
rect 670790 218864 670846 218920
rect 670606 217504 670662 217560
rect 670790 214104 670846 214160
rect 670790 197512 670846 197568
rect 671250 234504 671306 234560
rect 671250 225256 671306 225312
rect 672354 349288 672410 349344
rect 672170 333376 672226 333432
rect 672354 332696 672410 332752
rect 672998 394712 673054 394768
rect 672998 380976 673054 381032
rect 673918 401376 673974 401432
rect 673366 400424 673422 400480
rect 673182 357448 673238 357504
rect 676586 402872 676642 402928
rect 674838 402600 674894 402656
rect 674838 402056 674894 402112
rect 676586 400832 676642 400888
rect 676034 399336 676090 399392
rect 674746 397296 674802 397352
rect 674562 396616 674618 396672
rect 674102 395800 674158 395856
rect 679622 398384 679678 398440
rect 676218 397976 676274 398032
rect 676034 396092 676090 396128
rect 676034 396072 676036 396092
rect 676036 396072 676088 396092
rect 676088 396072 676090 396092
rect 678242 397568 678298 397624
rect 676218 394324 676274 394360
rect 676218 394304 676220 394324
rect 676220 394304 676272 394324
rect 676272 394304 676274 394324
rect 676678 393488 676734 393544
rect 676678 391176 676734 391232
rect 678242 387640 678298 387696
rect 675758 384920 675814 384976
rect 675206 382880 675262 382936
rect 675758 382200 675814 382256
rect 675390 380976 675446 381032
rect 675758 378664 675814 378720
rect 675758 377304 675814 377360
rect 675390 376216 675446 376272
rect 675758 373632 675814 373688
rect 675666 372952 675722 373008
rect 673918 358264 673974 358320
rect 673366 355816 673422 355872
rect 673366 355408 673422 355464
rect 672814 355000 672870 355056
rect 673182 354592 673238 354648
rect 672722 353368 672778 353424
rect 672906 348880 672962 348936
rect 672722 340720 672778 340776
rect 672906 331200 672962 331256
rect 672906 324944 672962 325000
rect 672538 312432 672594 312488
rect 672538 304272 672594 304328
rect 671894 262112 671950 262168
rect 671710 257216 671766 257272
rect 672538 287816 672594 287872
rect 672262 285676 672264 285696
rect 672264 285676 672316 285696
rect 672316 285676 672318 285696
rect 672262 285640 672318 285676
rect 672078 246200 672134 246256
rect 671894 245248 671950 245304
rect 671342 221040 671398 221096
rect 670606 170992 670662 171048
rect 670330 170720 670386 170776
rect 670422 169904 670478 169960
rect 670974 171128 671030 171184
rect 670422 155080 670478 155136
rect 671158 155352 671214 155408
rect 670790 154400 670846 154456
rect 670606 151680 670662 151736
rect 670790 149116 670846 149152
rect 670790 149096 670792 149116
rect 670792 149096 670844 149116
rect 670844 149096 670846 149116
rect 671526 149096 671582 149152
rect 672078 236272 672134 236328
rect 672262 227024 672318 227080
rect 672262 225836 672264 225856
rect 672264 225836 672316 225856
rect 672316 225836 672318 225856
rect 672262 225800 672318 225836
rect 672032 225392 672088 225448
rect 672154 225292 672156 225312
rect 672156 225292 672208 225312
rect 672208 225292 672210 225312
rect 672154 225256 672210 225292
rect 672262 224984 672318 225040
rect 672078 223896 672134 223952
rect 672262 223624 672318 223680
rect 672078 217776 672134 217832
rect 672078 217504 672134 217560
rect 672262 215872 672318 215928
rect 672078 213696 672134 213752
rect 672078 213288 672134 213344
rect 671894 145288 671950 145344
rect 670146 130872 670202 130928
rect 668582 128968 668638 129024
rect 668582 127744 668638 127800
rect 667202 122032 667258 122088
rect 589646 119856 589702 119912
rect 589462 116592 589518 116648
rect 590106 118224 590162 118280
rect 589462 113328 589518 113384
rect 590290 114960 590346 115016
rect 589462 111696 589518 111752
rect 589462 110064 589518 110120
rect 589462 108432 589518 108488
rect 589462 106800 589518 106856
rect 589830 105168 589886 105224
rect 666650 109316 666706 109372
rect 667938 107752 667994 107808
rect 668122 106120 668178 106176
rect 668398 106156 668400 106176
rect 668400 106156 668452 106176
rect 668452 106156 668454 106176
rect 668398 106120 668454 106156
rect 589462 101904 589518 101960
rect 591302 54440 591358 54496
rect 625434 94424 625490 94480
rect 635554 96872 635610 96928
rect 635738 95920 635794 95976
rect 637026 96872 637082 96928
rect 641994 96464 642050 96520
rect 644938 96092 644940 96112
rect 644940 96092 644992 96112
rect 644992 96092 644994 96112
rect 644938 96056 644994 96092
rect 647330 94968 647386 95024
rect 648066 96484 648122 96520
rect 648066 96464 648068 96484
rect 648068 96464 648120 96484
rect 648120 96464 648122 96484
rect 647882 95784 647938 95840
rect 626446 93608 626502 93664
rect 626262 92792 626318 92848
rect 625802 91976 625858 92032
rect 626446 91160 626502 91216
rect 626446 90344 626502 90400
rect 625250 89528 625306 89584
rect 625434 88712 625490 88768
rect 624974 88576 625030 88632
rect 625250 88576 625306 88632
rect 626446 87896 626502 87952
rect 626262 87080 626318 87136
rect 648250 89528 648306 89584
rect 648618 96076 648674 96112
rect 648618 96056 648620 96076
rect 648620 96056 648672 96076
rect 648672 96056 648674 96076
rect 648802 91976 648858 92032
rect 649262 96464 649318 96520
rect 626446 86300 626448 86320
rect 626448 86300 626500 86320
rect 626500 86300 626502 86320
rect 626446 86264 626502 86300
rect 626446 85484 626448 85504
rect 626448 85484 626500 85504
rect 626500 85484 626502 85504
rect 626446 85448 626502 85484
rect 625250 84632 625306 84688
rect 648618 84632 648674 84688
rect 626446 83816 626502 83872
rect 628746 83272 628802 83328
rect 650550 87080 650606 87136
rect 655242 94152 655298 94208
rect 654690 93336 654746 93392
rect 655426 91432 655482 91488
rect 655426 90616 655482 90672
rect 656346 95784 656402 95840
rect 655794 89800 655850 89856
rect 663798 93064 663854 93120
rect 663982 91704 664038 91760
rect 664350 90616 664406 90672
rect 664534 89800 664590 89856
rect 665362 93336 665418 93392
rect 665178 88984 665234 89040
rect 650274 82184 650330 82240
rect 629206 81640 629262 81696
rect 623042 77288 623098 77344
rect 633898 78512 633954 78568
rect 633898 77288 633954 77344
rect 639602 77560 639658 77616
rect 646502 74160 646558 74216
rect 646686 71712 646742 71768
rect 646318 69128 646374 69184
rect 646134 67088 646190 67144
rect 459834 53624 459890 53680
rect 460754 53624 460810 53680
rect 461674 53624 461730 53680
rect 462594 53624 462650 53680
rect 468298 53236 468354 53272
rect 468298 53216 468300 53236
rect 468300 53216 468352 53236
rect 468352 53216 468354 53236
rect 475198 53216 475254 53272
rect 308034 50224 308090 50280
rect 130566 44376 130622 44432
rect 458178 46960 458234 47016
rect 522946 47776 523002 47832
rect 132590 44416 132646 44432
rect 132590 44376 132592 44416
rect 132592 44376 132644 44416
rect 132644 44376 132646 44416
rect 458362 46688 458418 46744
rect 459190 44376 459246 44432
rect 142618 44240 142674 44296
rect 255870 44104 255926 44160
rect 307298 43832 307354 43888
rect 440238 43852 440294 43888
rect 440238 43832 440240 43852
rect 440240 43832 440292 43852
rect 440292 43832 440294 43852
rect 194322 42064 194378 42120
rect 441066 43852 441122 43888
rect 441066 43832 441068 43852
rect 441068 43832 441120 43852
rect 441120 43832 441122 43852
rect 416594 42336 416650 42392
rect 415766 42064 415822 42120
rect 405646 41792 405702 41848
rect 419906 41792 419962 41848
rect 446218 42200 446274 42256
rect 460110 44104 460166 44160
rect 460846 43424 460902 43480
rect 461950 44376 462006 44432
rect 462502 44376 462558 44432
rect 462318 43152 462374 43208
rect 461766 42880 461822 42936
rect 463882 44104 463938 44160
rect 463974 42880 464030 42936
rect 549994 48864 550050 48920
rect 553674 48048 553730 48104
rect 552018 47776 552074 47832
rect 547878 47504 547934 47560
rect 545670 47232 545726 47288
rect 465262 46960 465318 47016
rect 465078 46688 465134 46744
rect 647514 78104 647570 78160
rect 647330 64368 647386 64424
rect 648986 62056 649042 62112
rect 648618 59200 648674 59256
rect 647514 57296 647570 57352
rect 661590 48454 661646 48510
rect 661774 47733 661830 47789
rect 667938 102720 667994 102776
rect 668306 104352 668362 104408
rect 668950 126928 669006 126984
rect 668766 125704 668822 125760
rect 668950 120808 669006 120864
rect 668766 120536 668822 120592
rect 669042 116456 669098 116512
rect 669226 115776 669282 115832
rect 669226 114552 669282 114608
rect 669042 114280 669098 114336
rect 669226 114280 669282 114336
rect 669226 112648 669282 112704
rect 668766 111016 668822 111072
rect 671342 131688 671398 131744
rect 671526 129240 671582 129296
rect 672262 212064 672318 212120
rect 673734 351328 673790 351384
rect 674378 356496 674434 356552
rect 674102 356224 674158 356280
rect 673918 351056 673974 351112
rect 674654 352144 674710 352200
rect 673734 338000 673790 338056
rect 674470 350920 674526 350976
rect 674470 350512 674526 350568
rect 674286 349696 674342 349752
rect 675942 357856 675998 357912
rect 675942 356768 675998 356824
rect 676034 350104 676090 350160
rect 676034 346568 676090 346624
rect 675206 344936 675262 344992
rect 675114 340720 675170 340776
rect 675758 340312 675814 340368
rect 675482 339360 675538 339416
rect 674930 338680 674986 338736
rect 675114 338000 675170 338056
rect 675758 337864 675814 337920
rect 675298 335280 675354 335336
rect 675482 333376 675538 333432
rect 675482 332696 675538 332752
rect 675114 331200 675170 331256
rect 675022 327936 675078 327992
rect 674654 326848 674710 326904
rect 675390 327936 675446 327992
rect 675390 326848 675446 326904
rect 675206 325624 675262 325680
rect 675022 324944 675078 325000
rect 676034 313248 676090 313304
rect 674838 312840 674894 312896
rect 674378 311616 674434 311672
rect 673366 310800 673422 310856
rect 673918 310392 673974 310448
rect 673182 309984 673238 310040
rect 673366 309576 673422 309632
rect 673182 303864 673238 303920
rect 673182 286456 673238 286512
rect 672814 285640 672870 285696
rect 672998 266056 673054 266112
rect 673734 305904 673790 305960
rect 673734 291488 673790 291544
rect 673550 290400 673606 290456
rect 673642 268096 673698 268152
rect 675482 312044 675538 312080
rect 675482 312024 675484 312044
rect 675484 312024 675536 312044
rect 675536 312024 675538 312044
rect 674838 311888 674894 311944
rect 674746 311344 674802 311400
rect 675942 311072 675998 311128
rect 675022 309168 675078 309224
rect 674378 305496 674434 305552
rect 674470 303456 674526 303512
rect 674470 300736 674526 300792
rect 674470 293800 674526 293856
rect 674838 297336 674894 297392
rect 676678 308352 676734 308408
rect 675482 307944 675538 308000
rect 676034 307536 676090 307592
rect 676034 307128 676090 307184
rect 676402 304680 676458 304736
rect 676402 301552 676458 301608
rect 678242 306720 678298 306776
rect 676678 301416 676734 301472
rect 675206 296928 675262 296984
rect 678978 306312 679034 306368
rect 676862 297336 676918 297392
rect 676126 296928 676182 296984
rect 675942 296520 675998 296576
rect 675758 295704 675814 295760
rect 675390 292848 675446 292904
rect 675574 292168 675630 292224
rect 675482 291488 675538 291544
rect 675758 290944 675814 291000
rect 675114 287816 675170 287872
rect 675758 287000 675814 287056
rect 675390 286456 675446 286512
rect 674378 267416 674434 267472
rect 674470 267008 674526 267064
rect 673918 265784 673974 265840
rect 673918 265376 673974 265432
rect 673366 264968 673422 265024
rect 673550 261568 673606 261624
rect 673182 259256 673238 259312
rect 673734 258848 673790 258904
rect 673550 247016 673606 247072
rect 673182 242664 673238 242720
rect 673734 241440 673790 241496
rect 673182 236680 673238 236736
rect 673642 236272 673698 236328
rect 672722 226380 672724 226400
rect 672724 226380 672776 226400
rect 672776 226380 672778 226400
rect 672722 226344 672778 226380
rect 672602 226108 672604 226128
rect 672604 226108 672656 226128
rect 672656 226108 672658 226128
rect 672602 226072 672658 226108
rect 673458 230152 673514 230208
rect 674102 264560 674158 264616
rect 675758 283600 675814 283656
rect 675666 282648 675722 282704
rect 675666 281560 675722 281616
rect 676862 279384 676918 279440
rect 675114 278296 675170 278352
rect 676862 268504 676918 268560
rect 676218 268096 676274 268152
rect 676218 267688 676274 267744
rect 674654 266600 674710 266656
rect 675482 264016 675538 264072
rect 676218 263608 676274 263664
rect 674470 262520 674526 262576
rect 674286 260072 674342 260128
rect 674102 235184 674158 235240
rect 674102 230424 674158 230480
rect 674286 230424 674342 230480
rect 674470 230152 674526 230208
rect 673734 228520 673790 228576
rect 673090 221448 673146 221504
rect 673734 226516 673736 226536
rect 673736 226516 673788 226536
rect 673788 226516 673790 226536
rect 673734 226480 673790 226516
rect 673734 221856 673790 221912
rect 673550 220088 673606 220144
rect 673182 217504 673238 217560
rect 672446 206896 672502 206952
rect 672538 202952 672594 203008
rect 672538 182008 672594 182064
rect 672998 214512 673054 214568
rect 672998 200504 673054 200560
rect 673366 216960 673422 217016
rect 673182 195200 673238 195256
rect 673550 214920 673606 214976
rect 673550 197104 673606 197160
rect 673366 191120 673422 191176
rect 674470 229336 674526 229392
rect 674102 220632 674158 220688
rect 674102 220088 674158 220144
rect 672722 177656 672778 177712
rect 673642 177248 673698 177304
rect 673642 176840 673698 176896
rect 672538 175208 672594 175264
rect 673366 174392 673422 174448
rect 672998 169496 673054 169552
rect 672722 168272 672778 168328
rect 672538 130464 672594 130520
rect 672262 126928 672318 126984
rect 672078 124072 672134 124128
rect 672538 122848 672594 122904
rect 672078 121624 672134 121680
rect 673182 168680 673238 168736
rect 672998 155488 673054 155544
rect 673182 151000 673238 151056
rect 674286 213696 674342 213752
rect 679622 263200 679678 263256
rect 676402 262792 676458 262848
rect 676218 261160 676274 261216
rect 675022 255312 675078 255368
rect 675850 255312 675906 255368
rect 674838 249872 674894 249928
rect 675666 250688 675722 250744
rect 675758 250144 675814 250200
rect 675114 248920 675170 248976
rect 675114 247016 675170 247072
rect 675758 246608 675814 246664
rect 675114 245520 675170 245576
rect 675114 245248 675170 245304
rect 675390 242664 675446 242720
rect 675206 241440 675262 241496
rect 675206 240216 675262 240272
rect 674838 238584 674894 238640
rect 675022 238040 675078 238096
rect 675390 238584 675446 238640
rect 675390 238040 675446 238096
rect 675850 235184 675906 235240
rect 674930 228928 674986 228984
rect 675206 226480 675262 226536
rect 674838 226072 674894 226128
rect 674654 222264 674710 222320
rect 675022 225800 675078 225856
rect 674838 221176 674894 221232
rect 674654 220224 674710 220280
rect 675206 222672 675262 222728
rect 675022 219816 675078 219872
rect 676954 230424 677010 230480
rect 676218 230152 676274 230208
rect 675666 225256 675722 225312
rect 674930 219000 674986 219056
rect 674746 216144 674802 216200
rect 674470 213016 674526 213072
rect 675390 218592 675446 218648
rect 676034 223080 676090 223136
rect 676034 221040 676090 221096
rect 675298 218184 675354 218240
rect 675666 217912 675722 217968
rect 676034 217504 676090 217560
rect 675666 216416 675722 216472
rect 676034 215348 676090 215384
rect 676034 215328 676036 215348
rect 676036 215328 676088 215348
rect 676088 215328 676090 215348
rect 675666 215192 675722 215248
rect 676678 228520 676734 228576
rect 679254 223760 679310 223816
rect 683670 222672 683726 222728
rect 683302 219816 683358 219872
rect 675482 211384 675538 211440
rect 683118 212472 683174 212528
rect 683118 211384 683174 211440
rect 676586 211112 676642 211168
rect 675482 206896 675538 206952
rect 675758 204992 675814 205048
rect 675758 202680 675814 202736
rect 674746 201864 674802 201920
rect 675390 201864 675446 201920
rect 674286 196016 674342 196072
rect 675482 200504 675538 200560
rect 675114 198600 675170 198656
rect 675390 198328 675446 198384
rect 675482 197512 675538 197568
rect 675390 197104 675446 197160
rect 675114 196016 675170 196072
rect 675758 194520 675814 194576
rect 675758 193160 675814 193216
rect 675666 192752 675722 192808
rect 675114 191120 675170 191176
rect 676126 189080 676182 189136
rect 674102 178472 674158 178528
rect 675942 180240 675998 180296
rect 675942 178064 675998 178120
rect 674654 176024 674710 176080
rect 674470 175616 674526 175672
rect 674838 173984 674894 174040
rect 674562 171944 674618 172000
rect 674378 169088 674434 169144
rect 674102 166912 674158 166968
rect 674286 165552 674342 165608
rect 673826 160384 673882 160440
rect 674378 157528 674434 157584
rect 678242 173576 678298 173632
rect 676034 173168 676090 173224
rect 676034 167864 676090 167920
rect 675666 167456 675722 167512
rect 674746 157528 674802 157584
rect 676034 165552 676090 165608
rect 679622 171536 679678 171592
rect 678242 162152 678298 162208
rect 675942 161336 675998 161392
rect 675390 161064 675446 161120
rect 675666 159976 675722 160032
rect 674746 157120 674802 157176
rect 675758 156984 675814 157040
rect 673642 132096 673698 132152
rect 673366 129648 673422 129704
rect 673918 128288 673974 128344
rect 673366 126520 673422 126576
rect 673182 124752 673238 124808
rect 672998 123528 673054 123584
rect 672722 119176 672778 119232
rect 672538 116456 672594 116512
rect 672078 114280 672134 114336
rect 673182 106936 673238 106992
rect 672998 105984 673054 106040
rect 668582 102720 668638 102776
rect 674470 154808 674526 154864
rect 674470 152632 674526 152688
rect 675114 155488 675170 155544
rect 675022 155080 675078 155136
rect 675022 154400 675078 154456
rect 675114 152632 675170 152688
rect 675114 151680 675170 151736
rect 675114 151000 675170 151056
rect 674930 150320 674986 150376
rect 675758 150320 675814 150376
rect 675758 148416 675814 148472
rect 675390 147600 675446 147656
rect 674838 134544 674894 134600
rect 674838 133864 674894 133920
rect 676494 133048 676550 133104
rect 676494 132640 676550 132696
rect 674654 131280 674710 131336
rect 676218 130192 676274 130248
rect 675850 128832 675906 128888
rect 676218 127744 676274 127800
rect 676402 127744 676458 127800
rect 674654 125160 674710 125216
rect 674470 123936 674526 123992
rect 674286 117408 674342 117464
rect 674102 114552 674158 114608
rect 674470 107480 674526 107536
rect 678242 126112 678298 126168
rect 675022 122440 675078 122496
rect 675022 121624 675078 121680
rect 675114 116320 675170 116376
rect 675850 116320 675906 116376
rect 682382 125296 682438 125352
rect 682382 117272 682438 117328
rect 675114 116048 675170 116104
rect 676034 116048 676090 116104
rect 675482 115776 675538 115832
rect 675758 112376 675814 112432
rect 675758 111696 675814 111752
rect 675758 111288 675814 111344
rect 675758 110336 675814 110392
rect 675758 108160 675814 108216
rect 675390 107480 675446 107536
rect 675390 106936 675446 106992
rect 675390 105984 675446 106040
rect 675390 102584 675446 102640
rect 673366 100952 673422 101008
rect 675114 100952 675170 101008
rect 662418 47368 662474 47424
rect 471058 43424 471114 43480
rect 465814 43152 465870 43208
rect 461122 42200 461178 42256
rect 518806 42744 518862 42800
rect 515402 42064 515458 42120
rect 520922 42064 520978 42120
rect 522026 42064 522082 42120
rect 526442 42064 526498 42120
rect 529570 42064 529626 42120
rect 446218 41520 446274 41576
rect 141698 40296 141754 40352
<< metal3 >>
rect 676029 897154 676095 897157
rect 676029 897152 676292 897154
rect 676029 897096 676034 897152
rect 676090 897096 676292 897152
rect 676029 897094 676292 897096
rect 676029 897091 676095 897094
rect 675845 896746 675911 896749
rect 675845 896744 676292 896746
rect 675845 896688 675850 896744
rect 675906 896688 676292 896744
rect 675845 896686 676292 896688
rect 675845 896683 675911 896686
rect 676029 896338 676095 896341
rect 676029 896336 676292 896338
rect 676029 896280 676034 896336
rect 676090 896280 676292 896336
rect 676029 896278 676292 896280
rect 676029 896275 676095 896278
rect 675845 895522 675911 895525
rect 675845 895520 676292 895522
rect 675845 895464 675850 895520
rect 675906 895464 676292 895520
rect 675845 895462 676292 895464
rect 675845 895459 675911 895462
rect 676029 894706 676095 894709
rect 676029 894704 676292 894706
rect 676029 894648 676034 894704
rect 676090 894648 676292 894704
rect 676029 894646 676292 894648
rect 676029 894643 676095 894646
rect 675845 893890 675911 893893
rect 675845 893888 676292 893890
rect 675845 893832 675850 893888
rect 675906 893832 676292 893888
rect 675845 893830 676292 893832
rect 675845 893827 675911 893830
rect 676029 893074 676095 893077
rect 676029 893072 676292 893074
rect 676029 893016 676034 893072
rect 676090 893016 676292 893072
rect 676029 893014 676292 893016
rect 676029 893011 676095 893014
rect 676029 892666 676095 892669
rect 676029 892664 676292 892666
rect 676029 892608 676034 892664
rect 676090 892608 676292 892664
rect 676029 892606 676292 892608
rect 676029 892603 676095 892606
rect 675702 892196 675708 892260
rect 675772 892258 675778 892260
rect 675772 892198 676292 892258
rect 675772 892196 675778 892198
rect 679617 891850 679683 891853
rect 679604 891848 679683 891850
rect 679604 891792 679622 891848
rect 679678 891792 679683 891848
rect 679604 891790 679683 891792
rect 679617 891787 679683 891790
rect 676029 891442 676095 891445
rect 676029 891440 676292 891442
rect 676029 891384 676034 891440
rect 676090 891384 676292 891440
rect 676029 891382 676292 891384
rect 676029 891379 676095 891382
rect 675845 891034 675911 891037
rect 675845 891032 676292 891034
rect 675845 890976 675850 891032
rect 675906 890976 676292 891032
rect 675845 890974 676292 890976
rect 675845 890971 675911 890974
rect 676029 890626 676095 890629
rect 676029 890624 676292 890626
rect 676029 890568 676034 890624
rect 676090 890568 676292 890624
rect 676029 890566 676292 890568
rect 676029 890563 676095 890566
rect 676029 890218 676095 890221
rect 676029 890216 676292 890218
rect 676029 890160 676034 890216
rect 676090 890160 676292 890216
rect 676029 890158 676292 890160
rect 676029 890155 676095 890158
rect 678237 889810 678303 889813
rect 678237 889808 678316 889810
rect 678237 889752 678242 889808
rect 678298 889752 678316 889808
rect 678237 889750 678316 889752
rect 678237 889747 678303 889750
rect 683297 889402 683363 889405
rect 683284 889400 683363 889402
rect 683284 889344 683302 889400
rect 683358 889344 683363 889400
rect 683284 889342 683363 889344
rect 683297 889339 683363 889342
rect 676029 888994 676095 888997
rect 676029 888992 676292 888994
rect 676029 888936 676034 888992
rect 676090 888936 676292 888992
rect 676029 888934 676292 888936
rect 676029 888931 676095 888934
rect 676029 888586 676095 888589
rect 676029 888584 676292 888586
rect 676029 888528 676034 888584
rect 676090 888528 676292 888584
rect 676029 888526 676292 888528
rect 676029 888523 676095 888526
rect 676170 888118 676292 888178
rect 674465 888042 674531 888045
rect 676170 888042 676230 888118
rect 674465 888040 676230 888042
rect 674465 887984 674470 888040
rect 674526 887984 676230 888040
rect 674465 887982 676230 887984
rect 674465 887979 674531 887982
rect 676489 887770 676555 887773
rect 676476 887768 676555 887770
rect 676476 887712 676494 887768
rect 676550 887712 676555 887768
rect 676476 887710 676555 887712
rect 676489 887707 676555 887710
rect 675518 887436 675524 887500
rect 675588 887498 675594 887500
rect 676029 887498 676095 887501
rect 675588 887496 676095 887498
rect 675588 887440 676034 887496
rect 676090 887440 676095 887496
rect 675588 887438 676095 887440
rect 675588 887436 675594 887438
rect 676029 887435 676095 887438
rect 676305 887362 676371 887365
rect 676292 887360 676371 887362
rect 676292 887304 676310 887360
rect 676366 887304 676371 887360
rect 676292 887302 676371 887304
rect 676305 887299 676371 887302
rect 676029 886954 676095 886957
rect 676029 886952 676292 886954
rect 676029 886896 676034 886952
rect 676090 886896 676292 886952
rect 676029 886894 676292 886896
rect 676029 886891 676095 886894
rect 683070 886141 683130 886516
rect 683021 886136 683130 886141
rect 683021 886080 683026 886136
rect 683082 886108 683130 886136
rect 683082 886080 683100 886108
rect 683021 886078 683100 886080
rect 683021 886075 683087 886078
rect 676029 885730 676095 885733
rect 676029 885728 676292 885730
rect 676029 885672 676034 885728
rect 676090 885672 676292 885728
rect 676029 885670 676292 885672
rect 676029 885667 676095 885670
rect 676489 883420 676555 883421
rect 676438 883356 676444 883420
rect 676508 883418 676555 883420
rect 676508 883416 676600 883418
rect 676550 883360 676600 883416
rect 676508 883358 676600 883360
rect 676508 883356 676555 883358
rect 676489 883355 676555 883356
rect 676305 883284 676371 883285
rect 676254 883282 676260 883284
rect 676214 883222 676260 883282
rect 676324 883280 676371 883284
rect 676366 883224 676371 883280
rect 676254 883220 676260 883222
rect 676324 883220 676371 883224
rect 676305 883219 676371 883220
rect 675702 881860 675708 881924
rect 675772 881922 675778 881924
rect 683021 881922 683087 881925
rect 675772 881920 683087 881922
rect 675772 881864 683026 881920
rect 683082 881864 683087 881920
rect 675772 881862 683087 881864
rect 675772 881860 675778 881862
rect 683021 881859 683087 881862
rect 675753 878522 675819 878525
rect 675710 878520 675819 878522
rect 675710 878464 675758 878520
rect 675814 878464 675819 878520
rect 675710 878459 675819 878464
rect 675710 877845 675770 878459
rect 675661 877840 675770 877845
rect 675661 877784 675666 877840
rect 675722 877784 675770 877840
rect 675661 877782 675770 877784
rect 675661 877779 675727 877782
rect 674833 876618 674899 876621
rect 675150 876618 675156 876620
rect 674833 876616 675156 876618
rect 674833 876560 674838 876616
rect 674894 876560 675156 876616
rect 674833 876558 675156 876560
rect 674833 876555 674899 876558
rect 675150 876556 675156 876558
rect 675220 876556 675226 876620
rect 675150 874108 675156 874172
rect 675220 874170 675226 874172
rect 675477 874170 675543 874173
rect 675220 874168 675543 874170
rect 675220 874112 675482 874168
rect 675538 874112 675543 874168
rect 675220 874110 675543 874112
rect 675220 874108 675226 874110
rect 675477 874107 675543 874110
rect 675518 873564 675524 873628
rect 675588 873626 675594 873628
rect 676438 873626 676444 873628
rect 675588 873566 676444 873626
rect 675588 873564 675594 873566
rect 676438 873564 676444 873566
rect 676508 873564 676514 873628
rect 675201 872402 675267 872405
rect 676254 872402 676260 872404
rect 675201 872400 676260 872402
rect 675201 872344 675206 872400
rect 675262 872344 676260 872400
rect 675201 872342 676260 872344
rect 675201 872339 675267 872342
rect 676254 872340 676260 872342
rect 676324 872340 676330 872404
rect 674833 870498 674899 870501
rect 675477 870498 675543 870501
rect 674833 870496 675543 870498
rect 674833 870440 674838 870496
rect 674894 870440 675482 870496
rect 675538 870440 675543 870496
rect 674833 870438 675543 870440
rect 674833 870435 674899 870438
rect 675477 870435 675543 870438
rect 675569 869820 675635 869821
rect 675518 869756 675524 869820
rect 675588 869818 675635 869820
rect 675588 869816 675680 869818
rect 675630 869760 675680 869816
rect 675588 869758 675680 869760
rect 675588 869756 675635 869758
rect 675569 869755 675635 869756
rect 675017 869274 675083 869277
rect 675385 869274 675451 869277
rect 675017 869272 675451 869274
rect 675017 869216 675022 869272
rect 675078 869216 675390 869272
rect 675446 869216 675451 869272
rect 675017 869214 675451 869216
rect 675017 869211 675083 869214
rect 675385 869211 675451 869214
rect 651465 868594 651531 868597
rect 649950 868592 651531 868594
rect 649950 868536 651470 868592
rect 651526 868536 651531 868592
rect 649950 868534 651531 868536
rect 649950 868246 650010 868534
rect 651465 868531 651531 868534
rect 652017 867642 652083 867645
rect 649950 867640 652083 867642
rect 649950 867584 652022 867640
rect 652078 867584 652083 867640
rect 649950 867582 652083 867584
rect 649950 867064 650010 867582
rect 652017 867579 652083 867582
rect 675109 867234 675175 867237
rect 675702 867234 675708 867236
rect 675109 867232 675708 867234
rect 675109 867176 675114 867232
rect 675170 867176 675708 867232
rect 675109 867174 675708 867176
rect 675109 867171 675175 867174
rect 675702 867172 675708 867174
rect 675772 867172 675778 867236
rect 651465 866282 651531 866285
rect 649950 866280 651531 866282
rect 649950 866224 651470 866280
rect 651526 866224 651531 866280
rect 649950 866222 651531 866224
rect 649950 865882 650010 866222
rect 651465 866219 651531 866222
rect 674833 866282 674899 866285
rect 675385 866282 675451 866285
rect 674833 866280 675451 866282
rect 674833 866224 674838 866280
rect 674894 866224 675390 866280
rect 675446 866224 675451 866280
rect 674833 866222 675451 866224
rect 674833 866219 674899 866222
rect 675385 866219 675451 866222
rect 675109 865738 675175 865741
rect 675886 865738 675892 865740
rect 675109 865736 675892 865738
rect 675109 865680 675114 865736
rect 675170 865680 675892 865736
rect 675109 865678 675892 865680
rect 675109 865675 675175 865678
rect 675886 865676 675892 865678
rect 675956 865676 675962 865740
rect 675753 865466 675819 865469
rect 676070 865466 676076 865468
rect 675753 865464 676076 865466
rect 675753 865408 675758 865464
rect 675814 865408 676076 865464
rect 675753 865406 676076 865408
rect 675753 865403 675819 865406
rect 676070 865404 676076 865406
rect 676140 865404 676146 865468
rect 651373 865194 651439 865197
rect 649950 865192 651439 865194
rect 649950 865136 651378 865192
rect 651434 865136 651439 865192
rect 649950 865134 651439 865136
rect 649950 864700 650010 865134
rect 651373 865131 651439 865134
rect 651465 863834 651531 863837
rect 649766 863832 651531 863834
rect 649766 863776 651470 863832
rect 651526 863776 651531 863832
rect 649766 863774 651531 863776
rect 649766 863518 649826 863774
rect 651465 863771 651531 863774
rect 651465 862338 651531 862341
rect 649766 862336 651531 862338
rect 649766 862280 651470 862336
rect 651526 862280 651531 862336
rect 649766 862278 651531 862280
rect 651465 862275 651531 862278
rect 35617 818002 35683 818005
rect 35574 818000 35683 818002
rect 35574 817944 35622 818000
rect 35678 817944 35683 818000
rect 35574 817939 35683 817944
rect 35574 817700 35634 817939
rect 35801 817322 35867 817325
rect 35788 817320 35867 817322
rect 35788 817264 35806 817320
rect 35862 817264 35867 817320
rect 35788 817262 35867 817264
rect 35801 817259 35867 817262
rect 35617 816914 35683 816917
rect 35604 816912 35683 816914
rect 35604 816856 35622 816912
rect 35678 816856 35683 816912
rect 35604 816854 35683 816856
rect 35617 816851 35683 816854
rect 35801 816098 35867 816101
rect 35788 816096 35867 816098
rect 35788 816040 35806 816096
rect 35862 816040 35867 816096
rect 35788 816038 35867 816040
rect 35801 816035 35867 816038
rect 35617 815282 35683 815285
rect 35604 815280 35683 815282
rect 35604 815224 35622 815280
rect 35678 815224 35683 815280
rect 35604 815222 35683 815224
rect 35617 815219 35683 815222
rect 35801 814466 35867 814469
rect 35788 814464 35867 814466
rect 35788 814408 35806 814464
rect 35862 814408 35867 814464
rect 35788 814406 35867 814408
rect 35801 814403 35867 814406
rect 41321 813650 41387 813653
rect 41308 813648 41387 813650
rect 41308 813592 41326 813648
rect 41382 813592 41387 813648
rect 41308 813590 41387 813592
rect 41321 813587 41387 813590
rect 42006 813242 42012 813244
rect 41492 813182 42012 813242
rect 42006 813180 42012 813182
rect 42076 813180 42082 813244
rect 31661 812834 31727 812837
rect 31661 812832 31740 812834
rect 31661 812776 31666 812832
rect 31722 812776 31740 812832
rect 31661 812774 31740 812776
rect 31661 812771 31727 812774
rect 41321 812426 41387 812429
rect 41308 812424 41387 812426
rect 41308 812368 41326 812424
rect 41382 812368 41387 812424
rect 41308 812366 41387 812368
rect 41321 812363 41387 812366
rect 35157 812018 35223 812021
rect 35157 812016 35236 812018
rect 35157 811960 35162 812016
rect 35218 811960 35236 812016
rect 35157 811958 35236 811960
rect 35157 811955 35223 811958
rect 39297 811610 39363 811613
rect 39284 811608 39363 811610
rect 39284 811552 39302 811608
rect 39358 811552 39363 811608
rect 39284 811550 39363 811552
rect 39297 811547 39363 811550
rect 41781 811338 41847 811341
rect 42190 811338 42196 811340
rect 41781 811336 42196 811338
rect 41781 811280 41786 811336
rect 41842 811280 42196 811336
rect 41781 811278 42196 811280
rect 41781 811275 41847 811278
rect 42190 811276 42196 811278
rect 42260 811276 42266 811340
rect 32213 811202 32279 811205
rect 32213 811200 32292 811202
rect 32213 811144 32218 811200
rect 32274 811144 32292 811200
rect 32213 811142 32292 811144
rect 32213 811139 32279 811142
rect 41781 810794 41847 810797
rect 41492 810792 41847 810794
rect 41492 810736 41786 810792
rect 41842 810736 41847 810792
rect 41492 810734 41847 810736
rect 41781 810731 41847 810734
rect 42149 810386 42215 810389
rect 41492 810384 42215 810386
rect 41492 810328 42154 810384
rect 42210 810328 42215 810384
rect 41492 810326 42215 810328
rect 42149 810323 42215 810326
rect 31017 809978 31083 809981
rect 31004 809976 31083 809978
rect 31004 809920 31022 809976
rect 31078 809920 31083 809976
rect 31004 809918 31083 809920
rect 31017 809915 31083 809918
rect 33734 809403 33794 809540
rect 33734 809398 33843 809403
rect 33734 809342 33782 809398
rect 33838 809342 33843 809398
rect 33734 809340 33843 809342
rect 33777 809337 33843 809340
rect 30281 809162 30347 809165
rect 30268 809160 30347 809162
rect 30268 809104 30286 809160
rect 30342 809104 30347 809160
rect 30268 809102 30347 809104
rect 30281 809099 30347 809102
rect 41321 808754 41387 808757
rect 41308 808752 41387 808754
rect 41308 808696 41326 808752
rect 41382 808696 41387 808752
rect 41308 808694 41387 808696
rect 41321 808691 41387 808694
rect 41137 808346 41203 808349
rect 41124 808344 41203 808346
rect 41124 808288 41142 808344
rect 41198 808288 41203 808344
rect 41124 808286 41203 808288
rect 41137 808283 41203 808286
rect 41965 807938 42031 807941
rect 41492 807936 42031 807938
rect 41492 807880 41970 807936
rect 42026 807880 42031 807936
rect 41492 807878 42031 807880
rect 41965 807875 42031 807878
rect 41321 807530 41387 807533
rect 41308 807528 41387 807530
rect 41308 807472 41326 807528
rect 41382 807472 41387 807528
rect 41308 807470 41387 807472
rect 41321 807467 41387 807470
rect 41094 806717 41154 807092
rect 41094 806712 41203 806717
rect 41094 806684 41142 806712
rect 41124 806656 41142 806684
rect 41198 806656 41203 806712
rect 41124 806654 41203 806656
rect 41137 806651 41203 806654
rect 41321 806306 41387 806309
rect 41308 806304 41387 806306
rect 41308 806248 41326 806304
rect 41382 806248 41387 806304
rect 41308 806246 41387 806248
rect 41321 806243 41387 806246
rect 40534 805564 40540 805628
rect 40604 805626 40610 805628
rect 41781 805626 41847 805629
rect 40604 805624 41847 805626
rect 40604 805568 41786 805624
rect 41842 805568 41847 805624
rect 40604 805566 41847 805568
rect 40604 805564 40610 805566
rect 41781 805563 41847 805566
rect 40902 804748 40908 804812
rect 40972 804810 40978 804812
rect 41965 804810 42031 804813
rect 40972 804808 42031 804810
rect 40972 804752 41970 804808
rect 42026 804752 42031 804808
rect 40972 804750 42031 804752
rect 40972 804748 40978 804750
rect 41965 804747 42031 804750
rect 40718 804476 40724 804540
rect 40788 804538 40794 804540
rect 41965 804538 42031 804541
rect 40788 804536 42031 804538
rect 40788 804480 41970 804536
rect 42026 804480 42031 804536
rect 40788 804478 42031 804480
rect 40788 804476 40794 804478
rect 41965 804475 42031 804478
rect 35157 802498 35223 802501
rect 41822 802498 41828 802500
rect 35157 802496 41828 802498
rect 35157 802440 35162 802496
rect 35218 802440 41828 802496
rect 35157 802438 41828 802440
rect 35157 802435 35223 802438
rect 41822 802436 41828 802438
rect 41892 802436 41898 802500
rect 40493 800730 40559 800733
rect 41086 800730 41092 800732
rect 40493 800728 41092 800730
rect 40493 800672 40498 800728
rect 40554 800672 41092 800728
rect 40493 800670 41092 800672
rect 40493 800667 40559 800670
rect 41086 800668 41092 800670
rect 41156 800668 41162 800732
rect 39297 800594 39363 800597
rect 40350 800594 40356 800596
rect 39297 800592 40356 800594
rect 39297 800536 39302 800592
rect 39358 800536 40356 800592
rect 39297 800534 40356 800536
rect 39297 800531 39363 800534
rect 40350 800532 40356 800534
rect 40420 800532 40426 800596
rect 41781 800320 41847 800325
rect 41781 800264 41786 800320
rect 41842 800264 41847 800320
rect 41781 800259 41847 800264
rect 41784 799917 41844 800259
rect 41781 799912 41847 799917
rect 41781 799856 41786 799912
rect 41842 799856 41847 799912
rect 41781 799851 41847 799856
rect 42149 797330 42215 797333
rect 43621 797330 43687 797333
rect 42149 797328 43687 797330
rect 42149 797272 42154 797328
rect 42210 797272 43626 797328
rect 43682 797272 43687 797328
rect 42149 797270 43687 797272
rect 42149 797267 42215 797270
rect 43621 797267 43687 797270
rect 42149 795426 42215 795429
rect 45001 795426 45067 795429
rect 42149 795424 45067 795426
rect 42149 795368 42154 795424
rect 42210 795368 45006 795424
rect 45062 795368 45067 795424
rect 42149 795366 45067 795368
rect 42149 795363 42215 795366
rect 45001 795363 45067 795366
rect 40902 794820 40908 794884
rect 40972 794882 40978 794884
rect 41781 794882 41847 794885
rect 40972 794880 41847 794882
rect 40972 794824 41786 794880
rect 41842 794824 41847 794880
rect 40972 794822 41847 794824
rect 40972 794820 40978 794822
rect 41781 794819 41847 794822
rect 42057 793522 42123 793525
rect 42701 793522 42767 793525
rect 42057 793520 42767 793522
rect 42057 793464 42062 793520
rect 42118 793464 42706 793520
rect 42762 793464 42767 793520
rect 42057 793462 42767 793464
rect 42057 793459 42123 793462
rect 42701 793459 42767 793462
rect 40350 793052 40356 793116
rect 40420 793114 40426 793116
rect 41781 793114 41847 793117
rect 40420 793112 41847 793114
rect 40420 793056 41786 793112
rect 41842 793056 41847 793112
rect 40420 793054 41847 793056
rect 40420 793052 40426 793054
rect 41781 793051 41847 793054
rect 41086 792644 41092 792708
rect 41156 792706 41162 792708
rect 42425 792706 42491 792709
rect 41156 792704 42491 792706
rect 41156 792648 42430 792704
rect 42486 792648 42491 792704
rect 41156 792646 42491 792648
rect 41156 792644 41162 792646
rect 42425 792643 42491 792646
rect 41822 791556 41828 791620
rect 41892 791618 41898 791620
rect 42609 791618 42675 791621
rect 41892 791616 42675 791618
rect 41892 791560 42614 791616
rect 42670 791560 42675 791616
rect 41892 791558 42675 791560
rect 41892 791556 41898 791558
rect 42609 791555 42675 791558
rect 40718 791284 40724 791348
rect 40788 791346 40794 791348
rect 42241 791346 42307 791349
rect 40788 791344 42307 791346
rect 40788 791288 42246 791344
rect 42302 791288 42307 791344
rect 40788 791286 42307 791288
rect 40788 791284 40794 791286
rect 42241 791283 42307 791286
rect 42057 790666 42123 790669
rect 43069 790666 43135 790669
rect 42057 790664 43135 790666
rect 42057 790608 42062 790664
rect 42118 790608 43074 790664
rect 43130 790608 43135 790664
rect 42057 790606 43135 790608
rect 42057 790603 42123 790606
rect 43069 790603 43135 790606
rect 62205 790530 62271 790533
rect 62205 790528 64706 790530
rect 62205 790472 62210 790528
rect 62266 790472 64706 790528
rect 62205 790470 64706 790472
rect 62205 790467 62271 790470
rect 64646 790304 64706 790470
rect 62113 789170 62179 789173
rect 62113 789168 64706 789170
rect 62113 789112 62118 789168
rect 62174 789112 64706 789168
rect 62113 789110 64706 789112
rect 62113 789107 62179 789110
rect 41638 788156 41644 788220
rect 41708 788218 41714 788220
rect 42241 788218 42307 788221
rect 41708 788216 42307 788218
rect 41708 788160 42246 788216
rect 42302 788160 42307 788216
rect 41708 788158 42307 788160
rect 41708 788156 41714 788158
rect 42241 788155 42307 788158
rect 675753 788082 675819 788085
rect 676070 788082 676076 788084
rect 675753 788080 676076 788082
rect 675753 788024 675758 788080
rect 675814 788024 676076 788080
rect 675753 788022 676076 788024
rect 675753 788019 675819 788022
rect 676070 788020 676076 788022
rect 676140 788020 676146 788084
rect 62113 787402 62179 787405
rect 64646 787402 64706 787940
rect 62113 787400 64706 787402
rect 62113 787344 62118 787400
rect 62174 787344 64706 787400
rect 62113 787342 64706 787344
rect 62113 787339 62179 787342
rect 62757 787130 62823 787133
rect 62757 787128 64706 787130
rect 62757 787072 62762 787128
rect 62818 787072 64706 787128
rect 62757 787070 64706 787072
rect 62757 787067 62823 787070
rect 41454 786796 41460 786860
rect 41524 786858 41530 786860
rect 41781 786858 41847 786861
rect 41524 786856 41847 786858
rect 41524 786800 41786 786856
rect 41842 786800 41847 786856
rect 41524 786798 41847 786800
rect 41524 786796 41530 786798
rect 41781 786795 41847 786798
rect 64646 786758 64706 787070
rect 674414 786660 674420 786724
rect 674484 786722 674490 786724
rect 675109 786722 675175 786725
rect 674484 786720 675175 786722
rect 674484 786664 675114 786720
rect 675170 786664 675175 786720
rect 674484 786662 675175 786664
rect 674484 786660 674490 786662
rect 675109 786659 675175 786662
rect 40534 786116 40540 786180
rect 40604 786178 40610 786180
rect 41781 786178 41847 786181
rect 40604 786176 41847 786178
rect 40604 786120 41786 786176
rect 41842 786120 41847 786176
rect 40604 786118 41847 786120
rect 40604 786116 40610 786118
rect 41781 786115 41847 786118
rect 61377 786178 61443 786181
rect 61377 786176 64706 786178
rect 61377 786120 61382 786176
rect 61438 786120 64706 786176
rect 61377 786118 64706 786120
rect 61377 786115 61443 786118
rect 64646 785576 64706 786118
rect 62113 784954 62179 784957
rect 62113 784952 64706 784954
rect 62113 784896 62118 784952
rect 62174 784896 64706 784952
rect 62113 784894 64706 784896
rect 62113 784891 62179 784894
rect 64646 784394 64706 784894
rect 674598 784620 674604 784684
rect 674668 784682 674674 784684
rect 675109 784682 675175 784685
rect 674668 784680 675175 784682
rect 674668 784624 675114 784680
rect 675170 784624 675175 784680
rect 674668 784622 675175 784624
rect 674668 784620 674674 784622
rect 675109 784619 675175 784622
rect 675150 780540 675156 780604
rect 675220 780602 675226 780604
rect 675477 780602 675543 780605
rect 675220 780600 675543 780602
rect 675220 780544 675482 780600
rect 675538 780544 675543 780600
rect 675220 780542 675543 780544
rect 675220 780540 675226 780542
rect 675477 780539 675543 780542
rect 673729 780058 673795 780061
rect 675477 780058 675543 780061
rect 673729 780056 675543 780058
rect 673729 780000 673734 780056
rect 673790 780000 675482 780056
rect 675538 780000 675543 780056
rect 673729 779998 675543 780000
rect 673729 779995 673795 779998
rect 675477 779995 675543 779998
rect 674649 779242 674715 779245
rect 675385 779242 675451 779245
rect 674649 779240 675451 779242
rect 674649 779184 674654 779240
rect 674710 779184 675390 779240
rect 675446 779184 675451 779240
rect 674649 779182 675451 779184
rect 674649 779179 674715 779182
rect 675385 779179 675451 779182
rect 672993 778834 673059 778837
rect 675477 778834 675543 778837
rect 672993 778832 675543 778834
rect 649950 778426 650010 778824
rect 672993 778776 672998 778832
rect 673054 778776 675482 778832
rect 675538 778776 675543 778832
rect 672993 778774 675543 778776
rect 672993 778771 673059 778774
rect 675477 778771 675543 778774
rect 651465 778426 651531 778429
rect 649950 778424 651531 778426
rect 649950 778368 651470 778424
rect 651526 778368 651531 778424
rect 649950 778366 651531 778368
rect 651465 778363 651531 778366
rect 649950 777066 650010 777642
rect 652017 777066 652083 777069
rect 649950 777064 652083 777066
rect 649950 777008 652022 777064
rect 652078 777008 652083 777064
rect 649950 777006 652083 777008
rect 652017 777003 652083 777006
rect 649950 776114 650010 776460
rect 674833 776250 674899 776253
rect 674833 776248 676230 776250
rect 674833 776192 674838 776248
rect 674894 776192 676230 776248
rect 674833 776190 676230 776192
rect 674833 776187 674899 776190
rect 651465 776114 651531 776117
rect 649950 776112 651531 776114
rect 649950 776056 651470 776112
rect 651526 776056 651531 776112
rect 649950 776054 651531 776056
rect 676170 776114 676230 776190
rect 676806 776114 676812 776116
rect 676170 776054 676812 776114
rect 651465 776051 651531 776054
rect 676806 776052 676812 776054
rect 676876 776052 676882 776116
rect 669773 775842 669839 775845
rect 675477 775842 675543 775845
rect 669773 775840 675543 775842
rect 669773 775784 669778 775840
rect 669834 775784 675482 775840
rect 675538 775784 675543 775840
rect 669773 775782 675543 775784
rect 669773 775779 669839 775782
rect 675477 775779 675543 775782
rect 675109 775572 675175 775573
rect 675109 775570 675156 775572
rect 675064 775568 675156 775570
rect 675064 775512 675114 775568
rect 675064 775510 675156 775512
rect 675109 775508 675156 775510
rect 675220 775508 675226 775572
rect 675109 775507 675175 775508
rect 651373 775298 651439 775301
rect 649950 775296 651439 775298
rect 649950 775240 651378 775296
rect 651434 775240 651439 775296
rect 649950 775238 651439 775240
rect 651373 775235 651439 775238
rect 668393 775026 668459 775029
rect 675477 775026 675543 775029
rect 668393 775024 675543 775026
rect 668393 774968 668398 775024
rect 668454 774968 675482 775024
rect 675538 774968 675543 775024
rect 668393 774966 675543 774968
rect 668393 774963 668459 774966
rect 675477 774963 675543 774966
rect 35801 774754 35867 774757
rect 35758 774752 35867 774754
rect 35758 774696 35806 774752
rect 35862 774696 35867 774752
rect 35758 774691 35867 774696
rect 35758 774452 35818 774691
rect 674833 774618 674899 774621
rect 675477 774618 675543 774621
rect 674833 774616 675543 774618
rect 674833 774560 674838 774616
rect 674894 774560 675482 774616
rect 675538 774560 675543 774616
rect 674833 774558 675543 774560
rect 674833 774555 674899 774558
rect 675477 774555 675543 774558
rect 651465 774210 651531 774213
rect 649950 774208 651531 774210
rect 649950 774152 651470 774208
rect 651526 774152 651531 774208
rect 649950 774150 651531 774152
rect 649950 774096 650010 774150
rect 651465 774147 651531 774150
rect 35206 773941 35266 774044
rect 35206 773936 35315 773941
rect 35206 773880 35254 773936
rect 35310 773880 35315 773936
rect 35206 773878 35315 773880
rect 35249 773875 35315 773878
rect 35574 773533 35634 773636
rect 35574 773528 35683 773533
rect 35574 773472 35622 773528
rect 35678 773472 35683 773528
rect 35574 773470 35683 773472
rect 35617 773467 35683 773470
rect 651465 773394 651531 773397
rect 649950 773392 651531 773394
rect 649950 773336 651470 773392
rect 651526 773336 651531 773392
rect 649950 773334 651531 773336
rect 35758 773125 35818 773228
rect 35433 773122 35499 773125
rect 35390 773120 35499 773122
rect 35390 773064 35438 773120
rect 35494 773064 35499 773120
rect 35390 773059 35499 773064
rect 35758 773120 35867 773125
rect 35758 773064 35806 773120
rect 35862 773064 35867 773120
rect 35758 773062 35867 773064
rect 35801 773059 35867 773062
rect 41505 773122 41571 773125
rect 44909 773122 44975 773125
rect 41505 773120 44975 773122
rect 41505 773064 41510 773120
rect 41566 773064 44914 773120
rect 44970 773064 44975 773120
rect 41505 773062 44975 773064
rect 41505 773059 41571 773062
rect 44909 773059 44975 773062
rect 35390 772820 35450 773059
rect 649950 772914 650010 773334
rect 651465 773331 651531 773334
rect 35574 772309 35634 772412
rect 35574 772304 35683 772309
rect 35574 772248 35622 772304
rect 35678 772248 35683 772304
rect 35574 772246 35683 772248
rect 35617 772243 35683 772246
rect 35758 771901 35818 772004
rect 35758 771896 35867 771901
rect 35758 771840 35806 771896
rect 35862 771840 35867 771896
rect 35758 771838 35867 771840
rect 35801 771835 35867 771838
rect 35758 771493 35818 771596
rect 35758 771488 35867 771493
rect 35758 771432 35806 771488
rect 35862 771432 35867 771488
rect 35758 771430 35867 771432
rect 35801 771427 35867 771430
rect 35574 771085 35634 771188
rect 35574 771080 35683 771085
rect 35574 771024 35622 771080
rect 35678 771024 35683 771080
rect 35574 771022 35683 771024
rect 35617 771019 35683 771022
rect 35758 770677 35818 770780
rect 35758 770672 35867 770677
rect 35758 770616 35806 770672
rect 35862 770616 35867 770672
rect 35758 770614 35867 770616
rect 35801 770611 35867 770614
rect 39113 770674 39179 770677
rect 43253 770674 43319 770677
rect 39113 770672 43319 770674
rect 39113 770616 39118 770672
rect 39174 770616 43258 770672
rect 43314 770616 43319 770672
rect 39113 770614 43319 770616
rect 39113 770611 39179 770614
rect 43253 770611 43319 770614
rect 35758 770269 35818 770372
rect 35758 770264 35867 770269
rect 35758 770208 35806 770264
rect 35862 770208 35867 770264
rect 35758 770206 35867 770208
rect 35801 770203 35867 770206
rect 39481 770266 39547 770269
rect 43069 770266 43135 770269
rect 39481 770264 43135 770266
rect 39481 770208 39486 770264
rect 39542 770208 43074 770264
rect 43130 770208 43135 770264
rect 39481 770206 43135 770208
rect 39481 770203 39547 770206
rect 43069 770203 43135 770206
rect 41462 769860 41522 769964
rect 41454 769796 41460 769860
rect 41524 769796 41530 769860
rect 35758 769453 35818 769556
rect 35758 769448 35867 769453
rect 35758 769392 35806 769448
rect 35862 769392 35867 769448
rect 35758 769390 35867 769392
rect 35801 769387 35867 769390
rect 39849 769450 39915 769453
rect 44541 769450 44607 769453
rect 39849 769448 44607 769450
rect 39849 769392 39854 769448
rect 39910 769392 44546 769448
rect 44602 769392 44607 769448
rect 39849 769390 44607 769392
rect 39849 769387 39915 769390
rect 44541 769387 44607 769390
rect 35574 769045 35634 769148
rect 35574 769040 35683 769045
rect 35574 768984 35622 769040
rect 35678 768984 35683 769040
rect 35574 768982 35683 768984
rect 35617 768979 35683 768982
rect 35758 768637 35818 768740
rect 35758 768632 35867 768637
rect 35758 768576 35806 768632
rect 35862 768576 35867 768632
rect 35758 768574 35867 768576
rect 35801 768571 35867 768574
rect 35206 768229 35266 768332
rect 35157 768224 35266 768229
rect 35157 768168 35162 768224
rect 35218 768168 35266 768224
rect 35157 768166 35266 768168
rect 35157 768163 35223 768166
rect 32446 767821 32506 767924
rect 32397 767816 32506 767821
rect 32397 767760 32402 767816
rect 32458 767760 32506 767816
rect 32397 767758 32506 767760
rect 32397 767755 32463 767758
rect 35758 767413 35818 767516
rect 35758 767408 35867 767413
rect 35758 767352 35806 767408
rect 35862 767352 35867 767408
rect 35758 767350 35867 767352
rect 35801 767347 35867 767350
rect 33734 767005 33794 767108
rect 33734 767000 33843 767005
rect 33734 766944 33782 767000
rect 33838 766944 33843 767000
rect 33734 766942 33843 766944
rect 33777 766939 33843 766942
rect 40033 767002 40099 767005
rect 41638 767002 41644 767004
rect 40033 767000 41644 767002
rect 40033 766944 40038 767000
rect 40094 766944 41644 767000
rect 40033 766942 41644 766944
rect 40033 766939 40099 766942
rect 41638 766940 41644 766942
rect 41708 766940 41714 767004
rect 40726 766596 40786 766700
rect 40718 766532 40724 766596
rect 40788 766532 40794 766596
rect 35758 766189 35818 766292
rect 35758 766184 35867 766189
rect 35758 766128 35806 766184
rect 35862 766128 35867 766184
rect 35758 766126 35867 766128
rect 35801 766123 35867 766126
rect 35758 765781 35818 765884
rect 35758 765776 35867 765781
rect 35758 765720 35806 765776
rect 35862 765720 35867 765776
rect 35758 765718 35867 765720
rect 35801 765715 35867 765718
rect 40542 765372 40602 765476
rect 40534 765308 40540 765372
rect 40604 765308 40610 765372
rect 40910 764964 40970 765068
rect 40902 764900 40908 764964
rect 40972 764900 40978 764964
rect 35758 764557 35818 764660
rect 35758 764552 35867 764557
rect 35758 764496 35806 764552
rect 35862 764496 35867 764552
rect 35758 764494 35867 764496
rect 35801 764491 35867 764494
rect 39573 764554 39639 764557
rect 44357 764554 44423 764557
rect 39573 764552 44423 764554
rect 39573 764496 39578 764552
rect 39634 764496 44362 764552
rect 44418 764496 44423 764552
rect 39573 764494 44423 764496
rect 39573 764491 39639 764494
rect 44357 764491 44423 764494
rect 35574 764149 35634 764252
rect 35574 764144 35683 764149
rect 35574 764088 35622 764144
rect 35678 764088 35683 764144
rect 35574 764086 35683 764088
rect 35617 764083 35683 764086
rect 39757 764146 39823 764149
rect 42425 764146 42491 764149
rect 39757 764144 42491 764146
rect 39757 764088 39762 764144
rect 39818 764088 42430 764144
rect 42486 764088 42491 764144
rect 39757 764086 42491 764088
rect 39757 764083 39823 764086
rect 42425 764083 42491 764086
rect 35801 763738 35867 763741
rect 35758 763736 35867 763738
rect 35758 763680 35806 763736
rect 35862 763680 35867 763736
rect 35758 763675 35867 763680
rect 35758 763436 35818 763675
rect 37578 763432 37656 763932
rect 40493 763330 40559 763333
rect 45553 763330 45619 763333
rect 40493 763328 45619 763330
rect 40493 763272 40498 763328
rect 40554 763272 45558 763328
rect 45614 763272 45619 763328
rect 40493 763270 45619 763272
rect 40493 763267 40559 763270
rect 45553 763267 45619 763270
rect 35758 762925 35818 763028
rect 35758 762920 35867 762925
rect 35758 762864 35806 762920
rect 35862 762864 35867 762920
rect 35758 762862 35867 762864
rect 35801 762859 35867 762862
rect 40125 761834 40191 761837
rect 42609 761834 42675 761837
rect 40125 761832 42675 761834
rect 40125 761776 40130 761832
rect 40186 761776 42614 761832
rect 42670 761776 42675 761832
rect 40125 761774 42675 761776
rect 40125 761771 40191 761774
rect 42609 761771 42675 761774
rect 39941 758570 40007 758573
rect 43253 758570 43319 758573
rect 39941 758568 43319 758570
rect 39941 758512 39946 758568
rect 40002 758512 43258 758568
rect 43314 758512 43319 758568
rect 39941 758510 43319 758512
rect 39941 758507 40007 758510
rect 43253 758507 43319 758510
rect 36537 757754 36603 757757
rect 41822 757754 41828 757756
rect 36537 757752 41828 757754
rect 36537 757696 36542 757752
rect 36598 757696 41828 757752
rect 36537 757694 41828 757696
rect 36537 757691 36603 757694
rect 41822 757692 41828 757694
rect 41892 757692 41898 757756
rect 39849 757346 39915 757349
rect 40350 757346 40356 757348
rect 39849 757344 40356 757346
rect 39849 757288 39854 757344
rect 39910 757288 40356 757344
rect 39849 757286 40356 757288
rect 39849 757283 39915 757286
rect 40350 757284 40356 757286
rect 40420 757284 40426 757348
rect 41965 757212 42031 757213
rect 41965 757208 42012 757212
rect 42076 757210 42082 757212
rect 41965 757152 41970 757208
rect 41965 757148 42012 757152
rect 42076 757150 42122 757210
rect 42076 757148 42082 757150
rect 41965 757147 42031 757148
rect 41781 757074 41847 757077
rect 41781 757072 41890 757074
rect 41781 757016 41786 757072
rect 41842 757016 41890 757072
rect 41781 757011 41890 757016
rect 41830 756669 41890 757011
rect 41830 756664 41939 756669
rect 41830 756608 41878 756664
rect 41934 756608 41939 756664
rect 41830 756606 41939 756608
rect 41873 756603 41939 756606
rect 40902 754020 40908 754084
rect 40972 754082 40978 754084
rect 42241 754082 42307 754085
rect 40972 754080 42307 754082
rect 40972 754024 42246 754080
rect 42302 754024 42307 754080
rect 40972 754022 42307 754024
rect 40972 754020 40978 754022
rect 42241 754019 42307 754022
rect 40350 753612 40356 753676
rect 40420 753674 40426 753676
rect 42609 753674 42675 753677
rect 40420 753672 42675 753674
rect 40420 753616 42614 753672
rect 42670 753616 42675 753672
rect 40420 753614 42675 753616
rect 40420 753612 40426 753614
rect 42609 753611 42675 753614
rect 42149 753404 42215 753405
rect 42149 753400 42196 753404
rect 42260 753402 42266 753404
rect 42149 753344 42154 753400
rect 42149 753340 42196 753344
rect 42260 753342 42306 753402
rect 42260 753340 42266 753342
rect 42149 753339 42215 753340
rect 42057 752994 42123 752997
rect 44357 752994 44423 752997
rect 42057 752992 44423 752994
rect 42057 752936 42062 752992
rect 42118 752936 44362 752992
rect 44418 752936 44423 752992
rect 42057 752934 44423 752936
rect 42057 752931 42123 752934
rect 44357 752931 44423 752934
rect 44173 751906 44239 751909
rect 41876 751904 44239 751906
rect 41876 751848 44178 751904
rect 44234 751848 44239 751904
rect 41876 751846 44239 751848
rect 41876 751637 41936 751846
rect 44173 751843 44239 751846
rect 41873 751632 41939 751637
rect 41873 751576 41878 751632
rect 41934 751576 41939 751632
rect 41873 751571 41939 751576
rect 42057 751634 42123 751637
rect 45093 751634 45159 751637
rect 42057 751632 45159 751634
rect 42057 751576 42062 751632
rect 42118 751576 45098 751632
rect 45154 751576 45159 751632
rect 42057 751574 45159 751576
rect 42057 751571 42123 751574
rect 45093 751571 45159 751574
rect 41965 750546 42031 750549
rect 42190 750546 42196 750548
rect 41965 750544 42196 750546
rect 41965 750488 41970 750544
rect 42026 750488 42196 750544
rect 41965 750486 42196 750488
rect 41965 750483 42031 750486
rect 42190 750484 42196 750486
rect 42260 750484 42266 750548
rect 41965 749732 42031 749733
rect 41965 749728 42012 749732
rect 42076 749730 42082 749732
rect 41965 749672 41970 749728
rect 41965 749668 42012 749672
rect 42076 749670 42122 749730
rect 42076 749668 42082 749670
rect 41965 749667 42031 749668
rect 40534 749396 40540 749460
rect 40604 749458 40610 749460
rect 42241 749458 42307 749461
rect 40604 749456 42307 749458
rect 40604 749400 42246 749456
rect 42302 749400 42307 749456
rect 40604 749398 42307 749400
rect 40604 749396 40610 749398
rect 42241 749395 42307 749398
rect 62757 747690 62823 747693
rect 62757 747688 64706 747690
rect 62757 747632 62762 747688
rect 62818 747632 64706 747688
rect 62757 747630 64706 747632
rect 62757 747627 62823 747630
rect 64646 747082 64706 747630
rect 40718 746812 40724 746876
rect 40788 746874 40794 746876
rect 41781 746874 41847 746877
rect 40788 746872 41847 746874
rect 40788 746816 41786 746872
rect 41842 746816 41847 746872
rect 40788 746814 41847 746816
rect 40788 746812 40794 746814
rect 41781 746811 41847 746814
rect 62113 746194 62179 746197
rect 62113 746192 64706 746194
rect 62113 746136 62118 746192
rect 62174 746136 64706 746192
rect 62113 746134 64706 746136
rect 62113 746131 62179 746134
rect 64646 745900 64706 746134
rect 41965 745650 42031 745653
rect 42793 745650 42859 745653
rect 41965 745648 42859 745650
rect 41965 745592 41970 745648
rect 42026 745592 42798 745648
rect 42854 745592 42859 745648
rect 41965 745590 42859 745592
rect 41965 745587 42031 745590
rect 42793 745587 42859 745590
rect 41822 745316 41828 745380
rect 41892 745378 41898 745380
rect 42241 745378 42307 745381
rect 41892 745376 42307 745378
rect 41892 745320 42246 745376
rect 42302 745320 42307 745376
rect 41892 745318 42307 745320
rect 41892 745316 41898 745318
rect 42241 745315 42307 745318
rect 41638 744364 41644 744428
rect 41708 744426 41714 744428
rect 42517 744426 42583 744429
rect 41708 744424 42583 744426
rect 41708 744368 42522 744424
rect 42578 744368 42583 744424
rect 41708 744366 42583 744368
rect 41708 744364 41714 744366
rect 42517 744363 42583 744366
rect 62113 744154 62179 744157
rect 64646 744154 64706 744718
rect 62113 744152 64706 744154
rect 62113 744096 62118 744152
rect 62174 744096 64706 744152
rect 62113 744094 64706 744096
rect 62113 744091 62179 744094
rect 41454 743684 41460 743748
rect 41524 743746 41530 743748
rect 41781 743746 41847 743749
rect 41524 743744 41847 743746
rect 41524 743688 41786 743744
rect 41842 743688 41847 743744
rect 41524 743686 41847 743688
rect 41524 743684 41530 743686
rect 41781 743683 41847 743686
rect 62113 743746 62179 743749
rect 62113 743744 64706 743746
rect 62113 743688 62118 743744
rect 62174 743688 64706 743744
rect 62113 743686 64706 743688
rect 62113 743683 62179 743686
rect 64646 743536 64706 743686
rect 62113 742386 62179 742389
rect 62113 742384 64706 742386
rect 62113 742328 62118 742384
rect 62174 742328 64706 742384
rect 62113 742326 64706 742328
rect 62113 742323 62179 742326
rect 675385 742252 675451 742253
rect 675334 742250 675340 742252
rect 675294 742190 675340 742250
rect 675404 742248 675451 742252
rect 675446 742192 675451 742248
rect 675334 742188 675340 742190
rect 675404 742188 675451 742192
rect 675385 742187 675451 742188
rect 63033 741842 63099 741845
rect 63033 741840 64706 741842
rect 63033 741784 63038 741840
rect 63094 741784 64706 741840
rect 63033 741782 64706 741784
rect 63033 741779 63099 741782
rect 64646 741172 64706 741782
rect 672533 739938 672599 739941
rect 675477 739938 675543 739941
rect 672533 739936 675543 739938
rect 672533 739880 672538 739936
rect 672594 739880 675482 739936
rect 675538 739880 675543 739936
rect 672533 739878 675543 739880
rect 672533 739875 672599 739878
rect 675477 739875 675543 739878
rect 673545 738714 673611 738717
rect 675477 738714 675543 738717
rect 673545 738712 675543 738714
rect 673545 738656 673550 738712
rect 673606 738656 675482 738712
rect 675538 738656 675543 738712
rect 673545 738654 675543 738656
rect 673545 738651 673611 738654
rect 675477 738651 675543 738654
rect 674230 738108 674236 738172
rect 674300 738170 674306 738172
rect 675477 738170 675543 738173
rect 674300 738168 675543 738170
rect 674300 738112 675482 738168
rect 675538 738112 675543 738168
rect 674300 738110 675543 738112
rect 674300 738108 674306 738110
rect 675477 738107 675543 738110
rect 669589 735722 669655 735725
rect 675385 735722 675451 735725
rect 669589 735720 675451 735722
rect 669589 735664 669594 735720
rect 669650 735664 675390 735720
rect 675446 735664 675451 735720
rect 669589 735662 675451 735664
rect 669589 735659 669655 735662
rect 675385 735659 675451 735662
rect 674097 734906 674163 734909
rect 675477 734906 675543 734909
rect 674097 734904 675543 734906
rect 674097 734848 674102 734904
rect 674158 734848 675482 734904
rect 675538 734848 675543 734904
rect 674097 734846 675543 734848
rect 674097 734843 674163 734846
rect 675477 734843 675543 734846
rect 649950 734226 650010 734402
rect 651465 734226 651531 734229
rect 649950 734224 651531 734226
rect 649950 734168 651470 734224
rect 651526 734168 651531 734224
rect 649950 734166 651531 734168
rect 651465 734163 651531 734166
rect 673913 734226 673979 734229
rect 675477 734226 675543 734229
rect 673913 734224 675543 734226
rect 673913 734168 673918 734224
rect 673974 734168 675482 734224
rect 675538 734168 675543 734224
rect 673913 734166 675543 734168
rect 673913 734163 673979 734166
rect 675477 734163 675543 734166
rect 671613 733818 671679 733821
rect 675569 733818 675635 733821
rect 671613 733816 675635 733818
rect 671613 733760 671618 733816
rect 671674 733760 675574 733816
rect 675630 733760 675635 733816
rect 671613 733758 675635 733760
rect 671613 733755 671679 733758
rect 675569 733755 675635 733758
rect 649950 733002 650010 733220
rect 651465 733002 651531 733005
rect 649950 733000 651531 733002
rect 649950 732944 651470 733000
rect 651526 732944 651531 733000
rect 649950 732942 651531 732944
rect 651465 732939 651531 732942
rect 649950 731778 650010 732038
rect 651465 731778 651531 731781
rect 649950 731776 651531 731778
rect 649950 731720 651470 731776
rect 651526 731720 651531 731776
rect 649950 731718 651531 731720
rect 651465 731715 651531 731718
rect 43437 731370 43503 731373
rect 41492 731368 43503 731370
rect 41492 731312 43442 731368
rect 43498 731312 43503 731368
rect 41492 731310 43503 731312
rect 43437 731307 43503 731310
rect 651465 731098 651531 731101
rect 649950 731096 651531 731098
rect 649950 731040 651470 731096
rect 651526 731040 651531 731096
rect 649950 731038 651531 731040
rect 41137 730962 41203 730965
rect 41124 730960 41203 730962
rect 41124 730904 41142 730960
rect 41198 730904 41203 730960
rect 41124 730902 41203 730904
rect 41137 730899 41203 730902
rect 649950 730856 650010 731038
rect 651465 731035 651531 731038
rect 43621 730554 43687 730557
rect 41492 730552 43687 730554
rect 41492 730496 43626 730552
rect 43682 730496 43687 730552
rect 41492 730494 43687 730496
rect 43621 730491 43687 730494
rect 44909 730146 44975 730149
rect 41492 730144 44975 730146
rect 41492 730088 44914 730144
rect 44970 730088 44975 730144
rect 41492 730086 44975 730088
rect 44909 730083 44975 730086
rect 668945 730146 669011 730149
rect 675477 730146 675543 730149
rect 668945 730144 675543 730146
rect 668945 730088 668950 730144
rect 669006 730088 675482 730144
rect 675538 730088 675543 730144
rect 668945 730086 675543 730088
rect 668945 730083 669011 730086
rect 675477 730083 675543 730086
rect 651465 729874 651531 729877
rect 649950 729872 651531 729874
rect 649950 729816 651470 729872
rect 651526 729816 651531 729872
rect 649950 729814 651531 729816
rect 45185 729738 45251 729741
rect 41492 729736 45251 729738
rect 41492 729680 45190 729736
rect 45246 729680 45251 729736
rect 41492 729678 45251 729680
rect 45185 729675 45251 729678
rect 649950 729674 650010 729814
rect 651465 729811 651531 729814
rect 43069 729330 43135 729333
rect 41492 729328 43135 729330
rect 41492 729272 43074 729328
rect 43130 729272 43135 729328
rect 41492 729270 43135 729272
rect 43069 729267 43135 729270
rect 41278 728687 41338 728892
rect 670325 728786 670391 728789
rect 675477 728786 675543 728789
rect 670325 728784 675543 728786
rect 670325 728728 670330 728784
rect 670386 728728 675482 728784
rect 675538 728728 675543 728784
rect 670325 728726 675543 728728
rect 670325 728723 670391 728726
rect 675477 728723 675543 728726
rect 40769 728684 40835 728687
rect 40726 728682 40835 728684
rect 40726 728626 40774 728682
rect 40830 728626 40835 728682
rect 40726 728621 40835 728626
rect 41278 728682 41387 728687
rect 41278 728626 41326 728682
rect 41382 728626 41387 728682
rect 41278 728624 41387 728626
rect 41321 728621 41387 728624
rect 40726 728484 40786 728621
rect 651465 728514 651531 728517
rect 649950 728512 651531 728514
rect 649950 728456 651470 728512
rect 651526 728456 651531 728512
rect 649950 728454 651531 728456
rect 651465 728451 651531 728454
rect 44265 728106 44331 728109
rect 41492 728104 44331 728106
rect 41492 728048 44270 728104
rect 44326 728048 44331 728104
rect 41492 728046 44331 728048
rect 44265 728043 44331 728046
rect 44541 727698 44607 727701
rect 41492 727696 44607 727698
rect 41492 727640 44546 727696
rect 44602 727640 44607 727696
rect 41492 727638 44607 727640
rect 44541 727635 44607 727638
rect 41045 727460 41111 727463
rect 41045 727458 41154 727460
rect 41045 727402 41050 727458
rect 41106 727402 41154 727458
rect 41045 727397 41154 727402
rect 41094 727260 41154 727397
rect 674925 727290 674991 727293
rect 675334 727290 675340 727292
rect 674925 727288 675340 727290
rect 674925 727232 674930 727288
rect 674986 727232 675340 727288
rect 674925 727230 675340 727232
rect 674925 727227 674991 727230
rect 675334 727228 675340 727230
rect 675404 727228 675410 727292
rect 41137 726882 41203 726885
rect 41124 726880 41203 726882
rect 41124 726824 41142 726880
rect 41198 726824 41203 726880
rect 41124 726822 41203 726824
rect 41137 726819 41203 726822
rect 676070 726548 676076 726612
rect 676140 726610 676146 726612
rect 682377 726610 682443 726613
rect 676140 726608 682443 726610
rect 676140 726552 682382 726608
rect 682438 726552 682443 726608
rect 676140 726550 682443 726552
rect 676140 726548 676146 726550
rect 682377 726547 682443 726550
rect 41278 726239 41338 726444
rect 40953 726236 41019 726239
rect 40910 726234 41019 726236
rect 40910 726178 40958 726234
rect 41014 726178 41019 726234
rect 40910 726173 41019 726178
rect 41278 726234 41387 726239
rect 41278 726178 41326 726234
rect 41382 726178 41387 726234
rect 41278 726176 41387 726178
rect 41321 726173 41387 726176
rect 40910 726036 40970 726173
rect 41781 725796 41847 725797
rect 41781 725794 41828 725796
rect 41736 725792 41828 725794
rect 41736 725736 41786 725792
rect 41736 725734 41828 725736
rect 41781 725732 41828 725734
rect 41892 725732 41898 725796
rect 41781 725731 41847 725732
rect 41321 725658 41387 725661
rect 41308 725656 41387 725658
rect 41308 725600 41326 725656
rect 41382 725600 41387 725656
rect 41308 725598 41387 725600
rect 41321 725595 41387 725598
rect 41137 725250 41203 725253
rect 41124 725248 41203 725250
rect 41124 725192 41142 725248
rect 41198 725192 41203 725248
rect 41124 725190 41203 725192
rect 41137 725187 41203 725190
rect 35157 724842 35223 724845
rect 35157 724840 35236 724842
rect 35157 724784 35162 724840
rect 35218 724784 35236 724840
rect 35157 724782 35236 724784
rect 35157 724779 35223 724782
rect 33041 724434 33107 724437
rect 33028 724432 33107 724434
rect 33028 724376 33046 724432
rect 33102 724376 33107 724432
rect 33028 724374 33107 724376
rect 33041 724371 33107 724374
rect 33734 723791 33794 723996
rect 33734 723786 33843 723791
rect 33734 723730 33782 723786
rect 33838 723730 33843 723786
rect 33734 723728 33843 723730
rect 33777 723725 33843 723728
rect 43437 723618 43503 723621
rect 41492 723616 43503 723618
rect 41492 723560 43442 723616
rect 43498 723560 43503 723616
rect 41492 723558 43503 723560
rect 43437 723555 43503 723558
rect 39297 723210 39363 723213
rect 39284 723208 39363 723210
rect 39284 723152 39302 723208
rect 39358 723152 39363 723208
rect 39284 723150 39363 723152
rect 39297 723147 39363 723150
rect 44449 722802 44515 722805
rect 41492 722800 44515 722802
rect 41492 722744 44454 722800
rect 44510 722744 44515 722800
rect 41492 722742 44515 722744
rect 44449 722739 44515 722742
rect 41781 722394 41847 722397
rect 673821 722396 673887 722397
rect 673821 722394 673868 722396
rect 41492 722392 41847 722394
rect 41492 722336 41786 722392
rect 41842 722336 41847 722392
rect 41492 722334 41847 722336
rect 673776 722392 673868 722394
rect 673776 722336 673826 722392
rect 673776 722334 673868 722336
rect 41781 722331 41847 722334
rect 673821 722332 673868 722334
rect 673932 722332 673938 722396
rect 673821 722331 673887 722332
rect 41822 721986 41828 721988
rect 41492 721926 41828 721986
rect 41822 721924 41828 721926
rect 41892 721924 41898 721988
rect 674097 721852 674163 721853
rect 674046 721850 674052 721852
rect 674006 721790 674052 721850
rect 674116 721848 674163 721852
rect 674158 721792 674163 721848
rect 674046 721788 674052 721790
rect 674116 721788 674163 721792
rect 674097 721787 674163 721788
rect 674925 721714 674991 721717
rect 674925 721712 675034 721714
rect 674925 721656 674930 721712
rect 674986 721656 675034 721712
rect 674925 721651 675034 721656
rect 44633 721578 44699 721581
rect 41492 721576 44699 721578
rect 41492 721520 44638 721576
rect 44694 721520 44699 721576
rect 41492 721518 44699 721520
rect 674974 721578 675034 721651
rect 675334 721578 675340 721580
rect 674974 721518 675340 721578
rect 44633 721515 44699 721518
rect 675334 721516 675340 721518
rect 675404 721516 675410 721580
rect 47209 721170 47275 721173
rect 41492 721168 47275 721170
rect 41492 721112 47214 721168
rect 47270 721112 47275 721168
rect 41492 721110 47275 721112
rect 47209 721107 47275 721110
rect 41462 720354 41522 720732
rect 42057 720354 42123 720357
rect 41462 720352 42123 720354
rect 41462 720324 42062 720352
rect 41492 720296 42062 720324
rect 42118 720296 42123 720352
rect 41492 720294 42123 720296
rect 42057 720291 42123 720294
rect 673862 720020 673868 720084
rect 673932 720082 673938 720084
rect 674189 720082 674255 720085
rect 673932 720080 674255 720082
rect 673932 720024 674194 720080
rect 674250 720024 674255 720080
rect 673932 720022 674255 720024
rect 673932 720020 673938 720022
rect 674189 720019 674255 720022
rect 47025 719946 47091 719949
rect 41492 719944 47091 719946
rect 41492 719888 47030 719944
rect 47086 719888 47091 719944
rect 41492 719886 47091 719888
rect 47025 719883 47091 719886
rect 41321 718858 41387 718861
rect 42057 718858 42123 718861
rect 41321 718856 42123 718858
rect 41321 718800 41326 718856
rect 41382 718800 42062 718856
rect 42118 718800 42123 718856
rect 41321 718798 42123 718800
rect 41321 718795 41387 718798
rect 42057 718795 42123 718798
rect 40534 718524 40540 718588
rect 40604 718586 40610 718588
rect 41781 718586 41847 718589
rect 40604 718584 41847 718586
rect 40604 718528 41786 718584
rect 41842 718528 41847 718584
rect 40604 718526 41847 718528
rect 40604 718524 40610 718526
rect 41781 718523 41847 718526
rect 40718 718252 40724 718316
rect 40788 718314 40794 718316
rect 41822 718314 41828 718316
rect 40788 718254 41828 718314
rect 40788 718252 40794 718254
rect 41822 718252 41828 718254
rect 41892 718252 41898 718316
rect 40953 717634 41019 717637
rect 41638 717634 41644 717636
rect 40953 717632 41644 717634
rect 40953 717576 40958 717632
rect 41014 717576 41644 717632
rect 40953 717574 41644 717576
rect 40953 717571 41019 717574
rect 41638 717572 41644 717574
rect 41708 717572 41714 717636
rect 674005 717092 674071 717093
rect 674005 717090 674052 717092
rect 673960 717088 674052 717090
rect 673960 717032 674010 717088
rect 673960 717030 674052 717032
rect 674005 717028 674052 717030
rect 674116 717028 674122 717092
rect 674005 717027 674071 717028
rect 33041 716818 33107 716821
rect 41822 716818 41828 716820
rect 33041 716816 41828 716818
rect 33041 716760 33046 716816
rect 33102 716760 41828 716816
rect 33041 716758 41828 716760
rect 33041 716755 33107 716758
rect 41822 716756 41828 716758
rect 41892 716756 41898 716820
rect 673821 716546 673887 716549
rect 673821 716544 676292 716546
rect 673821 716488 673826 716544
rect 673882 716488 676292 716544
rect 673821 716486 676292 716488
rect 673821 716483 673887 716486
rect 673821 716138 673887 716141
rect 673821 716136 676292 716138
rect 673821 716080 673826 716136
rect 673882 716080 676292 716136
rect 673821 716078 676292 716080
rect 673821 716075 673887 716078
rect 672809 715730 672875 715733
rect 672809 715728 676292 715730
rect 672809 715672 672814 715728
rect 672870 715672 676292 715728
rect 672809 715670 676292 715672
rect 672809 715667 672875 715670
rect 40769 715322 40835 715325
rect 42425 715322 42491 715325
rect 40769 715320 42491 715322
rect 40769 715264 40774 715320
rect 40830 715264 42430 715320
rect 42486 715264 42491 715320
rect 40769 715262 42491 715264
rect 40769 715259 40835 715262
rect 42425 715259 42491 715262
rect 673361 715322 673427 715325
rect 673361 715320 676292 715322
rect 673361 715264 673366 715320
rect 673422 715264 676292 715320
rect 673361 715262 676292 715264
rect 673361 715259 673427 715262
rect 41137 714914 41203 714917
rect 42517 714914 42583 714917
rect 41137 714912 42583 714914
rect 41137 714856 41142 714912
rect 41198 714856 42522 714912
rect 42578 714856 42583 714912
rect 41137 714854 42583 714856
rect 41137 714851 41203 714854
rect 42517 714851 42583 714854
rect 673361 714914 673427 714917
rect 673361 714912 676292 714914
rect 673361 714856 673366 714912
rect 673422 714856 676292 714912
rect 673361 714854 676292 714856
rect 673361 714851 673427 714854
rect 42057 714644 42123 714645
rect 42006 714580 42012 714644
rect 42076 714642 42123 714644
rect 42076 714640 42168 714642
rect 42118 714584 42168 714640
rect 42076 714582 42168 714584
rect 42076 714580 42123 714582
rect 42057 714579 42123 714580
rect 673177 714506 673243 714509
rect 673177 714504 676292 714506
rect 673177 714448 673182 714504
rect 673238 714448 676292 714504
rect 673177 714446 676292 714448
rect 673177 714443 673243 714446
rect 39297 714234 39363 714237
rect 40350 714234 40356 714236
rect 39297 714232 40356 714234
rect 39297 714176 39302 714232
rect 39358 714176 40356 714232
rect 39297 714174 40356 714176
rect 39297 714171 39363 714174
rect 40350 714172 40356 714174
rect 40420 714172 40426 714236
rect 673821 714098 673887 714101
rect 673821 714096 676292 714098
rect 673821 714040 673826 714096
rect 673882 714040 676292 714096
rect 673821 714038 676292 714040
rect 673821 714035 673887 714038
rect 673821 713690 673887 713693
rect 673821 713688 676292 713690
rect 673821 713632 673826 713688
rect 673882 713632 676292 713688
rect 673821 713630 676292 713632
rect 673821 713627 673887 713630
rect 673821 713282 673887 713285
rect 673821 713280 676292 713282
rect 673821 713224 673826 713280
rect 673882 713224 676292 713280
rect 673821 713222 676292 713224
rect 673821 713219 673887 713222
rect 673821 712874 673887 712877
rect 673821 712872 676292 712874
rect 673821 712816 673826 712872
rect 673882 712816 676292 712872
rect 673821 712814 676292 712816
rect 673821 712811 673887 712814
rect 673821 712466 673887 712469
rect 673821 712464 676292 712466
rect 673821 712408 673826 712464
rect 673882 712408 676292 712464
rect 673821 712406 676292 712408
rect 673821 712403 673887 712406
rect 674414 711996 674420 712060
rect 674484 712058 674490 712060
rect 674484 711998 676292 712058
rect 674484 711996 674490 711998
rect 673821 711650 673887 711653
rect 673821 711648 676292 711650
rect 673821 711592 673826 711648
rect 673882 711592 676292 711648
rect 673821 711590 676292 711592
rect 673821 711587 673887 711590
rect 682377 711242 682443 711245
rect 682364 711240 682443 711242
rect 682364 711184 682382 711240
rect 682438 711184 682443 711240
rect 682364 711182 682443 711184
rect 682377 711179 682443 711182
rect 42149 710834 42215 710837
rect 43621 710834 43687 710837
rect 42149 710832 43687 710834
rect 42149 710776 42154 710832
rect 42210 710776 43626 710832
rect 43682 710776 43687 710832
rect 42149 710774 43687 710776
rect 42149 710771 42215 710774
rect 43621 710771 43687 710774
rect 675293 710834 675359 710837
rect 675293 710832 676292 710834
rect 675293 710776 675298 710832
rect 675354 710776 676292 710832
rect 675293 710774 676292 710776
rect 675293 710771 675359 710774
rect 678237 710426 678303 710429
rect 678237 710424 678316 710426
rect 678237 710368 678242 710424
rect 678298 710368 678316 710424
rect 678237 710366 678316 710368
rect 678237 710363 678303 710366
rect 673821 710018 673887 710021
rect 673821 710016 676292 710018
rect 673821 709960 673826 710016
rect 673882 709960 676292 710016
rect 673821 709958 676292 709960
rect 673821 709955 673887 709958
rect 40350 709820 40356 709884
rect 40420 709882 40426 709884
rect 41781 709882 41847 709885
rect 40420 709880 41847 709882
rect 40420 709824 41786 709880
rect 41842 709824 41847 709880
rect 40420 709822 41847 709824
rect 40420 709820 40426 709822
rect 41781 709819 41847 709822
rect 673821 709610 673887 709613
rect 673821 709608 676292 709610
rect 673821 709552 673826 709608
rect 673882 709552 676292 709608
rect 673821 709550 676292 709552
rect 673821 709547 673887 709550
rect 674598 709140 674604 709204
rect 674668 709202 674674 709204
rect 674668 709142 676292 709202
rect 674668 709140 674674 709142
rect 44633 708794 44699 708797
rect 683481 708794 683547 708797
rect 41830 708792 44699 708794
rect 41830 708736 44638 708792
rect 44694 708736 44699 708792
rect 41830 708734 44699 708736
rect 683468 708792 683547 708794
rect 683468 708736 683486 708792
rect 683542 708736 683547 708792
rect 683468 708734 683547 708736
rect 41830 708525 41890 708734
rect 44633 708731 44699 708734
rect 683481 708731 683547 708734
rect 41830 708520 41939 708525
rect 41830 708464 41878 708520
rect 41934 708464 41939 708520
rect 41830 708462 41939 708464
rect 41873 708459 41939 708462
rect 42057 708522 42123 708525
rect 44449 708522 44515 708525
rect 42057 708520 44515 708522
rect 42057 708464 42062 708520
rect 42118 708464 44454 708520
rect 44510 708464 44515 708520
rect 42057 708462 44515 708464
rect 42057 708459 42123 708462
rect 44449 708459 44515 708462
rect 684125 708386 684191 708389
rect 684125 708384 684204 708386
rect 684125 708328 684130 708384
rect 684186 708328 684204 708384
rect 684125 708326 684204 708328
rect 684125 708323 684191 708326
rect 683297 707978 683363 707981
rect 683284 707976 683363 707978
rect 683284 707920 683302 707976
rect 683358 707920 683363 707976
rect 683284 707918 683363 707920
rect 683297 707915 683363 707918
rect 42057 707842 42123 707845
rect 43621 707842 43687 707845
rect 42057 707840 43687 707842
rect 42057 707784 42062 707840
rect 42118 707784 43626 707840
rect 43682 707784 43687 707840
rect 42057 707782 43687 707784
rect 42057 707779 42123 707782
rect 43621 707779 43687 707782
rect 675886 707508 675892 707572
rect 675956 707570 675962 707572
rect 675956 707510 676292 707570
rect 675956 707508 675962 707510
rect 40718 707372 40724 707436
rect 40788 707434 40794 707436
rect 41781 707434 41847 707437
rect 40788 707432 41847 707434
rect 40788 707376 41786 707432
rect 41842 707376 41847 707432
rect 40788 707374 41847 707376
rect 40788 707372 40794 707374
rect 41781 707371 41847 707374
rect 676029 707162 676095 707165
rect 676029 707160 676292 707162
rect 676029 707104 676034 707160
rect 676090 707104 676292 707160
rect 676029 707102 676292 707104
rect 676029 707099 676095 707102
rect 672993 706754 673059 706757
rect 672993 706752 676292 706754
rect 672993 706696 672998 706752
rect 673054 706696 676292 706752
rect 672993 706694 676292 706696
rect 672993 706691 673059 706694
rect 42006 706420 42012 706484
rect 42076 706482 42082 706484
rect 42517 706482 42583 706485
rect 42076 706480 42583 706482
rect 42076 706424 42522 706480
rect 42578 706424 42583 706480
rect 42076 706422 42583 706424
rect 42076 706420 42082 706422
rect 42517 706419 42583 706422
rect 676029 706346 676095 706349
rect 676029 706344 676292 706346
rect 676029 706288 676034 706344
rect 676090 706288 676292 706344
rect 676029 706286 676292 706288
rect 676029 706283 676095 706286
rect 673361 705530 673427 705533
rect 674281 705530 674347 705533
rect 673361 705528 674347 705530
rect 673361 705472 673366 705528
rect 673422 705472 674286 705528
rect 674342 705472 674347 705528
rect 678470 705530 678530 705908
rect 683113 705530 683179 705533
rect 678470 705528 683179 705530
rect 678470 705500 683118 705528
rect 673361 705470 674347 705472
rect 678500 705472 683118 705500
rect 683174 705472 683179 705528
rect 678500 705470 683179 705472
rect 673361 705467 673427 705470
rect 674281 705467 674347 705470
rect 683113 705467 683179 705470
rect 673361 705258 673427 705261
rect 674465 705258 674531 705261
rect 673361 705256 674531 705258
rect 673361 705200 673366 705256
rect 673422 705200 674470 705256
rect 674526 705200 674531 705256
rect 673361 705198 674531 705200
rect 673361 705195 673427 705198
rect 674465 705195 674531 705198
rect 676029 705122 676095 705125
rect 676029 705120 676292 705122
rect 676029 705064 676034 705120
rect 676090 705064 676292 705120
rect 676029 705062 676292 705064
rect 676029 705059 676095 705062
rect 62113 704442 62179 704445
rect 62113 704440 64706 704442
rect 62113 704384 62118 704440
rect 62174 704384 64706 704440
rect 62113 704382 64706 704384
rect 62113 704379 62179 704382
rect 40534 704244 40540 704308
rect 40604 704306 40610 704308
rect 41781 704306 41847 704309
rect 40604 704304 41847 704306
rect 40604 704248 41786 704304
rect 41842 704248 41847 704304
rect 40604 704246 41847 704248
rect 40604 704244 40610 704246
rect 41781 704243 41847 704246
rect 64646 703860 64706 704382
rect 673177 703898 673243 703901
rect 674281 703898 674347 703901
rect 673177 703896 674347 703898
rect 673177 703840 673182 703896
rect 673238 703840 674286 703896
rect 674342 703840 674347 703896
rect 673177 703838 674347 703840
rect 673177 703835 673243 703838
rect 674281 703835 674347 703838
rect 41454 703564 41460 703628
rect 41524 703626 41530 703628
rect 42241 703626 42307 703629
rect 41524 703624 42307 703626
rect 41524 703568 42246 703624
rect 42302 703568 42307 703624
rect 41524 703566 42307 703568
rect 41524 703564 41530 703566
rect 42241 703563 42307 703566
rect 62113 703354 62179 703357
rect 62113 703352 64706 703354
rect 62113 703296 62118 703352
rect 62174 703296 64706 703352
rect 62113 703294 64706 703296
rect 62113 703291 62179 703294
rect 42057 703082 42123 703085
rect 42701 703082 42767 703085
rect 42057 703080 42767 703082
rect 42057 703024 42062 703080
rect 42118 703024 42706 703080
rect 42762 703024 42767 703080
rect 42057 703022 42767 703024
rect 42057 703019 42123 703022
rect 42701 703019 42767 703022
rect 64646 702678 64706 703294
rect 41965 702266 42031 702269
rect 42517 702266 42583 702269
rect 41965 702264 42583 702266
rect 41965 702208 41970 702264
rect 42026 702208 42522 702264
rect 42578 702208 42583 702264
rect 41965 702206 42583 702208
rect 41965 702203 42031 702206
rect 42517 702203 42583 702206
rect 41822 701796 41828 701860
rect 41892 701858 41898 701860
rect 42517 701858 42583 701861
rect 41892 701856 42583 701858
rect 41892 701800 42522 701856
rect 42578 701800 42583 701856
rect 41892 701798 42583 701800
rect 41892 701796 41898 701798
rect 42517 701795 42583 701798
rect 41638 701524 41644 701588
rect 41708 701586 41714 701588
rect 42517 701586 42583 701589
rect 41708 701584 42583 701586
rect 41708 701528 42522 701584
rect 42578 701528 42583 701584
rect 41708 701526 42583 701528
rect 41708 701524 41714 701526
rect 42517 701523 42583 701526
rect 62205 701314 62271 701317
rect 64646 701314 64706 701496
rect 675109 701450 675175 701453
rect 676806 701450 676812 701452
rect 675109 701448 676812 701450
rect 675109 701392 675114 701448
rect 675170 701392 676812 701448
rect 675109 701390 676812 701392
rect 675109 701387 675175 701390
rect 676806 701388 676812 701390
rect 676876 701388 676882 701452
rect 62205 701312 64706 701314
rect 62205 701256 62210 701312
rect 62266 701256 64706 701312
rect 62205 701254 64706 701256
rect 62205 701251 62271 701254
rect 673177 701178 673243 701181
rect 675109 701178 675175 701181
rect 673177 701176 675175 701178
rect 673177 701120 673182 701176
rect 673238 701120 675114 701176
rect 675170 701120 675175 701176
rect 673177 701118 675175 701120
rect 673177 701115 673243 701118
rect 675109 701115 675175 701118
rect 62757 700906 62823 700909
rect 672993 700906 673059 700909
rect 674925 700906 674991 700909
rect 62757 700904 64706 700906
rect 62757 700848 62762 700904
rect 62818 700848 64706 700904
rect 62757 700846 64706 700848
rect 62757 700843 62823 700846
rect 64646 700314 64706 700846
rect 672993 700904 674991 700906
rect 672993 700848 672998 700904
rect 673054 700848 674930 700904
rect 674986 700848 674991 700904
rect 672993 700846 674991 700848
rect 672993 700843 673059 700846
rect 674925 700843 674991 700846
rect 61377 699682 61443 699685
rect 61377 699680 64706 699682
rect 61377 699624 61382 699680
rect 61438 699624 64706 699680
rect 61377 699622 64706 699624
rect 61377 699619 61443 699622
rect 64646 699132 64706 699622
rect 62113 698186 62179 698189
rect 62113 698184 64706 698186
rect 62113 698128 62118 698184
rect 62174 698128 64706 698184
rect 62113 698126 64706 698128
rect 62113 698123 62179 698126
rect 64646 697950 64706 698126
rect 668393 696962 668459 696965
rect 675109 696962 675175 696965
rect 668393 696960 675175 696962
rect 668393 696904 668398 696960
rect 668454 696904 675114 696960
rect 675170 696904 675175 696960
rect 668393 696902 675175 696904
rect 668393 696899 668459 696902
rect 675109 696899 675175 696902
rect 675477 696828 675543 696829
rect 675477 696824 675524 696828
rect 675588 696826 675594 696828
rect 675477 696768 675482 696824
rect 675477 696764 675524 696768
rect 675588 696766 675634 696826
rect 675588 696764 675594 696766
rect 675477 696763 675543 696764
rect 670601 696146 670667 696149
rect 675109 696146 675175 696149
rect 670601 696144 675175 696146
rect 670601 696088 670606 696144
rect 670662 696088 675114 696144
rect 675170 696088 675175 696144
rect 670601 696086 675175 696088
rect 670601 696083 670667 696086
rect 675109 696083 675175 696086
rect 672993 695330 673059 695333
rect 672993 695328 675402 695330
rect 672993 695272 672998 695328
rect 673054 695272 675402 695328
rect 672993 695270 675402 695272
rect 672993 695267 673059 695270
rect 675342 695061 675402 695270
rect 672809 695058 672875 695061
rect 675109 695058 675175 695061
rect 672809 695056 675175 695058
rect 672809 695000 672814 695056
rect 672870 695000 675114 695056
rect 675170 695000 675175 695056
rect 672809 694998 675175 695000
rect 672809 694995 672875 694998
rect 675109 694995 675175 694998
rect 675293 695056 675402 695061
rect 675293 695000 675298 695056
rect 675354 695000 675402 695056
rect 675293 694998 675402 695000
rect 675293 694995 675359 694998
rect 673545 693290 673611 693293
rect 673862 693290 673868 693292
rect 673545 693288 673868 693290
rect 673545 693232 673550 693288
rect 673606 693232 673868 693288
rect 673545 693230 673868 693232
rect 673545 693227 673611 693230
rect 673862 693228 673868 693230
rect 673932 693228 673938 693292
rect 673545 693018 673611 693021
rect 675477 693018 675543 693021
rect 673545 693016 675543 693018
rect 673545 692960 673550 693016
rect 673606 692960 675482 693016
rect 675538 692960 675543 693016
rect 673545 692958 675543 692960
rect 673545 692955 673611 692958
rect 675477 692955 675543 692958
rect 674097 690434 674163 690437
rect 675293 690434 675359 690437
rect 674097 690432 675359 690434
rect 674097 690376 674102 690432
rect 674158 690376 675298 690432
rect 675354 690376 675359 690432
rect 674097 690374 675359 690376
rect 674097 690371 674163 690374
rect 675293 690371 675359 690374
rect 673177 690026 673243 690029
rect 674925 690026 674991 690029
rect 673177 690024 674991 690026
rect 649950 689482 650010 689980
rect 673177 689968 673182 690024
rect 673238 689968 674930 690024
rect 674986 689968 674991 690024
rect 673177 689966 674991 689968
rect 673177 689963 673243 689966
rect 674925 689963 674991 689966
rect 651465 689482 651531 689485
rect 649950 689480 651531 689482
rect 649950 689424 651470 689480
rect 651526 689424 651531 689480
rect 649950 689422 651531 689424
rect 651465 689419 651531 689422
rect 670969 689210 671035 689213
rect 675109 689210 675175 689213
rect 670969 689208 675175 689210
rect 670969 689152 670974 689208
rect 671030 689152 675114 689208
rect 675170 689152 675175 689208
rect 670969 689150 675175 689152
rect 670969 689147 671035 689150
rect 675109 689147 675175 689150
rect 649980 688802 650562 688828
rect 651649 688802 651715 688805
rect 649980 688800 651715 688802
rect 649980 688768 651654 688800
rect 650502 688744 651654 688768
rect 651710 688744 651715 688800
rect 650502 688742 651715 688744
rect 651649 688739 651715 688742
rect 673177 688802 673243 688805
rect 674649 688802 674715 688805
rect 673177 688800 674715 688802
rect 673177 688744 673182 688800
rect 673238 688744 674654 688800
rect 674710 688744 674715 688800
rect 673177 688742 674715 688744
rect 673177 688739 673243 688742
rect 674649 688739 674715 688742
rect 669405 688394 669471 688397
rect 675109 688394 675175 688397
rect 669405 688392 675175 688394
rect 669405 688336 669410 688392
rect 669466 688336 675114 688392
rect 675170 688336 675175 688392
rect 669405 688334 675175 688336
rect 669405 688331 669471 688334
rect 675109 688331 675175 688334
rect 42701 688122 42767 688125
rect 41492 688120 42767 688122
rect 41492 688064 42706 688120
rect 42762 688064 42767 688120
rect 41492 688062 42767 688064
rect 42701 688059 42767 688062
rect 673862 688060 673868 688124
rect 673932 688122 673938 688124
rect 674649 688122 674715 688125
rect 673932 688120 674715 688122
rect 673932 688064 674654 688120
rect 674710 688064 674715 688120
rect 673932 688062 674715 688064
rect 673932 688060 673938 688062
rect 674649 688059 674715 688062
rect 44817 687714 44883 687717
rect 41492 687712 44883 687714
rect 41492 687656 44822 687712
rect 44878 687656 44883 687712
rect 41492 687654 44883 687656
rect 44817 687651 44883 687654
rect 649950 687442 650010 687616
rect 651465 687442 651531 687445
rect 649950 687440 651531 687442
rect 649950 687384 651470 687440
rect 651526 687384 651531 687440
rect 649950 687382 651531 687384
rect 651465 687379 651531 687382
rect 43437 687306 43503 687309
rect 41492 687304 43503 687306
rect 41492 687248 43442 687304
rect 43498 687248 43503 687304
rect 41492 687246 43503 687248
rect 43437 687243 43503 687246
rect 40861 686898 40927 686901
rect 40861 686896 40940 686898
rect 40861 686840 40866 686896
rect 40922 686840 40940 686896
rect 40861 686838 40940 686840
rect 40861 686835 40927 686838
rect 651465 686762 651531 686765
rect 649950 686760 651531 686762
rect 649950 686704 651470 686760
rect 651526 686704 651531 686760
rect 649950 686702 651531 686704
rect 41137 686490 41203 686493
rect 41124 686488 41203 686490
rect 41124 686432 41142 686488
rect 41198 686432 41203 686488
rect 649950 686434 650010 686702
rect 651465 686699 651531 686702
rect 41124 686430 41203 686432
rect 41137 686427 41203 686430
rect 43069 686082 43135 686085
rect 41492 686080 43135 686082
rect 41492 686024 43074 686080
rect 43130 686024 43135 686080
rect 41492 686022 43135 686024
rect 43069 686019 43135 686022
rect 41045 685912 41111 685915
rect 41045 685910 41154 685912
rect 41045 685854 41050 685910
rect 41106 685854 41154 685910
rect 41045 685849 41154 685854
rect 41094 685644 41154 685849
rect 673637 685810 673703 685813
rect 675293 685810 675359 685813
rect 673637 685808 675359 685810
rect 673637 685752 673642 685808
rect 673698 685752 675298 685808
rect 675354 685752 675359 685808
rect 673637 685750 675359 685752
rect 673637 685747 673703 685750
rect 675293 685747 675359 685750
rect 44265 685266 44331 685269
rect 651465 685266 651531 685269
rect 41492 685264 44331 685266
rect 41492 685208 44270 685264
rect 44326 685208 44331 685264
rect 41492 685206 44331 685208
rect 649950 685264 651531 685266
rect 649950 685208 651470 685264
rect 651526 685208 651531 685264
rect 649950 685206 651531 685208
rect 44265 685203 44331 685206
rect 651465 685203 651531 685206
rect 672717 684994 672783 684997
rect 675477 684994 675543 684997
rect 672717 684992 675543 684994
rect 672717 684936 672722 684992
rect 672778 684936 675482 684992
rect 675538 684936 675543 684992
rect 672717 684934 675543 684936
rect 672717 684931 672783 684934
rect 675477 684931 675543 684934
rect 44633 684858 44699 684861
rect 41492 684856 44699 684858
rect 41492 684800 44638 684856
rect 44694 684800 44699 684856
rect 41492 684798 44699 684800
rect 44633 684795 44699 684798
rect 45001 684450 45067 684453
rect 652569 684450 652635 684453
rect 41492 684448 45067 684450
rect 41492 684392 45006 684448
rect 45062 684392 45067 684448
rect 41492 684390 45067 684392
rect 45001 684387 45067 684390
rect 649950 684448 652635 684450
rect 649950 684392 652574 684448
rect 652630 684392 652635 684448
rect 649950 684390 652635 684392
rect 649950 684070 650010 684390
rect 652569 684387 652635 684390
rect 44449 684042 44515 684045
rect 41492 684040 44515 684042
rect 41492 683984 44454 684040
rect 44510 683984 44515 684040
rect 41492 683982 44515 683984
rect 44449 683979 44515 683982
rect 42006 683634 42012 683636
rect 41492 683574 42012 683634
rect 42006 683572 42012 683574
rect 42076 683572 42082 683636
rect 41321 683464 41387 683467
rect 41278 683462 41387 683464
rect 41278 683406 41326 683462
rect 41382 683406 41387 683462
rect 41278 683401 41387 683406
rect 41278 683196 41338 683401
rect 42190 682818 42196 682820
rect 41492 682758 42196 682818
rect 42190 682756 42196 682758
rect 42260 682756 42266 682820
rect 42701 682410 42767 682413
rect 41492 682408 42767 682410
rect 41492 682352 42706 682408
rect 42762 682352 42767 682408
rect 41492 682350 42767 682352
rect 42701 682347 42767 682350
rect 674230 682348 674236 682412
rect 674300 682410 674306 682412
rect 683389 682410 683455 682413
rect 674300 682408 683455 682410
rect 674300 682352 683394 682408
rect 683450 682352 683455 682408
rect 674300 682350 683455 682352
rect 674300 682348 674306 682350
rect 683389 682347 683455 682350
rect 35157 682002 35223 682005
rect 35157 682000 35236 682002
rect 35157 681944 35162 682000
rect 35218 681944 35236 682000
rect 35157 681942 35236 681944
rect 35157 681939 35223 681942
rect 31661 681594 31727 681597
rect 31661 681592 31740 681594
rect 31661 681536 31666 681592
rect 31722 681536 31740 681592
rect 31661 681534 31740 681536
rect 31661 681531 31727 681534
rect 675518 681396 675524 681460
rect 675588 681458 675594 681460
rect 675753 681458 675819 681461
rect 675588 681456 675819 681458
rect 675588 681400 675758 681456
rect 675814 681400 675819 681456
rect 675588 681398 675819 681400
rect 675588 681396 675594 681398
rect 675753 681395 675819 681398
rect 32446 681019 32506 681156
rect 41689 681050 41755 681053
rect 44265 681050 44331 681053
rect 675385 681052 675451 681053
rect 41689 681048 44331 681050
rect 32397 681014 32506 681019
rect 33777 681016 33843 681019
rect 32397 680958 32402 681014
rect 32458 680958 32506 681014
rect 32397 680956 32506 680958
rect 33734 681014 33843 681016
rect 33734 680958 33782 681014
rect 33838 680958 33843 681014
rect 41689 680992 41694 681048
rect 41750 680992 44270 681048
rect 44326 680992 44331 681048
rect 41689 680990 44331 680992
rect 41689 680987 41755 680990
rect 44265 680987 44331 680990
rect 675334 680988 675340 681052
rect 675404 681050 675451 681052
rect 675404 681048 675496 681050
rect 675446 680992 675496 681048
rect 675404 680990 675496 680992
rect 675404 680988 675451 680990
rect 675385 680987 675451 680988
rect 32397 680953 32463 680956
rect 33734 680953 33843 680958
rect 33734 680748 33794 680953
rect 43069 680370 43135 680373
rect 41492 680368 43135 680370
rect 41492 680312 43074 680368
rect 43130 680312 43135 680368
rect 41492 680310 43135 680312
rect 43069 680307 43135 680310
rect 45001 679962 45067 679965
rect 41492 679960 45067 679962
rect 41492 679904 45006 679960
rect 45062 679904 45067 679960
rect 41492 679902 45067 679904
rect 45001 679899 45067 679902
rect 43621 679554 43687 679557
rect 41492 679552 43687 679554
rect 41492 679496 43626 679552
rect 43682 679496 43687 679552
rect 41492 679494 43687 679496
rect 43621 679491 43687 679494
rect 40542 678992 40602 679116
rect 40534 678928 40540 678992
rect 40604 678928 40610 678992
rect 40718 678928 40724 678992
rect 40788 678928 40794 678992
rect 40726 678708 40786 678928
rect 41822 678330 41828 678332
rect 41492 678270 41828 678330
rect 41822 678268 41828 678270
rect 41892 678268 41898 678332
rect 43989 677922 44055 677925
rect 41492 677920 44055 677922
rect 41492 677864 43994 677920
rect 44050 677864 44055 677920
rect 41492 677862 44055 677864
rect 43989 677859 44055 677862
rect 41094 677109 41154 677484
rect 41094 677104 41203 677109
rect 41094 677076 41142 677104
rect 41124 677048 41142 677076
rect 41198 677048 41203 677104
rect 41124 677046 41203 677048
rect 41137 677043 41203 677046
rect 43437 676698 43503 676701
rect 41492 676696 43503 676698
rect 41492 676640 43442 676696
rect 43498 676640 43503 676696
rect 41492 676638 43503 676640
rect 43437 676635 43503 676638
rect 674833 676426 674899 676429
rect 675150 676426 675156 676428
rect 674833 676424 675156 676426
rect 674833 676368 674838 676424
rect 674894 676368 675156 676424
rect 674833 676366 675156 676368
rect 674833 676363 674899 676366
rect 675150 676364 675156 676366
rect 675220 676364 675226 676428
rect 675753 676426 675819 676429
rect 676070 676426 676076 676428
rect 675753 676424 676076 676426
rect 675753 676368 675758 676424
rect 675814 676368 676076 676424
rect 675753 676366 676076 676368
rect 675753 676363 675819 676366
rect 676070 676364 676076 676366
rect 676140 676364 676146 676428
rect 673729 674386 673795 674389
rect 674649 674386 674715 674389
rect 673729 674384 674715 674386
rect 673729 674328 673734 674384
rect 673790 674328 674654 674384
rect 674710 674328 674715 674384
rect 673729 674326 674715 674328
rect 673729 674323 673795 674326
rect 674649 674323 674715 674326
rect 32397 672754 32463 672757
rect 41822 672754 41828 672756
rect 32397 672752 41828 672754
rect 32397 672696 32402 672752
rect 32458 672696 41828 672752
rect 32397 672694 41828 672696
rect 32397 672691 32463 672694
rect 41822 672692 41828 672694
rect 41892 672692 41898 672756
rect 42006 671604 42012 671668
rect 42076 671666 42082 671668
rect 42333 671666 42399 671669
rect 42076 671664 42399 671666
rect 42076 671608 42338 671664
rect 42394 671608 42399 671664
rect 42076 671606 42399 671608
rect 42076 671604 42082 671606
rect 42333 671603 42399 671606
rect 673729 671394 673795 671397
rect 673729 671392 676292 671394
rect 673729 671336 673734 671392
rect 673790 671336 676292 671392
rect 673729 671334 676292 671336
rect 673729 671331 673795 671334
rect 673729 670986 673795 670989
rect 673729 670984 676292 670986
rect 673729 670928 673734 670984
rect 673790 670928 676292 670984
rect 673729 670926 676292 670928
rect 673729 670923 673795 670926
rect 673545 670578 673611 670581
rect 673545 670576 676292 670578
rect 673545 670520 673550 670576
rect 673606 670520 676292 670576
rect 673545 670518 676292 670520
rect 673545 670515 673611 670518
rect 672165 670170 672231 670173
rect 672165 670168 676292 670170
rect 672165 670112 672170 670168
rect 672226 670112 676292 670168
rect 672165 670110 676292 670112
rect 672165 670107 672231 670110
rect 672165 669762 672231 669765
rect 672165 669760 676292 669762
rect 672165 669704 672170 669760
rect 672226 669704 676292 669760
rect 672165 669702 676292 669704
rect 672165 669699 672231 669702
rect 673545 669218 673611 669221
rect 676262 669218 676322 669330
rect 673545 669216 676322 669218
rect 673545 669160 673550 669216
rect 673606 669160 676322 669216
rect 673545 669158 676322 669160
rect 673545 669155 673611 669158
rect 673545 668946 673611 668949
rect 673545 668944 676292 668946
rect 673545 668888 673550 668944
rect 673606 668888 676292 668944
rect 673545 668886 676292 668888
rect 673545 668883 673611 668886
rect 42057 668540 42123 668541
rect 42006 668476 42012 668540
rect 42076 668538 42123 668540
rect 673545 668538 673611 668541
rect 42076 668536 42168 668538
rect 42118 668480 42168 668536
rect 42076 668478 42168 668480
rect 673545 668536 676292 668538
rect 673545 668480 673550 668536
rect 673606 668480 676292 668536
rect 673545 668478 676292 668480
rect 42076 668476 42123 668478
rect 42057 668475 42123 668476
rect 673545 668475 673611 668478
rect 673545 668130 673611 668133
rect 673545 668128 676292 668130
rect 673545 668072 673550 668128
rect 673606 668072 676292 668128
rect 673545 668070 676292 668072
rect 673545 668067 673611 668070
rect 673545 667722 673611 667725
rect 673545 667720 676292 667722
rect 673545 667664 673550 667720
rect 673606 667664 676292 667720
rect 673545 667662 676292 667664
rect 673545 667659 673611 667662
rect 676262 667042 676322 667284
rect 673548 666982 676322 667042
rect 673548 666773 673608 666982
rect 673545 666768 673611 666773
rect 673545 666712 673550 666768
rect 673606 666712 673611 666768
rect 673545 666707 673611 666712
rect 676029 666770 676095 666773
rect 676262 666770 676322 666876
rect 676029 666768 676322 666770
rect 676029 666712 676034 666768
rect 676090 666712 676322 666768
rect 676029 666710 676322 666712
rect 676029 666707 676095 666710
rect 42057 666634 42123 666637
rect 45001 666634 45067 666637
rect 42057 666632 45067 666634
rect 42057 666576 42062 666632
rect 42118 666576 45006 666632
rect 45062 666576 45067 666632
rect 42057 666574 45067 666576
rect 42057 666571 42123 666574
rect 45001 666571 45067 666574
rect 676806 666572 676812 666636
rect 676876 666572 676882 666636
rect 676814 666468 676874 666572
rect 673545 666090 673611 666093
rect 673545 666088 676292 666090
rect 673545 666032 673550 666088
rect 673606 666032 676292 666088
rect 673545 666030 676292 666032
rect 673545 666027 673611 666030
rect 672533 665546 672599 665549
rect 676262 665546 676322 665652
rect 672533 665544 676322 665546
rect 672533 665488 672538 665544
rect 672594 665488 676322 665544
rect 672533 665486 676322 665488
rect 672533 665483 672599 665486
rect 673545 665274 673611 665277
rect 673545 665272 676292 665274
rect 673545 665216 673550 665272
rect 673606 665216 676292 665272
rect 673545 665214 676292 665216
rect 673545 665211 673611 665214
rect 40902 665076 40908 665140
rect 40972 665138 40978 665140
rect 41781 665138 41847 665141
rect 40972 665136 41847 665138
rect 40972 665080 41786 665136
rect 41842 665080 41847 665136
rect 40972 665078 41847 665080
rect 40972 665076 40978 665078
rect 41781 665075 41847 665078
rect 673545 664866 673611 664869
rect 673545 664864 676292 664866
rect 673545 664808 673550 664864
rect 673606 664808 676292 664864
rect 673545 664806 676292 664808
rect 673545 664803 673611 664806
rect 672349 664186 672415 664189
rect 676262 664186 676322 664428
rect 672349 664184 676322 664186
rect 672349 664128 672354 664184
rect 672410 664128 676322 664184
rect 672349 664126 676322 664128
rect 672349 664123 672415 664126
rect 40718 663988 40724 664052
rect 40788 664050 40794 664052
rect 41781 664050 41847 664053
rect 40788 664048 41847 664050
rect 40788 663992 41786 664048
rect 41842 663992 41847 664048
rect 40788 663990 41847 663992
rect 40788 663988 40794 663990
rect 41781 663987 41847 663990
rect 676262 663781 676322 664020
rect 676213 663776 676322 663781
rect 676213 663720 676218 663776
rect 676274 663720 676322 663776
rect 676213 663718 676322 663720
rect 683205 663778 683271 663781
rect 683205 663776 683314 663778
rect 683205 663720 683210 663776
rect 683266 663720 683314 663776
rect 676213 663715 676279 663718
rect 683205 663715 683314 663720
rect 673545 663642 673611 663645
rect 674833 663642 674899 663645
rect 673545 663640 674899 663642
rect 673545 663584 673550 663640
rect 673606 663584 674838 663640
rect 674894 663584 674899 663640
rect 683254 663612 683314 663715
rect 673545 663582 674899 663584
rect 673545 663579 673611 663582
rect 674833 663579 674899 663582
rect 674606 663174 676292 663234
rect 673913 663098 673979 663101
rect 674606 663098 674666 663174
rect 673913 663096 674666 663098
rect 673913 663040 673918 663096
rect 673974 663040 674666 663096
rect 673913 663038 674666 663040
rect 673913 663035 673979 663038
rect 676213 662962 676279 662965
rect 676213 662960 676322 662962
rect 676213 662904 676218 662960
rect 676274 662904 676322 662960
rect 676213 662899 676322 662904
rect 40534 662764 40540 662828
rect 40604 662826 40610 662828
rect 42241 662826 42307 662829
rect 40604 662824 42307 662826
rect 40604 662768 42246 662824
rect 42302 662768 42307 662824
rect 676262 662796 676322 662899
rect 40604 662766 42307 662768
rect 40604 662764 40610 662766
rect 42241 662763 42307 662766
rect 683389 662554 683455 662557
rect 683389 662552 683498 662554
rect 683389 662496 683394 662552
rect 683450 662496 683498 662552
rect 683389 662491 683498 662496
rect 683438 662388 683498 662491
rect 673545 662010 673611 662013
rect 673545 662008 676292 662010
rect 673545 661952 673550 662008
rect 673606 661952 676292 662008
rect 673545 661950 676292 661952
rect 673545 661947 673611 661950
rect 673913 661602 673979 661605
rect 673913 661600 676292 661602
rect 673913 661544 673918 661600
rect 673974 661544 676292 661600
rect 673913 661542 676292 661544
rect 673913 661539 673979 661542
rect 673913 661194 673979 661197
rect 673913 661192 676292 661194
rect 673913 661136 673918 661192
rect 673974 661136 676292 661192
rect 673913 661134 676292 661136
rect 673913 661131 673979 661134
rect 62113 660922 62179 660925
rect 62113 660920 64706 660922
rect 62113 660864 62118 660920
rect 62174 660864 64706 660920
rect 62113 660862 64706 660864
rect 62113 660859 62179 660862
rect 64646 660638 64706 660862
rect 683070 660109 683130 660756
rect 673913 660106 673979 660109
rect 674649 660106 674715 660109
rect 673913 660104 674715 660106
rect 673913 660048 673918 660104
rect 673974 660048 674654 660104
rect 674710 660048 674715 660104
rect 673913 660046 674715 660048
rect 683070 660104 683179 660109
rect 683070 660048 683118 660104
rect 683174 660048 683179 660104
rect 683070 660046 683179 660048
rect 673913 660043 673979 660046
rect 674649 660043 674715 660046
rect 683113 660043 683179 660046
rect 672809 659698 672875 659701
rect 676262 659698 676322 659940
rect 672809 659696 676322 659698
rect 672809 659640 672814 659696
rect 672870 659640 676322 659696
rect 672809 659638 676322 659640
rect 672809 659635 672875 659638
rect 62113 659562 62179 659565
rect 62113 659560 64706 659562
rect 62113 659504 62118 659560
rect 62174 659504 64706 659560
rect 62113 659502 64706 659504
rect 62113 659499 62179 659502
rect 64646 659456 64706 659502
rect 41638 658548 41644 658612
rect 41708 658610 41714 658612
rect 42517 658610 42583 658613
rect 41708 658608 42583 658610
rect 41708 658552 42522 658608
rect 42578 658552 42583 658608
rect 41708 658550 42583 658552
rect 41708 658548 41714 658550
rect 42517 658547 42583 658550
rect 41781 658340 41847 658341
rect 41781 658336 41828 658340
rect 41892 658338 41898 658340
rect 62113 658338 62179 658341
rect 41781 658280 41786 658336
rect 41781 658276 41828 658280
rect 41892 658278 41938 658338
rect 62113 658336 64706 658338
rect 62113 658280 62118 658336
rect 62174 658280 64706 658336
rect 62113 658278 64706 658280
rect 41892 658276 41898 658278
rect 41781 658275 41847 658276
rect 62113 658275 62179 658278
rect 64646 658274 64706 658278
rect 62757 657658 62823 657661
rect 62757 657656 64706 657658
rect 62757 657600 62762 657656
rect 62818 657600 64706 657656
rect 62757 657598 64706 657600
rect 62757 657595 62823 657598
rect 41454 657188 41460 657252
rect 41524 657250 41530 657252
rect 41781 657250 41847 657253
rect 41524 657248 41847 657250
rect 41524 657192 41786 657248
rect 41842 657192 41847 657248
rect 41524 657190 41847 657192
rect 41524 657188 41530 657190
rect 41781 657187 41847 657190
rect 64646 657092 64706 657598
rect 61377 656570 61443 656573
rect 61377 656568 64706 656570
rect 61377 656512 61382 656568
rect 61438 656512 64706 656568
rect 61377 656510 64706 656512
rect 61377 656507 61443 656510
rect 64646 655910 64706 656510
rect 673913 655618 673979 655621
rect 675109 655618 675175 655621
rect 673913 655616 675175 655618
rect 673913 655560 673918 655616
rect 673974 655560 675114 655616
rect 675170 655560 675175 655616
rect 673913 655558 675175 655560
rect 673913 655555 673979 655558
rect 675109 655555 675175 655558
rect 62113 655346 62179 655349
rect 62113 655344 64706 655346
rect 62113 655288 62118 655344
rect 62174 655288 64706 655344
rect 62113 655286 64706 655288
rect 62113 655283 62179 655286
rect 64646 654728 64706 655286
rect 674414 652836 674420 652900
rect 674484 652898 674490 652900
rect 675385 652898 675451 652901
rect 674484 652896 675451 652898
rect 674484 652840 675390 652896
rect 675446 652840 675451 652896
rect 674484 652838 675451 652840
rect 674484 652836 674490 652838
rect 675385 652835 675451 652838
rect 671981 652490 672047 652493
rect 675109 652490 675175 652493
rect 671981 652488 675175 652490
rect 671981 652432 671986 652488
rect 672042 652432 675114 652488
rect 675170 652432 675175 652488
rect 671981 652430 675175 652432
rect 671981 652427 672047 652430
rect 675109 652427 675175 652430
rect 675201 650180 675267 650181
rect 675150 650178 675156 650180
rect 675110 650118 675156 650178
rect 675220 650176 675267 650180
rect 675262 650120 675267 650176
rect 675150 650116 675156 650118
rect 675220 650116 675267 650120
rect 675201 650115 675267 650116
rect 671797 649770 671863 649773
rect 675385 649770 675451 649773
rect 671797 649768 675451 649770
rect 671797 649712 671802 649768
rect 671858 649712 675390 649768
rect 675446 649712 675451 649768
rect 671797 649710 675451 649712
rect 671797 649707 671863 649710
rect 675385 649707 675451 649710
rect 672533 649226 672599 649229
rect 675385 649226 675451 649229
rect 672533 649224 675451 649226
rect 672533 649168 672538 649224
rect 672594 649168 675390 649224
rect 675446 649168 675451 649224
rect 672533 649166 675451 649168
rect 672533 649163 672599 649166
rect 675385 649163 675451 649166
rect 675753 648682 675819 648685
rect 677174 648682 677180 648684
rect 675753 648680 677180 648682
rect 675753 648624 675758 648680
rect 675814 648624 677180 648680
rect 675753 648622 677180 648624
rect 675753 648619 675819 648622
rect 677174 648620 677180 648622
rect 677244 648620 677250 648684
rect 671613 647866 671679 647869
rect 675385 647866 675451 647869
rect 671613 647864 675451 647866
rect 671613 647808 671618 647864
rect 671674 647808 675390 647864
rect 675446 647808 675451 647864
rect 671613 647806 675451 647808
rect 671613 647803 671679 647806
rect 675385 647803 675451 647806
rect 674005 647322 674071 647325
rect 675201 647322 675267 647325
rect 674005 647320 675267 647322
rect 674005 647264 674010 647320
rect 674066 647264 675206 647320
rect 675262 647264 675267 647320
rect 674005 647262 675267 647264
rect 674005 647259 674071 647262
rect 675201 647259 675267 647262
rect 674005 645554 674071 645557
rect 675201 645554 675267 645557
rect 674005 645552 675267 645554
rect 674005 645496 674010 645552
rect 674066 645496 675206 645552
rect 675262 645496 675267 645552
rect 674005 645494 675267 645496
rect 674005 645491 674071 645494
rect 675201 645491 675267 645494
rect 35758 644741 35818 644912
rect 673545 644874 673611 644877
rect 675385 644874 675451 644877
rect 673545 644872 675451 644874
rect 673545 644816 673550 644872
rect 673606 644816 675390 644872
rect 675446 644816 675451 644872
rect 673545 644814 675451 644816
rect 673545 644811 673611 644814
rect 675385 644811 675451 644814
rect 35758 644736 35867 644741
rect 35758 644680 35806 644736
rect 35862 644680 35867 644736
rect 35758 644678 35867 644680
rect 35801 644675 35867 644678
rect 39481 644738 39547 644741
rect 44265 644738 44331 644741
rect 39481 644736 44331 644738
rect 39481 644680 39486 644736
rect 39542 644680 44270 644736
rect 44326 644680 44331 644736
rect 39481 644678 44331 644680
rect 39481 644675 39547 644678
rect 44265 644675 44331 644678
rect 675753 644738 675819 644741
rect 676806 644738 676812 644740
rect 675753 644736 676812 644738
rect 675753 644680 675758 644736
rect 675814 644680 676812 644736
rect 675753 644678 676812 644680
rect 675753 644675 675819 644678
rect 676806 644676 676812 644678
rect 676876 644676 676882 644740
rect 38518 644333 38578 644504
rect 38518 644328 38627 644333
rect 38518 644272 38566 644328
rect 38622 644272 38627 644328
rect 38518 644270 38627 644272
rect 38561 644267 38627 644270
rect 35390 643925 35450 644096
rect 35341 643920 35450 643925
rect 35341 643864 35346 643920
rect 35402 643864 35450 643920
rect 35341 643862 35450 643864
rect 35341 643859 35407 643862
rect 35574 643517 35634 643688
rect 674741 643650 674807 643653
rect 675385 643650 675451 643653
rect 674741 643648 675451 643650
rect 674741 643592 674746 643648
rect 674802 643592 675390 643648
rect 675446 643592 675451 643648
rect 674741 643590 675451 643592
rect 674741 643587 674807 643590
rect 675385 643587 675451 643590
rect 35525 643512 35634 643517
rect 35801 643514 35867 643517
rect 35525 643456 35530 643512
rect 35586 643456 35634 643512
rect 35525 643454 35634 643456
rect 35758 643512 35867 643514
rect 35758 643456 35806 643512
rect 35862 643456 35867 643512
rect 35525 643451 35591 643454
rect 35758 643451 35867 643456
rect 40493 643514 40559 643517
rect 45001 643514 45067 643517
rect 40493 643512 45067 643514
rect 40493 643456 40498 643512
rect 40554 643456 45006 643512
rect 45062 643456 45067 643512
rect 40493 643454 45067 643456
rect 40493 643451 40559 643454
rect 45001 643451 45067 643454
rect 35758 643280 35818 643451
rect 649950 643242 650010 643558
rect 651465 643242 651531 643245
rect 649950 643240 651531 643242
rect 649950 643184 651470 643240
rect 651526 643184 651531 643240
rect 649950 643182 651531 643184
rect 651465 643179 651531 643182
rect 674005 643106 674071 643109
rect 675293 643106 675359 643109
rect 674005 643104 675359 643106
rect 674005 643048 674010 643104
rect 674066 643048 675298 643104
rect 675354 643048 675359 643104
rect 674005 643046 675359 643048
rect 674005 643043 674071 643046
rect 675293 643043 675359 643046
rect 35574 642701 35634 642872
rect 35574 642696 35683 642701
rect 35574 642640 35622 642696
rect 35678 642640 35683 642696
rect 35574 642638 35683 642640
rect 35617 642635 35683 642638
rect 35801 642290 35867 642293
rect 35758 642288 35867 642290
rect 35758 642232 35806 642288
rect 35862 642232 35867 642288
rect 35758 642227 35867 642232
rect 41462 642290 41522 642464
rect 44214 642290 44220 642292
rect 41462 642230 44220 642290
rect 44214 642228 44220 642230
rect 44284 642228 44290 642292
rect 35758 642056 35818 642227
rect 649950 641882 650010 642376
rect 652017 641882 652083 641885
rect 649950 641880 652083 641882
rect 649950 641824 652022 641880
rect 652078 641824 652083 641880
rect 649950 641822 652083 641824
rect 652017 641819 652083 641822
rect 673913 641746 673979 641749
rect 675293 641746 675359 641749
rect 673913 641744 675359 641746
rect 673913 641688 673918 641744
rect 673974 641688 675298 641744
rect 675354 641688 675359 641744
rect 673913 641686 675359 641688
rect 673913 641683 673979 641686
rect 675293 641683 675359 641686
rect 35574 641477 35634 641648
rect 35574 641472 35683 641477
rect 35574 641416 35622 641472
rect 35678 641416 35683 641472
rect 35574 641414 35683 641416
rect 35617 641411 35683 641414
rect 35758 641069 35818 641240
rect 35758 641064 35867 641069
rect 35758 641008 35806 641064
rect 35862 641008 35867 641064
rect 35758 641006 35867 641008
rect 35801 641003 35867 641006
rect 39573 641066 39639 641069
rect 44449 641066 44515 641069
rect 39573 641064 44515 641066
rect 39573 641008 39578 641064
rect 39634 641008 44454 641064
rect 44510 641008 44515 641064
rect 39573 641006 44515 641008
rect 39573 641003 39639 641006
rect 44449 641003 44515 641006
rect 35758 640661 35818 640832
rect 649950 640794 650010 641194
rect 651465 640794 651531 640797
rect 649950 640792 651531 640794
rect 649950 640736 651470 640792
rect 651526 640736 651531 640792
rect 649950 640734 651531 640736
rect 651465 640731 651531 640734
rect 35758 640656 35867 640661
rect 35758 640600 35806 640656
rect 35862 640600 35867 640656
rect 35758 640598 35867 640600
rect 35801 640595 35867 640598
rect 41454 640596 41460 640660
rect 41524 640596 41530 640660
rect 41462 640424 41522 640596
rect 39941 640250 40007 640253
rect 45185 640250 45251 640253
rect 39941 640248 45251 640250
rect 39941 640192 39946 640248
rect 40002 640192 45190 640248
rect 45246 640192 45251 640248
rect 39941 640190 45251 640192
rect 39941 640187 40007 640190
rect 45185 640187 45251 640190
rect 651373 640114 651439 640117
rect 649950 640112 651439 640114
rect 649950 640056 651378 640112
rect 651434 640056 651439 640112
rect 649950 640054 651439 640056
rect 35390 639845 35450 640016
rect 649950 640012 650010 640054
rect 651373 640051 651439 640054
rect 35341 639840 35450 639845
rect 35341 639784 35346 639840
rect 35402 639784 35450 639840
rect 35341 639782 35450 639784
rect 667657 639842 667723 639845
rect 675477 639842 675543 639845
rect 667657 639840 675543 639842
rect 667657 639784 667662 639840
rect 667718 639784 675482 639840
rect 675538 639784 675543 639840
rect 667657 639782 675543 639784
rect 35341 639779 35407 639782
rect 667657 639779 667723 639782
rect 675477 639779 675543 639782
rect 35574 639437 35634 639608
rect 35525 639432 35634 639437
rect 35801 639434 35867 639437
rect 35525 639376 35530 639432
rect 35586 639376 35634 639432
rect 35525 639374 35634 639376
rect 35758 639432 35867 639434
rect 35758 639376 35806 639432
rect 35862 639376 35867 639432
rect 35525 639371 35591 639374
rect 35758 639371 35867 639376
rect 35758 639200 35818 639371
rect 35574 638621 35634 638792
rect 35574 638616 35683 638621
rect 35574 638560 35622 638616
rect 35678 638560 35683 638616
rect 35574 638558 35683 638560
rect 649766 638618 649826 638830
rect 670417 638754 670483 638757
rect 675477 638754 675543 638757
rect 670417 638752 675543 638754
rect 670417 638696 670422 638752
rect 670478 638696 675482 638752
rect 675538 638696 675543 638752
rect 670417 638694 675543 638696
rect 670417 638691 670483 638694
rect 675477 638691 675543 638694
rect 651465 638618 651531 638621
rect 649766 638616 651531 638618
rect 649766 638560 651470 638616
rect 651526 638560 651531 638616
rect 649766 638558 651531 638560
rect 35617 638555 35683 638558
rect 651465 638555 651531 638558
rect 35758 638213 35818 638384
rect 35758 638208 35867 638213
rect 651649 638210 651715 638213
rect 35758 638152 35806 638208
rect 35862 638152 35867 638208
rect 35758 638150 35867 638152
rect 35801 638147 35867 638150
rect 649950 638208 651715 638210
rect 649950 638152 651654 638208
rect 651710 638152 651715 638208
rect 649950 638150 651715 638152
rect 32446 637805 32506 637976
rect 32397 637800 32506 637805
rect 32397 637744 32402 637800
rect 32458 637744 32506 637800
rect 32397 637742 32506 637744
rect 32397 637739 32463 637742
rect 649950 637648 650010 638150
rect 651649 638147 651715 638150
rect 35206 637397 35266 637568
rect 35157 637392 35266 637397
rect 35157 637336 35162 637392
rect 35218 637336 35266 637392
rect 35157 637334 35266 637336
rect 35157 637331 35223 637334
rect 35574 636989 35634 637160
rect 35574 636984 35683 636989
rect 35574 636928 35622 636984
rect 35678 636928 35683 636984
rect 35574 636926 35683 636928
rect 35617 636923 35683 636926
rect 35801 636578 35867 636581
rect 40910 636580 40970 636752
rect 35758 636576 35867 636578
rect 35758 636520 35806 636576
rect 35862 636520 35867 636576
rect 35758 636515 35867 636520
rect 40902 636516 40908 636580
rect 40972 636516 40978 636580
rect 35758 636344 35818 636515
rect 39021 636170 39087 636173
rect 44633 636170 44699 636173
rect 39021 636168 44699 636170
rect 39021 636112 39026 636168
rect 39082 636112 44638 636168
rect 44694 636112 44699 636168
rect 39021 636110 44699 636112
rect 39021 636107 39087 636110
rect 44633 636107 44699 636110
rect 676070 636108 676076 636172
rect 676140 636170 676146 636172
rect 682377 636170 682443 636173
rect 676140 636168 682443 636170
rect 676140 636112 682382 636168
rect 682438 636112 682443 636168
rect 676140 636110 682443 636112
rect 676140 636108 676146 636110
rect 682377 636107 682443 636110
rect 35758 635765 35818 635936
rect 35758 635760 35867 635765
rect 35758 635704 35806 635760
rect 35862 635704 35867 635760
rect 35758 635702 35867 635704
rect 35801 635699 35867 635702
rect 39849 635762 39915 635765
rect 43069 635762 43135 635765
rect 39849 635760 43135 635762
rect 39849 635704 39854 635760
rect 39910 635704 43074 635760
rect 43130 635704 43135 635760
rect 39849 635702 43135 635704
rect 39849 635699 39915 635702
rect 43069 635699 43135 635702
rect 40542 635356 40602 635528
rect 673729 635490 673795 635493
rect 674281 635490 674347 635493
rect 673729 635488 674347 635490
rect 673729 635432 673734 635488
rect 673790 635432 674286 635488
rect 674342 635432 674347 635488
rect 673729 635430 674347 635432
rect 673729 635427 673795 635430
rect 674281 635427 674347 635430
rect 40534 635292 40540 635356
rect 40604 635292 40610 635356
rect 40726 634948 40786 635120
rect 40718 634884 40724 634948
rect 40788 634884 40794 634948
rect 35758 634541 35818 634712
rect 35758 634536 35867 634541
rect 35758 634480 35806 634536
rect 35862 634480 35867 634536
rect 35758 634478 35867 634480
rect 35801 634475 35867 634478
rect 39481 634538 39547 634541
rect 44265 634538 44331 634541
rect 39481 634536 44331 634538
rect 39481 634480 39486 634536
rect 39542 634480 44270 634536
rect 44326 634480 44331 634536
rect 39481 634478 44331 634480
rect 39481 634475 39547 634478
rect 44265 634475 44331 634478
rect 35574 633725 35634 634304
rect 35574 633720 35683 633725
rect 35574 633664 35622 633720
rect 35678 633664 35683 633720
rect 35574 633662 35683 633664
rect 35617 633659 35683 633662
rect 40125 633722 40191 633725
rect 43621 633722 43687 633725
rect 40125 633720 43687 633722
rect 40125 633664 40130 633720
rect 40186 633664 43626 633720
rect 43682 633664 43687 633720
rect 40125 633662 43687 633664
rect 40125 633659 40191 633662
rect 43621 633659 43687 633662
rect 35758 633317 35818 633488
rect 35758 633312 35867 633317
rect 35758 633256 35806 633312
rect 35862 633256 35867 633312
rect 35758 633254 35867 633256
rect 35801 633251 35867 633254
rect 41597 633314 41663 633317
rect 42057 633314 42123 633317
rect 41597 633312 42123 633314
rect 41597 633256 41602 633312
rect 41658 633256 42062 633312
rect 42118 633256 42123 633312
rect 41597 633254 42123 633256
rect 41597 633251 41663 633254
rect 42057 633251 42123 633254
rect 39757 632906 39823 632909
rect 44817 632906 44883 632909
rect 39757 632904 44883 632906
rect 39757 632848 39762 632904
rect 39818 632848 44822 632904
rect 44878 632848 44883 632904
rect 39757 632846 44883 632848
rect 39757 632843 39823 632846
rect 44817 632843 44883 632846
rect 40401 632634 40467 632637
rect 42701 632634 42767 632637
rect 40401 632632 42767 632634
rect 40401 632576 40406 632632
rect 40462 632576 42706 632632
rect 42762 632576 42767 632632
rect 40401 632574 42767 632576
rect 40401 632571 40467 632574
rect 42701 632571 42767 632574
rect 674925 631410 674991 631413
rect 676070 631410 676076 631412
rect 674925 631408 676076 631410
rect 674925 631352 674930 631408
rect 674986 631352 676076 631408
rect 674925 631350 676076 631352
rect 674925 631347 674991 631350
rect 676070 631348 676076 631350
rect 676140 631348 676146 631412
rect 32397 629914 32463 629917
rect 41638 629914 41644 629916
rect 32397 629912 41644 629914
rect 32397 629856 32402 629912
rect 32458 629856 41644 629912
rect 32397 629854 41644 629856
rect 32397 629851 32463 629854
rect 41638 629852 41644 629854
rect 41708 629852 41714 629916
rect 37917 629234 37983 629237
rect 41822 629234 41828 629236
rect 37917 629232 41828 629234
rect 37917 629176 37922 629232
rect 37978 629176 41828 629232
rect 37917 629174 41828 629176
rect 37917 629171 37983 629174
rect 41822 629172 41828 629174
rect 41892 629172 41898 629236
rect 40493 628690 40559 628693
rect 42333 628690 42399 628693
rect 40493 628688 42399 628690
rect 40493 628632 40498 628688
rect 40554 628632 42338 628688
rect 42394 628632 42399 628688
rect 40493 628630 42399 628632
rect 40493 628627 40559 628630
rect 42333 628627 42399 628630
rect 41781 627464 41847 627469
rect 41781 627408 41786 627464
rect 41842 627408 41847 627464
rect 41781 627403 41847 627408
rect 41784 627197 41844 627403
rect 41781 627192 41847 627197
rect 41781 627136 41786 627192
rect 41842 627136 41847 627192
rect 41781 627131 41847 627136
rect 676262 626109 676322 626348
rect 676213 626104 676322 626109
rect 676213 626048 676218 626104
rect 676274 626048 676322 626104
rect 676213 626046 676322 626048
rect 676213 626043 676279 626046
rect 676262 625701 676322 625940
rect 676213 625696 676322 625701
rect 676213 625640 676218 625696
rect 676274 625640 676322 625696
rect 676213 625638 676322 625640
rect 676213 625635 676279 625638
rect 676262 625293 676322 625532
rect 676213 625288 676322 625293
rect 676489 625290 676555 625293
rect 676213 625232 676218 625288
rect 676274 625232 676322 625288
rect 676213 625230 676322 625232
rect 676446 625288 676555 625290
rect 676446 625232 676494 625288
rect 676550 625232 676555 625288
rect 676213 625227 676279 625230
rect 676446 625227 676555 625232
rect 676446 625124 676506 625227
rect 676029 624746 676095 624749
rect 676029 624744 676292 624746
rect 676029 624688 676034 624744
rect 676090 624688 676292 624744
rect 676029 624686 676292 624688
rect 676029 624683 676095 624686
rect 42057 624474 42123 624477
rect 44449 624474 44515 624477
rect 42057 624472 44515 624474
rect 42057 624416 42062 624472
rect 42118 624416 44454 624472
rect 44510 624416 44515 624472
rect 42057 624414 44515 624416
rect 42057 624411 42123 624414
rect 44449 624411 44515 624414
rect 676213 624474 676279 624477
rect 676213 624472 676322 624474
rect 676213 624416 676218 624472
rect 676274 624416 676322 624472
rect 676213 624411 676322 624416
rect 676262 624308 676322 624411
rect 674005 623930 674071 623933
rect 674005 623928 676292 623930
rect 674005 623872 674010 623928
rect 674066 623872 676292 623928
rect 674005 623870 676292 623872
rect 674005 623867 674071 623870
rect 676213 623658 676279 623661
rect 676213 623656 676322 623658
rect 676213 623600 676218 623656
rect 676274 623600 676322 623656
rect 676213 623595 676322 623600
rect 676262 623492 676322 623595
rect 40902 623324 40908 623388
rect 40972 623386 40978 623388
rect 41781 623386 41847 623389
rect 40972 623384 41847 623386
rect 40972 623328 41786 623384
rect 41842 623328 41847 623384
rect 40972 623326 41847 623328
rect 40972 623324 40978 623326
rect 41781 623323 41847 623326
rect 674005 623114 674071 623117
rect 674005 623112 676292 623114
rect 674005 623056 674010 623112
rect 674066 623056 676292 623112
rect 674005 623054 676292 623056
rect 674005 623051 674071 623054
rect 676213 622842 676279 622845
rect 676213 622840 676322 622842
rect 676213 622784 676218 622840
rect 676274 622784 676322 622840
rect 676213 622779 676322 622784
rect 676262 622676 676322 622779
rect 674005 622298 674071 622301
rect 674005 622296 676292 622298
rect 674005 622240 674010 622296
rect 674066 622240 676292 622296
rect 674005 622238 676292 622240
rect 674005 622235 674071 622238
rect 40718 621964 40724 622028
rect 40788 622026 40794 622028
rect 41781 622026 41847 622029
rect 40788 622024 41847 622026
rect 40788 621968 41786 622024
rect 41842 621968 41847 622024
rect 40788 621966 41847 621968
rect 40788 621964 40794 621966
rect 41781 621963 41847 621966
rect 42149 622026 42215 622029
rect 44725 622026 44791 622029
rect 682377 622026 682443 622029
rect 42149 622024 44791 622026
rect 42149 621968 42154 622024
rect 42210 621968 44730 622024
rect 44786 621968 44791 622024
rect 42149 621966 44791 621968
rect 42149 621963 42215 621966
rect 44725 621963 44791 621966
rect 682334 622024 682443 622026
rect 682334 621968 682382 622024
rect 682438 621968 682443 622024
rect 682334 621963 682443 621968
rect 682334 621860 682394 621963
rect 675293 621482 675359 621485
rect 675293 621480 676292 621482
rect 675293 621424 675298 621480
rect 675354 621424 676292 621480
rect 675293 621422 676292 621424
rect 675293 621419 675359 621422
rect 676213 621210 676279 621213
rect 676213 621208 676322 621210
rect 676213 621152 676218 621208
rect 676274 621152 676322 621208
rect 676213 621147 676322 621152
rect 676262 621044 676322 621147
rect 40534 620740 40540 620804
rect 40604 620802 40610 620804
rect 41781 620802 41847 620805
rect 40604 620800 41847 620802
rect 40604 620744 41786 620800
rect 41842 620744 41847 620800
rect 40604 620742 41847 620744
rect 40604 620740 40610 620742
rect 41781 620739 41847 620742
rect 676213 620802 676279 620805
rect 676213 620800 676322 620802
rect 676213 620744 676218 620800
rect 676274 620744 676322 620800
rect 676213 620739 676322 620744
rect 676262 620636 676322 620739
rect 683941 620394 684007 620397
rect 683941 620392 684050 620394
rect 683941 620336 683946 620392
rect 684002 620336 684050 620392
rect 683941 620331 684050 620336
rect 683990 620228 684050 620331
rect 676029 619850 676095 619853
rect 676029 619848 676292 619850
rect 676029 619792 676034 619848
rect 676090 619792 676292 619848
rect 676029 619790 676292 619792
rect 676029 619787 676095 619790
rect 676262 619173 676322 619412
rect 676213 619168 676322 619173
rect 676489 619170 676555 619173
rect 676213 619112 676218 619168
rect 676274 619112 676322 619168
rect 676213 619110 676322 619112
rect 676446 619168 676555 619170
rect 676446 619112 676494 619168
rect 676550 619112 676555 619168
rect 676213 619107 676279 619110
rect 676446 619107 676555 619112
rect 676446 619004 676506 619107
rect 672993 618626 673059 618629
rect 672993 618624 676292 618626
rect 672993 618568 672998 618624
rect 673054 618568 676292 618624
rect 672993 618566 676292 618568
rect 672993 618563 673059 618566
rect 676029 618218 676095 618221
rect 676029 618216 676292 618218
rect 676029 618160 676034 618216
rect 676090 618160 676292 618216
rect 676029 618158 676292 618160
rect 676029 618155 676095 618158
rect 63125 618082 63191 618085
rect 63125 618080 64706 618082
rect 63125 618024 63130 618080
rect 63186 618024 64706 618080
rect 63125 618022 64706 618024
rect 63125 618019 63191 618022
rect 64646 617416 64706 618022
rect 676213 617946 676279 617949
rect 676213 617944 676322 617946
rect 676213 617888 676218 617944
rect 676274 617888 676322 617944
rect 676213 617883 676322 617888
rect 676262 617780 676322 617883
rect 683113 617538 683179 617541
rect 683070 617536 683179 617538
rect 683070 617480 683118 617536
rect 683174 617480 683179 617536
rect 683070 617475 683179 617480
rect 683070 617372 683130 617475
rect 683297 617130 683363 617133
rect 683254 617128 683363 617130
rect 683254 617072 683302 617128
rect 683358 617072 683363 617128
rect 683254 617067 683363 617072
rect 683254 616964 683314 617067
rect 676213 616722 676279 616725
rect 676213 616720 676322 616722
rect 676213 616664 676218 616720
rect 676274 616664 676322 616720
rect 676213 616659 676322 616664
rect 62113 616586 62179 616589
rect 62113 616584 64706 616586
rect 62113 616528 62118 616584
rect 62174 616528 64706 616584
rect 676262 616556 676322 616659
rect 62113 616526 64706 616528
rect 62113 616523 62179 616526
rect 64646 616234 64706 616526
rect 673862 616116 673868 616180
rect 673932 616178 673938 616180
rect 673932 616118 676292 616178
rect 673932 616116 673938 616118
rect 41454 615980 41460 616044
rect 41524 616042 41530 616044
rect 41873 616042 41939 616045
rect 41524 616040 41939 616042
rect 41524 615984 41878 616040
rect 41934 615984 41939 616040
rect 41524 615982 41939 615984
rect 41524 615980 41530 615982
rect 41873 615979 41939 615982
rect 42057 615906 42123 615909
rect 42701 615906 42767 615909
rect 42057 615904 42767 615906
rect 42057 615848 42062 615904
rect 42118 615848 42706 615904
rect 42762 615848 42767 615904
rect 42057 615846 42767 615848
rect 42057 615843 42123 615846
rect 42701 615843 42767 615846
rect 683070 615501 683130 615740
rect 41822 615436 41828 615500
rect 41892 615498 41898 615500
rect 42609 615498 42675 615501
rect 41892 615496 42675 615498
rect 41892 615440 42614 615496
rect 42670 615440 42675 615496
rect 41892 615438 42675 615440
rect 41892 615436 41898 615438
rect 42609 615435 42675 615438
rect 683070 615498 683179 615501
rect 683070 615496 683260 615498
rect 683070 615440 683118 615496
rect 683174 615440 683260 615496
rect 683070 615438 683260 615440
rect 683070 615435 683179 615438
rect 683070 615332 683130 615435
rect 62113 614682 62179 614685
rect 64646 614682 64706 615052
rect 674005 614954 674071 614957
rect 674005 614952 676292 614954
rect 674005 614896 674010 614952
rect 674066 614896 676292 614952
rect 674005 614894 676292 614896
rect 674005 614891 674071 614894
rect 62113 614680 64706 614682
rect 62113 614624 62118 614680
rect 62174 614624 64706 614680
rect 62113 614622 64706 614624
rect 62113 614619 62179 614622
rect 61377 613866 61443 613869
rect 64646 613866 64706 613870
rect 61377 613864 64706 613866
rect 61377 613808 61382 613864
rect 61438 613808 64706 613864
rect 61377 613806 64706 613808
rect 61377 613803 61443 613806
rect 41873 613460 41939 613461
rect 41822 613458 41828 613460
rect 41782 613398 41828 613458
rect 41892 613456 41939 613460
rect 41934 613400 41939 613456
rect 41822 613396 41828 613398
rect 41892 613396 41939 613400
rect 41873 613395 41939 613396
rect 62113 612642 62179 612645
rect 64646 612642 64706 612688
rect 62113 612640 64706 612642
rect 62113 612584 62118 612640
rect 62174 612584 64706 612640
rect 62113 612582 64706 612584
rect 62113 612579 62179 612582
rect 43253 612234 43319 612237
rect 43759 612234 43825 612237
rect 43253 612232 43825 612234
rect 43253 612176 43258 612232
rect 43314 612176 43764 612232
rect 43820 612176 43825 612232
rect 43253 612174 43825 612176
rect 43253 612171 43319 612174
rect 43759 612171 43825 612174
rect 43868 612098 43934 612101
rect 45553 612098 45619 612101
rect 43868 612096 45619 612098
rect 43868 612040 43873 612096
rect 43929 612040 45558 612096
rect 45614 612040 45619 612096
rect 43868 612038 45619 612040
rect 43868 612035 43934 612038
rect 45553 612035 45619 612038
rect 62941 612098 63007 612101
rect 62941 612096 64706 612098
rect 62941 612040 62946 612096
rect 63002 612040 64706 612096
rect 62941 612038 64706 612040
rect 62941 612035 63007 612038
rect 64646 611506 64706 612038
rect 673177 608154 673243 608157
rect 675109 608154 675175 608157
rect 673177 608152 675175 608154
rect 673177 608096 673182 608152
rect 673238 608096 675114 608152
rect 675170 608096 675175 608152
rect 673177 608094 675175 608096
rect 673177 608091 673243 608094
rect 675109 608091 675175 608094
rect 671153 607338 671219 607341
rect 675109 607338 675175 607341
rect 671153 607336 675175 607338
rect 671153 607280 671158 607336
rect 671214 607280 675114 607336
rect 675170 607280 675175 607336
rect 671153 607278 675175 607280
rect 671153 607275 671219 607278
rect 675109 607275 675175 607278
rect 674833 607066 674899 607069
rect 675886 607066 675892 607068
rect 674833 607064 675892 607066
rect 674833 607008 674838 607064
rect 674894 607008 675892 607064
rect 674833 607006 675892 607008
rect 674833 607003 674899 607006
rect 675886 607004 675892 607006
rect 675956 607004 675962 607068
rect 672349 604346 672415 604349
rect 675385 604346 675451 604349
rect 672349 604344 675451 604346
rect 672349 604288 672354 604344
rect 672410 604288 675390 604344
rect 675446 604288 675451 604344
rect 672349 604286 675451 604288
rect 672349 604283 672415 604286
rect 675385 604283 675451 604286
rect 672993 604074 673059 604077
rect 675477 604074 675543 604077
rect 672993 604072 675543 604074
rect 672993 604016 672998 604072
rect 673054 604016 675482 604072
rect 675538 604016 675543 604072
rect 672993 604014 675543 604016
rect 672993 604011 673059 604014
rect 675477 604011 675543 604014
rect 673729 603802 673795 603805
rect 674465 603802 674531 603805
rect 673729 603800 674531 603802
rect 673729 603744 673734 603800
rect 673790 603744 674470 603800
rect 674526 603744 674531 603800
rect 673729 603742 674531 603744
rect 673729 603739 673795 603742
rect 674465 603739 674531 603742
rect 674230 602788 674236 602852
rect 674300 602850 674306 602852
rect 675385 602850 675451 602853
rect 674300 602848 675451 602850
rect 674300 602792 675390 602848
rect 675446 602792 675451 602848
rect 674300 602790 675451 602792
rect 674300 602788 674306 602790
rect 675385 602787 675451 602790
rect 33777 601762 33843 601765
rect 33764 601760 33843 601762
rect 33764 601704 33782 601760
rect 33838 601704 33843 601760
rect 33764 601702 33843 601704
rect 33777 601699 33843 601702
rect 38561 601354 38627 601357
rect 38548 601352 38627 601354
rect 38548 601296 38566 601352
rect 38622 601296 38627 601352
rect 38548 601294 38627 601296
rect 38561 601291 38627 601294
rect 39941 600946 40007 600949
rect 668945 600946 669011 600949
rect 675477 600946 675543 600949
rect 39941 600944 40020 600946
rect 39941 600888 39946 600944
rect 40002 600888 40020 600944
rect 39941 600886 40020 600888
rect 668945 600944 675543 600946
rect 668945 600888 668950 600944
rect 669006 600888 675482 600944
rect 675538 600888 675543 600944
rect 668945 600886 675543 600888
rect 39941 600883 40007 600886
rect 668945 600883 669011 600886
rect 675477 600883 675543 600886
rect 45001 600538 45067 600541
rect 41492 600536 45067 600538
rect 41492 600480 45006 600536
rect 45062 600480 45067 600536
rect 41492 600478 45067 600480
rect 45001 600475 45067 600478
rect 670877 600402 670943 600405
rect 675385 600402 675451 600405
rect 670877 600400 675451 600402
rect 670877 600344 670882 600400
rect 670938 600344 675390 600400
rect 675446 600344 675451 600400
rect 670877 600342 675451 600344
rect 670877 600339 670943 600342
rect 675385 600339 675451 600342
rect 44633 600130 44699 600133
rect 41492 600128 44699 600130
rect 41492 600072 44638 600128
rect 44694 600072 44699 600128
rect 41492 600070 44699 600072
rect 44633 600067 44699 600070
rect 673729 599858 673795 599861
rect 675477 599858 675543 599861
rect 673729 599856 675543 599858
rect 673729 599800 673734 599856
rect 673790 599800 675482 599856
rect 675538 599800 675543 599856
rect 673729 599798 675543 599800
rect 673729 599795 673795 599798
rect 675477 599795 675543 599798
rect 44214 599722 44220 599724
rect 41492 599662 44220 599722
rect 44214 599660 44220 599662
rect 44284 599660 44290 599724
rect 43110 599314 43116 599316
rect 41492 599254 43116 599314
rect 43110 599252 43116 599254
rect 43180 599252 43186 599316
rect 670785 599178 670851 599181
rect 674097 599178 674163 599181
rect 670785 599176 674163 599178
rect 670785 599120 670790 599176
rect 670846 599120 674102 599176
rect 674158 599120 674163 599176
rect 670785 599118 674163 599120
rect 670785 599115 670851 599118
rect 674097 599115 674163 599118
rect 674281 599178 674347 599181
rect 675385 599178 675451 599181
rect 674281 599176 675451 599178
rect 674281 599120 674286 599176
rect 674342 599120 675390 599176
rect 675446 599120 675451 599176
rect 674281 599118 675451 599120
rect 674281 599115 674347 599118
rect 675385 599115 675451 599118
rect 675886 599116 675892 599180
rect 675956 599116 675962 599180
rect 675894 598950 675954 599116
rect 45369 598906 45435 598909
rect 41492 598904 45435 598906
rect 41492 598848 45374 598904
rect 45430 598848 45435 598904
rect 41492 598846 45435 598848
rect 675710 598906 675954 598950
rect 676990 598906 676996 598908
rect 675710 598846 676996 598906
rect 45369 598843 45435 598846
rect 676990 598844 676996 598846
rect 677060 598844 677066 598908
rect 674465 598634 674531 598637
rect 675477 598634 675543 598637
rect 674465 598632 675543 598634
rect 674465 598576 674470 598632
rect 674526 598576 675482 598632
rect 675538 598576 675543 598632
rect 674465 598574 675543 598576
rect 674465 598571 674531 598574
rect 675477 598571 675543 598574
rect 44909 598498 44975 598501
rect 41492 598496 44975 598498
rect 41492 598440 44914 598496
rect 44970 598440 44975 598496
rect 41492 598438 44975 598440
rect 44909 598435 44975 598438
rect 45185 598090 45251 598093
rect 41492 598088 45251 598090
rect 41492 598032 45190 598088
rect 45246 598032 45251 598088
rect 41492 598030 45251 598032
rect 45185 598027 45251 598030
rect 649950 597954 650010 598336
rect 674005 598090 674071 598093
rect 675293 598090 675359 598093
rect 674005 598088 675359 598090
rect 674005 598032 674010 598088
rect 674066 598032 675298 598088
rect 675354 598032 675359 598088
rect 674005 598030 675359 598032
rect 674005 598027 674071 598030
rect 675293 598027 675359 598030
rect 651465 597954 651531 597957
rect 649950 597952 651531 597954
rect 649950 597896 651470 597952
rect 651526 597896 651531 597952
rect 649950 597894 651531 597896
rect 651465 597891 651531 597894
rect 42885 597682 42951 597685
rect 41492 597680 42951 597682
rect 41492 597624 42890 597680
rect 42946 597624 42951 597680
rect 41492 597622 42951 597624
rect 42885 597619 42951 597622
rect 674097 597410 674163 597413
rect 675477 597410 675543 597413
rect 674097 597408 675543 597410
rect 674097 597352 674102 597408
rect 674158 597352 675482 597408
rect 675538 597352 675543 597408
rect 674097 597350 675543 597352
rect 674097 597347 674163 597350
rect 675477 597347 675543 597350
rect 41094 597038 41154 597244
rect 41086 596974 41092 597038
rect 41156 596974 41162 597038
rect 43069 597004 43135 597005
rect 43069 597000 43116 597004
rect 43180 597002 43186 597004
rect 43069 596944 43074 597000
rect 43069 596940 43116 596944
rect 43180 596942 43226 597002
rect 43180 596940 43186 596942
rect 43069 596939 43135 596940
rect 42149 596866 42215 596869
rect 41492 596864 42215 596866
rect 41492 596808 42154 596864
rect 42210 596808 42215 596864
rect 41492 596806 42215 596808
rect 42149 596803 42215 596806
rect 649950 596730 650010 597154
rect 651465 596730 651531 596733
rect 649950 596728 651531 596730
rect 649950 596672 651470 596728
rect 651526 596672 651531 596728
rect 649950 596670 651531 596672
rect 651465 596667 651531 596670
rect 41822 596458 41828 596460
rect 41492 596398 41828 596458
rect 41822 596396 41828 596398
rect 41892 596396 41898 596460
rect 42701 596050 42767 596053
rect 41492 596048 42767 596050
rect 41492 595992 42706 596048
rect 42762 595992 42767 596048
rect 41492 595990 42767 595992
rect 42701 595987 42767 595990
rect 35433 595812 35499 595815
rect 35390 595810 35499 595812
rect 35390 595754 35438 595810
rect 35494 595754 35499 595810
rect 35390 595749 35499 595754
rect 41689 595778 41755 595781
rect 62665 595778 62731 595781
rect 41689 595776 62731 595778
rect 35390 595612 35450 595749
rect 41689 595720 41694 595776
rect 41750 595720 62670 595776
rect 62726 595720 62731 595776
rect 41689 595718 62731 595720
rect 41689 595715 41755 595718
rect 62665 595715 62731 595718
rect 649950 595370 650010 595972
rect 651465 595370 651531 595373
rect 649950 595368 651531 595370
rect 649950 595312 651470 595368
rect 651526 595312 651531 595368
rect 649950 595310 651531 595312
rect 651465 595307 651531 595310
rect 32397 595234 32463 595237
rect 32397 595232 32476 595234
rect 32397 595176 32402 595232
rect 32458 595176 32476 595232
rect 32397 595174 32476 595176
rect 32397 595171 32463 595174
rect 651649 595098 651715 595101
rect 649950 595096 651715 595098
rect 649950 595040 651654 595096
rect 651710 595040 651715 595096
rect 649950 595038 651715 595040
rect 39297 594826 39363 594829
rect 39284 594824 39363 594826
rect 39284 594768 39302 594824
rect 39358 594768 39363 594824
rect 649950 594790 650010 595038
rect 651649 595035 651715 595038
rect 668761 594826 668827 594829
rect 675477 594826 675543 594829
rect 668761 594824 675543 594826
rect 39284 594766 39363 594768
rect 39297 594763 39363 594766
rect 668761 594768 668766 594824
rect 668822 594768 675482 594824
rect 675538 594768 675543 594824
rect 668761 594766 675543 594768
rect 668761 594763 668827 594766
rect 675477 594763 675543 594766
rect 31017 594418 31083 594421
rect 31004 594416 31083 594418
rect 31004 594360 31022 594416
rect 31078 594360 31083 594416
rect 31004 594358 31083 594360
rect 31017 594355 31083 594358
rect 40534 594118 40540 594182
rect 40604 594118 40610 594182
rect 41689 594146 41755 594149
rect 63125 594146 63191 594149
rect 651465 594146 651531 594149
rect 41689 594144 63191 594146
rect 40542 593980 40602 594118
rect 41689 594088 41694 594144
rect 41750 594088 63130 594144
rect 63186 594088 63191 594144
rect 41689 594086 63191 594088
rect 41689 594083 41755 594086
rect 63125 594083 63191 594086
rect 649950 594144 651531 594146
rect 649950 594088 651470 594144
rect 651526 594088 651531 594144
rect 649950 594086 651531 594088
rect 649950 593608 650010 594086
rect 651465 594083 651531 594086
rect 36537 593602 36603 593605
rect 36524 593600 36603 593602
rect 36524 593544 36542 593600
rect 36598 593544 36603 593600
rect 36524 593542 36603 593544
rect 36537 593539 36603 593542
rect 670969 593602 671035 593605
rect 675477 593602 675543 593605
rect 670969 593600 675543 593602
rect 670969 593544 670974 593600
rect 671030 593544 675482 593600
rect 675538 593544 675543 593600
rect 670969 593542 675543 593544
rect 670969 593539 671035 593542
rect 675477 593539 675543 593542
rect 44357 593194 44423 593197
rect 41492 593192 44423 593194
rect 41492 593136 44362 593192
rect 44418 593136 44423 593192
rect 41492 593134 44423 593136
rect 44357 593131 44423 593134
rect 677174 592860 677180 592924
rect 677244 592922 677250 592924
rect 677501 592922 677567 592925
rect 677244 592920 677567 592922
rect 677244 592864 677506 592920
rect 677562 592864 677567 592920
rect 677244 592862 677567 592864
rect 677244 592860 677250 592862
rect 677501 592859 677567 592862
rect 41965 592786 42031 592789
rect 651465 592786 651531 592789
rect 41492 592784 42031 592786
rect 41492 592728 41970 592784
rect 42026 592728 42031 592784
rect 41492 592726 42031 592728
rect 41965 592723 42031 592726
rect 649950 592784 651531 592786
rect 649950 592728 651470 592784
rect 651526 592728 651531 592784
rect 649950 592726 651531 592728
rect 649950 592426 650010 592726
rect 651465 592723 651531 592726
rect 676070 592588 676076 592652
rect 676140 592650 676146 592652
rect 678237 592650 678303 592653
rect 676140 592648 678303 592650
rect 676140 592592 678242 592648
rect 678298 592592 678303 592648
rect 676140 592590 678303 592592
rect 676140 592588 676146 592590
rect 678237 592587 678303 592590
rect 41781 592378 41847 592381
rect 41492 592376 41847 592378
rect 41492 592320 41786 592376
rect 41842 592320 41847 592376
rect 41492 592318 41847 592320
rect 41781 592315 41847 592318
rect 44173 591970 44239 591973
rect 41492 591968 44239 591970
rect 41492 591912 44178 591968
rect 44234 591912 44239 591968
rect 41492 591910 44239 591912
rect 44173 591907 44239 591910
rect 43345 591562 43411 591565
rect 41492 591560 43411 591562
rect 41492 591504 43350 591560
rect 43406 591504 43411 591560
rect 41492 591502 43411 591504
rect 43345 591499 43411 591502
rect 674414 591228 674420 591292
rect 674484 591290 674490 591292
rect 684217 591290 684283 591293
rect 674484 591288 684283 591290
rect 674484 591232 684222 591288
rect 684278 591232 684283 591288
rect 674484 591230 684283 591232
rect 674484 591228 674490 591230
rect 684217 591227 684283 591230
rect 41462 590746 41522 591124
rect 62941 590746 63007 590749
rect 41462 590744 63007 590746
rect 41462 590716 62946 590744
rect 41492 590688 62946 590716
rect 63002 590688 63007 590744
rect 41492 590686 63007 590688
rect 62941 590683 63007 590686
rect 41781 590338 41847 590341
rect 41492 590336 41847 590338
rect 41492 590280 41786 590336
rect 41842 590280 41847 590336
rect 41492 590278 41847 590280
rect 41781 590275 41847 590278
rect 62849 590066 62915 590069
rect 51030 590064 62915 590066
rect 51030 590008 62854 590064
rect 62910 590008 62915 590064
rect 51030 590006 62915 590008
rect 40718 589596 40724 589660
rect 40788 589658 40794 589660
rect 41965 589658 42031 589661
rect 40788 589656 42031 589658
rect 40788 589600 41970 589656
rect 42026 589600 42031 589656
rect 40788 589598 42031 589600
rect 40788 589596 40794 589598
rect 41965 589595 42031 589598
rect 33777 589386 33843 589389
rect 51030 589386 51090 590006
rect 62849 590003 62915 590006
rect 33777 589384 51090 589386
rect 33777 589328 33782 589384
rect 33838 589328 51090 589384
rect 33777 589326 51090 589328
rect 33777 589323 33843 589326
rect 40902 589052 40908 589116
rect 40972 589114 40978 589116
rect 41505 589114 41571 589117
rect 40972 589112 41571 589114
rect 40972 589056 41510 589112
rect 41566 589056 41571 589112
rect 40972 589054 41571 589056
rect 40972 589052 40978 589054
rect 41505 589051 41571 589054
rect 41689 589114 41755 589117
rect 43621 589114 43687 589117
rect 41689 589112 43687 589114
rect 41689 589056 41694 589112
rect 41750 589056 43626 589112
rect 43682 589056 43687 589112
rect 41689 589054 43687 589056
rect 41689 589051 41755 589054
rect 43621 589051 43687 589054
rect 673545 588570 673611 588573
rect 675569 588570 675635 588573
rect 673545 588568 675635 588570
rect 673545 588512 673550 588568
rect 673606 588512 675574 588568
rect 675630 588512 675635 588568
rect 673545 588510 675635 588512
rect 673545 588507 673611 588510
rect 675569 588507 675635 588510
rect 41505 586938 41571 586941
rect 42793 586938 42859 586941
rect 41505 586936 42859 586938
rect 41505 586880 41510 586936
rect 41566 586880 42798 586936
rect 42854 586880 42859 586936
rect 41505 586878 42859 586880
rect 41505 586875 41571 586878
rect 42793 586875 42859 586878
rect 674925 586532 674991 586533
rect 674925 586530 674972 586532
rect 674880 586528 674972 586530
rect 674880 586472 674930 586528
rect 674880 586470 674972 586472
rect 674925 586468 674972 586470
rect 675036 586468 675042 586532
rect 674925 586467 674991 586468
rect 675109 586258 675175 586261
rect 676070 586258 676076 586260
rect 675109 586256 676076 586258
rect 675109 586200 675114 586256
rect 675170 586200 676076 586256
rect 675109 586198 676076 586200
rect 675109 586195 675175 586198
rect 676070 586196 676076 586198
rect 676140 586196 676146 586260
rect 39665 586122 39731 586125
rect 40350 586122 40356 586124
rect 39665 586120 40356 586122
rect 39665 586064 39670 586120
rect 39726 586064 40356 586120
rect 39665 586062 40356 586064
rect 39665 586059 39731 586062
rect 40350 586060 40356 586062
rect 40420 586060 40426 586124
rect 39297 585170 39363 585173
rect 41822 585170 41828 585172
rect 39297 585168 41828 585170
rect 39297 585112 39302 585168
rect 39358 585112 41828 585168
rect 39297 585110 41828 585112
rect 39297 585107 39363 585110
rect 41822 585108 41828 585110
rect 41892 585108 41898 585172
rect 39757 584626 39823 584629
rect 42609 584626 42675 584629
rect 39757 584624 42675 584626
rect 39757 584568 39762 584624
rect 39818 584568 42614 584624
rect 42670 584568 42675 584624
rect 39757 584566 42675 584568
rect 39757 584563 39823 584566
rect 42609 584563 42675 584566
rect 42333 581226 42399 581229
rect 44173 581226 44239 581229
rect 42333 581224 44239 581226
rect 42333 581168 42338 581224
rect 42394 581168 44178 581224
rect 44234 581168 44239 581224
rect 42333 581166 44239 581168
rect 42333 581163 42399 581166
rect 44173 581163 44239 581166
rect 673913 581090 673979 581093
rect 673913 581088 676292 581090
rect 673913 581032 673918 581088
rect 673974 581032 676292 581088
rect 673913 581030 676292 581032
rect 673913 581027 673979 581030
rect 42057 580682 42123 580685
rect 45093 580682 45159 580685
rect 42057 580680 45159 580682
rect 42057 580624 42062 580680
rect 42118 580624 45098 580680
rect 45154 580624 45159 580680
rect 42057 580622 45159 580624
rect 42057 580619 42123 580622
rect 45093 580619 45159 580622
rect 673545 580682 673611 580685
rect 673545 580680 676292 580682
rect 673545 580624 673550 580680
rect 673606 580624 676292 580680
rect 673545 580622 676292 580624
rect 673545 580619 673611 580622
rect 40350 580212 40356 580276
rect 40420 580274 40426 580276
rect 41781 580274 41847 580277
rect 40420 580272 41847 580274
rect 40420 580216 41786 580272
rect 41842 580216 41847 580272
rect 40420 580214 41847 580216
rect 40420 580212 40426 580214
rect 41781 580211 41847 580214
rect 673913 580274 673979 580277
rect 673913 580272 676292 580274
rect 673913 580216 673918 580272
rect 673974 580216 676292 580272
rect 673913 580214 676292 580216
rect 673913 580211 673979 580214
rect 673913 579866 673979 579869
rect 673913 579864 676292 579866
rect 673913 579808 673918 579864
rect 673974 579808 676292 579864
rect 673913 579806 676292 579808
rect 673913 579803 673979 579806
rect 673913 579458 673979 579461
rect 673913 579456 676292 579458
rect 673913 579400 673918 579456
rect 673974 579400 676292 579456
rect 673913 579398 676292 579400
rect 673913 579395 673979 579398
rect 673913 579050 673979 579053
rect 673913 579048 676292 579050
rect 673913 578992 673918 579048
rect 673974 578992 676292 579048
rect 673913 578990 676292 578992
rect 673913 578987 673979 578990
rect 42241 578914 42307 578917
rect 45553 578914 45619 578917
rect 42241 578912 45619 578914
rect 42241 578856 42246 578912
rect 42302 578856 45558 578912
rect 45614 578856 45619 578912
rect 42241 578854 45619 578856
rect 42241 578851 42307 578854
rect 45553 578851 45619 578854
rect 673913 578642 673979 578645
rect 673913 578640 676292 578642
rect 673913 578584 673918 578640
rect 673974 578584 676292 578640
rect 673913 578582 676292 578584
rect 673913 578579 673979 578582
rect 673913 578234 673979 578237
rect 673913 578232 676292 578234
rect 673913 578176 673918 578232
rect 673974 578176 676292 578232
rect 673913 578174 676292 578176
rect 673913 578171 673979 578174
rect 42241 578098 42307 578101
rect 44357 578098 44423 578101
rect 42241 578096 44423 578098
rect 42241 578040 42246 578096
rect 42302 578040 44362 578096
rect 44418 578040 44423 578096
rect 42241 578038 44423 578040
rect 42241 578035 42307 578038
rect 44357 578035 44423 578038
rect 40902 577764 40908 577828
rect 40972 577826 40978 577828
rect 41781 577826 41847 577829
rect 40972 577824 41847 577826
rect 40972 577768 41786 577824
rect 41842 577768 41847 577824
rect 40972 577766 41847 577768
rect 40972 577764 40978 577766
rect 41781 577763 41847 577766
rect 673913 577826 673979 577829
rect 673913 577824 676292 577826
rect 673913 577768 673918 577824
rect 673974 577768 676292 577824
rect 673913 577766 676292 577768
rect 673913 577763 673979 577766
rect 42793 577418 42859 577421
rect 42014 577416 42859 577418
rect 42014 577360 42798 577416
rect 42854 577360 42859 577416
rect 42014 577358 42859 577360
rect 42014 577149 42074 577358
rect 42793 577355 42859 577358
rect 673913 577418 673979 577421
rect 673913 577416 676292 577418
rect 673913 577360 673918 577416
rect 673974 577360 676292 577416
rect 673913 577358 676292 577360
rect 673913 577355 673979 577358
rect 41965 577144 42074 577149
rect 41965 577088 41970 577144
rect 42026 577088 42074 577144
rect 41965 577086 42074 577088
rect 41965 577083 42031 577086
rect 673913 577010 673979 577013
rect 673913 577008 676292 577010
rect 673913 576952 673918 577008
rect 673974 576952 676292 577008
rect 673913 576950 676292 576952
rect 673913 576947 673979 576950
rect 678237 576874 678303 576877
rect 678237 576872 678346 576874
rect 678237 576816 678242 576872
rect 678298 576816 678346 576872
rect 678237 576811 678346 576816
rect 678286 576572 678346 576811
rect 676990 576404 676996 576468
rect 677060 576404 677066 576468
rect 676998 576164 677058 576404
rect 684217 576058 684283 576061
rect 684174 576056 684283 576058
rect 684174 576000 684222 576056
rect 684278 576000 684283 576056
rect 684174 575995 684283 576000
rect 684174 575756 684234 575995
rect 673913 575378 673979 575381
rect 673913 575376 676292 575378
rect 673913 575320 673918 575376
rect 673974 575320 676292 575376
rect 673913 575318 676292 575320
rect 673913 575315 673979 575318
rect 673913 574970 673979 574973
rect 673913 574968 676292 574970
rect 673913 574912 673918 574968
rect 673974 574912 676292 574968
rect 673913 574910 676292 574912
rect 673913 574907 673979 574910
rect 62389 574834 62455 574837
rect 62389 574832 64706 574834
rect 62389 574776 62394 574832
rect 62450 574776 64706 574832
rect 62389 574774 64706 574776
rect 62389 574771 62455 574774
rect 40718 574636 40724 574700
rect 40788 574698 40794 574700
rect 41781 574698 41847 574701
rect 40788 574696 41847 574698
rect 40788 574640 41786 574696
rect 41842 574640 41847 574696
rect 40788 574638 41847 574640
rect 40788 574636 40794 574638
rect 41781 574635 41847 574638
rect 64646 574194 64706 574774
rect 673545 574562 673611 574565
rect 673545 574560 676292 574562
rect 673545 574504 673550 574560
rect 673606 574504 676292 574560
rect 673545 574502 676292 574504
rect 673545 574499 673611 574502
rect 673545 574154 673611 574157
rect 673545 574152 676292 574154
rect 673545 574096 673550 574152
rect 673606 574096 676292 574152
rect 673545 574094 676292 574096
rect 673545 574091 673611 574094
rect 40534 573820 40540 573884
rect 40604 573882 40610 573884
rect 41781 573882 41847 573885
rect 40604 573880 41847 573882
rect 40604 573824 41786 573880
rect 41842 573824 41847 573880
rect 40604 573822 41847 573824
rect 40604 573820 40610 573822
rect 41781 573819 41847 573822
rect 673913 573746 673979 573749
rect 673913 573744 676292 573746
rect 673913 573688 673918 573744
rect 673974 573688 676292 573744
rect 673913 573686 676292 573688
rect 673913 573683 673979 573686
rect 62389 573610 62455 573613
rect 677501 573610 677567 573613
rect 62389 573608 64706 573610
rect 62389 573552 62394 573608
rect 62450 573552 64706 573608
rect 62389 573550 64706 573552
rect 62389 573547 62455 573550
rect 64646 573012 64706 573550
rect 677501 573608 677610 573610
rect 677501 573552 677506 573608
rect 677562 573552 677610 573608
rect 677501 573547 677610 573552
rect 677550 573308 677610 573547
rect 683389 573202 683455 573205
rect 683389 573200 683498 573202
rect 683389 573144 683394 573200
rect 683450 573144 683498 573200
rect 683389 573139 683498 573144
rect 683438 572900 683498 573139
rect 676806 572732 676812 572796
rect 676876 572732 676882 572796
rect 676814 572492 676874 572732
rect 41822 572188 41828 572252
rect 41892 572250 41898 572252
rect 42241 572250 42307 572253
rect 41892 572248 42307 572250
rect 41892 572192 42246 572248
rect 42302 572192 42307 572248
rect 41892 572190 42307 572192
rect 41892 572188 41898 572190
rect 42241 572187 42307 572190
rect 673913 572114 673979 572117
rect 673913 572112 676292 572114
rect 673913 572056 673918 572112
rect 673974 572056 676292 572112
rect 673913 572054 676292 572056
rect 673913 572051 673979 572054
rect 41638 571916 41644 571980
rect 41708 571978 41714 571980
rect 42609 571978 42675 571981
rect 684033 571978 684099 571981
rect 41708 571976 42675 571978
rect 41708 571920 42614 571976
rect 42670 571920 42675 571976
rect 41708 571918 42675 571920
rect 41708 571916 41714 571918
rect 42609 571915 42675 571918
rect 683990 571976 684099 571978
rect 683990 571920 684038 571976
rect 684094 571920 684099 571976
rect 683990 571915 684099 571920
rect 42425 571434 42491 571437
rect 64646 571434 64706 571830
rect 683990 571676 684050 571915
rect 676213 571570 676279 571573
rect 676213 571568 676322 571570
rect 676213 571512 676218 571568
rect 676274 571512 676322 571568
rect 676213 571507 676322 571512
rect 42425 571432 64706 571434
rect 42425 571376 42430 571432
rect 42486 571376 64706 571432
rect 42425 571374 64706 571376
rect 42425 571371 42491 571374
rect 676262 571268 676322 571507
rect 62389 571162 62455 571165
rect 62389 571160 64706 571162
rect 62389 571104 62394 571160
rect 62450 571104 64706 571160
rect 62389 571102 64706 571104
rect 62389 571099 62455 571102
rect 41454 570828 41460 570892
rect 41524 570890 41530 570892
rect 41781 570890 41847 570893
rect 41524 570888 41847 570890
rect 41524 570832 41786 570888
rect 41842 570832 41847 570888
rect 41524 570830 41847 570832
rect 41524 570828 41530 570830
rect 41781 570827 41847 570830
rect 64646 570648 64706 571102
rect 673913 570890 673979 570893
rect 673913 570888 676292 570890
rect 673913 570832 673918 570888
rect 673974 570832 676292 570888
rect 673913 570830 676292 570832
rect 673913 570827 673979 570830
rect 682886 570346 682946 570452
rect 683113 570346 683179 570349
rect 682886 570344 683179 570346
rect 682886 570288 683118 570344
rect 683174 570288 683179 570344
rect 682886 570286 683179 570288
rect 673913 570210 673979 570213
rect 674649 570210 674715 570213
rect 673913 570208 674715 570210
rect 673913 570152 673918 570208
rect 673974 570152 674654 570208
rect 674710 570152 674715 570208
rect 673913 570150 674715 570152
rect 673913 570147 673979 570150
rect 674649 570147 674715 570150
rect 682886 570044 682946 570286
rect 683113 570283 683179 570286
rect 62573 569938 62639 569941
rect 62573 569936 64706 569938
rect 62573 569880 62578 569936
rect 62634 569880 64706 569936
rect 62573 569878 64706 569880
rect 62573 569875 62639 569878
rect 64646 569466 64706 569878
rect 673545 569666 673611 569669
rect 673545 569664 676292 569666
rect 673545 569608 673550 569664
rect 673606 569608 676292 569664
rect 673545 569606 676292 569608
rect 673545 569603 673611 569606
rect 63125 568578 63191 568581
rect 63125 568576 64706 568578
rect 63125 568520 63130 568576
rect 63186 568520 64706 568576
rect 63125 568518 64706 568520
rect 63125 568515 63191 568518
rect 64646 568284 64706 568518
rect 673545 565858 673611 565861
rect 675385 565858 675451 565861
rect 673545 565856 675451 565858
rect 673545 565800 673550 565856
rect 673606 565800 675390 565856
rect 675446 565800 675451 565856
rect 673545 565798 675451 565800
rect 673545 565795 673611 565798
rect 675385 565795 675451 565798
rect 673913 565178 673979 565181
rect 674281 565178 674347 565181
rect 673913 565176 674347 565178
rect 673913 565120 673918 565176
rect 673974 565120 674286 565176
rect 674342 565120 674347 565176
rect 673913 565118 674347 565120
rect 673913 565115 673979 565118
rect 674281 565115 674347 565118
rect 671797 562458 671863 562461
rect 675109 562458 675175 562461
rect 671797 562456 675175 562458
rect 671797 562400 671802 562456
rect 671858 562400 675114 562456
rect 675170 562400 675175 562456
rect 671797 562398 675175 562400
rect 671797 562395 671863 562398
rect 675109 562395 675175 562398
rect 667013 562186 667079 562189
rect 675385 562186 675451 562189
rect 667013 562184 675451 562186
rect 667013 562128 667018 562184
rect 667074 562128 675390 562184
rect 675446 562128 675451 562184
rect 667013 562126 675451 562128
rect 667013 562123 667079 562126
rect 675385 562123 675451 562126
rect 675385 561916 675451 561917
rect 675334 561914 675340 561916
rect 675294 561854 675340 561914
rect 675404 561912 675451 561916
rect 675446 561856 675451 561912
rect 675334 561852 675340 561854
rect 675404 561852 675451 561856
rect 675385 561851 675451 561852
rect 675150 559404 675156 559468
rect 675220 559466 675226 559468
rect 675477 559466 675543 559469
rect 675220 559464 675543 559466
rect 675220 559408 675482 559464
rect 675538 559408 675543 559464
rect 675220 559406 675543 559408
rect 675220 559404 675226 559406
rect 675477 559403 675543 559406
rect 673545 559058 673611 559061
rect 675201 559058 675267 559061
rect 673545 559056 675267 559058
rect 673545 559000 673550 559056
rect 673606 559000 675206 559056
rect 675262 559000 675267 559056
rect 673545 558998 675267 559000
rect 673545 558995 673611 558998
rect 675201 558995 675267 558998
rect 41086 558724 41092 558788
rect 41156 558786 41162 558788
rect 44633 558786 44699 558789
rect 41156 558784 44699 558786
rect 41156 558728 44638 558784
rect 44694 558728 44699 558784
rect 41156 558726 44699 558728
rect 41156 558724 41162 558726
rect 44633 558723 44699 558726
rect 54477 558514 54543 558517
rect 41492 558512 54543 558514
rect 41492 558456 54482 558512
rect 54538 558456 54543 558512
rect 41492 558454 54543 558456
rect 54477 558451 54543 558454
rect 41137 558106 41203 558109
rect 41124 558104 41203 558106
rect 41124 558048 41142 558104
rect 41198 558048 41203 558104
rect 41124 558046 41203 558048
rect 41137 558043 41203 558046
rect 41086 557488 41092 557552
rect 41156 557488 41162 557552
rect 41278 557550 41338 557668
rect 41278 557490 41890 557550
rect 41094 557260 41154 557488
rect 41830 557426 41890 557490
rect 41830 557366 51090 557426
rect 44541 556882 44607 556885
rect 41492 556880 44607 556882
rect 41492 556824 44546 556880
rect 44602 556824 44607 556880
rect 41492 556822 44607 556824
rect 44541 556819 44607 556822
rect 51030 556746 51090 557366
rect 62205 556746 62271 556749
rect 51030 556744 62271 556746
rect 51030 556688 62210 556744
rect 62266 556688 62271 556744
rect 51030 556686 62271 556688
rect 62205 556683 62271 556686
rect 43069 556474 43135 556477
rect 41492 556472 43135 556474
rect 41492 556416 43074 556472
rect 43130 556416 43135 556472
rect 41492 556414 43135 556416
rect 43069 556411 43135 556414
rect 44725 556066 44791 556069
rect 41492 556064 44791 556066
rect 41492 556008 44730 556064
rect 44786 556008 44791 556064
rect 41492 556006 44791 556008
rect 44725 556003 44791 556006
rect 44909 555658 44975 555661
rect 41492 555656 44975 555658
rect 41492 555600 44914 555656
rect 44970 555600 44975 555656
rect 41492 555598 44975 555600
rect 44909 555595 44975 555598
rect 674925 555524 674991 555525
rect 674925 555522 674972 555524
rect 674880 555520 674972 555522
rect 674880 555464 674930 555520
rect 674880 555462 674972 555464
rect 674925 555460 674972 555462
rect 675036 555460 675042 555524
rect 674925 555459 674991 555460
rect 45829 555250 45895 555253
rect 41492 555248 45895 555250
rect 41492 555192 45834 555248
rect 45890 555192 45895 555248
rect 41492 555190 45895 555192
rect 45829 555187 45895 555190
rect 672257 555250 672323 555253
rect 675385 555250 675451 555253
rect 672257 555248 675451 555250
rect 672257 555192 672262 555248
rect 672318 555192 675390 555248
rect 675446 555192 675451 555248
rect 672257 555190 675451 555192
rect 672257 555187 672323 555190
rect 675385 555187 675451 555190
rect 42793 554842 42859 554845
rect 41492 554840 42859 554842
rect 41492 554784 42798 554840
rect 42854 554784 42859 554840
rect 41492 554782 42859 554784
rect 42793 554779 42859 554782
rect 668393 554706 668459 554709
rect 675109 554706 675175 554709
rect 668393 554704 675175 554706
rect 668393 554648 668398 554704
rect 668454 554648 675114 554704
rect 675170 554648 675175 554704
rect 668393 554646 675175 554648
rect 668393 554643 668459 554646
rect 675109 554643 675175 554646
rect 45645 554434 45711 554437
rect 41492 554432 45711 554434
rect 41492 554376 45650 554432
rect 45706 554376 45711 554432
rect 41492 554374 45711 554376
rect 45645 554371 45711 554374
rect 674005 554434 674071 554437
rect 675293 554434 675359 554437
rect 674005 554432 675359 554434
rect 674005 554376 674010 554432
rect 674066 554376 675298 554432
rect 675354 554376 675359 554432
rect 674005 554374 675359 554376
rect 674005 554371 674071 554374
rect 675293 554371 675359 554374
rect 42190 554026 42196 554028
rect 41492 553966 42196 554026
rect 42190 553964 42196 553966
rect 42260 553964 42266 554028
rect 675753 554026 675819 554029
rect 676438 554026 676444 554028
rect 675753 554024 676444 554026
rect 675753 553968 675758 554024
rect 675814 553968 676444 554024
rect 675753 553966 676444 553968
rect 675753 553963 675819 553966
rect 676438 553964 676444 553966
rect 676508 553964 676514 554028
rect 39990 553413 40050 553588
rect 649950 553482 650010 553914
rect 667565 553890 667631 553893
rect 675477 553890 675543 553893
rect 667565 553888 675543 553890
rect 667565 553832 667570 553888
rect 667626 553832 675482 553888
rect 675538 553832 675543 553888
rect 667565 553830 675543 553832
rect 667565 553827 667631 553830
rect 675477 553827 675543 553830
rect 651465 553482 651531 553485
rect 649950 553480 651531 553482
rect 649950 553424 651470 553480
rect 651526 553424 651531 553480
rect 649950 553422 651531 553424
rect 651465 553419 651531 553422
rect 674005 553482 674071 553485
rect 675109 553482 675175 553485
rect 674005 553480 675175 553482
rect 674005 553424 674010 553480
rect 674066 553424 675114 553480
rect 675170 553424 675175 553480
rect 674005 553422 675175 553424
rect 674005 553419 674071 553422
rect 675109 553419 675175 553422
rect 39990 553408 40099 553413
rect 39990 553352 40038 553408
rect 40094 553352 40099 553408
rect 39990 553350 40099 553352
rect 40033 553347 40099 553350
rect 41362 553348 41368 553412
rect 41432 553348 41438 553412
rect 41370 553210 41430 553348
rect 41370 553150 41492 553210
rect 41321 552802 41387 552805
rect 41308 552800 41387 552802
rect 41308 552744 41326 552800
rect 41382 552744 41387 552800
rect 41308 552742 41387 552744
rect 41321 552739 41387 552742
rect 37917 552394 37983 552397
rect 37917 552392 37996 552394
rect 37917 552336 37922 552392
rect 37978 552336 37996 552392
rect 37917 552334 37996 552336
rect 37917 552331 37983 552334
rect 649950 552122 650010 552732
rect 652017 552122 652083 552125
rect 649950 552120 652083 552122
rect 649950 552064 652022 552120
rect 652078 552064 652083 552120
rect 649950 552062 652083 552064
rect 652017 552059 652083 552062
rect 675753 552122 675819 552125
rect 676990 552122 676996 552124
rect 675753 552120 676996 552122
rect 675753 552064 675758 552120
rect 675814 552064 676996 552120
rect 675753 552062 676996 552064
rect 675753 552059 675819 552062
rect 676990 552060 676996 552062
rect 677060 552060 677066 552124
rect 29637 551986 29703 551989
rect 29637 551984 29716 551986
rect 29637 551928 29642 551984
rect 29698 551928 29716 551984
rect 29637 551926 29716 551928
rect 29637 551923 29703 551926
rect 41689 551850 41755 551853
rect 42374 551850 42380 551852
rect 41689 551848 42380 551850
rect 41689 551792 41694 551848
rect 41750 551792 42380 551848
rect 41689 551790 42380 551792
rect 41689 551787 41755 551790
rect 42374 551788 42380 551790
rect 42444 551788 42450 551852
rect 673913 551850 673979 551853
rect 674741 551850 674807 551853
rect 673913 551848 674807 551850
rect 673913 551792 673918 551848
rect 673974 551792 674746 551848
rect 674802 551792 674807 551848
rect 673913 551790 674807 551792
rect 673913 551787 673979 551790
rect 674741 551787 674807 551790
rect 44357 551578 44423 551581
rect 41492 551576 44423 551578
rect 41492 551520 44362 551576
rect 44418 551520 44423 551576
rect 41492 551518 44423 551520
rect 44357 551515 44423 551518
rect 42793 551170 42859 551173
rect 41492 551168 42859 551170
rect 41492 551112 42798 551168
rect 42854 551112 42859 551168
rect 41492 551110 42859 551112
rect 649950 551170 650010 551550
rect 651465 551170 651531 551173
rect 649950 551168 651531 551170
rect 649950 551112 651470 551168
rect 651526 551112 651531 551168
rect 649950 551110 651531 551112
rect 42793 551107 42859 551110
rect 651465 551107 651531 551110
rect 45093 550762 45159 550765
rect 41492 550760 45159 550762
rect 41492 550704 45098 550760
rect 45154 550704 45159 550760
rect 41492 550702 45159 550704
rect 45093 550699 45159 550702
rect 675150 550428 675156 550492
rect 675220 550490 675226 550492
rect 675385 550490 675451 550493
rect 675220 550488 675451 550490
rect 675220 550432 675390 550488
rect 675446 550432 675451 550488
rect 675220 550430 675451 550432
rect 675220 550428 675226 550430
rect 675385 550427 675451 550430
rect 41965 550354 42031 550357
rect 41492 550352 42031 550354
rect 41492 550296 41970 550352
rect 42026 550296 42031 550352
rect 41492 550294 42031 550296
rect 649950 550354 650010 550368
rect 651373 550354 651439 550357
rect 649950 550352 651439 550354
rect 649950 550296 651378 550352
rect 651434 550296 651439 550352
rect 649950 550294 651439 550296
rect 41965 550291 42031 550294
rect 651373 550291 651439 550294
rect 42149 550218 42215 550221
rect 62665 550218 62731 550221
rect 42149 550216 62731 550218
rect 42149 550160 42154 550216
rect 42210 550160 62670 550216
rect 62726 550160 62731 550216
rect 42149 550158 62731 550160
rect 42149 550155 42215 550158
rect 62665 550155 62731 550158
rect 41781 549946 41847 549949
rect 41492 549944 41847 549946
rect 41492 549888 41786 549944
rect 41842 549888 41847 549944
rect 41492 549886 41847 549888
rect 41781 549883 41847 549886
rect 670417 549810 670483 549813
rect 675293 549810 675359 549813
rect 670417 549808 675359 549810
rect 670417 549752 670422 549808
rect 670478 549752 675298 549808
rect 675354 549752 675359 549808
rect 670417 549750 675359 549752
rect 670417 549747 670483 549750
rect 675293 549747 675359 549750
rect 42977 549538 43043 549541
rect 41492 549536 43043 549538
rect 41492 549480 42982 549536
rect 43038 549480 43043 549536
rect 41492 549478 43043 549480
rect 42977 549475 43043 549478
rect 674966 549476 674972 549540
rect 675036 549538 675042 549540
rect 675293 549538 675359 549541
rect 675036 549536 675359 549538
rect 675036 549480 675298 549536
rect 675354 549480 675359 549536
rect 675036 549478 675359 549480
rect 675036 549476 675042 549478
rect 675293 549475 675359 549478
rect 651465 549266 651531 549269
rect 649950 549264 651531 549266
rect 649950 549208 651470 549264
rect 651526 549208 651531 549264
rect 649950 549206 651531 549208
rect 649950 549186 650010 549206
rect 651465 549203 651531 549206
rect 44173 549130 44239 549133
rect 41492 549128 44239 549130
rect 41492 549072 44178 549128
rect 44234 549072 44239 549128
rect 41492 549070 44239 549072
rect 44173 549067 44239 549070
rect 45277 548722 45343 548725
rect 41492 548720 45343 548722
rect 41492 548664 45282 548720
rect 45338 548664 45343 548720
rect 41492 548662 45343 548664
rect 45277 548659 45343 548662
rect 651465 548450 651531 548453
rect 649950 548448 651531 548450
rect 649950 548392 651470 548448
rect 651526 548392 651531 548448
rect 649950 548390 651531 548392
rect 43805 548314 43871 548317
rect 41492 548312 43871 548314
rect 41492 548256 43810 548312
rect 43866 548256 43871 548312
rect 41492 548254 43871 548256
rect 43805 548251 43871 548254
rect 649950 548004 650010 548390
rect 651465 548387 651531 548390
rect 674833 548450 674899 548453
rect 675334 548450 675340 548452
rect 674833 548448 675340 548450
rect 674833 548392 674838 548448
rect 674894 548392 675340 548448
rect 674833 548390 675340 548392
rect 674833 548387 674899 548390
rect 675334 548388 675340 548390
rect 675404 548388 675410 548452
rect 675753 548314 675819 548317
rect 676806 548314 676812 548316
rect 675753 548312 676812 548314
rect 675753 548256 675758 548312
rect 675814 548256 676812 548312
rect 675753 548254 676812 548256
rect 675753 548251 675819 548254
rect 676806 548252 676812 548254
rect 676876 548252 676882 548316
rect 41462 547498 41522 547876
rect 676438 547572 676444 547636
rect 676508 547634 676514 547636
rect 677409 547634 677475 547637
rect 676508 547632 677475 547634
rect 676508 547576 677414 547632
rect 677470 547576 677475 547632
rect 676508 547574 677475 547576
rect 676508 547572 676514 547574
rect 677409 547571 677475 547574
rect 47577 547498 47643 547501
rect 41462 547496 47643 547498
rect 41462 547468 47582 547496
rect 41492 547440 47582 547468
rect 47638 547440 47643 547496
rect 41492 547438 47643 547440
rect 47577 547435 47643 547438
rect 674230 547300 674236 547364
rect 674300 547362 674306 547364
rect 683389 547362 683455 547365
rect 674300 547360 683455 547362
rect 674300 547304 683394 547360
rect 683450 547304 683455 547360
rect 674300 547302 683455 547304
rect 674300 547300 674306 547302
rect 683389 547299 683455 547302
rect 43989 547090 44055 547093
rect 41492 547088 44055 547090
rect 41492 547032 43994 547088
rect 44050 547032 44055 547088
rect 41492 547030 44055 547032
rect 43989 547027 44055 547030
rect 675886 547028 675892 547092
rect 675956 547090 675962 547092
rect 680997 547090 681063 547093
rect 675956 547088 681063 547090
rect 675956 547032 681002 547088
rect 681058 547032 681063 547088
rect 675956 547030 681063 547032
rect 675956 547028 675962 547030
rect 680997 547027 681063 547030
rect 676070 546756 676076 546820
rect 676140 546818 676146 546820
rect 679617 546818 679683 546821
rect 676140 546816 679683 546818
rect 676140 546760 679622 546816
rect 679678 546760 679683 546816
rect 676140 546758 679683 546760
rect 676140 546756 676146 546758
rect 679617 546755 679683 546758
rect 41638 546348 41644 546412
rect 41708 546410 41714 546412
rect 42374 546410 42380 546412
rect 41708 546350 42380 546410
rect 41708 546348 41714 546350
rect 42374 546348 42380 546350
rect 42444 546348 42450 546412
rect 40902 545668 40908 545732
rect 40972 545730 40978 545732
rect 41965 545730 42031 545733
rect 40972 545728 42031 545730
rect 40972 545672 41970 545728
rect 42026 545672 42031 545728
rect 40972 545670 42031 545672
rect 40972 545668 40978 545670
rect 41965 545667 42031 545670
rect 40718 545396 40724 545460
rect 40788 545458 40794 545460
rect 41781 545458 41847 545461
rect 40788 545456 41847 545458
rect 40788 545400 41786 545456
rect 41842 545400 41847 545456
rect 40788 545398 41847 545400
rect 40788 545396 40794 545398
rect 41781 545395 41847 545398
rect 37917 542330 37983 542333
rect 41454 542330 41460 542332
rect 37917 542328 41460 542330
rect 37917 542272 37922 542328
rect 37978 542272 41460 542328
rect 37917 542270 41460 542272
rect 37917 542267 37983 542270
rect 41454 542268 41460 542270
rect 41524 542268 41530 542332
rect 675201 541244 675267 541245
rect 675150 541242 675156 541244
rect 675110 541182 675156 541242
rect 675220 541240 675267 541244
rect 675262 541184 675267 541240
rect 675150 541180 675156 541182
rect 675220 541180 675267 541184
rect 675201 541179 675267 541180
rect 42425 539610 42491 539613
rect 53097 539610 53163 539613
rect 675109 539612 675175 539613
rect 675109 539610 675156 539612
rect 42425 539608 53163 539610
rect 42425 539552 42430 539608
rect 42486 539552 53102 539608
rect 53158 539552 53163 539608
rect 42425 539550 53163 539552
rect 675064 539608 675156 539610
rect 675064 539552 675114 539608
rect 675064 539550 675156 539552
rect 42425 539547 42491 539550
rect 53097 539547 53163 539550
rect 675109 539548 675156 539550
rect 675220 539548 675226 539612
rect 675109 539547 675175 539548
rect 42517 537570 42583 537573
rect 44173 537570 44239 537573
rect 42517 537568 44239 537570
rect 42517 537512 42522 537568
rect 42578 537512 44178 537568
rect 44234 537512 44239 537568
rect 42517 537510 44239 537512
rect 42517 537507 42583 537510
rect 44173 537507 44239 537510
rect 40718 537236 40724 537300
rect 40788 537298 40794 537300
rect 42333 537298 42399 537301
rect 40788 537296 42399 537298
rect 40788 537240 42338 537296
rect 42394 537240 42399 537296
rect 40788 537238 42399 537240
rect 40788 537236 40794 537238
rect 42333 537235 42399 537238
rect 40902 536964 40908 537028
rect 40972 537026 40978 537028
rect 41781 537026 41847 537029
rect 40972 537024 41847 537026
rect 40972 536968 41786 537024
rect 41842 536968 41847 537024
rect 40972 536966 41847 536968
rect 40972 536964 40978 536966
rect 41781 536963 41847 536966
rect 673729 536346 673795 536349
rect 674281 536346 674347 536349
rect 673729 536344 674347 536346
rect 673729 536288 673734 536344
rect 673790 536288 674286 536344
rect 674342 536288 674347 536344
rect 673729 536286 674347 536288
rect 673729 536283 673795 536286
rect 674281 536283 674347 536286
rect 673729 536074 673795 536077
rect 676262 536074 676322 536112
rect 673729 536072 676322 536074
rect 673729 536016 673734 536072
rect 673790 536016 676322 536072
rect 673729 536014 676322 536016
rect 673729 536011 673795 536014
rect 42057 535802 42123 535805
rect 44725 535802 44791 535805
rect 42057 535800 44791 535802
rect 42057 535744 42062 535800
rect 42118 535744 44730 535800
rect 44786 535744 44791 535800
rect 42057 535742 44791 535744
rect 42057 535739 42123 535742
rect 44725 535739 44791 535742
rect 673729 535802 673795 535805
rect 673729 535800 676322 535802
rect 673729 535744 673734 535800
rect 673790 535744 676322 535800
rect 673729 535742 676322 535744
rect 673729 535739 673795 535742
rect 676262 535704 676322 535742
rect 42149 535530 42215 535533
rect 45277 535530 45343 535533
rect 42149 535528 45343 535530
rect 42149 535472 42154 535528
rect 42210 535472 45282 535528
rect 45338 535472 45343 535528
rect 42149 535470 45343 535472
rect 42149 535467 42215 535470
rect 45277 535467 45343 535470
rect 673729 535258 673795 535261
rect 676262 535258 676322 535296
rect 673729 535256 676322 535258
rect 673729 535200 673734 535256
rect 673790 535200 676322 535256
rect 673729 535198 676322 535200
rect 673729 535195 673795 535198
rect 672625 534986 672691 534989
rect 672625 534984 676322 534986
rect 672625 534928 672630 534984
rect 672686 534928 676322 534984
rect 672625 534926 676322 534928
rect 672625 534923 672691 534926
rect 676262 534888 676322 534926
rect 676262 534309 676322 534480
rect 676213 534304 676322 534309
rect 676213 534248 676218 534304
rect 676274 534248 676322 534304
rect 676213 534246 676322 534248
rect 676213 534243 676279 534246
rect 672625 534170 672691 534173
rect 672625 534168 675770 534170
rect 672625 534112 672630 534168
rect 672686 534112 675770 534168
rect 672625 534110 675770 534112
rect 672625 534107 672691 534110
rect 675710 534102 675770 534110
rect 675710 534042 676292 534102
rect 42425 533898 42491 533901
rect 45093 533898 45159 533901
rect 42425 533896 45159 533898
rect 42425 533840 42430 533896
rect 42486 533840 45098 533896
rect 45154 533840 45159 533896
rect 42425 533838 45159 533840
rect 42425 533835 42491 533838
rect 45093 533835 45159 533838
rect 670785 533898 670851 533901
rect 674281 533898 674347 533901
rect 670785 533896 674347 533898
rect 670785 533840 670790 533896
rect 670846 533840 674286 533896
rect 674342 533840 674347 533896
rect 670785 533838 674347 533840
rect 670785 533835 670851 533838
rect 674281 533835 674347 533838
rect 41454 533700 41460 533764
rect 41524 533762 41530 533764
rect 41781 533762 41847 533765
rect 41524 533760 41847 533762
rect 41524 533704 41786 533760
rect 41842 533704 41847 533760
rect 41524 533702 41847 533704
rect 41524 533700 41530 533702
rect 41781 533699 41847 533702
rect 676029 533694 676095 533697
rect 676029 533692 676292 533694
rect 676029 533636 676034 533692
rect 676090 533636 676292 533692
rect 676029 533634 676292 533636
rect 676029 533631 676095 533634
rect 672625 533354 672691 533357
rect 672625 533352 676322 533354
rect 672625 533296 672630 533352
rect 672686 533296 676322 533352
rect 672625 533294 676322 533296
rect 672625 533291 672691 533294
rect 676262 533256 676322 533294
rect 671521 533082 671587 533085
rect 671521 533080 676322 533082
rect 671521 533024 671526 533080
rect 671582 533024 676322 533080
rect 671521 533022 676322 533024
rect 671521 533019 671587 533022
rect 40534 532884 40540 532948
rect 40604 532946 40610 532948
rect 42609 532946 42675 532949
rect 40604 532944 42675 532946
rect 40604 532888 42614 532944
rect 42670 532888 42675 532944
rect 40604 532886 42675 532888
rect 40604 532884 40610 532886
rect 42609 532883 42675 532886
rect 676262 532848 676322 533022
rect 672533 532810 672599 532813
rect 674281 532810 674347 532813
rect 672533 532808 674347 532810
rect 672533 532752 672538 532808
rect 672594 532752 674286 532808
rect 674342 532752 674347 532808
rect 672533 532750 674347 532752
rect 672533 532747 672599 532750
rect 674281 532747 674347 532750
rect 671337 532266 671403 532269
rect 676262 532266 676322 532440
rect 671337 532264 676322 532266
rect 671337 532208 671342 532264
rect 671398 532208 676322 532264
rect 671337 532206 676322 532208
rect 671337 532203 671403 532206
rect 676262 531858 676322 532032
rect 673686 531798 676322 531858
rect 680997 531858 681063 531861
rect 680997 531856 681106 531858
rect 680997 531800 681002 531856
rect 681058 531800 681106 531856
rect 671337 531586 671403 531589
rect 673686 531586 673746 531798
rect 680997 531795 681106 531800
rect 681046 531624 681106 531795
rect 671337 531584 673746 531586
rect 671337 531528 671342 531584
rect 671398 531528 673746 531584
rect 671337 531526 673746 531528
rect 671337 531523 671403 531526
rect 682377 531450 682443 531453
rect 682334 531448 682443 531450
rect 682334 531392 682382 531448
rect 682438 531392 682443 531448
rect 682334 531387 682443 531392
rect 682334 531216 682394 531387
rect 62113 531178 62179 531181
rect 62113 531176 64706 531178
rect 62113 531120 62118 531176
rect 62174 531120 64706 531176
rect 62113 531118 64706 531120
rect 62113 531115 62179 531118
rect 673729 530770 673795 530773
rect 676262 530770 676322 530808
rect 673729 530768 676322 530770
rect 673729 530712 673734 530768
rect 673790 530712 676322 530768
rect 673729 530710 676322 530712
rect 673729 530707 673795 530710
rect 62297 530634 62363 530637
rect 679617 530634 679683 530637
rect 62297 530632 64706 530634
rect 62297 530576 62302 530632
rect 62358 530576 64706 530632
rect 62297 530574 64706 530576
rect 62297 530571 62363 530574
rect 42057 530226 42123 530229
rect 42701 530226 42767 530229
rect 42057 530224 42767 530226
rect 42057 530168 42062 530224
rect 42118 530168 42706 530224
rect 42762 530168 42767 530224
rect 42057 530166 42767 530168
rect 42057 530163 42123 530166
rect 42701 530163 42767 530166
rect 64646 529990 64706 530574
rect 679574 530632 679683 530634
rect 679574 530576 679622 530632
rect 679678 530576 679683 530632
rect 679574 530571 679683 530576
rect 679574 530400 679634 530571
rect 41822 529892 41828 529956
rect 41892 529954 41898 529956
rect 42333 529954 42399 529957
rect 41892 529952 42399 529954
rect 41892 529896 42338 529952
rect 42394 529896 42399 529952
rect 41892 529894 42399 529896
rect 41892 529892 41898 529894
rect 42333 529891 42399 529894
rect 673729 529954 673795 529957
rect 676262 529954 676322 529992
rect 673729 529952 676322 529954
rect 673729 529896 673734 529952
rect 673790 529896 676322 529952
rect 673729 529894 676322 529896
rect 673729 529891 673795 529894
rect 673729 529546 673795 529549
rect 676262 529546 676322 529584
rect 673729 529544 676322 529546
rect 673729 529488 673734 529544
rect 673790 529488 676322 529544
rect 673729 529486 676322 529488
rect 673729 529483 673795 529486
rect 41873 529412 41939 529413
rect 41822 529410 41828 529412
rect 41782 529350 41828 529410
rect 41892 529408 41939 529412
rect 41934 529352 41939 529408
rect 41822 529348 41828 529350
rect 41892 529348 41939 529352
rect 41873 529347 41939 529348
rect 673729 529274 673795 529277
rect 673729 529272 676322 529274
rect 673729 529216 673734 529272
rect 673790 529216 676322 529272
rect 673729 529214 676322 529216
rect 673729 529211 673795 529214
rect 676262 529176 676322 529214
rect 42425 529002 42491 529005
rect 44357 529002 44423 529005
rect 42425 529000 44423 529002
rect 42425 528944 42430 529000
rect 42486 528944 44362 529000
rect 44418 528944 44423 529000
rect 42425 528942 44423 528944
rect 42425 528939 42491 528942
rect 44357 528939 44423 528942
rect 673729 528866 673795 528869
rect 673729 528864 676322 528866
rect 673729 528808 673734 528864
rect 673790 528808 676322 528864
rect 62113 528594 62179 528597
rect 64646 528594 64706 528808
rect 673729 528806 676322 528808
rect 673729 528803 673795 528806
rect 676262 528768 676322 528806
rect 62113 528592 64706 528594
rect 62113 528536 62118 528592
rect 62174 528536 64706 528592
rect 62113 528534 64706 528536
rect 62113 528531 62179 528534
rect 676262 528189 676322 528360
rect 676213 528184 676322 528189
rect 676213 528128 676218 528184
rect 676274 528128 676322 528184
rect 676213 528126 676322 528128
rect 683205 528186 683271 528189
rect 683205 528184 683314 528186
rect 683205 528128 683210 528184
rect 683266 528128 683314 528184
rect 676213 528123 676279 528126
rect 683205 528123 683314 528128
rect 62481 528050 62547 528053
rect 62481 528048 64706 528050
rect 62481 527992 62486 528048
rect 62542 527992 64706 528048
rect 62481 527990 64706 527992
rect 62481 527987 62547 527990
rect 64646 527626 64706 527990
rect 683254 527952 683314 528123
rect 683573 527778 683639 527781
rect 683573 527776 683682 527778
rect 683573 527720 683578 527776
rect 683634 527720 683682 527776
rect 683573 527715 683682 527720
rect 683622 527544 683682 527715
rect 683389 527370 683455 527373
rect 683389 527368 683498 527370
rect 683389 527312 683394 527368
rect 683450 527312 683498 527368
rect 683389 527307 683498 527312
rect 42701 527234 42767 527237
rect 45093 527234 45159 527237
rect 42701 527232 45159 527234
rect 42701 527176 42706 527232
rect 42762 527176 45098 527232
rect 45154 527176 45159 527232
rect 42701 527174 45159 527176
rect 42701 527171 42767 527174
rect 45093 527171 45159 527174
rect 673177 527234 673243 527237
rect 674373 527234 674439 527237
rect 673177 527232 674439 527234
rect 673177 527176 673182 527232
rect 673238 527176 674378 527232
rect 674434 527176 674439 527232
rect 673177 527174 674439 527176
rect 673177 527171 673243 527174
rect 674373 527171 674439 527174
rect 683438 527136 683498 527307
rect 62113 527098 62179 527101
rect 62113 527096 64706 527098
rect 62113 527040 62118 527096
rect 62174 527040 64706 527096
rect 62113 527038 64706 527040
rect 62113 527035 62179 527038
rect 64646 526444 64706 527038
rect 676029 526758 676095 526761
rect 676029 526756 676292 526758
rect 676029 526700 676034 526756
rect 676090 526700 676292 526756
rect 676029 526698 676292 526700
rect 676029 526695 676095 526698
rect 676029 526350 676095 526353
rect 676029 526348 676292 526350
rect 676029 526292 676034 526348
rect 676090 526292 676292 526348
rect 676029 526290 676292 526292
rect 676029 526287 676095 526290
rect 679022 525741 679082 525912
rect 62665 525738 62731 525741
rect 62665 525736 64706 525738
rect 62665 525680 62670 525736
rect 62726 525680 64706 525736
rect 62665 525678 64706 525680
rect 62665 525675 62731 525678
rect 64646 525262 64706 525678
rect 678973 525736 679082 525741
rect 678973 525680 678978 525736
rect 679034 525680 679082 525736
rect 678973 525678 679082 525680
rect 678973 525675 679039 525678
rect 683070 524925 683130 525504
rect 683070 524920 683179 524925
rect 683070 524864 683118 524920
rect 683174 524864 683179 524920
rect 683070 524862 683179 524864
rect 683113 524859 683179 524862
rect 680310 524517 680370 524688
rect 680310 524512 680419 524517
rect 680310 524456 680358 524512
rect 680414 524456 680419 524512
rect 680310 524454 680419 524456
rect 680353 524451 680419 524454
rect 676806 503644 676812 503708
rect 676876 503706 676882 503708
rect 683205 503706 683271 503709
rect 676876 503704 683271 503706
rect 676876 503648 683210 503704
rect 683266 503648 683271 503704
rect 676876 503646 683271 503648
rect 676876 503644 676882 503646
rect 683205 503643 683271 503646
rect 673177 492146 673243 492149
rect 673177 492144 676292 492146
rect 673177 492088 673182 492144
rect 673238 492088 676292 492144
rect 673177 492086 676292 492088
rect 673177 492083 673243 492086
rect 676029 491738 676095 491741
rect 676029 491736 676292 491738
rect 676029 491680 676034 491736
rect 676090 491680 676292 491736
rect 676029 491678 676292 491680
rect 676029 491675 676095 491678
rect 673821 491330 673887 491333
rect 673821 491328 676292 491330
rect 673821 491272 673826 491328
rect 673882 491272 676292 491328
rect 673821 491270 676292 491272
rect 673821 491267 673887 491270
rect 674005 490922 674071 490925
rect 674005 490920 676292 490922
rect 674005 490864 674010 490920
rect 674066 490864 676292 490920
rect 674005 490862 676292 490864
rect 674005 490859 674071 490862
rect 673177 490514 673243 490517
rect 673177 490512 676292 490514
rect 673177 490456 673182 490512
rect 673238 490456 676292 490512
rect 673177 490454 676292 490456
rect 673177 490451 673243 490454
rect 674005 490106 674071 490109
rect 674005 490104 676292 490106
rect 674005 490048 674010 490104
rect 674066 490048 676292 490104
rect 674005 490046 676292 490048
rect 674005 490043 674071 490046
rect 674005 489698 674071 489701
rect 674005 489696 676292 489698
rect 674005 489640 674010 489696
rect 674066 489640 676292 489696
rect 674005 489638 676292 489640
rect 674005 489635 674071 489638
rect 674005 489290 674071 489293
rect 674005 489288 676292 489290
rect 674005 489232 674010 489288
rect 674066 489232 676292 489288
rect 674005 489230 676292 489232
rect 674005 489227 674071 489230
rect 676029 488882 676095 488885
rect 676029 488880 676292 488882
rect 676029 488824 676034 488880
rect 676090 488824 676292 488880
rect 676029 488822 676292 488824
rect 676029 488819 676095 488822
rect 674005 488474 674071 488477
rect 674005 488472 676292 488474
rect 674005 488416 674010 488472
rect 674066 488416 676292 488472
rect 674005 488414 676292 488416
rect 674005 488411 674071 488414
rect 675702 488004 675708 488068
rect 675772 488066 675778 488068
rect 675772 488006 676292 488066
rect 675772 488004 675778 488006
rect 678237 487658 678303 487661
rect 678237 487656 678316 487658
rect 678237 487600 678242 487656
rect 678298 487600 678316 487656
rect 678237 487598 678316 487600
rect 678237 487595 678303 487598
rect 679617 487250 679683 487253
rect 679604 487248 679683 487250
rect 679604 487192 679622 487248
rect 679678 487192 679683 487248
rect 679604 487190 679683 487192
rect 679617 487187 679683 487190
rect 674005 486842 674071 486845
rect 674005 486840 676292 486842
rect 674005 486784 674010 486840
rect 674066 486784 676292 486840
rect 674005 486782 676292 486784
rect 674005 486779 674071 486782
rect 680997 486434 681063 486437
rect 680997 486432 681076 486434
rect 680997 486376 681002 486432
rect 681058 486376 681076 486432
rect 680997 486374 681076 486376
rect 680997 486371 681063 486374
rect 674005 486026 674071 486029
rect 674005 486024 676292 486026
rect 674005 485968 674010 486024
rect 674066 485968 676292 486024
rect 674005 485966 676292 485968
rect 674005 485963 674071 485966
rect 683205 485618 683271 485621
rect 683205 485616 683284 485618
rect 683205 485560 683210 485616
rect 683266 485560 683284 485616
rect 683205 485558 683284 485560
rect 683205 485555 683271 485558
rect 676029 485210 676095 485213
rect 676029 485208 676292 485210
rect 676029 485152 676034 485208
rect 676090 485152 676292 485208
rect 676029 485150 676292 485152
rect 676029 485147 676095 485150
rect 673545 484802 673611 484805
rect 673545 484800 676292 484802
rect 673545 484744 673550 484800
rect 673606 484744 676292 484800
rect 673545 484742 676292 484744
rect 673545 484739 673611 484742
rect 674649 484394 674715 484397
rect 674649 484392 676292 484394
rect 674649 484336 674654 484392
rect 674710 484336 676292 484392
rect 674649 484334 676292 484336
rect 674649 484331 674715 484334
rect 675886 483924 675892 483988
rect 675956 483986 675962 483988
rect 675956 483926 676292 483986
rect 675956 483924 675962 483926
rect 676029 483578 676095 483581
rect 676029 483576 676292 483578
rect 676029 483520 676034 483576
rect 676090 483520 676292 483576
rect 676029 483518 676292 483520
rect 676029 483515 676095 483518
rect 675845 483170 675911 483173
rect 675845 483168 676292 483170
rect 675845 483112 675850 483168
rect 675906 483112 676292 483168
rect 675845 483110 676292 483112
rect 675845 483107 675911 483110
rect 676029 482762 676095 482765
rect 676029 482760 676292 482762
rect 676029 482704 676034 482760
rect 676090 482704 676292 482760
rect 676029 482702 676292 482704
rect 676029 482699 676095 482702
rect 677133 482526 677199 482527
rect 677133 482522 677180 482526
rect 677244 482524 677250 482526
rect 677133 482466 677138 482522
rect 677133 482462 677180 482466
rect 677244 482464 677290 482524
rect 677244 482462 677250 482464
rect 677133 482461 677199 482462
rect 676029 482354 676095 482357
rect 676029 482352 676292 482354
rect 676029 482296 676034 482352
rect 676090 482296 676292 482352
rect 676029 482294 676292 482296
rect 676029 482291 676095 482294
rect 680353 481946 680419 481949
rect 680340 481944 680419 481946
rect 680340 481888 680358 481944
rect 680414 481888 680419 481944
rect 680340 481886 680419 481888
rect 680353 481883 680419 481886
rect 677182 481130 677242 481508
rect 683113 481130 683179 481133
rect 677182 481128 683179 481130
rect 677182 481100 683118 481128
rect 677212 481072 683118 481100
rect 683174 481072 683179 481128
rect 677212 481070 683179 481072
rect 683113 481067 683179 481070
rect 675845 480722 675911 480725
rect 675845 480720 676292 480722
rect 675845 480664 675850 480720
rect 675906 480664 676292 480720
rect 675845 480662 676292 480664
rect 675845 480659 675911 480662
rect 669773 455426 669839 455429
rect 673269 455426 673335 455429
rect 669773 455424 673335 455426
rect 669773 455368 669778 455424
rect 669834 455368 673274 455424
rect 673330 455368 673335 455424
rect 669773 455366 673335 455368
rect 669773 455363 669839 455366
rect 673269 455363 673335 455366
rect 673381 455290 673447 455293
rect 673862 455290 673868 455292
rect 673381 455288 673868 455290
rect 673381 455232 673386 455288
rect 673442 455232 673868 455288
rect 673381 455230 673868 455232
rect 673381 455227 673447 455230
rect 673862 455228 673868 455230
rect 673932 455228 673938 455292
rect 670601 455018 670667 455021
rect 673499 455018 673565 455021
rect 670601 455016 673565 455018
rect 670601 454960 670606 455016
rect 670662 454960 673504 455016
rect 673560 454960 673565 455016
rect 670601 454958 673565 454960
rect 670601 454955 670667 454958
rect 673499 454955 673565 454958
rect 673039 454746 673105 454749
rect 674281 454746 674347 454749
rect 673039 454744 674347 454746
rect 673039 454688 673044 454744
rect 673100 454688 674286 454744
rect 674342 454688 674347 454744
rect 673039 454686 674347 454688
rect 673039 454683 673105 454686
rect 674281 454683 674347 454686
rect 672947 454474 673013 454477
rect 674281 454474 674347 454477
rect 672947 454472 674347 454474
rect 672947 454416 672952 454472
rect 673008 454416 674286 454472
rect 674342 454416 674347 454472
rect 672947 454414 674347 454416
rect 672947 454411 673013 454414
rect 674281 454411 674347 454414
rect 672809 454202 672875 454205
rect 674281 454202 674347 454205
rect 672809 454200 674347 454202
rect 672809 454144 672814 454200
rect 672870 454144 674286 454200
rect 674342 454144 674347 454200
rect 672809 454142 674347 454144
rect 672809 454139 672875 454142
rect 674281 454139 674347 454142
rect 672257 453930 672323 453933
rect 674281 453930 674347 453933
rect 672257 453928 674347 453930
rect 672257 453872 672262 453928
rect 672318 453872 674286 453928
rect 674342 453872 674347 453928
rect 672257 453870 674347 453872
rect 672257 453867 672323 453870
rect 674281 453867 674347 453870
rect 47945 430946 48011 430949
rect 41492 430944 48011 430946
rect 41492 430888 47950 430944
rect 48006 430888 48011 430944
rect 41492 430886 48011 430888
rect 47945 430883 48011 430886
rect 54477 430538 54543 430541
rect 41492 430536 54543 430538
rect 41492 430480 54482 430536
rect 54538 430480 54543 430536
rect 41492 430478 54543 430480
rect 54477 430475 54543 430478
rect 35801 430130 35867 430133
rect 35788 430128 35867 430130
rect 35788 430072 35806 430128
rect 35862 430072 35867 430128
rect 35788 430070 35867 430072
rect 35801 430067 35867 430070
rect 44541 429722 44607 429725
rect 41492 429720 44607 429722
rect 41492 429664 44546 429720
rect 44602 429664 44607 429720
rect 41492 429662 44607 429664
rect 44541 429659 44607 429662
rect 44265 429314 44331 429317
rect 41492 429312 44331 429314
rect 41492 429256 44270 429312
rect 44326 429256 44331 429312
rect 41492 429254 44331 429256
rect 44265 429251 44331 429254
rect 44909 428906 44975 428909
rect 41492 428904 44975 428906
rect 41492 428848 44914 428904
rect 44970 428848 44975 428904
rect 41492 428846 44975 428848
rect 44909 428843 44975 428846
rect 44633 428498 44699 428501
rect 41492 428496 44699 428498
rect 41492 428440 44638 428496
rect 44694 428440 44699 428496
rect 41492 428438 44699 428440
rect 44633 428435 44699 428438
rect 45829 428090 45895 428093
rect 41492 428088 45895 428090
rect 41492 428032 45834 428088
rect 45890 428032 45895 428088
rect 41492 428030 45895 428032
rect 45829 428027 45895 428030
rect 45553 427682 45619 427685
rect 41492 427680 45619 427682
rect 41492 427624 45558 427680
rect 45614 427624 45619 427680
rect 41492 427622 45619 427624
rect 45553 427619 45619 427622
rect 45737 427274 45803 427277
rect 41492 427272 45803 427274
rect 41492 427216 45742 427272
rect 45798 427216 45803 427272
rect 41492 427214 45803 427216
rect 45737 427211 45803 427214
rect 45921 426866 45987 426869
rect 41492 426864 45987 426866
rect 41492 426808 45926 426864
rect 45982 426808 45987 426864
rect 41492 426806 45987 426808
rect 45921 426803 45987 426806
rect 45737 426458 45803 426461
rect 41492 426456 45803 426458
rect 41492 426400 45742 426456
rect 45798 426400 45803 426456
rect 41492 426398 45803 426400
rect 45737 426395 45803 426398
rect 41137 426050 41203 426053
rect 41124 426048 41203 426050
rect 41124 425992 41142 426048
rect 41198 425992 41203 426048
rect 41124 425990 41203 425992
rect 41137 425987 41203 425990
rect 39254 425407 39314 425612
rect 35157 425404 35223 425407
rect 35157 425402 35266 425404
rect 35157 425346 35162 425402
rect 35218 425346 35266 425402
rect 35157 425341 35266 425346
rect 39254 425402 39363 425407
rect 39254 425346 39302 425402
rect 39358 425346 39363 425402
rect 39254 425344 39363 425346
rect 39297 425341 39363 425344
rect 35206 425204 35266 425341
rect 33041 424826 33107 424829
rect 33028 424824 33107 424826
rect 33028 424768 33046 424824
rect 33102 424768 33107 424824
rect 33028 424766 33107 424768
rect 33041 424763 33107 424766
rect 40953 424418 41019 424421
rect 40940 424416 41019 424418
rect 40940 424360 40958 424416
rect 41014 424360 41019 424416
rect 40940 424358 41019 424360
rect 40953 424355 41019 424358
rect 33777 424010 33843 424013
rect 33764 424008 33843 424010
rect 33764 423952 33782 424008
rect 33838 423952 33843 424008
rect 33764 423950 33843 423952
rect 33777 423947 33843 423950
rect 41781 424010 41847 424013
rect 42149 424010 42215 424013
rect 41781 424008 42215 424010
rect 41781 423952 41786 424008
rect 41842 423952 42154 424008
rect 42210 423952 42215 424008
rect 41781 423950 42215 423952
rect 41781 423947 41847 423950
rect 42149 423947 42215 423950
rect 42793 423602 42859 423605
rect 41492 423600 42859 423602
rect 41492 423544 42798 423600
rect 42854 423544 42859 423600
rect 41492 423542 42859 423544
rect 42793 423539 42859 423542
rect 44909 423194 44975 423197
rect 41492 423192 44975 423194
rect 41492 423136 44914 423192
rect 44970 423136 44975 423192
rect 41492 423134 44975 423136
rect 44909 423131 44975 423134
rect 42149 422922 42215 422925
rect 62389 422922 62455 422925
rect 42149 422920 62455 422922
rect 42149 422864 42154 422920
rect 42210 422864 62394 422920
rect 62450 422864 62455 422920
rect 42149 422862 62455 422864
rect 42149 422859 42215 422862
rect 62389 422859 62455 422862
rect 41492 422726 41844 422786
rect 41784 422650 41844 422726
rect 45093 422650 45159 422653
rect 41784 422648 45159 422650
rect 41784 422592 45098 422648
rect 45154 422592 45159 422648
rect 41784 422590 45159 422592
rect 45093 422587 45159 422590
rect 41822 422378 41828 422380
rect 41492 422318 41828 422378
rect 41822 422316 41828 422318
rect 41892 422316 41898 422380
rect 41781 421970 41847 421973
rect 41492 421968 41847 421970
rect 41492 421912 41786 421968
rect 41842 421912 41847 421968
rect 41492 421910 41847 421912
rect 41781 421907 41847 421910
rect 44449 421562 44515 421565
rect 41492 421560 44515 421562
rect 41492 421504 44454 421560
rect 44510 421504 44515 421560
rect 41492 421502 44515 421504
rect 44449 421499 44515 421502
rect 45277 421154 45343 421157
rect 41492 421152 45343 421154
rect 41492 421096 45282 421152
rect 45338 421096 45343 421152
rect 41492 421094 45343 421096
rect 45277 421091 45343 421094
rect 43253 420746 43319 420749
rect 41492 420744 43319 420746
rect 41492 420688 43258 420744
rect 43314 420688 43319 420744
rect 41492 420686 43319 420688
rect 43253 420683 43319 420686
rect 41462 419930 41522 420308
rect 47761 419930 47827 419933
rect 41462 419928 47827 419930
rect 41462 419900 47766 419928
rect 41492 419872 47766 419900
rect 47822 419872 47827 419928
rect 41492 419870 47827 419872
rect 47761 419867 47827 419870
rect 43069 419522 43135 419525
rect 41492 419520 43135 419522
rect 41492 419464 43074 419520
rect 43130 419464 43135 419520
rect 41492 419462 43135 419464
rect 43069 419459 43135 419462
rect 40534 418644 40540 418708
rect 40604 418706 40610 418708
rect 41505 418706 41571 418709
rect 40604 418704 41571 418706
rect 40604 418648 41510 418704
rect 41566 418648 41571 418704
rect 40604 418646 41571 418648
rect 40604 418644 40610 418646
rect 41505 418643 41571 418646
rect 40585 415986 40651 415989
rect 42609 415986 42675 415989
rect 40585 415984 42675 415986
rect 40585 415928 40590 415984
rect 40646 415928 42614 415984
rect 42670 415928 42675 415984
rect 40585 415926 42675 415928
rect 40585 415923 40651 415926
rect 42609 415923 42675 415926
rect 39297 415306 39363 415309
rect 41454 415306 41460 415308
rect 39297 415304 41460 415306
rect 39297 415248 39302 415304
rect 39358 415248 41460 415304
rect 39297 415246 41460 415248
rect 39297 415243 39363 415246
rect 41454 415244 41460 415246
rect 41524 415244 41530 415308
rect 35157 414898 35223 414901
rect 41822 414898 41828 414900
rect 35157 414896 41828 414898
rect 35157 414840 35162 414896
rect 35218 414840 41828 414896
rect 35157 414838 41828 414840
rect 35157 414835 35223 414838
rect 41822 414836 41828 414838
rect 41892 414836 41898 414900
rect 33777 414626 33843 414629
rect 41638 414626 41644 414628
rect 33777 414624 41644 414626
rect 33777 414568 33782 414624
rect 33838 414568 41644 414624
rect 33777 414566 41644 414568
rect 33777 414563 33843 414566
rect 41638 414564 41644 414566
rect 41708 414564 41714 414628
rect 42241 409866 42307 409869
rect 45093 409866 45159 409869
rect 42241 409864 45159 409866
rect 42241 409808 42246 409864
rect 42302 409808 45098 409864
rect 45154 409808 45159 409864
rect 42241 409806 45159 409808
rect 42241 409803 42307 409806
rect 45093 409803 45159 409806
rect 42057 408098 42123 408101
rect 45277 408098 45343 408101
rect 42057 408096 45343 408098
rect 42057 408040 42062 408096
rect 42118 408040 45282 408096
rect 45338 408040 45343 408096
rect 42057 408038 45343 408040
rect 42057 408035 42123 408038
rect 45277 408035 45343 408038
rect 42425 407282 42491 407285
rect 45093 407282 45159 407285
rect 42425 407280 45159 407282
rect 42425 407224 42430 407280
rect 42486 407224 45098 407280
rect 45154 407224 45159 407280
rect 42425 407222 45159 407224
rect 42425 407219 42491 407222
rect 45093 407219 45159 407222
rect 40718 406948 40724 407012
rect 40788 407010 40794 407012
rect 41781 407010 41847 407013
rect 40788 407008 41847 407010
rect 40788 406952 41786 407008
rect 41842 406952 41847 407008
rect 40788 406950 41847 406952
rect 40788 406948 40794 406950
rect 41781 406947 41847 406950
rect 42057 406738 42123 406741
rect 44449 406738 44515 406741
rect 42057 406736 44515 406738
rect 42057 406680 42062 406736
rect 42118 406680 44454 406736
rect 44510 406680 44515 406736
rect 42057 406678 44515 406680
rect 42057 406675 42123 406678
rect 44449 406675 44515 406678
rect 42241 404562 42307 404565
rect 46105 404562 46171 404565
rect 42241 404560 46171 404562
rect 42241 404504 42246 404560
rect 42302 404504 46110 404560
rect 46166 404504 46171 404560
rect 42241 404502 46171 404504
rect 42241 404499 42307 404502
rect 46105 404499 46171 404502
rect 62113 404154 62179 404157
rect 62113 404152 64706 404154
rect 62113 404096 62118 404152
rect 62174 404096 64706 404152
rect 62113 404094 64706 404096
rect 62113 404091 62179 404094
rect 40534 403820 40540 403884
rect 40604 403882 40610 403884
rect 41781 403882 41847 403885
rect 40604 403880 41847 403882
rect 40604 403824 41786 403880
rect 41842 403824 41847 403880
rect 40604 403822 41847 403824
rect 40604 403820 40610 403822
rect 41781 403819 41847 403822
rect 64646 403550 64706 404094
rect 676262 403746 676322 403852
rect 663750 403686 676322 403746
rect 657537 403338 657603 403341
rect 663750 403338 663810 403686
rect 676262 403341 676322 403444
rect 657537 403336 663810 403338
rect 657537 403280 657542 403336
rect 657598 403280 663810 403336
rect 657537 403278 663810 403280
rect 676213 403336 676322 403341
rect 676213 403280 676218 403336
rect 676274 403280 676322 403336
rect 676213 403278 676322 403280
rect 657537 403275 657603 403278
rect 676213 403275 676279 403278
rect 676630 402933 676690 403036
rect 42333 402930 42399 402933
rect 44909 402930 44975 402933
rect 42333 402928 44975 402930
rect 42333 402872 42338 402928
rect 42394 402872 44914 402928
rect 44970 402872 44975 402928
rect 42333 402870 44975 402872
rect 42333 402867 42399 402870
rect 44909 402867 44975 402870
rect 676581 402928 676690 402933
rect 676581 402872 676586 402928
rect 676642 402872 676690 402928
rect 676581 402870 676690 402872
rect 676581 402867 676647 402870
rect 62113 402658 62179 402661
rect 674833 402658 674899 402661
rect 62113 402656 64706 402658
rect 62113 402600 62118 402656
rect 62174 402600 64706 402656
rect 62113 402598 64706 402600
rect 62113 402595 62179 402598
rect 64646 402368 64706 402598
rect 674833 402656 676292 402658
rect 674833 402600 674838 402656
rect 674894 402600 676292 402656
rect 674833 402598 676292 402600
rect 674833 402595 674899 402598
rect 673177 402386 673243 402389
rect 673177 402384 676322 402386
rect 673177 402328 673182 402384
rect 673238 402328 676322 402384
rect 673177 402326 676322 402328
rect 673177 402323 673243 402326
rect 676262 402220 676322 402326
rect 672625 402114 672691 402117
rect 674833 402114 674899 402117
rect 672625 402112 674899 402114
rect 672625 402056 672630 402112
rect 672686 402056 674838 402112
rect 674894 402056 674899 402112
rect 672625 402054 674899 402056
rect 672625 402051 672691 402054
rect 674833 402051 674899 402054
rect 41781 401980 41847 401981
rect 41781 401976 41828 401980
rect 41892 401978 41898 401980
rect 41781 401920 41786 401976
rect 41781 401916 41828 401920
rect 41892 401918 41938 401978
rect 41892 401916 41898 401918
rect 41781 401915 41847 401916
rect 672441 401706 672507 401709
rect 676262 401706 676322 401812
rect 672441 401704 676322 401706
rect 672441 401648 672446 401704
rect 672502 401648 676322 401704
rect 672441 401646 676322 401648
rect 672441 401643 672507 401646
rect 673913 401434 673979 401437
rect 673913 401432 676292 401434
rect 673913 401376 673918 401432
rect 673974 401376 676292 401432
rect 673913 401374 676292 401376
rect 673913 401371 673979 401374
rect 677174 401236 677180 401300
rect 677244 401236 677250 401300
rect 62113 400618 62179 400621
rect 64646 400618 64706 401186
rect 677182 400996 677242 401236
rect 652017 400890 652083 400893
rect 676581 400890 676647 400893
rect 652017 400888 676647 400890
rect 652017 400832 652022 400888
rect 652078 400832 676586 400888
rect 676642 400832 676647 400888
rect 652017 400830 676647 400832
rect 652017 400827 652083 400830
rect 676581 400827 676647 400830
rect 62113 400616 64706 400618
rect 62113 400560 62118 400616
rect 62174 400560 64706 400616
rect 62113 400558 64706 400560
rect 62113 400555 62179 400558
rect 673361 400482 673427 400485
rect 676262 400482 676322 400588
rect 673361 400480 676322 400482
rect 673361 400424 673366 400480
rect 673422 400424 676322 400480
rect 673361 400422 676322 400424
rect 673361 400419 673427 400422
rect 676806 400420 676812 400484
rect 676876 400420 676882 400484
rect 62389 400210 62455 400213
rect 62389 400208 64706 400210
rect 62389 400152 62394 400208
rect 62450 400152 64706 400208
rect 676814 400180 676874 400420
rect 62389 400150 64706 400152
rect 62389 400147 62455 400150
rect 64646 400004 64706 400150
rect 42425 399802 42491 399805
rect 45737 399802 45803 399805
rect 42425 399800 45803 399802
rect 42425 399744 42430 399800
rect 42486 399744 45742 399800
rect 45798 399744 45803 399800
rect 42425 399742 45803 399744
rect 42425 399739 42491 399742
rect 45737 399739 45803 399742
rect 672809 399666 672875 399669
rect 676262 399666 676322 399772
rect 672809 399664 676322 399666
rect 672809 399608 672814 399664
rect 672870 399608 676322 399664
rect 672809 399606 676322 399608
rect 672809 399603 672875 399606
rect 41781 399396 41847 399397
rect 41781 399392 41828 399396
rect 41892 399394 41898 399396
rect 62113 399394 62179 399397
rect 676029 399394 676095 399397
rect 41781 399336 41786 399392
rect 41781 399332 41828 399336
rect 41892 399334 41938 399394
rect 62113 399392 64706 399394
rect 62113 399336 62118 399392
rect 62174 399336 64706 399392
rect 62113 399334 64706 399336
rect 41892 399332 41898 399334
rect 41781 399331 41847 399332
rect 62113 399331 62179 399334
rect 41454 398788 41460 398852
rect 41524 398850 41530 398852
rect 41781 398850 41847 398853
rect 41524 398848 41847 398850
rect 41524 398792 41786 398848
rect 41842 398792 41847 398848
rect 64646 398822 64706 399334
rect 676029 399392 676292 399394
rect 676029 399336 676034 399392
rect 676090 399336 676292 399392
rect 676029 399334 676292 399336
rect 676029 399331 676095 399334
rect 41524 398790 41847 398792
rect 41524 398788 41530 398790
rect 41781 398787 41847 398790
rect 676070 398788 676076 398852
rect 676140 398850 676146 398852
rect 676262 398850 676322 398956
rect 676140 398790 676322 398850
rect 676140 398788 676146 398790
rect 679574 398445 679634 398548
rect 679574 398440 679683 398445
rect 679574 398384 679622 398440
rect 679678 398384 679683 398440
rect 679574 398382 679683 398384
rect 679617 398379 679683 398382
rect 62113 398306 62179 398309
rect 62113 398304 64706 398306
rect 62113 398248 62118 398304
rect 62174 398248 64706 398304
rect 62113 398246 64706 398248
rect 62113 398243 62179 398246
rect 64646 397640 64706 398246
rect 676262 398037 676322 398140
rect 676213 398032 676322 398037
rect 676213 397976 676218 398032
rect 676274 397976 676322 398032
rect 676213 397974 676322 397976
rect 676213 397971 676279 397974
rect 678286 397629 678346 397732
rect 678237 397624 678346 397629
rect 678237 397568 678242 397624
rect 678298 397568 678346 397624
rect 678237 397566 678346 397568
rect 678237 397563 678303 397566
rect 674741 397354 674807 397357
rect 674741 397352 676292 397354
rect 674741 397296 674746 397352
rect 674802 397296 676292 397352
rect 674741 397294 676292 397296
rect 674741 397291 674807 397294
rect 676630 396812 676690 396916
rect 676622 396748 676628 396812
rect 676692 396748 676698 396812
rect 652201 396674 652267 396677
rect 674557 396674 674623 396677
rect 652201 396672 674623 396674
rect 652201 396616 652206 396672
rect 652262 396616 674562 396672
rect 674618 396616 674623 396672
rect 652201 396614 674623 396616
rect 652201 396611 652267 396614
rect 674557 396611 674623 396614
rect 676446 396404 676506 396508
rect 676438 396340 676444 396404
rect 676508 396340 676514 396404
rect 676029 396130 676095 396133
rect 676029 396128 676292 396130
rect 676029 396072 676034 396128
rect 676090 396072 676292 396128
rect 676029 396070 676292 396072
rect 676029 396067 676095 396070
rect 674097 395858 674163 395861
rect 674097 395856 676322 395858
rect 674097 395800 674102 395856
rect 674158 395800 676322 395856
rect 674097 395798 676322 395800
rect 674097 395795 674163 395798
rect 42149 395722 42215 395725
rect 51073 395722 51139 395725
rect 42149 395720 51139 395722
rect 42149 395664 42154 395720
rect 42210 395664 51078 395720
rect 51134 395664 51139 395720
rect 676262 395692 676322 395798
rect 42149 395662 51139 395664
rect 42149 395659 42215 395662
rect 51073 395659 51139 395662
rect 676262 395180 676322 395284
rect 676254 395116 676260 395180
rect 676324 395116 676330 395180
rect 672993 394770 673059 394773
rect 676262 394770 676322 394876
rect 672993 394768 676322 394770
rect 672993 394712 672998 394768
rect 673054 394712 676322 394768
rect 672993 394710 676322 394712
rect 672993 394707 673059 394710
rect 676262 394365 676322 394468
rect 676213 394360 676322 394365
rect 676213 394304 676218 394360
rect 676274 394304 676322 394360
rect 676213 394302 676322 394304
rect 676213 394299 676279 394302
rect 672625 393954 672691 393957
rect 676262 393954 676322 394060
rect 672625 393952 676322 393954
rect 672625 393896 672630 393952
rect 672686 393896 676322 393952
rect 672625 393894 676322 393896
rect 672625 393891 672691 393894
rect 676630 393549 676690 393652
rect 676630 393544 676739 393549
rect 676630 393488 676678 393544
rect 676734 393488 676739 393544
rect 676630 393486 676739 393488
rect 676673 393483 676739 393486
rect 675886 392804 675892 392868
rect 675956 392866 675962 392868
rect 676262 392866 676322 393244
rect 675956 392836 676322 392866
rect 675956 392806 676292 392836
rect 675956 392804 675962 392806
rect 671337 392594 671403 392597
rect 671337 392592 676322 392594
rect 671337 392536 671342 392592
rect 671398 392536 676322 392592
rect 671337 392534 676322 392536
rect 671337 392531 671403 392534
rect 676262 392428 676322 392534
rect 668577 391234 668643 391237
rect 676673 391234 676739 391237
rect 668577 391232 676739 391234
rect 668577 391176 668582 391232
rect 668638 391176 676678 391232
rect 676734 391176 676739 391232
rect 668577 391174 676739 391176
rect 668577 391171 668643 391174
rect 676673 391171 676739 391174
rect 47945 387698 48011 387701
rect 41492 387696 48011 387698
rect 41492 387640 47950 387696
rect 48006 387640 48011 387696
rect 41492 387638 48011 387640
rect 47945 387635 48011 387638
rect 675702 387636 675708 387700
rect 675772 387698 675778 387700
rect 678237 387698 678303 387701
rect 675772 387696 678303 387698
rect 675772 387640 678242 387696
rect 678298 387640 678303 387696
rect 675772 387638 678303 387640
rect 675772 387636 675778 387638
rect 678237 387635 678303 387638
rect 41094 387157 41154 387260
rect 41094 387152 41203 387157
rect 41094 387096 41142 387152
rect 41198 387096 41203 387152
rect 41094 387094 41203 387096
rect 41137 387091 41203 387094
rect 41278 386749 41338 386852
rect 41278 386744 41387 386749
rect 41278 386688 41326 386744
rect 41382 386688 41387 386744
rect 41278 386686 41387 386688
rect 41321 386683 41387 386686
rect 44265 386474 44331 386477
rect 41492 386472 44331 386474
rect 41492 386416 44270 386472
rect 44326 386416 44331 386472
rect 41492 386414 44331 386416
rect 44265 386411 44331 386414
rect 40910 385933 40970 386036
rect 40910 385928 41019 385933
rect 40910 385872 40958 385928
rect 41014 385872 41019 385928
rect 40910 385870 41019 385872
rect 40953 385867 41019 385870
rect 41321 385930 41387 385933
rect 62205 385930 62271 385933
rect 41321 385928 62271 385930
rect 41321 385872 41326 385928
rect 41382 385872 62210 385928
rect 62266 385872 62271 385928
rect 41321 385870 62271 385872
rect 41321 385867 41387 385870
rect 62205 385867 62271 385870
rect 44633 385658 44699 385661
rect 41492 385656 44699 385658
rect 41492 385600 44638 385656
rect 44694 385600 44699 385656
rect 41492 385598 44699 385600
rect 44633 385595 44699 385598
rect 45093 385250 45159 385253
rect 41492 385248 45159 385250
rect 41492 385192 45098 385248
rect 45154 385192 45159 385248
rect 41492 385190 45159 385192
rect 45093 385187 45159 385190
rect 675753 384978 675819 384981
rect 676622 384978 676628 384980
rect 675753 384976 676628 384978
rect 675753 384920 675758 384976
rect 675814 384920 676628 384976
rect 675753 384918 676628 384920
rect 675753 384915 675819 384918
rect 676622 384916 676628 384918
rect 676692 384916 676698 384980
rect 45553 384842 45619 384845
rect 41492 384840 45619 384842
rect 41492 384784 45558 384840
rect 45614 384784 45619 384840
rect 41492 384782 45619 384784
rect 45553 384779 45619 384782
rect 45553 384434 45619 384437
rect 41492 384432 45619 384434
rect 41492 384376 45558 384432
rect 45614 384376 45619 384432
rect 41492 384374 45619 384376
rect 45553 384371 45619 384374
rect 45921 384026 45987 384029
rect 41492 384024 45987 384026
rect 41492 383968 45926 384024
rect 45982 383968 45987 384024
rect 41492 383966 45987 383968
rect 45921 383963 45987 383966
rect 46197 383618 46263 383621
rect 41492 383616 46263 383618
rect 41492 383560 46202 383616
rect 46258 383560 46263 383616
rect 41492 383558 46263 383560
rect 46197 383555 46263 383558
rect 41462 383076 41522 383180
rect 41454 383012 41460 383076
rect 41524 383012 41530 383076
rect 654777 382938 654843 382941
rect 675201 382938 675267 382941
rect 654777 382936 675267 382938
rect 654777 382880 654782 382936
rect 654838 382880 675206 382936
rect 675262 382880 675267 382936
rect 654777 382878 675267 382880
rect 654777 382875 654843 382878
rect 675201 382875 675267 382878
rect 41278 382669 41338 382772
rect 41278 382664 41387 382669
rect 41278 382608 41326 382664
rect 41382 382608 41387 382664
rect 41278 382606 41387 382608
rect 41321 382603 41387 382606
rect 40174 382261 40234 382364
rect 40174 382256 40283 382261
rect 40174 382200 40222 382256
rect 40278 382200 40283 382256
rect 40174 382198 40283 382200
rect 40217 382195 40283 382198
rect 40953 382258 41019 382261
rect 44909 382258 44975 382261
rect 40953 382256 44975 382258
rect 40953 382200 40958 382256
rect 41014 382200 44914 382256
rect 44970 382200 44975 382256
rect 40953 382198 44975 382200
rect 40953 382195 41019 382198
rect 44909 382195 44975 382198
rect 675753 382258 675819 382261
rect 676438 382258 676444 382260
rect 675753 382256 676444 382258
rect 675753 382200 675758 382256
rect 675814 382200 676444 382256
rect 675753 382198 676444 382200
rect 675753 382195 675819 382198
rect 676438 382196 676444 382198
rect 676508 382196 676514 382260
rect 39990 381853 40050 381956
rect 39990 381848 40099 381853
rect 39990 381792 40038 381848
rect 40094 381792 40099 381848
rect 39990 381790 40099 381792
rect 40033 381787 40099 381790
rect 41137 381850 41203 381853
rect 62665 381850 62731 381853
rect 41137 381848 62731 381850
rect 41137 381792 41142 381848
rect 41198 381792 62670 381848
rect 62726 381792 62731 381848
rect 41137 381790 62731 381792
rect 41137 381787 41203 381790
rect 62665 381787 62731 381790
rect 32446 381445 32506 381548
rect 32397 381440 32506 381445
rect 32397 381384 32402 381440
rect 32458 381384 32506 381440
rect 32397 381382 32506 381384
rect 32397 381379 32463 381382
rect 37966 381037 38026 381140
rect 37917 381032 38026 381037
rect 37917 380976 37922 381032
rect 37978 380976 38026 381032
rect 37917 380974 38026 380976
rect 672993 381034 673059 381037
rect 675385 381034 675451 381037
rect 672993 381032 675451 381034
rect 672993 380976 672998 381032
rect 673054 380976 675390 381032
rect 675446 380976 675451 381032
rect 672993 380974 675451 380976
rect 37917 380971 37983 380974
rect 672993 380971 673059 380974
rect 675385 380971 675451 380974
rect 46013 380762 46079 380765
rect 41492 380760 46079 380762
rect 41492 380704 46018 380760
rect 46074 380704 46079 380760
rect 41492 380702 46079 380704
rect 46013 380699 46079 380702
rect 44449 380354 44515 380357
rect 41492 380352 44515 380354
rect 41492 380296 44454 380352
rect 44510 380296 44515 380352
rect 41492 380294 44515 380296
rect 44449 380291 44515 380294
rect 42793 379946 42859 379949
rect 41492 379944 42859 379946
rect 41492 379888 42798 379944
rect 42854 379888 42859 379944
rect 41492 379886 42859 379888
rect 42793 379883 42859 379886
rect 40726 379404 40786 379530
rect 40718 379340 40724 379404
rect 40788 379340 40794 379404
rect 44633 379402 44699 379405
rect 41278 379400 44699 379402
rect 41278 379344 44638 379400
rect 44694 379344 44699 379400
rect 41278 379342 44699 379344
rect 41278 379100 41338 379342
rect 44633 379339 44699 379342
rect 40217 378994 40283 378997
rect 41638 378994 41644 378996
rect 40217 378992 41644 378994
rect 40217 378936 40222 378992
rect 40278 378936 41644 378992
rect 40217 378934 41644 378936
rect 40217 378931 40283 378934
rect 41638 378932 41644 378934
rect 41708 378932 41714 378996
rect 46473 378722 46539 378725
rect 675753 378724 675819 378725
rect 675702 378722 675708 378724
rect 41492 378720 46539 378722
rect 41492 378664 46478 378720
rect 46534 378664 46539 378720
rect 41492 378662 46539 378664
rect 675662 378662 675708 378722
rect 675772 378720 675819 378724
rect 675814 378664 675819 378720
rect 46473 378659 46539 378662
rect 675702 378660 675708 378662
rect 675772 378660 675819 378664
rect 675753 378659 675819 378660
rect 40542 378180 40602 378284
rect 40534 378116 40540 378180
rect 40604 378116 40610 378180
rect 40910 377772 40970 377876
rect 40902 377708 40908 377772
rect 40972 377708 40978 377772
rect 44173 377498 44239 377501
rect 41492 377496 44239 377498
rect 41492 377440 44178 377496
rect 44234 377440 44239 377496
rect 41492 377438 44239 377440
rect 44173 377435 44239 377438
rect 675753 377362 675819 377365
rect 676254 377362 676260 377364
rect 675753 377360 676260 377362
rect 675753 377304 675758 377360
rect 675814 377304 676260 377360
rect 675753 377302 676260 377304
rect 675753 377299 675819 377302
rect 676254 377300 676260 377302
rect 676324 377300 676330 377364
rect 35758 376549 35818 377060
rect 40033 376954 40099 376957
rect 41822 376954 41828 376956
rect 40033 376952 41828 376954
rect 40033 376896 40038 376952
rect 40094 376896 41828 376952
rect 40033 376894 41828 376896
rect 40033 376891 40099 376894
rect 41822 376892 41828 376894
rect 41892 376892 41898 376956
rect 47577 376682 47643 376685
rect 39100 376680 47643 376682
rect 39100 376652 47582 376680
rect 39070 376624 47582 376652
rect 47638 376624 47643 376680
rect 39070 376622 47643 376624
rect 39070 376549 39130 376622
rect 47577 376619 47643 376622
rect 35758 376544 35867 376549
rect 35758 376488 35806 376544
rect 35862 376488 35867 376544
rect 35758 376486 35867 376488
rect 35801 376483 35867 376486
rect 39021 376544 39130 376549
rect 39021 376488 39026 376544
rect 39082 376488 39130 376544
rect 39021 376486 39130 376488
rect 39021 376483 39087 376486
rect 45829 376274 45895 376277
rect 41492 376272 45895 376274
rect 41492 376216 45834 376272
rect 45890 376216 45895 376272
rect 41492 376214 45895 376216
rect 45829 376211 45895 376214
rect 672625 376274 672691 376277
rect 675385 376274 675451 376277
rect 672625 376272 675451 376274
rect 672625 376216 672630 376272
rect 672686 376216 675390 376272
rect 675446 376216 675451 376272
rect 672625 376214 675451 376216
rect 672625 376211 672691 376214
rect 675385 376211 675451 376214
rect 35801 376138 35867 376141
rect 39021 376138 39087 376141
rect 35801 376136 39087 376138
rect 35801 376080 35806 376136
rect 35862 376080 39026 376136
rect 39082 376080 39087 376136
rect 35801 376078 39087 376080
rect 35801 376075 35867 376078
rect 39021 376075 39087 376078
rect 652201 373962 652267 373965
rect 649950 373960 652267 373962
rect 649950 373904 652206 373960
rect 652262 373904 652267 373960
rect 649950 373902 652267 373904
rect 649950 373892 650010 373902
rect 652201 373899 652267 373902
rect 675753 373690 675819 373693
rect 676070 373690 676076 373692
rect 675753 373688 676076 373690
rect 675753 373632 675758 373688
rect 675814 373632 676076 373688
rect 675753 373630 676076 373632
rect 675753 373627 675819 373630
rect 676070 373628 676076 373630
rect 676140 373628 676146 373692
rect 651465 373282 651531 373285
rect 649950 373280 651531 373282
rect 649950 373224 651470 373280
rect 651526 373224 651531 373280
rect 649950 373222 651531 373224
rect 649950 372710 650010 373222
rect 651465 373219 651531 373222
rect 675661 373012 675727 373013
rect 675661 373008 675708 373012
rect 675772 373010 675778 373012
rect 675661 372952 675666 373008
rect 675661 372948 675708 372952
rect 675772 372950 675818 373010
rect 675772 372948 675778 372950
rect 675661 372947 675727 372948
rect 652017 372194 652083 372197
rect 649950 372192 652083 372194
rect 649950 372136 652022 372192
rect 652078 372136 652083 372192
rect 649950 372134 652083 372136
rect 649950 371528 650010 372134
rect 652017 372131 652083 372134
rect 651465 370698 651531 370701
rect 649950 370696 651531 370698
rect 649950 370640 651470 370696
rect 651526 370640 651531 370696
rect 649950 370638 651531 370640
rect 649950 370346 650010 370638
rect 651465 370635 651531 370638
rect 40718 365604 40724 365668
rect 40788 365666 40794 365668
rect 41781 365666 41847 365669
rect 40788 365664 41847 365666
rect 40788 365608 41786 365664
rect 41842 365608 41847 365664
rect 40788 365606 41847 365608
rect 40788 365604 40794 365606
rect 41781 365603 41847 365606
rect 40902 364244 40908 364308
rect 40972 364306 40978 364308
rect 41781 364306 41847 364309
rect 40972 364304 41847 364306
rect 40972 364248 41786 364304
rect 41842 364248 41847 364304
rect 40972 364246 41847 364248
rect 40972 364244 40978 364246
rect 41781 364243 41847 364246
rect 42149 364306 42215 364309
rect 44633 364306 44699 364309
rect 42149 364304 44699 364306
rect 42149 364248 42154 364304
rect 42210 364248 44638 364304
rect 44694 364248 44699 364304
rect 42149 364246 44699 364248
rect 42149 364243 42215 364246
rect 44633 364243 44699 364246
rect 40534 363700 40540 363764
rect 40604 363762 40610 363764
rect 41781 363762 41847 363765
rect 40604 363760 41847 363762
rect 40604 363704 41786 363760
rect 41842 363704 41847 363760
rect 40604 363702 41847 363704
rect 40604 363700 40610 363702
rect 41781 363699 41847 363702
rect 42425 363082 42491 363085
rect 45369 363082 45435 363085
rect 42425 363080 45435 363082
rect 42425 363024 42430 363080
rect 42486 363024 45374 363080
rect 45430 363024 45435 363080
rect 42425 363022 45435 363024
rect 42425 363019 42491 363022
rect 45369 363019 45435 363022
rect 42241 362946 42307 362949
rect 42198 362944 42307 362946
rect 42198 362888 42246 362944
rect 42302 362888 42307 362944
rect 42198 362883 42307 362888
rect 42198 362674 42258 362883
rect 46749 362674 46815 362677
rect 42198 362672 46815 362674
rect 42198 362616 46754 362672
rect 46810 362616 46815 362672
rect 42198 362614 46815 362616
rect 46749 362611 46815 362614
rect 62113 360906 62179 360909
rect 62113 360904 64706 360906
rect 62113 360848 62118 360904
rect 62174 360848 64706 360904
rect 62113 360846 64706 360848
rect 62113 360843 62179 360846
rect 64646 360328 64706 360846
rect 62113 359818 62179 359821
rect 62113 359816 64706 359818
rect 62113 359760 62118 359816
rect 62174 359760 64706 359816
rect 62113 359758 64706 359760
rect 62113 359755 62179 359758
rect 42057 359274 42123 359277
rect 44449 359274 44515 359277
rect 42057 359272 44515 359274
rect 42057 359216 42062 359272
rect 42118 359216 44454 359272
rect 44510 359216 44515 359272
rect 42057 359214 44515 359216
rect 42057 359211 42123 359214
rect 44449 359211 44515 359214
rect 64646 359146 64706 359758
rect 41873 358732 41939 358733
rect 41822 358730 41828 358732
rect 41782 358670 41828 358730
rect 41892 358728 41939 358732
rect 41934 358672 41939 358728
rect 41822 358668 41828 358670
rect 41892 358668 41939 358672
rect 41873 358667 41939 358668
rect 42425 358730 42491 358733
rect 46473 358730 46539 358733
rect 42425 358728 46539 358730
rect 42425 358672 42430 358728
rect 42486 358672 46478 358728
rect 46534 358672 46539 358728
rect 42425 358670 46539 358672
rect 42425 358667 42491 358670
rect 46473 358667 46539 358670
rect 667381 358730 667447 358733
rect 667381 358728 676292 358730
rect 667381 358672 667386 358728
rect 667442 358672 676292 358728
rect 667381 358670 676292 358672
rect 667381 358667 667447 358670
rect 673913 358322 673979 358325
rect 673913 358320 676292 358322
rect 673913 358264 673918 358320
rect 673974 358264 676292 358320
rect 673913 358262 676292 358264
rect 673913 358259 673979 358262
rect 62113 357778 62179 357781
rect 64646 357778 64706 357964
rect 675937 357914 676003 357917
rect 675937 357912 676292 357914
rect 675937 357856 675942 357912
rect 675998 357856 676292 357912
rect 675937 357854 676292 357856
rect 675937 357851 676003 357854
rect 62113 357776 64706 357778
rect 62113 357720 62118 357776
rect 62174 357720 64706 357776
rect 62113 357718 64706 357720
rect 62113 357715 62179 357718
rect 673177 357506 673243 357509
rect 673177 357504 676292 357506
rect 673177 357448 673182 357504
rect 673238 357448 676292 357504
rect 673177 357446 676292 357448
rect 673177 357443 673243 357446
rect 62297 357370 62363 357373
rect 62297 357368 64706 357370
rect 62297 357312 62302 357368
rect 62358 357312 64706 357368
rect 62297 357310 64706 357312
rect 62297 357307 62363 357310
rect 41454 356900 41460 356964
rect 41524 356962 41530 356964
rect 41781 356962 41847 356965
rect 41524 356960 41847 356962
rect 41524 356904 41786 356960
rect 41842 356904 41847 356960
rect 41524 356902 41847 356904
rect 41524 356900 41530 356902
rect 41781 356899 41847 356902
rect 64646 356782 64706 357310
rect 672533 357098 672599 357101
rect 672533 357096 676292 357098
rect 672533 357040 672538 357096
rect 672594 357040 676292 357096
rect 672533 357038 676292 357040
rect 672533 357035 672599 357038
rect 675937 356826 676003 356829
rect 669270 356824 676003 356826
rect 669270 356768 675942 356824
rect 675998 356768 676003 356824
rect 669270 356766 676003 356768
rect 652017 356690 652083 356693
rect 669270 356690 669330 356766
rect 675937 356763 676003 356766
rect 652017 356688 669330 356690
rect 652017 356632 652022 356688
rect 652078 356632 669330 356688
rect 652017 356630 669330 356632
rect 676170 356630 676292 356690
rect 652017 356627 652083 356630
rect 674373 356554 674439 356557
rect 676170 356554 676230 356630
rect 674373 356552 676230 356554
rect 674373 356496 674378 356552
rect 674434 356496 676230 356552
rect 674373 356494 676230 356496
rect 674373 356491 674439 356494
rect 674097 356282 674163 356285
rect 674097 356280 676292 356282
rect 674097 356224 674102 356280
rect 674158 356224 676292 356280
rect 674097 356222 676292 356224
rect 674097 356219 674163 356222
rect 62113 356010 62179 356013
rect 62113 356008 64706 356010
rect 62113 355952 62118 356008
rect 62174 355952 64706 356008
rect 62113 355950 64706 355952
rect 62113 355947 62179 355950
rect 41873 355604 41939 355605
rect 41822 355602 41828 355604
rect 41782 355542 41828 355602
rect 41892 355600 41939 355604
rect 64646 355600 64706 355950
rect 673361 355874 673427 355877
rect 673361 355872 676292 355874
rect 673361 355816 673366 355872
rect 673422 355816 676292 355872
rect 673361 355814 676292 355816
rect 673361 355811 673427 355814
rect 41934 355544 41939 355600
rect 41822 355540 41828 355542
rect 41892 355540 41939 355544
rect 41873 355539 41939 355540
rect 673361 355466 673427 355469
rect 673361 355464 676292 355466
rect 673361 355408 673366 355464
rect 673422 355408 676292 355464
rect 673361 355406 676292 355408
rect 673361 355403 673427 355406
rect 672809 355058 672875 355061
rect 672809 355056 676292 355058
rect 672809 355000 672814 355056
rect 672870 355000 676292 355056
rect 672809 354998 676292 355000
rect 672809 354995 672875 354998
rect 43897 354922 43963 354925
rect 45185 354922 45251 354925
rect 43897 354920 45251 354922
rect 43897 354864 43902 354920
rect 43958 354864 45190 354920
rect 45246 354864 45251 354920
rect 43897 354862 45251 354864
rect 43897 354859 43963 354862
rect 45185 354859 45251 354862
rect 673177 354650 673243 354653
rect 673177 354648 676292 354650
rect 673177 354592 673182 354648
rect 673238 354592 676292 354648
rect 673177 354590 676292 354592
rect 673177 354587 673243 354590
rect 62665 354514 62731 354517
rect 62665 354512 64706 354514
rect 62665 354456 62670 354512
rect 62726 354456 64706 354512
rect 62665 354454 64706 354456
rect 62665 354451 62731 354454
rect 64646 354418 64706 354454
rect 675518 354180 675524 354244
rect 675588 354242 675594 354244
rect 675588 354182 676292 354242
rect 675588 354180 675594 354182
rect 43069 353970 43135 353973
rect 45277 353970 45343 353973
rect 43069 353968 45343 353970
rect 43069 353912 43074 353968
rect 43130 353912 45282 353968
rect 45338 353912 45343 353968
rect 43069 353910 45343 353912
rect 43069 353907 43135 353910
rect 45277 353907 45343 353910
rect 675886 353908 675892 353972
rect 675956 353970 675962 353972
rect 675956 353910 676230 353970
rect 675956 353908 675962 353910
rect 676170 353834 676230 353910
rect 676170 353774 676292 353834
rect 43253 353698 43319 353701
rect 45277 353698 45343 353701
rect 43253 353696 45343 353698
rect 43253 353640 43258 353696
rect 43314 353640 45282 353696
rect 45338 353640 45343 353696
rect 43253 353638 45343 353640
rect 43253 353635 43319 353638
rect 45277 353635 45343 353638
rect 672717 353426 672783 353429
rect 672717 353424 676292 353426
rect 672717 353368 672722 353424
rect 672778 353368 676292 353424
rect 672717 353366 676292 353368
rect 672717 353363 672783 353366
rect 42149 353290 42215 353293
rect 51717 353290 51783 353293
rect 42149 353288 51783 353290
rect 42149 353232 42154 353288
rect 42210 353232 51722 353288
rect 51778 353232 51783 353288
rect 42149 353230 51783 353232
rect 42149 353227 42215 353230
rect 51717 353227 51783 353230
rect 42425 353018 42491 353021
rect 45921 353018 45987 353021
rect 42425 353016 45987 353018
rect 42425 352960 42430 353016
rect 42486 352960 45926 353016
rect 45982 352960 45987 353016
rect 42425 352958 45987 352960
rect 42425 352955 42491 352958
rect 45921 352955 45987 352958
rect 675702 352956 675708 353020
rect 675772 353018 675778 353020
rect 675772 352958 676292 353018
rect 675772 352956 675778 352958
rect 672165 352610 672231 352613
rect 672165 352608 676292 352610
rect 672165 352552 672170 352608
rect 672226 352552 676292 352608
rect 672165 352550 676292 352552
rect 672165 352547 672231 352550
rect 674649 352202 674715 352205
rect 674649 352200 676292 352202
rect 674649 352144 674654 352200
rect 674710 352144 676292 352200
rect 674649 352142 676292 352144
rect 674649 352139 674715 352142
rect 676170 351734 676292 351794
rect 675886 351596 675892 351660
rect 675956 351658 675962 351660
rect 676170 351658 676230 351734
rect 675956 351598 676230 351658
rect 675956 351596 675962 351598
rect 673729 351386 673795 351389
rect 673729 351384 676292 351386
rect 673729 351328 673734 351384
rect 673790 351328 676292 351384
rect 673729 351326 676292 351328
rect 673729 351323 673795 351326
rect 652385 351114 652451 351117
rect 673913 351114 673979 351117
rect 652385 351112 673979 351114
rect 652385 351056 652390 351112
rect 652446 351056 673918 351112
rect 673974 351056 673979 351112
rect 652385 351054 673979 351056
rect 652385 351051 652451 351054
rect 673913 351051 673979 351054
rect 674465 350978 674531 350981
rect 674465 350976 676292 350978
rect 674465 350920 674470 350976
rect 674526 350920 676292 350976
rect 674465 350918 676292 350920
rect 674465 350915 674531 350918
rect 674465 350570 674531 350573
rect 674465 350568 676292 350570
rect 674465 350512 674470 350568
rect 674526 350512 676292 350568
rect 674465 350510 676292 350512
rect 674465 350507 674531 350510
rect 676029 350162 676095 350165
rect 676029 350160 676292 350162
rect 676029 350104 676034 350160
rect 676090 350104 676292 350160
rect 676029 350102 676292 350104
rect 676029 350099 676095 350102
rect 674281 349754 674347 349757
rect 674281 349752 676292 349754
rect 674281 349696 674286 349752
rect 674342 349696 676292 349752
rect 674281 349694 676292 349696
rect 674281 349691 674347 349694
rect 672349 349346 672415 349349
rect 672349 349344 676292 349346
rect 672349 349288 672354 349344
rect 672410 349288 676292 349344
rect 672349 349286 676292 349288
rect 672349 349283 672415 349286
rect 672901 348938 672967 348941
rect 672901 348936 676292 348938
rect 672901 348880 672906 348936
rect 672962 348880 676292 348936
rect 672901 348878 676292 348880
rect 672901 348875 672967 348878
rect 671521 348530 671587 348533
rect 671521 348528 676292 348530
rect 671521 348472 671526 348528
rect 671582 348472 676292 348528
rect 671521 348470 676292 348472
rect 671521 348467 671587 348470
rect 675334 347652 675340 347716
rect 675404 347714 675410 347716
rect 683070 347714 683130 348092
rect 675404 347684 683130 347714
rect 675404 347654 683100 347684
rect 675404 347652 675410 347654
rect 670601 347306 670667 347309
rect 670601 347304 676292 347306
rect 670601 347248 670606 347304
rect 670662 347248 676292 347304
rect 670601 347246 676292 347248
rect 670601 347243 670667 347246
rect 676029 346626 676095 346629
rect 676438 346626 676444 346628
rect 676029 346624 676444 346626
rect 676029 346568 676034 346624
rect 676090 346568 676444 346624
rect 676029 346566 676444 346568
rect 676029 346563 676095 346566
rect 676438 346564 676444 346566
rect 676508 346564 676514 346628
rect 669313 344994 669379 344997
rect 675201 344994 675267 344997
rect 669313 344992 675267 344994
rect 669313 344936 669318 344992
rect 669374 344936 675206 344992
rect 675262 344936 675267 344992
rect 669313 344934 675267 344936
rect 669313 344931 669379 344934
rect 675201 344931 675267 344934
rect 35574 344317 35634 344556
rect 35525 344312 35634 344317
rect 35801 344314 35867 344317
rect 35525 344256 35530 344312
rect 35586 344256 35634 344312
rect 35525 344254 35634 344256
rect 35758 344312 35867 344314
rect 35758 344256 35806 344312
rect 35862 344256 35867 344312
rect 35525 344251 35591 344254
rect 35758 344251 35867 344256
rect 39665 344314 39731 344317
rect 45553 344314 45619 344317
rect 39665 344312 45619 344314
rect 39665 344256 39670 344312
rect 39726 344256 45558 344312
rect 45614 344256 45619 344312
rect 39665 344254 45619 344256
rect 39665 344251 39731 344254
rect 45553 344251 45619 344254
rect 35758 344148 35818 344251
rect 35758 343501 35818 343740
rect 35758 343496 35867 343501
rect 35758 343440 35806 343496
rect 35862 343440 35867 343496
rect 35758 343438 35867 343440
rect 35801 343435 35867 343438
rect 44909 343362 44975 343365
rect 41492 343360 44975 343362
rect 41492 343304 44914 343360
rect 44970 343304 44975 343360
rect 41492 343302 44975 343304
rect 44909 343299 44975 343302
rect 44214 342954 44220 342956
rect 41492 342894 44220 342954
rect 44214 342892 44220 342894
rect 44284 342892 44290 342956
rect 45093 342546 45159 342549
rect 41492 342544 45159 342546
rect 41492 342488 45098 342544
rect 45154 342488 45159 342544
rect 41492 342486 45159 342488
rect 45093 342483 45159 342486
rect 40217 342274 40283 342277
rect 45461 342274 45527 342277
rect 40217 342272 45527 342274
rect 40217 342216 40222 342272
rect 40278 342216 45466 342272
rect 45522 342216 45527 342272
rect 40217 342214 45527 342216
rect 40217 342211 40283 342214
rect 45461 342211 45527 342214
rect 39438 341869 39498 342108
rect 39438 341864 39547 341869
rect 39438 341808 39486 341864
rect 39542 341808 39547 341864
rect 39438 341806 39547 341808
rect 39481 341803 39547 341806
rect 40033 341866 40099 341869
rect 40033 341864 45570 341866
rect 40033 341808 40038 341864
rect 40094 341808 45570 341864
rect 40033 341806 45570 341808
rect 40033 341803 40099 341806
rect 45510 341730 45570 341806
rect 62665 341730 62731 341733
rect 45510 341728 62731 341730
rect 35574 341461 35634 341700
rect 45510 341672 62670 341728
rect 62726 341672 62731 341728
rect 45510 341670 62731 341672
rect 62665 341667 62731 341670
rect 35574 341456 35683 341461
rect 35574 341400 35622 341456
rect 35678 341400 35683 341456
rect 35574 341398 35683 341400
rect 35617 341395 35683 341398
rect 39849 341458 39915 341461
rect 62481 341458 62547 341461
rect 39849 341456 62547 341458
rect 39849 341400 39854 341456
rect 39910 341400 62486 341456
rect 62542 341400 62547 341456
rect 39849 341398 62547 341400
rect 39849 341395 39915 341398
rect 62481 341395 62547 341398
rect 35801 341050 35867 341053
rect 35758 341048 35867 341050
rect 35758 340992 35806 341048
rect 35862 340992 35867 341048
rect 35758 340987 35867 340992
rect 40217 341050 40283 341053
rect 41462 341050 41522 341292
rect 44582 341050 44588 341052
rect 40217 341048 40602 341050
rect 40217 340992 40222 341048
rect 40278 340992 40602 341048
rect 40217 340990 40602 340992
rect 41462 340990 44588 341050
rect 40217 340987 40283 340990
rect 35758 340884 35818 340987
rect 40542 340778 40602 340990
rect 44582 340988 44588 340990
rect 44652 340988 44658 341052
rect 46105 340778 46171 340781
rect 40542 340776 46171 340778
rect 40542 340720 46110 340776
rect 46166 340720 46171 340776
rect 40542 340718 46171 340720
rect 46105 340715 46171 340718
rect 672717 340778 672783 340781
rect 675109 340778 675175 340781
rect 672717 340776 675175 340778
rect 672717 340720 672722 340776
rect 672778 340720 675114 340776
rect 675170 340720 675175 340776
rect 672717 340718 675175 340720
rect 672717 340715 672783 340718
rect 675109 340715 675175 340718
rect 42742 340506 42748 340508
rect 41492 340446 42748 340506
rect 42742 340444 42748 340446
rect 42812 340444 42818 340508
rect 675753 340370 675819 340373
rect 676254 340370 676260 340372
rect 675753 340368 676260 340370
rect 675753 340312 675758 340368
rect 675814 340312 676260 340368
rect 675753 340310 676260 340312
rect 675753 340307 675819 340310
rect 676254 340308 676260 340310
rect 676324 340308 676330 340372
rect 39481 340234 39547 340237
rect 44398 340234 44404 340236
rect 39481 340232 44404 340234
rect 39481 340176 39486 340232
rect 39542 340176 44404 340232
rect 39481 340174 44404 340176
rect 39481 340171 39547 340174
rect 44398 340172 44404 340174
rect 44468 340172 44474 340236
rect 35574 339829 35634 340068
rect 35525 339824 35634 339829
rect 35801 339826 35867 339829
rect 35525 339768 35530 339824
rect 35586 339768 35634 339824
rect 35525 339766 35634 339768
rect 35758 339824 35867 339826
rect 35758 339768 35806 339824
rect 35862 339768 35867 339824
rect 35525 339763 35591 339766
rect 35758 339763 35867 339768
rect 35758 339660 35818 339763
rect 675477 339420 675543 339421
rect 675477 339416 675524 339420
rect 675588 339418 675594 339420
rect 675477 339360 675482 339416
rect 675477 339356 675524 339360
rect 675588 339358 675634 339418
rect 675588 339356 675594 339358
rect 675477 339355 675543 339356
rect 45645 339282 45711 339285
rect 41492 339280 45711 339282
rect 41492 339224 45650 339280
rect 45706 339224 45711 339280
rect 41492 339222 45711 339224
rect 45645 339219 45711 339222
rect 35206 338605 35266 338844
rect 653397 338738 653463 338741
rect 674925 338738 674991 338741
rect 653397 338736 674991 338738
rect 653397 338680 653402 338736
rect 653458 338680 674930 338736
rect 674986 338680 674991 338736
rect 653397 338678 674991 338680
rect 653397 338675 653463 338678
rect 674925 338675 674991 338678
rect 35157 338600 35266 338605
rect 35157 338544 35162 338600
rect 35218 338544 35266 338600
rect 35157 338542 35266 338544
rect 35157 338539 35223 338542
rect 46933 338466 46999 338469
rect 41492 338464 46999 338466
rect 41492 338408 46938 338464
rect 46994 338408 46999 338464
rect 41492 338406 46999 338408
rect 46933 338403 46999 338406
rect 45461 338058 45527 338061
rect 41492 338056 45527 338058
rect 41492 338000 45466 338056
rect 45522 338000 45527 338056
rect 41492 337998 45527 338000
rect 45461 337995 45527 337998
rect 673729 338058 673795 338061
rect 675109 338058 675175 338061
rect 673729 338056 675175 338058
rect 673729 338000 673734 338056
rect 673790 338000 675114 338056
rect 675170 338000 675175 338056
rect 673729 337998 675175 338000
rect 673729 337995 673795 337998
rect 675109 337995 675175 337998
rect 675753 337922 675819 337925
rect 676070 337922 676076 337924
rect 675753 337920 676076 337922
rect 675753 337864 675758 337920
rect 675814 337864 676076 337920
rect 675753 337862 676076 337864
rect 675753 337859 675819 337862
rect 676070 337860 676076 337862
rect 676140 337860 676146 337924
rect 42926 337650 42932 337652
rect 41492 337590 42932 337650
rect 42926 337588 42932 337590
rect 42996 337588 43002 337652
rect 40542 336972 40602 337212
rect 40534 336908 40540 336972
rect 40604 336908 40610 336972
rect 40726 336564 40786 336804
rect 40718 336500 40724 336564
rect 40788 336500 40794 336564
rect 40910 336156 40970 336396
rect 40902 336092 40908 336156
rect 40972 336092 40978 336156
rect 35574 335749 35634 335988
rect 35525 335744 35634 335749
rect 35801 335746 35867 335749
rect 35525 335688 35530 335744
rect 35586 335688 35634 335744
rect 35525 335686 35634 335688
rect 35758 335744 35867 335746
rect 35758 335688 35806 335744
rect 35862 335688 35867 335744
rect 35525 335683 35591 335686
rect 35758 335683 35867 335688
rect 38561 335746 38627 335749
rect 41822 335746 41828 335748
rect 38561 335744 41828 335746
rect 38561 335688 38566 335744
rect 38622 335688 41828 335744
rect 38561 335686 41828 335688
rect 38561 335683 38627 335686
rect 41822 335684 41828 335686
rect 41892 335684 41898 335748
rect 35758 335580 35818 335683
rect 675293 335338 675359 335341
rect 676438 335338 676444 335340
rect 675293 335336 676444 335338
rect 675293 335280 675298 335336
rect 675354 335280 676444 335336
rect 675293 335278 676444 335280
rect 675293 335275 675359 335278
rect 676438 335276 676444 335278
rect 676508 335276 676514 335340
rect 41462 334930 41522 335172
rect 41462 334870 42074 334930
rect 35758 334525 35818 334764
rect 42014 334658 42074 334870
rect 44173 334658 44239 334661
rect 42014 334656 44239 334658
rect 42014 334600 44178 334656
rect 44234 334600 44239 334656
rect 42014 334598 44239 334600
rect 44173 334595 44239 334598
rect 35758 334520 35867 334525
rect 35758 334464 35806 334520
rect 35862 334464 35867 334520
rect 35758 334462 35867 334464
rect 35801 334459 35867 334462
rect 40033 334522 40099 334525
rect 40033 334520 41890 334522
rect 40033 334464 40038 334520
rect 40094 334464 41890 334520
rect 40033 334462 41890 334464
rect 40033 334459 40099 334462
rect 41830 334386 41890 334462
rect 42793 334386 42859 334389
rect 41830 334384 42859 334386
rect 41462 334114 41522 334356
rect 41830 334328 42798 334384
rect 42854 334328 42859 334384
rect 41830 334326 42859 334328
rect 42793 334323 42859 334326
rect 51717 334114 51783 334117
rect 41462 334112 51783 334114
rect 41462 334056 51722 334112
rect 51778 334056 51783 334112
rect 41462 334054 51783 334056
rect 51717 334051 51783 334054
rect 41278 333570 41338 333948
rect 41278 333540 41492 333570
rect 41308 333510 41522 333540
rect 41462 333298 41522 333510
rect 672165 333434 672231 333437
rect 675477 333434 675543 333437
rect 672165 333432 675543 333434
rect 672165 333376 672170 333432
rect 672226 333376 675482 333432
rect 675538 333376 675543 333432
rect 672165 333374 675543 333376
rect 672165 333371 672231 333374
rect 675477 333371 675543 333374
rect 41462 333238 51090 333298
rect 35758 332893 35818 333132
rect 35758 332888 35867 332893
rect 35758 332832 35806 332888
rect 35862 332832 35867 332888
rect 35758 332830 35867 332832
rect 35801 332827 35867 332830
rect 39757 332890 39823 332893
rect 42977 332890 43043 332893
rect 39757 332888 43043 332890
rect 39757 332832 39762 332888
rect 39818 332832 42982 332888
rect 43038 332832 43043 332888
rect 39757 332830 43043 332832
rect 39757 332827 39823 332830
rect 42977 332827 43043 332830
rect 51030 332618 51090 333238
rect 672349 332754 672415 332757
rect 675477 332754 675543 332757
rect 672349 332752 675543 332754
rect 672349 332696 672354 332752
rect 672410 332696 675482 332752
rect 675538 332696 675543 332752
rect 672349 332694 675543 332696
rect 672349 332691 672415 332694
rect 675477 332691 675543 332694
rect 63217 332618 63283 332621
rect 51030 332616 63283 332618
rect 51030 332560 63222 332616
rect 63278 332560 63283 332616
rect 51030 332558 63283 332560
rect 63217 332555 63283 332558
rect 40217 332482 40283 332485
rect 43161 332482 43227 332485
rect 40217 332480 43227 332482
rect 40217 332424 40222 332480
rect 40278 332424 43166 332480
rect 43222 332424 43227 332480
rect 40217 332422 43227 332424
rect 40217 332419 40283 332422
rect 43161 332419 43227 332422
rect 35801 331802 35867 331805
rect 50337 331802 50403 331805
rect 35801 331800 50403 331802
rect 35801 331744 35806 331800
rect 35862 331744 50342 331800
rect 50398 331744 50403 331800
rect 35801 331742 50403 331744
rect 35801 331739 35867 331742
rect 50337 331739 50403 331742
rect 36537 331258 36603 331261
rect 41454 331258 41460 331260
rect 36537 331256 41460 331258
rect 36537 331200 36542 331256
rect 36598 331200 41460 331256
rect 36537 331198 41460 331200
rect 36537 331195 36603 331198
rect 41454 331196 41460 331198
rect 41524 331196 41530 331260
rect 672901 331258 672967 331261
rect 675109 331258 675175 331261
rect 672901 331256 675175 331258
rect 672901 331200 672906 331256
rect 672962 331200 675114 331256
rect 675170 331200 675175 331256
rect 672901 331198 675175 331200
rect 672901 331195 672967 331198
rect 675109 331195 675175 331198
rect 35157 330442 35223 330445
rect 41638 330442 41644 330444
rect 35157 330440 41644 330442
rect 35157 330384 35162 330440
rect 35218 330384 41644 330440
rect 35157 330382 41644 330384
rect 35157 330379 35223 330382
rect 41638 330380 41644 330382
rect 41708 330380 41714 330444
rect 652385 329762 652451 329765
rect 649950 329760 652451 329762
rect 649950 329704 652390 329760
rect 652446 329704 652451 329760
rect 649950 329702 652451 329704
rect 649950 329234 650010 329702
rect 652385 329699 652451 329702
rect 651465 328266 651531 328269
rect 649950 328264 651531 328266
rect 649950 328208 651470 328264
rect 651526 328208 651531 328264
rect 649950 328206 651531 328208
rect 649950 328052 650010 328206
rect 651465 328203 651531 328206
rect 675017 327994 675083 327997
rect 675385 327996 675451 327997
rect 675334 327994 675340 327996
rect 675017 327992 675340 327994
rect 675404 327994 675451 327996
rect 675404 327992 675496 327994
rect 675017 327936 675022 327992
rect 675078 327936 675340 327992
rect 675446 327936 675496 327992
rect 675017 327934 675340 327936
rect 675017 327931 675083 327934
rect 675334 327932 675340 327934
rect 675404 327934 675496 327936
rect 675404 327932 675451 327934
rect 675385 327931 675451 327932
rect 42425 327042 42491 327045
rect 45277 327042 45343 327045
rect 42425 327040 45343 327042
rect 42425 326984 42430 327040
rect 42486 326984 45282 327040
rect 45338 326984 45343 327040
rect 42425 326982 45343 326984
rect 42425 326979 42491 326982
rect 45277 326979 45343 326982
rect 652017 326906 652083 326909
rect 650502 326904 652083 326906
rect 650502 326900 652022 326904
rect 649980 326848 652022 326900
rect 652078 326848 652083 326904
rect 649980 326846 652083 326848
rect 649980 326840 650562 326846
rect 652017 326843 652083 326846
rect 674649 326906 674715 326909
rect 675385 326906 675451 326909
rect 674649 326904 675451 326906
rect 674649 326848 674654 326904
rect 674710 326848 675390 326904
rect 675446 326848 675451 326904
rect 674649 326846 675451 326848
rect 674649 326843 674715 326846
rect 675385 326843 675451 326846
rect 649950 325682 650010 325710
rect 651373 325682 651439 325685
rect 649950 325680 651439 325682
rect 649950 325624 651378 325680
rect 651434 325624 651439 325680
rect 649950 325622 651439 325624
rect 651373 325619 651439 325622
rect 675201 325682 675267 325685
rect 676622 325682 676628 325684
rect 675201 325680 676628 325682
rect 675201 325624 675206 325680
rect 675262 325624 676628 325680
rect 675201 325622 676628 325624
rect 675201 325619 675267 325622
rect 676622 325620 676628 325622
rect 676692 325620 676698 325684
rect 672901 325002 672967 325005
rect 675017 325002 675083 325005
rect 672901 325000 675083 325002
rect 672901 324944 672906 325000
rect 672962 324944 675022 325000
rect 675078 324944 675083 325000
rect 672901 324942 675083 324944
rect 672901 324939 672967 324942
rect 675017 324939 675083 324942
rect 41781 324868 41847 324869
rect 41781 324864 41828 324868
rect 41892 324866 41898 324868
rect 41781 324808 41786 324864
rect 41781 324804 41828 324808
rect 41892 324806 41938 324866
rect 41892 324804 41898 324806
rect 41781 324803 41847 324804
rect 40902 322764 40908 322828
rect 40972 322826 40978 322828
rect 41781 322826 41847 322829
rect 40972 322824 41847 322826
rect 40972 322768 41786 322824
rect 41842 322768 41847 322824
rect 40972 322766 41847 322768
rect 40972 322764 40978 322766
rect 41781 322763 41847 322766
rect 42057 321194 42123 321197
rect 42977 321194 43043 321197
rect 42057 321192 43043 321194
rect 42057 321136 42062 321192
rect 42118 321136 42982 321192
rect 43038 321136 43043 321192
rect 42057 321134 43043 321136
rect 42057 321131 42123 321134
rect 42977 321131 43043 321134
rect 42425 320786 42491 320789
rect 53833 320786 53899 320789
rect 42425 320784 53899 320786
rect 42425 320728 42430 320784
rect 42486 320728 53838 320784
rect 53894 320728 53899 320784
rect 42425 320726 53899 320728
rect 42425 320723 42491 320726
rect 53833 320723 53899 320726
rect 42149 320514 42215 320517
rect 43161 320514 43227 320517
rect 42149 320512 43227 320514
rect 42149 320456 42154 320512
rect 42210 320456 43166 320512
rect 43222 320456 43227 320512
rect 42149 320454 43227 320456
rect 42149 320451 42215 320454
rect 43161 320451 43227 320454
rect 42333 320106 42399 320109
rect 53097 320106 53163 320109
rect 42333 320104 53163 320106
rect 42333 320048 42338 320104
rect 42394 320048 53102 320104
rect 53158 320048 53163 320104
rect 42333 320046 53163 320048
rect 42333 320043 42399 320046
rect 53097 320043 53163 320046
rect 42425 319698 42491 319701
rect 46933 319698 46999 319701
rect 42425 319696 46999 319698
rect 42425 319640 42430 319696
rect 42486 319640 46938 319696
rect 46994 319640 46999 319696
rect 42425 319638 46999 319640
rect 42425 319635 42491 319638
rect 46933 319635 46999 319638
rect 62113 317386 62179 317389
rect 62113 317384 64706 317386
rect 62113 317328 62118 317384
rect 62174 317328 64706 317384
rect 62113 317326 64706 317328
rect 62113 317323 62179 317326
rect 64646 317106 64706 317326
rect 40718 316780 40724 316844
rect 40788 316842 40794 316844
rect 41781 316842 41847 316845
rect 40788 316840 41847 316842
rect 40788 316784 41786 316840
rect 41842 316784 41847 316840
rect 40788 316782 41847 316784
rect 40788 316780 40794 316782
rect 41781 316779 41847 316782
rect 40534 315964 40540 316028
rect 40604 316026 40610 316028
rect 41781 316026 41847 316029
rect 40604 316024 41847 316026
rect 40604 315968 41786 316024
rect 41842 315968 41847 316024
rect 40604 315966 41847 315968
rect 40604 315964 40610 315966
rect 41781 315963 41847 315966
rect 62113 316026 62179 316029
rect 62113 316024 64706 316026
rect 62113 315968 62118 316024
rect 62174 315968 64706 316024
rect 62113 315966 64706 315968
rect 62113 315963 62179 315966
rect 64646 315924 64706 315966
rect 41781 315620 41847 315621
rect 41781 315616 41828 315620
rect 41892 315618 41898 315620
rect 41781 315560 41786 315616
rect 41781 315556 41828 315560
rect 41892 315558 41938 315618
rect 41892 315556 41898 315558
rect 41781 315555 41847 315556
rect 62113 314802 62179 314805
rect 62113 314800 64706 314802
rect 62113 314744 62118 314800
rect 62174 314744 64706 314800
rect 62113 314742 64706 314744
rect 62113 314739 62179 314742
rect 62297 314122 62363 314125
rect 62297 314120 64706 314122
rect 62297 314064 62302 314120
rect 62358 314064 64706 314120
rect 62297 314062 64706 314064
rect 62297 314059 62363 314062
rect 41454 313652 41460 313716
rect 41524 313714 41530 313716
rect 41781 313714 41847 313717
rect 41524 313712 41847 313714
rect 41524 313656 41786 313712
rect 41842 313656 41847 313712
rect 41524 313654 41847 313656
rect 41524 313652 41530 313654
rect 41781 313651 41847 313654
rect 64646 313560 64706 314062
rect 667381 313714 667447 313717
rect 667381 313712 676292 313714
rect 667381 313656 667386 313712
rect 667442 313656 676292 313712
rect 667381 313654 676292 313656
rect 667381 313651 667447 313654
rect 676029 313306 676095 313309
rect 676029 313304 676292 313306
rect 676029 313248 676034 313304
rect 676090 313248 676292 313304
rect 676029 313246 676292 313248
rect 676029 313243 676095 313246
rect 62481 313034 62547 313037
rect 62481 313032 64706 313034
rect 62481 312976 62486 313032
rect 62542 312976 64706 313032
rect 62481 312974 64706 312976
rect 62481 312971 62547 312974
rect 42425 312762 42491 312765
rect 42926 312762 42932 312764
rect 42425 312760 42932 312762
rect 42425 312704 42430 312760
rect 42486 312704 42932 312760
rect 42425 312702 42932 312704
rect 42425 312699 42491 312702
rect 42926 312700 42932 312702
rect 42996 312700 43002 312764
rect 64646 312378 64706 312974
rect 674833 312898 674899 312901
rect 674833 312896 676292 312898
rect 674833 312840 674838 312896
rect 674894 312840 676292 312896
rect 674833 312838 676292 312840
rect 674833 312835 674899 312838
rect 672533 312490 672599 312493
rect 672533 312488 676292 312490
rect 672533 312432 672538 312488
rect 672594 312432 676292 312488
rect 672533 312430 676292 312432
rect 672533 312427 672599 312430
rect 42149 312354 42215 312357
rect 45553 312354 45619 312357
rect 42149 312352 45619 312354
rect 42149 312296 42154 312352
rect 42210 312296 45558 312352
rect 45614 312296 45619 312352
rect 42149 312294 45619 312296
rect 42149 312291 42215 312294
rect 45553 312291 45619 312294
rect 675477 312082 675543 312085
rect 675477 312080 676292 312082
rect 675477 312024 675482 312080
rect 675538 312024 676292 312080
rect 675477 312022 676292 312024
rect 675477 312019 675543 312022
rect 660297 311946 660363 311949
rect 674833 311946 674899 311949
rect 660297 311944 674899 311946
rect 660297 311888 660302 311944
rect 660358 311888 674838 311944
rect 674894 311888 674899 311944
rect 660297 311886 674899 311888
rect 660297 311883 660363 311886
rect 674833 311883 674899 311886
rect 62665 311810 62731 311813
rect 62665 311808 64706 311810
rect 62665 311752 62670 311808
rect 62726 311752 64706 311808
rect 62665 311750 64706 311752
rect 62665 311747 62731 311750
rect 64646 311196 64706 311750
rect 674373 311674 674439 311677
rect 674373 311672 676292 311674
rect 674373 311616 674378 311672
rect 674434 311616 676292 311672
rect 674373 311614 676292 311616
rect 674373 311611 674439 311614
rect 674741 311402 674807 311405
rect 674741 311400 676230 311402
rect 674741 311344 674746 311400
rect 674802 311344 676230 311400
rect 674741 311342 676230 311344
rect 674741 311339 674807 311342
rect 676170 311266 676230 311342
rect 676170 311206 676292 311266
rect 652201 311130 652267 311133
rect 675937 311130 676003 311133
rect 652201 311128 676003 311130
rect 652201 311072 652206 311128
rect 652262 311072 675942 311128
rect 675998 311072 676003 311128
rect 652201 311070 676003 311072
rect 652201 311067 652267 311070
rect 675937 311067 676003 311070
rect 673361 310858 673427 310861
rect 673361 310856 676292 310858
rect 673361 310800 673366 310856
rect 673422 310800 676292 310856
rect 673361 310798 676292 310800
rect 673361 310795 673427 310798
rect 42057 310450 42123 310453
rect 53833 310450 53899 310453
rect 42057 310448 53899 310450
rect 42057 310392 42062 310448
rect 42118 310392 53838 310448
rect 53894 310392 53899 310448
rect 42057 310390 53899 310392
rect 42057 310387 42123 310390
rect 53833 310387 53899 310390
rect 673913 310450 673979 310453
rect 673913 310448 676292 310450
rect 673913 310392 673918 310448
rect 673974 310392 676292 310448
rect 673913 310390 676292 310392
rect 673913 310387 673979 310390
rect 673177 310042 673243 310045
rect 673177 310040 676292 310042
rect 673177 309984 673182 310040
rect 673238 309984 676292 310040
rect 673177 309982 676292 309984
rect 673177 309979 673243 309982
rect 673361 309634 673427 309637
rect 673361 309632 676292 309634
rect 673361 309576 673366 309632
rect 673422 309576 676292 309632
rect 673361 309574 676292 309576
rect 673361 309571 673427 309574
rect 675017 309226 675083 309229
rect 675017 309224 676292 309226
rect 675017 309168 675022 309224
rect 675078 309168 676292 309224
rect 675017 309166 676292 309168
rect 675017 309163 675083 309166
rect 675886 308756 675892 308820
rect 675956 308818 675962 308820
rect 675956 308758 676292 308818
rect 675956 308756 675962 308758
rect 676673 308410 676739 308413
rect 676660 308408 676739 308410
rect 676660 308352 676678 308408
rect 676734 308352 676739 308408
rect 676660 308350 676739 308352
rect 676673 308347 676739 308350
rect 675477 308002 675543 308005
rect 675477 308000 676292 308002
rect 675477 307944 675482 308000
rect 675538 307944 676292 308000
rect 675477 307942 676292 307944
rect 675477 307939 675543 307942
rect 676029 307594 676095 307597
rect 676029 307592 676292 307594
rect 676029 307536 676034 307592
rect 676090 307536 676292 307592
rect 676029 307534 676292 307536
rect 676029 307531 676095 307534
rect 676029 307186 676095 307189
rect 676029 307184 676292 307186
rect 676029 307128 676034 307184
rect 676090 307128 676292 307184
rect 676029 307126 676292 307128
rect 676029 307123 676095 307126
rect 678237 306778 678303 306781
rect 678237 306776 678316 306778
rect 678237 306720 678242 306776
rect 678298 306720 678316 306776
rect 678237 306718 678316 306720
rect 678237 306715 678303 306718
rect 678973 306370 679039 306373
rect 678973 306368 679052 306370
rect 678973 306312 678978 306368
rect 679034 306312 679052 306368
rect 678973 306310 679052 306312
rect 678973 306307 679039 306310
rect 673729 305962 673795 305965
rect 673729 305960 676292 305962
rect 673729 305904 673734 305960
rect 673790 305904 676292 305960
rect 673729 305902 676292 305904
rect 673729 305899 673795 305902
rect 674373 305554 674439 305557
rect 674373 305552 676292 305554
rect 674373 305496 674378 305552
rect 674434 305496 676292 305552
rect 674373 305494 676292 305496
rect 674373 305491 674439 305494
rect 675894 305086 676292 305146
rect 675894 304602 675954 305086
rect 676397 304738 676463 304741
rect 676397 304736 676476 304738
rect 676397 304680 676402 304736
rect 676458 304680 676476 304736
rect 676397 304678 676476 304680
rect 676397 304675 676463 304678
rect 676070 304602 676076 304604
rect 675894 304542 676076 304602
rect 676070 304540 676076 304542
rect 676140 304540 676146 304604
rect 672533 304330 672599 304333
rect 672533 304328 676292 304330
rect 672533 304272 672538 304328
rect 672594 304272 676292 304328
rect 672533 304270 676292 304272
rect 672533 304267 672599 304270
rect 673177 303922 673243 303925
rect 673177 303920 676292 303922
rect 673177 303864 673182 303920
rect 673238 303864 676292 303920
rect 673177 303862 676292 303864
rect 673177 303859 673243 303862
rect 674465 303514 674531 303517
rect 674465 303512 676292 303514
rect 674465 303456 674470 303512
rect 674526 303456 676292 303512
rect 674465 303454 676292 303456
rect 674465 303451 674531 303454
rect 652201 303378 652267 303381
rect 649950 303376 652267 303378
rect 649950 303320 652206 303376
rect 652262 303320 652267 303376
rect 649950 303318 652267 303320
rect 649950 302776 650010 303318
rect 652201 303315 652267 303318
rect 675886 302636 675892 302700
rect 675956 302698 675962 302700
rect 676262 302698 676322 303076
rect 675956 302668 676322 302698
rect 675956 302638 676292 302668
rect 675956 302636 675962 302638
rect 676262 302250 676322 302260
rect 676078 302190 676322 302250
rect 669957 302154 670023 302157
rect 676078 302154 676138 302190
rect 669957 302152 676138 302154
rect 669957 302096 669962 302152
rect 670018 302096 676138 302152
rect 669957 302094 676138 302096
rect 669957 302091 670023 302094
rect 651465 301882 651531 301885
rect 649950 301880 651531 301882
rect 649950 301824 651470 301880
rect 651526 301824 651531 301880
rect 649950 301822 651531 301824
rect 649950 301594 650010 301822
rect 651465 301819 651531 301822
rect 676397 301612 676463 301613
rect 676397 301608 676444 301612
rect 676508 301610 676514 301612
rect 676397 301552 676402 301608
rect 676397 301548 676444 301552
rect 676508 301550 676554 301610
rect 676508 301548 676514 301550
rect 676397 301547 676463 301548
rect 676673 301476 676739 301477
rect 676622 301412 676628 301476
rect 676692 301474 676739 301476
rect 676692 301472 676784 301474
rect 676734 301416 676784 301472
rect 676692 301414 676784 301416
rect 676692 301412 676739 301414
rect 676673 301411 676739 301412
rect 41492 301278 51090 301338
rect 35617 300930 35683 300933
rect 35604 300928 35683 300930
rect 35604 300872 35622 300928
rect 35678 300872 35683 300928
rect 35604 300870 35683 300872
rect 51030 300930 51090 301278
rect 59997 300930 60063 300933
rect 51030 300928 60063 300930
rect 51030 300872 60002 300928
rect 60058 300872 60063 300928
rect 51030 300870 60063 300872
rect 35617 300867 35683 300870
rect 59997 300867 60063 300870
rect 668761 300794 668827 300797
rect 674465 300794 674531 300797
rect 668761 300792 674531 300794
rect 668761 300736 668766 300792
rect 668822 300736 674470 300792
rect 674526 300736 674531 300792
rect 668761 300734 674531 300736
rect 668761 300731 668827 300734
rect 674465 300731 674531 300734
rect 651465 300658 651531 300661
rect 649950 300656 651531 300658
rect 649950 300600 651470 300656
rect 651526 300600 651531 300656
rect 649950 300598 651531 300600
rect 46197 300522 46263 300525
rect 41492 300520 46263 300522
rect 41492 300464 46202 300520
rect 46258 300464 46263 300520
rect 41492 300462 46263 300464
rect 46197 300459 46263 300462
rect 649950 300412 650010 300598
rect 651465 300595 651531 300598
rect 44214 300114 44220 300116
rect 41492 300054 44220 300114
rect 44214 300052 44220 300054
rect 44284 300052 44290 300116
rect 44173 299706 44239 299709
rect 41492 299704 44239 299706
rect 41492 299648 44178 299704
rect 44234 299648 44239 299704
rect 41492 299646 44239 299648
rect 44173 299643 44239 299646
rect 44398 299298 44404 299300
rect 41492 299238 44404 299298
rect 44398 299236 44404 299238
rect 44468 299236 44474 299300
rect 35801 298890 35867 298893
rect 35788 298888 35867 298890
rect 35788 298832 35806 298888
rect 35862 298832 35867 298888
rect 35788 298830 35867 298832
rect 35801 298827 35867 298830
rect 41781 298754 41847 298757
rect 62665 298754 62731 298757
rect 41781 298752 62731 298754
rect 41781 298696 41786 298752
rect 41842 298696 62670 298752
rect 62726 298696 62731 298752
rect 41781 298694 62731 298696
rect 41781 298691 41847 298694
rect 62665 298691 62731 298694
rect 649950 298618 650010 299230
rect 652569 298618 652635 298621
rect 649950 298616 652635 298618
rect 649950 298560 652574 298616
rect 652630 298560 652635 298616
rect 649950 298558 652635 298560
rect 652569 298555 652635 298558
rect 44582 298482 44588 298484
rect 41492 298422 44588 298482
rect 44582 298420 44588 298422
rect 44652 298420 44658 298484
rect 44633 298074 44699 298077
rect 41492 298072 44699 298074
rect 41492 298016 44638 298072
rect 44694 298016 44699 298072
rect 41492 298014 44699 298016
rect 44633 298011 44699 298014
rect 42742 297666 42748 297668
rect 41492 297606 42748 297666
rect 42742 297604 42748 297606
rect 42812 297604 42818 297668
rect 649950 297530 650010 298048
rect 651741 297530 651807 297533
rect 649950 297528 651807 297530
rect 649950 297472 651746 297528
rect 651802 297472 651807 297528
rect 649950 297470 651807 297472
rect 651741 297467 651807 297470
rect 41781 297394 41847 297397
rect 42793 297394 42859 297397
rect 674833 297396 674899 297397
rect 41781 297392 42859 297394
rect 41781 297336 41786 297392
rect 41842 297336 42798 297392
rect 42854 297336 42859 297392
rect 41781 297334 42859 297336
rect 41781 297331 41847 297334
rect 42793 297331 42859 297334
rect 674782 297332 674788 297396
rect 674852 297394 674899 297396
rect 674852 297392 674944 297394
rect 674894 297336 674944 297392
rect 674852 297334 674944 297336
rect 674852 297332 674899 297334
rect 675702 297332 675708 297396
rect 675772 297394 675778 297396
rect 676857 297394 676923 297397
rect 675772 297392 676923 297394
rect 675772 297336 676862 297392
rect 676918 297336 676923 297392
rect 675772 297334 676923 297336
rect 675772 297332 675778 297334
rect 674833 297331 674899 297332
rect 676857 297331 676923 297334
rect 35801 297258 35867 297261
rect 35788 297256 35867 297258
rect 35788 297200 35806 297256
rect 35862 297200 35867 297256
rect 35788 297198 35867 297200
rect 35801 297195 35867 297198
rect 675201 296986 675267 296989
rect 676121 296986 676187 296989
rect 675201 296984 676187 296986
rect 675201 296928 675206 296984
rect 675262 296928 676126 296984
rect 676182 296928 676187 296984
rect 675201 296926 676187 296928
rect 675201 296923 675267 296926
rect 676121 296923 676187 296926
rect 42006 296850 42012 296852
rect 41492 296790 42012 296850
rect 42006 296788 42012 296790
rect 42076 296788 42082 296852
rect 649950 296850 650010 296866
rect 651741 296850 651807 296853
rect 649950 296848 651807 296850
rect 649950 296792 651746 296848
rect 651802 296792 651807 296848
rect 649950 296790 651807 296792
rect 651741 296787 651807 296790
rect 41781 296578 41847 296581
rect 43161 296578 43227 296581
rect 41781 296576 43227 296578
rect 41781 296520 41786 296576
rect 41842 296520 43166 296576
rect 43222 296520 43227 296576
rect 41781 296518 43227 296520
rect 41781 296515 41847 296518
rect 43161 296515 43227 296518
rect 675518 296516 675524 296580
rect 675588 296578 675594 296580
rect 675937 296578 676003 296581
rect 675588 296576 676003 296578
rect 675588 296520 675942 296576
rect 675998 296520 676003 296576
rect 675588 296518 676003 296520
rect 675588 296516 675594 296518
rect 675937 296515 676003 296518
rect 35433 296442 35499 296445
rect 35420 296440 35499 296442
rect 35420 296384 35438 296440
rect 35494 296384 35499 296440
rect 35420 296382 35499 296384
rect 35433 296379 35499 296382
rect 35617 296034 35683 296037
rect 35604 296032 35683 296034
rect 35604 295976 35622 296032
rect 35678 295976 35683 296032
rect 35604 295974 35683 295976
rect 35617 295971 35683 295974
rect 675753 295762 675819 295765
rect 676622 295762 676628 295764
rect 675753 295760 676628 295762
rect 675753 295704 675758 295760
rect 675814 295704 676628 295760
rect 675753 295702 676628 295704
rect 675753 295699 675819 295702
rect 676622 295700 676628 295702
rect 676692 295700 676698 295764
rect 35801 295626 35867 295629
rect 35788 295624 35867 295626
rect 35788 295568 35806 295624
rect 35862 295568 35867 295624
rect 35788 295566 35867 295568
rect 35801 295563 35867 295566
rect 61561 295354 61627 295357
rect 64646 295354 64706 295684
rect 61561 295352 64706 295354
rect 61561 295296 61566 295352
rect 61622 295296 64706 295352
rect 61561 295294 64706 295296
rect 649950 295354 650010 295684
rect 651649 295354 651715 295357
rect 649950 295352 651715 295354
rect 649950 295296 651654 295352
rect 651710 295296 651715 295352
rect 649950 295294 651715 295296
rect 61561 295291 61627 295294
rect 651649 295291 651715 295294
rect 35801 295218 35867 295221
rect 35788 295216 35867 295218
rect 35788 295160 35806 295216
rect 35862 295160 35867 295216
rect 35788 295158 35867 295160
rect 35801 295155 35867 295158
rect 31017 294810 31083 294813
rect 31004 294808 31083 294810
rect 31004 294752 31022 294808
rect 31078 294752 31083 294808
rect 31004 294750 31083 294752
rect 31017 294747 31083 294750
rect 44357 294402 44423 294405
rect 41492 294400 44423 294402
rect 41492 294344 44362 294400
rect 44418 294344 44423 294400
rect 41492 294342 44423 294344
rect 44357 294339 44423 294342
rect 62205 294266 62271 294269
rect 64646 294266 64706 294502
rect 62205 294264 64706 294266
rect 62205 294208 62210 294264
rect 62266 294208 64706 294264
rect 62205 294206 64706 294208
rect 649950 294266 650010 294502
rect 651465 294266 651531 294269
rect 649950 294264 651531 294266
rect 649950 294208 651470 294264
rect 651526 294208 651531 294264
rect 649950 294206 651531 294208
rect 62205 294203 62271 294206
rect 651465 294203 651531 294206
rect 44817 293994 44883 293997
rect 41492 293992 44883 293994
rect 41492 293936 44822 293992
rect 44878 293936 44883 293992
rect 41492 293934 44883 293936
rect 44817 293931 44883 293934
rect 652845 293858 652911 293861
rect 674465 293858 674531 293861
rect 652845 293856 674531 293858
rect 652845 293800 652850 293856
rect 652906 293800 674470 293856
rect 674526 293800 674531 293856
rect 652845 293798 674531 293800
rect 652845 293795 652911 293798
rect 674465 293795 674531 293798
rect 35801 293586 35867 293589
rect 35788 293584 35867 293586
rect 35788 293528 35806 293584
rect 35862 293528 35867 293584
rect 35788 293526 35867 293528
rect 35801 293523 35867 293526
rect 41822 293178 41828 293180
rect 41492 293118 41828 293178
rect 41822 293116 41828 293118
rect 41892 293116 41898 293180
rect 35801 292770 35867 292773
rect 35788 292768 35867 292770
rect 35788 292712 35806 292768
rect 35862 292712 35867 292768
rect 35788 292710 35867 292712
rect 35801 292707 35867 292710
rect 62297 292770 62363 292773
rect 64646 292770 64706 293320
rect 62297 292768 64706 292770
rect 62297 292712 62302 292768
rect 62358 292712 64706 292768
rect 62297 292710 64706 292712
rect 649950 292770 650010 293320
rect 674782 292844 674788 292908
rect 674852 292906 674858 292908
rect 675385 292906 675451 292909
rect 674852 292904 675451 292906
rect 674852 292848 675390 292904
rect 675446 292848 675451 292904
rect 674852 292846 675451 292848
rect 674852 292844 674858 292846
rect 675385 292843 675451 292846
rect 652385 292770 652451 292773
rect 649950 292768 652451 292770
rect 649950 292712 652390 292768
rect 652446 292712 652451 292768
rect 649950 292710 652451 292712
rect 62297 292707 62363 292710
rect 652385 292707 652451 292710
rect 40769 292592 40835 292593
rect 40534 292528 40540 292592
rect 40604 292528 40610 292592
rect 40718 292528 40724 292592
rect 40788 292590 40835 292592
rect 40788 292588 40880 292590
rect 40830 292532 40880 292588
rect 40788 292530 40880 292532
rect 40788 292528 40835 292530
rect 40542 292332 40602 292528
rect 40769 292527 40835 292528
rect 41781 292500 41847 292501
rect 41781 292496 41828 292500
rect 41892 292498 41898 292500
rect 62113 292498 62179 292501
rect 41781 292440 41786 292496
rect 41781 292436 41828 292440
rect 41892 292438 41938 292498
rect 62113 292496 64706 292498
rect 62113 292440 62118 292496
rect 62174 292440 64706 292496
rect 62113 292438 64706 292440
rect 41892 292436 41898 292438
rect 41781 292435 41847 292436
rect 62113 292435 62179 292438
rect 41781 292226 41847 292229
rect 42977 292226 43043 292229
rect 41781 292224 43043 292226
rect 41781 292168 41786 292224
rect 41842 292168 42982 292224
rect 43038 292168 43043 292224
rect 41781 292166 43043 292168
rect 41781 292163 41847 292166
rect 42977 292163 43043 292166
rect 64646 292138 64706 292438
rect 675569 292228 675635 292229
rect 675518 292164 675524 292228
rect 675588 292226 675635 292228
rect 675588 292224 675680 292226
rect 675630 292168 675680 292224
rect 675588 292166 675680 292168
rect 675588 292164 675635 292166
rect 675569 292163 675635 292164
rect 41781 291954 41847 291957
rect 41492 291952 41847 291954
rect 41492 291896 41786 291952
rect 41842 291896 41847 291952
rect 41492 291894 41847 291896
rect 41781 291891 41847 291894
rect 45001 291546 45067 291549
rect 41492 291544 45067 291546
rect 41492 291488 45006 291544
rect 45062 291488 45067 291544
rect 41492 291486 45067 291488
rect 649950 291546 650010 292138
rect 652201 291546 652267 291549
rect 649950 291544 652267 291546
rect 649950 291488 652206 291544
rect 652262 291488 652267 291544
rect 649950 291486 652267 291488
rect 45001 291483 45067 291486
rect 652201 291483 652267 291486
rect 673729 291546 673795 291549
rect 675477 291546 675543 291549
rect 673729 291544 675543 291546
rect 673729 291488 673734 291544
rect 673790 291488 675482 291544
rect 675538 291488 675543 291544
rect 673729 291486 675543 291488
rect 673729 291483 673795 291486
rect 675477 291483 675543 291486
rect 42149 291376 42215 291379
rect 41462 291374 42215 291376
rect 41462 291318 42154 291374
rect 42210 291318 42215 291374
rect 41462 291316 42215 291318
rect 41462 291108 41522 291316
rect 42149 291313 42215 291316
rect 41781 291138 41847 291141
rect 43621 291138 43687 291141
rect 41781 291136 43687 291138
rect 41781 291080 41786 291136
rect 41842 291080 43626 291136
rect 43682 291080 43687 291136
rect 41781 291078 43687 291080
rect 41781 291075 41847 291078
rect 43621 291075 43687 291078
rect 62297 291002 62363 291005
rect 675753 291002 675819 291005
rect 676438 291002 676444 291004
rect 62297 291000 64154 291002
rect 62297 290944 62302 291000
rect 62358 290986 64154 291000
rect 675753 291000 676444 291002
rect 62358 290944 64676 290986
rect 62297 290942 64676 290944
rect 62297 290939 62363 290942
rect 64094 290926 64676 290942
rect 50521 290730 50587 290733
rect 41492 290728 50587 290730
rect 41492 290672 50526 290728
rect 50582 290672 50587 290728
rect 41492 290670 50587 290672
rect 50521 290667 50587 290670
rect 649950 290458 650010 290956
rect 675753 290944 675758 291000
rect 675814 290944 676444 291000
rect 675753 290942 676444 290944
rect 675753 290939 675819 290942
rect 676438 290940 676444 290942
rect 676508 290940 676514 291004
rect 651465 290458 651531 290461
rect 649950 290456 651531 290458
rect 649950 290400 651470 290456
rect 651526 290400 651531 290456
rect 649950 290398 651531 290400
rect 651465 290395 651531 290398
rect 651649 290458 651715 290461
rect 673545 290458 673611 290461
rect 651649 290456 673611 290458
rect 651649 290400 651654 290456
rect 651710 290400 673550 290456
rect 673606 290400 673611 290456
rect 651649 290398 673611 290400
rect 651649 290395 651715 290398
rect 673545 290395 673611 290398
rect 35801 290322 35867 290325
rect 35788 290320 35867 290322
rect 35788 290264 35806 290320
rect 35862 290264 35867 290320
rect 35788 290262 35867 290264
rect 35801 290259 35867 290262
rect 48957 289914 49023 289917
rect 41492 289912 49023 289914
rect 41492 289856 48962 289912
rect 49018 289856 49023 289912
rect 41492 289854 49023 289856
rect 48957 289851 49023 289854
rect 62665 289778 62731 289781
rect 62665 289776 64706 289778
rect 62665 289720 62670 289776
rect 62726 289720 64706 289776
rect 62665 289718 64706 289720
rect 62665 289715 62731 289718
rect 649950 289234 650010 289774
rect 651649 289234 651715 289237
rect 649950 289232 651715 289234
rect 649950 289176 651654 289232
rect 651710 289176 651715 289232
rect 649950 289174 651715 289176
rect 651649 289171 651715 289174
rect 651465 288690 651531 288693
rect 649950 288688 651531 288690
rect 649950 288632 651470 288688
rect 651526 288632 651531 288688
rect 649950 288630 651531 288632
rect 649950 288592 650010 288630
rect 651465 288627 651531 288630
rect 62113 288554 62179 288557
rect 64646 288554 64706 288592
rect 62113 288552 64706 288554
rect 62113 288496 62118 288552
rect 62174 288496 64706 288552
rect 62113 288494 64706 288496
rect 62113 288491 62179 288494
rect 672533 287874 672599 287877
rect 675109 287874 675175 287877
rect 672533 287872 675175 287874
rect 672533 287816 672538 287872
rect 672594 287816 675114 287872
rect 675170 287816 675175 287872
rect 672533 287814 675175 287816
rect 672533 287811 672599 287814
rect 675109 287811 675175 287814
rect 62389 287194 62455 287197
rect 64646 287194 64706 287410
rect 62389 287192 64706 287194
rect 62389 287136 62394 287192
rect 62450 287136 64706 287192
rect 62389 287134 64706 287136
rect 649950 287194 650010 287410
rect 652017 287194 652083 287197
rect 649950 287192 652083 287194
rect 649950 287136 652022 287192
rect 652078 287136 652083 287192
rect 649950 287134 652083 287136
rect 62389 287131 62455 287134
rect 652017 287131 652083 287134
rect 675753 287058 675819 287061
rect 676254 287058 676260 287060
rect 675753 287056 676260 287058
rect 675753 287000 675758 287056
rect 675814 287000 676260 287056
rect 675753 286998 676260 287000
rect 675753 286995 675819 286998
rect 676254 286996 676260 286998
rect 676324 286996 676330 287060
rect 673177 286514 673243 286517
rect 675385 286514 675451 286517
rect 673177 286512 675451 286514
rect 673177 286456 673182 286512
rect 673238 286456 675390 286512
rect 675446 286456 675451 286512
rect 673177 286454 675451 286456
rect 673177 286451 673243 286454
rect 675385 286451 675451 286454
rect 62113 285970 62179 285973
rect 64646 285970 64706 286228
rect 62113 285968 64706 285970
rect 62113 285912 62118 285968
rect 62174 285912 64706 285968
rect 62113 285910 64706 285912
rect 649950 285970 650010 286228
rect 651465 285970 651531 285973
rect 649950 285968 651531 285970
rect 649950 285912 651470 285968
rect 651526 285912 651531 285968
rect 649950 285910 651531 285912
rect 62113 285907 62179 285910
rect 651465 285907 651531 285910
rect 672257 285698 672323 285701
rect 672809 285698 672875 285701
rect 672257 285696 672875 285698
rect 672257 285640 672262 285696
rect 672318 285640 672814 285696
rect 672870 285640 672875 285696
rect 672257 285638 672875 285640
rect 672257 285635 672323 285638
rect 672809 285635 672875 285638
rect 62941 284610 63007 284613
rect 64646 284610 64706 285046
rect 649950 284746 650010 285046
rect 651465 284746 651531 284749
rect 649950 284744 651531 284746
rect 649950 284688 651470 284744
rect 651526 284688 651531 284744
rect 649950 284686 651531 284688
rect 651465 284683 651531 284686
rect 62941 284608 64706 284610
rect 62941 284552 62946 284608
rect 63002 284552 64706 284608
rect 62941 284550 64706 284552
rect 62941 284547 63007 284550
rect 39297 284338 39363 284341
rect 42006 284338 42012 284340
rect 39297 284336 42012 284338
rect 39297 284280 39302 284336
rect 39358 284280 42012 284336
rect 39297 284278 42012 284280
rect 39297 284275 39363 284278
rect 42006 284276 42012 284278
rect 42076 284276 42082 284340
rect 62665 283250 62731 283253
rect 64646 283250 64706 283864
rect 649950 283522 650010 283864
rect 675753 283658 675819 283661
rect 676070 283658 676076 283660
rect 675753 283656 676076 283658
rect 675753 283600 675758 283656
rect 675814 283600 676076 283656
rect 675753 283598 676076 283600
rect 675753 283595 675819 283598
rect 676070 283596 676076 283598
rect 676140 283596 676146 283660
rect 651465 283522 651531 283525
rect 649950 283520 651531 283522
rect 649950 283464 651470 283520
rect 651526 283464 651531 283520
rect 649950 283462 651531 283464
rect 651465 283459 651531 283462
rect 62665 283248 64706 283250
rect 62665 283192 62670 283248
rect 62726 283192 64706 283248
rect 62665 283190 64706 283192
rect 62665 283187 62731 283190
rect 675661 282706 675727 282709
rect 675886 282706 675892 282708
rect 675661 282704 675892 282706
rect 62205 282162 62271 282165
rect 64646 282162 64706 282682
rect 62205 282160 64706 282162
rect 62205 282104 62210 282160
rect 62266 282104 64706 282160
rect 62205 282102 64706 282104
rect 649950 282162 650010 282682
rect 675661 282648 675666 282704
rect 675722 282648 675892 282704
rect 675661 282646 675892 282648
rect 675661 282643 675727 282646
rect 675886 282644 675892 282646
rect 675956 282644 675962 282708
rect 651465 282162 651531 282165
rect 649950 282160 651531 282162
rect 649950 282104 651470 282160
rect 651526 282104 651531 282160
rect 649950 282102 651531 282104
rect 62205 282099 62271 282102
rect 651465 282099 651531 282102
rect 675661 281620 675727 281621
rect 675661 281616 675708 281620
rect 675772 281618 675778 281620
rect 675661 281560 675666 281616
rect 675661 281556 675708 281560
rect 675772 281558 675818 281618
rect 675772 281556 675778 281558
rect 675661 281555 675727 281556
rect 62113 280938 62179 280941
rect 64646 280938 64706 281500
rect 62113 280936 64706 280938
rect 62113 280880 62118 280936
rect 62174 280880 64706 280936
rect 62113 280878 64706 280880
rect 649950 280938 650010 281500
rect 651465 280938 651531 280941
rect 649950 280936 651531 280938
rect 649950 280880 651470 280936
rect 651526 280880 651531 280936
rect 649950 280878 651531 280880
rect 62113 280875 62179 280878
rect 651465 280875 651531 280878
rect 61377 280394 61443 280397
rect 652569 280394 652635 280397
rect 61377 280392 64706 280394
rect 61377 280336 61382 280392
rect 61438 280336 64706 280392
rect 61377 280334 64706 280336
rect 61377 280331 61443 280334
rect 64646 280318 64706 280334
rect 649950 280392 652635 280394
rect 649950 280336 652574 280392
rect 652630 280336 652635 280392
rect 649950 280334 652635 280336
rect 649950 280318 650010 280334
rect 652569 280331 652635 280334
rect 40902 279788 40908 279852
rect 40972 279850 40978 279852
rect 41781 279850 41847 279853
rect 40972 279848 41847 279850
rect 40972 279792 41786 279848
rect 41842 279792 41847 279848
rect 40972 279790 41847 279792
rect 40972 279788 40978 279790
rect 41781 279787 41847 279790
rect 651833 279442 651899 279445
rect 676857 279442 676923 279445
rect 651833 279440 676923 279442
rect 651833 279384 651838 279440
rect 651894 279384 676862 279440
rect 676918 279384 676923 279440
rect 651833 279382 676923 279384
rect 651833 279379 651899 279382
rect 676857 279379 676923 279382
rect 42425 278762 42491 278765
rect 61561 278762 61627 278765
rect 42425 278760 61627 278762
rect 42425 278704 42430 278760
rect 42486 278704 61566 278760
rect 61622 278704 61627 278760
rect 42425 278702 61627 278704
rect 42425 278699 42491 278702
rect 61561 278699 61627 278702
rect 63401 278762 63467 278765
rect 63401 278760 663810 278762
rect 63401 278704 63406 278760
rect 63462 278704 663810 278760
rect 63401 278702 663810 278704
rect 63401 278699 63467 278702
rect 42057 278490 42123 278493
rect 45001 278490 45067 278493
rect 42057 278488 45067 278490
rect 42057 278432 42062 278488
rect 42118 278432 45006 278488
rect 45062 278432 45067 278488
rect 42057 278430 45067 278432
rect 42057 278427 42123 278430
rect 45001 278427 45067 278430
rect 663750 278354 663810 278702
rect 675109 278354 675175 278357
rect 663750 278352 675175 278354
rect 663750 278296 675114 278352
rect 675170 278296 675175 278352
rect 663750 278294 675175 278296
rect 675109 278291 675175 278294
rect 42057 277946 42123 277949
rect 42977 277946 43043 277949
rect 42057 277944 43043 277946
rect 42057 277888 42062 277944
rect 42118 277888 42982 277944
rect 43038 277888 43043 277944
rect 42057 277886 43043 277888
rect 42057 277883 42123 277886
rect 42977 277883 43043 277886
rect 40718 277068 40724 277132
rect 40788 277130 40794 277132
rect 41781 277130 41847 277133
rect 40788 277128 41847 277130
rect 40788 277072 41786 277128
rect 41842 277072 41847 277128
rect 40788 277070 41847 277072
rect 40788 277068 40794 277070
rect 41781 277067 41847 277070
rect 42057 276722 42123 276725
rect 42609 276722 42675 276725
rect 42057 276720 42675 276722
rect 42057 276664 42062 276720
rect 42118 276664 42614 276720
rect 42670 276664 42675 276720
rect 42057 276662 42675 276664
rect 42057 276659 42123 276662
rect 42609 276659 42675 276662
rect 42241 275906 42307 275909
rect 53097 275906 53163 275909
rect 42241 275904 53163 275906
rect 42241 275848 42246 275904
rect 42302 275848 53102 275904
rect 53158 275848 53163 275904
rect 42241 275846 53163 275848
rect 42241 275843 42307 275846
rect 53097 275843 53163 275846
rect 40534 274212 40540 274276
rect 40604 274274 40610 274276
rect 41781 274274 41847 274277
rect 40604 274272 41847 274274
rect 40604 274216 41786 274272
rect 41842 274216 41847 274272
rect 40604 274214 41847 274216
rect 40604 274212 40610 274214
rect 41781 274211 41847 274214
rect 539317 274002 539383 274005
rect 545941 274002 546007 274005
rect 539317 274000 546007 274002
rect 539317 273944 539322 274000
rect 539378 273944 545946 274000
rect 546002 273944 546007 274000
rect 539317 273942 546007 273944
rect 539317 273939 539383 273942
rect 545941 273939 546007 273942
rect 42333 273186 42399 273189
rect 43621 273186 43687 273189
rect 42333 273184 43687 273186
rect 42333 273128 42338 273184
rect 42394 273128 43626 273184
rect 43682 273128 43687 273184
rect 42333 273126 43687 273128
rect 42333 273123 42399 273126
rect 43621 273123 43687 273126
rect 499481 273050 499547 273053
rect 503345 273050 503411 273053
rect 499481 273048 503411 273050
rect 499481 272992 499486 273048
rect 499542 272992 503350 273048
rect 503406 272992 503411 273048
rect 499481 272990 503411 272992
rect 499481 272987 499547 272990
rect 503345 272987 503411 272990
rect 42425 272914 42491 272917
rect 44817 272914 44883 272917
rect 42425 272912 44883 272914
rect 42425 272856 42430 272912
rect 42486 272856 44822 272912
rect 44878 272856 44883 272912
rect 42425 272854 44883 272856
rect 42425 272851 42491 272854
rect 44817 272851 44883 272854
rect 461025 272914 461091 272917
rect 466269 272914 466335 272917
rect 461025 272912 466335 272914
rect 461025 272856 461030 272912
rect 461086 272856 466274 272912
rect 466330 272856 466335 272912
rect 461025 272854 466335 272856
rect 461025 272851 461091 272854
rect 466269 272851 466335 272854
rect 460841 272642 460907 272645
rect 461853 272642 461919 272645
rect 460841 272640 461919 272642
rect 460841 272584 460846 272640
rect 460902 272584 461858 272640
rect 461914 272584 461919 272640
rect 460841 272582 461919 272584
rect 460841 272579 460907 272582
rect 461853 272579 461919 272582
rect 489913 272642 489979 272645
rect 499665 272642 499731 272645
rect 489913 272640 499731 272642
rect 489913 272584 489918 272640
rect 489974 272584 499670 272640
rect 499726 272584 499731 272640
rect 489913 272582 499731 272584
rect 489913 272579 489979 272582
rect 499665 272579 499731 272582
rect 464705 272506 464771 272509
rect 470685 272506 470751 272509
rect 464705 272504 470751 272506
rect 464705 272448 464710 272504
rect 464766 272448 470690 272504
rect 470746 272448 470751 272504
rect 464705 272446 470751 272448
rect 464705 272443 464771 272446
rect 470685 272443 470751 272446
rect 536557 272506 536623 272509
rect 547689 272506 547755 272509
rect 536557 272504 547755 272506
rect 536557 272448 536562 272504
rect 536618 272448 547694 272504
rect 547750 272448 547755 272504
rect 536557 272446 547755 272448
rect 536557 272443 536623 272446
rect 547689 272443 547755 272446
rect 41781 272372 41847 272373
rect 41781 272368 41828 272372
rect 41892 272370 41898 272372
rect 480253 272370 480319 272373
rect 484853 272370 484919 272373
rect 41781 272312 41786 272368
rect 41781 272308 41828 272312
rect 41892 272310 41938 272370
rect 480253 272368 484919 272370
rect 480253 272312 480258 272368
rect 480314 272312 484858 272368
rect 484914 272312 484919 272368
rect 480253 272310 484919 272312
rect 41892 272308 41898 272310
rect 41781 272307 41847 272308
rect 480253 272307 480319 272310
rect 484853 272307 484919 272310
rect 470547 271962 470613 271965
rect 478045 271962 478111 271965
rect 470547 271960 478111 271962
rect 470547 271904 470552 271960
rect 470608 271904 478050 271960
rect 478106 271904 478111 271960
rect 470547 271902 478111 271904
rect 470547 271899 470613 271902
rect 478045 271899 478111 271902
rect 547505 271962 547571 271965
rect 547873 271962 547939 271965
rect 547505 271960 547939 271962
rect 547505 271904 547510 271960
rect 547566 271904 547878 271960
rect 547934 271904 547939 271960
rect 547505 271902 547939 271904
rect 547505 271899 547571 271902
rect 547873 271899 547939 271902
rect 479517 271826 479583 271829
rect 483197 271826 483263 271829
rect 479517 271824 483263 271826
rect 479517 271768 479522 271824
rect 479578 271768 483202 271824
rect 483258 271768 483263 271824
rect 479517 271766 483263 271768
rect 479517 271763 479583 271766
rect 483197 271763 483263 271766
rect 41454 270404 41460 270468
rect 41524 270466 41530 270468
rect 41781 270466 41847 270469
rect 41524 270464 41847 270466
rect 41524 270408 41786 270464
rect 41842 270408 41847 270464
rect 41524 270406 41847 270408
rect 41524 270404 41530 270406
rect 41781 270403 41847 270406
rect 42425 270466 42491 270469
rect 44357 270466 44423 270469
rect 42425 270464 44423 270466
rect 42425 270408 42430 270464
rect 42486 270408 44362 270464
rect 44418 270408 44423 270464
rect 42425 270406 44423 270408
rect 42425 270403 42491 270406
rect 44357 270403 44423 270406
rect 532233 270194 532299 270197
rect 534073 270194 534139 270197
rect 532233 270192 534139 270194
rect 532233 270136 532238 270192
rect 532294 270136 534078 270192
rect 534134 270136 534139 270192
rect 532233 270134 534139 270136
rect 532233 270131 532299 270134
rect 534073 270131 534139 270134
rect 509233 269922 509299 269925
rect 516501 269922 516567 269925
rect 509233 269920 516567 269922
rect 509233 269864 509238 269920
rect 509294 269864 516506 269920
rect 516562 269864 516567 269920
rect 509233 269862 516567 269864
rect 509233 269859 509299 269862
rect 516501 269859 516567 269862
rect 538029 269786 538095 269789
rect 541801 269786 541867 269789
rect 538029 269784 541867 269786
rect 538029 269728 538034 269784
rect 538090 269728 541806 269784
rect 541862 269728 541867 269784
rect 538029 269726 541867 269728
rect 538029 269723 538095 269726
rect 541801 269723 541867 269726
rect 509141 269514 509207 269517
rect 509877 269514 509943 269517
rect 509141 269512 509943 269514
rect 509141 269456 509146 269512
rect 509202 269456 509882 269512
rect 509938 269456 509943 269512
rect 509141 269454 509943 269456
rect 509141 269451 509207 269454
rect 509877 269451 509943 269454
rect 42057 269108 42123 269109
rect 42006 269106 42012 269108
rect 41966 269046 42012 269106
rect 42076 269104 42123 269108
rect 42118 269048 42123 269104
rect 42006 269044 42012 269046
rect 42076 269044 42123 269048
rect 42057 269043 42123 269044
rect 665817 268562 665883 268565
rect 676262 268562 676322 268668
rect 676857 268562 676923 268565
rect 665817 268560 676322 268562
rect 665817 268504 665822 268560
rect 665878 268504 676322 268560
rect 665817 268502 676322 268504
rect 676814 268560 676923 268562
rect 676814 268504 676862 268560
rect 676918 268504 676923 268560
rect 665817 268499 665883 268502
rect 676814 268499 676923 268504
rect 676814 268260 676874 268499
rect 673637 268154 673703 268157
rect 676213 268154 676279 268157
rect 673637 268152 676279 268154
rect 673637 268096 673642 268152
rect 673698 268096 676218 268152
rect 676274 268096 676279 268152
rect 673637 268094 676279 268096
rect 673637 268091 673703 268094
rect 676213 268091 676279 268094
rect 676262 267749 676322 267852
rect 676213 267744 676322 267749
rect 676213 267688 676218 267744
rect 676274 267688 676322 267744
rect 676213 267686 676322 267688
rect 676213 267683 676279 267686
rect 674373 267474 674439 267477
rect 674373 267472 676292 267474
rect 674373 267416 674378 267472
rect 674434 267416 676292 267472
rect 674373 267414 676292 267416
rect 674373 267411 674439 267414
rect 40677 267066 40743 267069
rect 62389 267066 62455 267069
rect 40677 267064 62455 267066
rect 40677 267008 40682 267064
rect 40738 267008 62394 267064
rect 62450 267008 62455 267064
rect 40677 267006 62455 267008
rect 40677 267003 40743 267006
rect 62389 267003 62455 267006
rect 674465 267066 674531 267069
rect 674465 267064 676292 267066
rect 674465 267008 674470 267064
rect 674526 267008 676292 267064
rect 674465 267006 676292 267008
rect 674465 267003 674531 267006
rect 674649 266658 674715 266661
rect 674649 266656 676292 266658
rect 674649 266600 674654 266656
rect 674710 266600 676292 266656
rect 674649 266598 676292 266600
rect 674649 266595 674715 266598
rect 42149 266250 42215 266253
rect 54477 266250 54543 266253
rect 42149 266248 54543 266250
rect 42149 266192 42154 266248
rect 42210 266192 54482 266248
rect 54538 266192 54543 266248
rect 42149 266190 54543 266192
rect 42149 266187 42215 266190
rect 54477 266187 54543 266190
rect 672993 266114 673059 266117
rect 676262 266114 676322 266220
rect 672993 266112 676322 266114
rect 672993 266056 672998 266112
rect 673054 266056 676322 266112
rect 672993 266054 676322 266056
rect 672993 266051 673059 266054
rect 673913 265842 673979 265845
rect 673913 265840 676292 265842
rect 673913 265784 673918 265840
rect 673974 265784 676292 265840
rect 673913 265782 676292 265784
rect 673913 265779 673979 265782
rect 673913 265434 673979 265437
rect 673913 265432 676292 265434
rect 673913 265376 673918 265432
rect 673974 265376 676292 265432
rect 673913 265374 676292 265376
rect 673913 265371 673979 265374
rect 673361 265026 673427 265029
rect 673361 265024 676292 265026
rect 673361 264968 673366 265024
rect 673422 264968 676292 265024
rect 673361 264966 676292 264968
rect 673361 264963 673427 264966
rect 674097 264618 674163 264621
rect 674097 264616 676292 264618
rect 674097 264560 674102 264616
rect 674158 264560 676292 264616
rect 674097 264558 676292 264560
rect 674097 264555 674163 264558
rect 55857 264210 55923 264213
rect 675334 264210 675340 264212
rect 55857 264208 675340 264210
rect 55857 264152 55862 264208
rect 55918 264152 675340 264208
rect 55857 264150 675340 264152
rect 55857 264147 55923 264150
rect 675334 264148 675340 264150
rect 675404 264148 675410 264212
rect 675477 264074 675543 264077
rect 676262 264074 676322 264180
rect 675477 264072 676322 264074
rect 675477 264016 675482 264072
rect 675538 264016 676322 264072
rect 675477 264014 676322 264016
rect 675477 264011 675543 264014
rect 676262 263669 676322 263772
rect 676213 263664 676322 263669
rect 676213 263608 676218 263664
rect 676274 263608 676322 263664
rect 676213 263606 676322 263608
rect 676213 263603 676279 263606
rect 679574 263261 679634 263364
rect 679574 263256 679683 263261
rect 679574 263200 679622 263256
rect 679678 263200 679683 263256
rect 679574 263198 679683 263200
rect 679617 263195 679683 263198
rect 676446 262853 676506 262956
rect 676397 262848 676506 262853
rect 676397 262792 676402 262848
rect 676458 262792 676506 262848
rect 676397 262790 676506 262792
rect 676397 262787 676463 262790
rect 674465 262578 674531 262581
rect 674465 262576 676292 262578
rect 674465 262520 674470 262576
rect 674526 262520 676292 262576
rect 674465 262518 676292 262520
rect 674465 262515 674531 262518
rect 554405 262170 554471 262173
rect 552460 262168 554471 262170
rect 552460 262112 554410 262168
rect 554466 262112 554471 262168
rect 552460 262110 554471 262112
rect 554405 262107 554471 262110
rect 671889 262170 671955 262173
rect 671889 262168 676292 262170
rect 671889 262112 671894 262168
rect 671950 262112 676292 262168
rect 671889 262110 676292 262112
rect 671889 262107 671955 262110
rect 673545 261626 673611 261629
rect 676998 261628 677058 261732
rect 673545 261624 676506 261626
rect 673545 261568 673550 261624
rect 673606 261568 676506 261624
rect 673545 261566 676506 261568
rect 673545 261563 673611 261566
rect 676446 261324 676506 261566
rect 676990 261564 676996 261628
rect 677060 261564 677066 261628
rect 675886 261156 675892 261220
rect 675956 261218 675962 261220
rect 676213 261218 676279 261221
rect 675956 261216 676279 261218
rect 675956 261160 676218 261216
rect 676274 261160 676279 261216
rect 675956 261158 676279 261160
rect 675956 261156 675962 261158
rect 676213 261155 676279 261158
rect 676814 260812 676874 260916
rect 676806 260748 676812 260812
rect 676876 260748 676882 260812
rect 670417 260538 670483 260541
rect 670417 260536 676292 260538
rect 670417 260480 670422 260536
rect 670478 260480 676292 260536
rect 670417 260478 676292 260480
rect 670417 260475 670483 260478
rect 674281 260130 674347 260133
rect 674281 260128 676292 260130
rect 674281 260072 674286 260128
rect 674342 260072 676292 260128
rect 674281 260070 676292 260072
rect 674281 260067 674347 260070
rect 554313 259994 554379 259997
rect 552460 259992 554379 259994
rect 552460 259936 554318 259992
rect 554374 259936 554379 259992
rect 552460 259934 554379 259936
rect 554313 259931 554379 259934
rect 671153 259722 671219 259725
rect 671153 259720 676292 259722
rect 671153 259664 671158 259720
rect 671214 259664 676292 259720
rect 671153 259662 676292 259664
rect 671153 259659 671219 259662
rect 673177 259314 673243 259317
rect 673177 259312 676292 259314
rect 673177 259256 673182 259312
rect 673238 259256 676292 259312
rect 673177 259254 676292 259256
rect 673177 259251 673243 259254
rect 673729 258906 673795 258909
rect 673729 258904 676292 258906
rect 673729 258848 673734 258904
rect 673790 258848 676292 258904
rect 673729 258846 676292 258848
rect 673729 258843 673795 258846
rect 670141 258498 670207 258501
rect 670141 258496 676292 258498
rect 670141 258440 670146 258496
rect 670202 258440 676292 258496
rect 670141 258438 676292 258440
rect 670141 258435 670207 258438
rect 46197 258090 46263 258093
rect 41492 258088 46263 258090
rect 41492 258032 46202 258088
rect 46258 258032 46263 258088
rect 41492 258030 46263 258032
rect 46197 258027 46263 258030
rect 675334 258028 675340 258092
rect 675404 258090 675410 258092
rect 675404 258060 676292 258090
rect 675404 258030 676322 258060
rect 675404 258028 675410 258030
rect 553945 257818 554011 257821
rect 552460 257816 554011 257818
rect 552460 257760 553950 257816
rect 554006 257760 554011 257816
rect 552460 257758 554011 257760
rect 553945 257755 554011 257758
rect 47577 257682 47643 257685
rect 41492 257680 47643 257682
rect 41492 257624 47582 257680
rect 47638 257624 47643 257680
rect 676262 257652 676322 258030
rect 41492 257622 47643 257624
rect 47577 257619 47643 257622
rect 671705 257274 671771 257277
rect 671705 257272 676292 257274
rect 35758 257141 35818 257244
rect 671705 257216 671710 257272
rect 671766 257216 676292 257272
rect 671705 257214 676292 257216
rect 671705 257211 671771 257214
rect 35758 257136 35867 257141
rect 35758 257080 35806 257136
rect 35862 257080 35867 257136
rect 35758 257078 35867 257080
rect 35801 257075 35867 257078
rect 44173 256866 44239 256869
rect 41492 256864 44239 256866
rect 41492 256808 44178 256864
rect 44234 256808 44239 256864
rect 41492 256806 44239 256808
rect 44173 256803 44239 256806
rect 44357 256458 44423 256461
rect 41492 256456 44423 256458
rect 41492 256400 44362 256456
rect 44418 256400 44423 256456
rect 41492 256398 44423 256400
rect 44357 256395 44423 256398
rect 35758 255917 35818 256020
rect 35758 255912 35867 255917
rect 35758 255856 35806 255912
rect 35862 255856 35867 255912
rect 35758 255854 35867 255856
rect 35801 255851 35867 255854
rect 39389 255914 39455 255917
rect 42793 255914 42859 255917
rect 39389 255912 42859 255914
rect 39389 255856 39394 255912
rect 39450 255856 42798 255912
rect 42854 255856 42859 255912
rect 39389 255854 42859 255856
rect 39389 255851 39455 255854
rect 42793 255851 42859 255854
rect 44909 255642 44975 255645
rect 553485 255642 553551 255645
rect 41492 255640 44975 255642
rect 41492 255584 44914 255640
rect 44970 255584 44975 255640
rect 41492 255582 44975 255584
rect 552460 255640 553551 255642
rect 552460 255584 553490 255640
rect 553546 255584 553551 255640
rect 552460 255582 553551 255584
rect 44909 255579 44975 255582
rect 553485 255579 553551 255582
rect 675017 255370 675083 255373
rect 675845 255370 675911 255373
rect 675017 255368 675911 255370
rect 675017 255312 675022 255368
rect 675078 255312 675850 255368
rect 675906 255312 675911 255368
rect 675017 255310 675911 255312
rect 675017 255307 675083 255310
rect 675845 255307 675911 255310
rect 44633 255234 44699 255237
rect 41492 255232 44699 255234
rect 41492 255176 44638 255232
rect 44694 255176 44699 255232
rect 41492 255174 44699 255176
rect 44633 255171 44699 255174
rect 44173 254826 44239 254829
rect 41492 254824 44239 254826
rect 41492 254768 44178 254824
rect 44234 254768 44239 254824
rect 41492 254766 44239 254768
rect 44173 254763 44239 254766
rect 35574 254285 35634 254388
rect 35525 254280 35634 254285
rect 35801 254282 35867 254285
rect 35525 254224 35530 254280
rect 35586 254224 35634 254280
rect 35525 254222 35634 254224
rect 35758 254280 35867 254282
rect 35758 254224 35806 254280
rect 35862 254224 35867 254280
rect 35525 254219 35591 254222
rect 35758 254219 35867 254224
rect 35758 253980 35818 254219
rect 39389 253874 39455 253877
rect 42885 253874 42951 253877
rect 39389 253872 42951 253874
rect 39389 253816 39394 253872
rect 39450 253816 42890 253872
rect 42946 253816 42951 253872
rect 39389 253814 42951 253816
rect 39389 253811 39455 253814
rect 42885 253811 42951 253814
rect 45553 253602 45619 253605
rect 41492 253600 45619 253602
rect 41492 253544 45558 253600
rect 45614 253544 45619 253600
rect 41492 253542 45619 253544
rect 45553 253539 45619 253542
rect 554405 253466 554471 253469
rect 552460 253464 554471 253466
rect 552460 253408 554410 253464
rect 554466 253408 554471 253464
rect 552460 253406 554471 253408
rect 554405 253403 554471 253406
rect 35758 253061 35818 253164
rect 35758 253056 35867 253061
rect 35758 253000 35806 253056
rect 35862 253000 35867 253056
rect 35758 252998 35867 253000
rect 35801 252995 35867 252998
rect 35758 252653 35818 252756
rect 35758 252648 35867 252653
rect 35758 252592 35806 252648
rect 35862 252592 35867 252648
rect 35758 252590 35867 252592
rect 35801 252587 35867 252590
rect 47209 252378 47275 252381
rect 41492 252376 47275 252378
rect 41492 252320 47214 252376
rect 47270 252320 47275 252376
rect 41492 252318 47275 252320
rect 47209 252315 47275 252318
rect 45921 251970 45987 251973
rect 41492 251968 45987 251970
rect 41492 251912 45926 251968
rect 45982 251912 45987 251968
rect 41492 251910 45987 251912
rect 45921 251907 45987 251910
rect 44541 251562 44607 251565
rect 41492 251560 44607 251562
rect 41492 251504 44546 251560
rect 44602 251504 44607 251560
rect 41492 251502 44607 251504
rect 44541 251499 44607 251502
rect 554129 251290 554195 251293
rect 552460 251288 554195 251290
rect 552460 251232 554134 251288
rect 554190 251232 554195 251288
rect 552460 251230 554195 251232
rect 554129 251227 554195 251230
rect 47025 251154 47091 251157
rect 41492 251152 47091 251154
rect 41492 251096 47030 251152
rect 47086 251096 47091 251152
rect 41492 251094 47091 251096
rect 47025 251091 47091 251094
rect 670969 250746 671035 250749
rect 675661 250746 675727 250749
rect 670969 250744 675727 250746
rect 40542 250612 40602 250716
rect 670969 250688 670974 250744
rect 671030 250688 675666 250744
rect 675722 250688 675727 250744
rect 670969 250686 675727 250688
rect 670969 250683 671035 250686
rect 675661 250683 675727 250686
rect 40534 250548 40540 250612
rect 40604 250548 40610 250612
rect 35758 250205 35818 250308
rect 35758 250200 35867 250205
rect 35758 250144 35806 250200
rect 35862 250144 35867 250200
rect 35758 250142 35867 250144
rect 35801 250139 35867 250142
rect 675753 250202 675819 250205
rect 676990 250202 676996 250204
rect 675753 250200 676996 250202
rect 675753 250144 675758 250200
rect 675814 250144 676996 250200
rect 675753 250142 676996 250144
rect 675753 250139 675819 250142
rect 676990 250140 676996 250142
rect 677060 250140 677066 250204
rect 674833 249930 674899 249933
rect 676070 249930 676076 249932
rect 674833 249928 676076 249930
rect 40726 249796 40786 249900
rect 674833 249872 674838 249928
rect 674894 249872 676076 249928
rect 674833 249870 676076 249872
rect 674833 249867 674899 249870
rect 676070 249868 676076 249870
rect 676140 249868 676146 249932
rect 40718 249732 40724 249796
rect 40788 249732 40794 249796
rect 675334 249596 675340 249660
rect 675404 249596 675410 249660
rect 46105 249522 46171 249525
rect 41492 249520 46171 249522
rect 41492 249464 46110 249520
rect 46166 249464 46171 249520
rect 41492 249462 46171 249464
rect 46105 249459 46171 249462
rect 45737 249114 45803 249117
rect 554037 249114 554103 249117
rect 41492 249112 45803 249114
rect 41492 249056 45742 249112
rect 45798 249056 45803 249112
rect 41492 249054 45803 249056
rect 552460 249112 554103 249114
rect 552460 249056 554042 249112
rect 554098 249056 554103 249112
rect 552460 249054 554103 249056
rect 45737 249051 45803 249054
rect 554037 249051 554103 249054
rect 675109 248978 675175 248981
rect 675342 248978 675402 249596
rect 675109 248976 675402 248978
rect 675109 248920 675114 248976
rect 675170 248920 675402 248976
rect 675109 248918 675402 248920
rect 675109 248915 675175 248918
rect 35758 248573 35818 248676
rect 35758 248568 35867 248573
rect 35758 248512 35806 248568
rect 35862 248512 35867 248568
rect 35758 248510 35867 248512
rect 35801 248507 35867 248510
rect 44725 248298 44791 248301
rect 41492 248296 44791 248298
rect 41492 248240 44730 248296
rect 44786 248240 44791 248296
rect 41492 248238 44791 248240
rect 44725 248235 44791 248238
rect 664437 248298 664503 248301
rect 670969 248298 671035 248301
rect 664437 248296 671035 248298
rect 664437 248240 664442 248296
rect 664498 248240 670974 248296
rect 671030 248240 671035 248296
rect 664437 248238 671035 248240
rect 664437 248235 664503 248238
rect 670969 248235 671035 248238
rect 35758 247757 35818 247860
rect 35758 247752 35867 247757
rect 35758 247696 35806 247752
rect 35862 247696 35867 247752
rect 35758 247694 35867 247696
rect 35801 247691 35867 247694
rect 40953 247754 41019 247757
rect 43345 247754 43411 247757
rect 40953 247752 43411 247754
rect 40953 247696 40958 247752
rect 41014 247696 43350 247752
rect 43406 247696 43411 247752
rect 40953 247694 43411 247696
rect 40953 247691 41019 247694
rect 43345 247691 43411 247694
rect 49141 247482 49207 247485
rect 41492 247480 49207 247482
rect 41492 247424 49146 247480
rect 49202 247424 49207 247480
rect 41492 247422 49207 247424
rect 49141 247419 49207 247422
rect 673545 247074 673611 247077
rect 675109 247074 675175 247077
rect 673545 247072 675175 247074
rect 35758 246941 35818 247044
rect 673545 247016 673550 247072
rect 673606 247016 675114 247072
rect 675170 247016 675175 247072
rect 673545 247014 675175 247016
rect 673545 247011 673611 247014
rect 675109 247011 675175 247014
rect 35758 246936 35867 246941
rect 553853 246938 553919 246941
rect 35758 246880 35806 246936
rect 35862 246880 35867 246936
rect 35758 246878 35867 246880
rect 552460 246936 553919 246938
rect 552460 246880 553858 246936
rect 553914 246880 553919 246936
rect 552460 246878 553919 246880
rect 35801 246875 35867 246878
rect 553853 246875 553919 246878
rect 47577 246666 47643 246669
rect 41492 246664 47643 246666
rect 41492 246608 47582 246664
rect 47638 246608 47643 246664
rect 41492 246606 47643 246608
rect 47577 246603 47643 246606
rect 675753 246666 675819 246669
rect 676806 246666 676812 246668
rect 675753 246664 676812 246666
rect 675753 246608 675758 246664
rect 675814 246608 676812 246664
rect 675753 246606 676812 246608
rect 675753 246603 675819 246606
rect 676806 246604 676812 246606
rect 676876 246604 676882 246668
rect 672073 246258 672139 246261
rect 673310 246258 673316 246260
rect 672073 246256 673316 246258
rect 672073 246200 672078 246256
rect 672134 246200 673316 246256
rect 672073 246198 673316 246200
rect 672073 246195 672139 246198
rect 673310 246196 673316 246198
rect 673380 246196 673386 246260
rect 40309 245714 40375 245717
rect 43161 245714 43227 245717
rect 40309 245712 43227 245714
rect 40309 245656 40314 245712
rect 40370 245656 43166 245712
rect 43222 245656 43227 245712
rect 40309 245654 43227 245656
rect 40309 245651 40375 245654
rect 43161 245651 43227 245654
rect 671153 245578 671219 245581
rect 675109 245578 675175 245581
rect 671153 245576 675175 245578
rect 671153 245520 671158 245576
rect 671214 245520 675114 245576
rect 675170 245520 675175 245576
rect 671153 245518 675175 245520
rect 671153 245515 671219 245518
rect 675109 245515 675175 245518
rect 671889 245306 671955 245309
rect 675109 245306 675175 245309
rect 671889 245304 675175 245306
rect 671889 245248 671894 245304
rect 671950 245248 675114 245304
rect 675170 245248 675175 245304
rect 671889 245246 675175 245248
rect 671889 245243 671955 245246
rect 675109 245243 675175 245246
rect 39389 244762 39455 244765
rect 42517 244762 42583 244765
rect 554497 244762 554563 244765
rect 39389 244760 42583 244762
rect 39389 244704 39394 244760
rect 39450 244704 42522 244760
rect 42578 244704 42583 244760
rect 39389 244702 42583 244704
rect 552460 244760 554563 244762
rect 552460 244704 554502 244760
rect 554558 244704 554563 244760
rect 552460 244702 554563 244704
rect 39389 244699 39455 244702
rect 42517 244699 42583 244702
rect 554497 244699 554563 244702
rect 39573 244082 39639 244085
rect 43069 244082 43135 244085
rect 39573 244080 43135 244082
rect 39573 244024 39578 244080
rect 39634 244024 43074 244080
rect 43130 244024 43135 244080
rect 39573 244022 43135 244024
rect 39573 244019 39639 244022
rect 43069 244019 43135 244022
rect 673177 242722 673243 242725
rect 675385 242722 675451 242725
rect 673177 242720 675451 242722
rect 673177 242664 673182 242720
rect 673238 242664 675390 242720
rect 675446 242664 675451 242720
rect 673177 242662 675451 242664
rect 673177 242659 673243 242662
rect 675385 242659 675451 242662
rect 553669 242586 553735 242589
rect 552460 242584 553735 242586
rect 552460 242528 553674 242584
rect 553730 242528 553735 242584
rect 552460 242526 553735 242528
rect 553669 242523 553735 242526
rect 673729 241498 673795 241501
rect 675201 241498 675267 241501
rect 673729 241496 675267 241498
rect 673729 241440 673734 241496
rect 673790 241440 675206 241496
rect 675262 241440 675267 241496
rect 673729 241438 675267 241440
rect 673729 241435 673795 241438
rect 675201 241435 675267 241438
rect 554497 240410 554563 240413
rect 552460 240408 554563 240410
rect 552460 240352 554502 240408
rect 554558 240352 554563 240408
rect 552460 240350 554563 240352
rect 554497 240347 554563 240350
rect 670417 240274 670483 240277
rect 675201 240274 675267 240277
rect 670417 240272 675267 240274
rect 670417 240216 670422 240272
rect 670478 240216 675206 240272
rect 675262 240216 675267 240272
rect 670417 240214 675267 240216
rect 670417 240211 670483 240214
rect 675201 240211 675267 240214
rect 42057 240138 42123 240141
rect 44541 240138 44607 240141
rect 42057 240136 44607 240138
rect 42057 240080 42062 240136
rect 42118 240080 44546 240136
rect 44602 240080 44607 240136
rect 42057 240078 44607 240080
rect 42057 240075 42123 240078
rect 44541 240075 44607 240078
rect 42241 238914 42307 238917
rect 42198 238912 42307 238914
rect 42198 238856 42246 238912
rect 42302 238856 42307 238912
rect 42198 238851 42307 238856
rect 42006 238036 42012 238100
rect 42076 238098 42082 238100
rect 42198 238098 42258 238851
rect 674833 238642 674899 238645
rect 675385 238642 675451 238645
rect 674833 238640 675451 238642
rect 674833 238584 674838 238640
rect 674894 238584 675390 238640
rect 675446 238584 675451 238640
rect 674833 238582 675451 238584
rect 674833 238579 674899 238582
rect 675385 238579 675451 238582
rect 554313 238234 554379 238237
rect 552460 238232 554379 238234
rect 552460 238176 554318 238232
rect 554374 238176 554379 238232
rect 552460 238174 554379 238176
rect 554313 238171 554379 238174
rect 42076 238038 42258 238098
rect 675017 238098 675083 238101
rect 675385 238098 675451 238101
rect 675017 238096 675451 238098
rect 675017 238040 675022 238096
rect 675078 238040 675390 238096
rect 675446 238040 675451 238096
rect 675017 238038 675451 238040
rect 42076 238036 42082 238038
rect 675017 238035 675083 238038
rect 675385 238035 675451 238038
rect 43805 237962 43871 237965
rect 62205 237962 62271 237965
rect 43805 237960 62271 237962
rect 43805 237904 43810 237960
rect 43866 237904 62210 237960
rect 62266 237904 62271 237960
rect 43805 237902 62271 237904
rect 43805 237899 43871 237902
rect 62205 237899 62271 237902
rect 673177 236738 673243 236741
rect 674230 236738 674236 236740
rect 673177 236736 674236 236738
rect 673177 236680 673182 236736
rect 673238 236680 674236 236736
rect 673177 236678 674236 236680
rect 673177 236675 673243 236678
rect 674230 236676 674236 236678
rect 674300 236676 674306 236740
rect 40718 236540 40724 236604
rect 40788 236602 40794 236604
rect 41781 236602 41847 236605
rect 40788 236600 41847 236602
rect 40788 236544 41786 236600
rect 41842 236544 41847 236600
rect 40788 236542 41847 236544
rect 40788 236540 40794 236542
rect 41781 236539 41847 236542
rect 672073 236330 672139 236333
rect 673637 236330 673703 236333
rect 672073 236328 673703 236330
rect 672073 236272 672078 236328
rect 672134 236272 673642 236328
rect 673698 236272 673703 236328
rect 672073 236270 673703 236272
rect 672073 236267 672139 236270
rect 673637 236267 673703 236270
rect 554497 236058 554563 236061
rect 552460 236056 554563 236058
rect 552460 236000 554502 236056
rect 554558 236000 554563 236056
rect 552460 235998 554563 236000
rect 554497 235995 554563 235998
rect 42425 235922 42491 235925
rect 44725 235922 44791 235925
rect 42425 235920 44791 235922
rect 42425 235864 42430 235920
rect 42486 235864 44730 235920
rect 44786 235864 44791 235920
rect 42425 235862 44791 235864
rect 42425 235859 42491 235862
rect 44725 235859 44791 235862
rect 674097 235242 674163 235245
rect 675845 235242 675911 235245
rect 674097 235240 675911 235242
rect 674097 235184 674102 235240
rect 674158 235184 675850 235240
rect 675906 235184 675911 235240
rect 674097 235182 675911 235184
rect 674097 235179 674163 235182
rect 675845 235179 675911 235182
rect 668945 234562 669011 234565
rect 671245 234562 671311 234565
rect 668945 234560 671311 234562
rect 668945 234504 668950 234560
rect 669006 234504 671250 234560
rect 671306 234504 671311 234560
rect 668945 234502 671311 234504
rect 668945 234499 669011 234502
rect 671245 234499 671311 234502
rect 554405 233882 554471 233885
rect 552460 233880 554471 233882
rect 552460 233824 554410 233880
rect 554466 233824 554471 233880
rect 552460 233822 554471 233824
rect 554405 233819 554471 233822
rect 42425 233338 42491 233341
rect 46105 233338 46171 233341
rect 42425 233336 46171 233338
rect 42425 233280 42430 233336
rect 42486 233280 46110 233336
rect 46166 233280 46171 233336
rect 42425 233278 46171 233280
rect 42425 233275 42491 233278
rect 46105 233275 46171 233278
rect 42425 231978 42491 231981
rect 45921 231978 45987 231981
rect 42425 231976 45987 231978
rect 42425 231920 42430 231976
rect 42486 231920 45926 231976
rect 45982 231920 45987 231976
rect 42425 231918 45987 231920
rect 42425 231915 42491 231918
rect 45921 231915 45987 231918
rect 43989 230618 44055 230621
rect 43486 230616 44055 230618
rect 43486 230560 43994 230616
rect 44050 230560 44055 230616
rect 43486 230558 44055 230560
rect 43486 230493 43546 230558
rect 43989 230555 44055 230558
rect 43437 230488 43546 230493
rect 43437 230432 43442 230488
rect 43498 230432 43546 230488
rect 43437 230430 43546 230432
rect 142613 230482 142679 230485
rect 144085 230482 144151 230485
rect 142613 230480 144151 230482
rect 43437 230427 43503 230430
rect 142613 230424 142618 230480
rect 142674 230424 144090 230480
rect 144146 230424 144151 230480
rect 142613 230422 144151 230424
rect 142613 230419 142679 230422
rect 144085 230419 144151 230422
rect 659561 230482 659627 230485
rect 674097 230482 674163 230485
rect 659561 230480 674163 230482
rect 659561 230424 659566 230480
rect 659622 230424 674102 230480
rect 674158 230424 674163 230480
rect 659561 230422 674163 230424
rect 659561 230419 659627 230422
rect 674097 230419 674163 230422
rect 674281 230482 674347 230485
rect 676949 230482 677015 230485
rect 674281 230480 677015 230482
rect 674281 230424 674286 230480
rect 674342 230424 676954 230480
rect 677010 230424 677015 230480
rect 674281 230422 677015 230424
rect 674281 230419 674347 230422
rect 676949 230419 677015 230422
rect 665173 230210 665239 230213
rect 673453 230210 673519 230213
rect 665173 230208 673519 230210
rect 665173 230152 665178 230208
rect 665234 230152 673458 230208
rect 673514 230152 673519 230208
rect 665173 230150 673519 230152
rect 665173 230147 665239 230150
rect 673453 230147 673519 230150
rect 674465 230210 674531 230213
rect 676213 230210 676279 230213
rect 674465 230208 676279 230210
rect 674465 230152 674470 230208
rect 674526 230152 676218 230208
rect 676274 230152 676279 230208
rect 674465 230150 676279 230152
rect 674465 230147 674531 230150
rect 676213 230147 676279 230150
rect 156689 229938 156755 229941
rect 157425 229938 157491 229941
rect 156689 229936 157491 229938
rect 156689 229880 156694 229936
rect 156750 229880 157430 229936
rect 157486 229880 157491 229936
rect 156689 229878 157491 229880
rect 156689 229875 156755 229878
rect 157425 229875 157491 229878
rect 40534 229604 40540 229668
rect 40604 229666 40610 229668
rect 41781 229666 41847 229669
rect 40604 229664 41847 229666
rect 40604 229608 41786 229664
rect 41842 229608 41847 229664
rect 40604 229606 41847 229608
rect 40604 229604 40610 229606
rect 41781 229603 41847 229606
rect 157701 229666 157767 229669
rect 158713 229666 158779 229669
rect 157701 229664 158779 229666
rect 157701 229608 157706 229664
rect 157762 229608 158718 229664
rect 158774 229608 158779 229664
rect 157701 229606 158779 229608
rect 157701 229603 157767 229606
rect 158713 229603 158779 229606
rect 150341 229394 150407 229397
rect 156321 229394 156387 229397
rect 150341 229392 156387 229394
rect 150341 229336 150346 229392
rect 150402 229336 156326 229392
rect 156382 229336 156387 229392
rect 150341 229334 156387 229336
rect 150341 229331 150407 229334
rect 156321 229331 156387 229334
rect 663701 229394 663767 229397
rect 674465 229394 674531 229397
rect 663701 229392 674531 229394
rect 663701 229336 663706 229392
rect 663762 229336 674470 229392
rect 674526 229336 674531 229392
rect 663701 229334 674531 229336
rect 663701 229331 663767 229334
rect 674465 229331 674531 229334
rect 140037 229258 140103 229261
rect 145833 229258 145899 229261
rect 140037 229256 145899 229258
rect 140037 229200 140042 229256
rect 140098 229200 145838 229256
rect 145894 229200 145899 229256
rect 140037 229198 145899 229200
rect 140037 229195 140103 229198
rect 145833 229195 145899 229198
rect 147121 229258 147187 229261
rect 149973 229258 150039 229261
rect 147121 229256 150039 229258
rect 147121 229200 147126 229256
rect 147182 229200 149978 229256
rect 150034 229200 150039 229256
rect 147121 229198 150039 229200
rect 147121 229195 147187 229198
rect 149973 229195 150039 229198
rect 202873 229122 202939 229125
rect 205173 229122 205239 229125
rect 202873 229120 205239 229122
rect 202873 229064 202878 229120
rect 202934 229064 205178 229120
rect 205234 229064 205239 229120
rect 202873 229062 205239 229064
rect 202873 229059 202939 229062
rect 205173 229059 205239 229062
rect 42425 228986 42491 228989
rect 45737 228986 45803 228989
rect 42425 228984 45803 228986
rect 42425 228928 42430 228984
rect 42486 228928 45742 228984
rect 45798 228928 45803 228984
rect 42425 228926 45803 228928
rect 42425 228923 42491 228926
rect 45737 228923 45803 228926
rect 146477 228986 146543 228989
rect 149237 228986 149303 228989
rect 146477 228984 149303 228986
rect 146477 228928 146482 228984
rect 146538 228928 149242 228984
rect 149298 228928 149303 228984
rect 146477 228926 149303 228928
rect 146477 228923 146543 228926
rect 149237 228923 149303 228926
rect 166809 228986 166875 228989
rect 167361 228986 167427 228989
rect 674925 228988 674991 228989
rect 674925 228986 674972 228988
rect 166809 228984 167427 228986
rect 166809 228928 166814 228984
rect 166870 228928 167366 228984
rect 167422 228928 167427 228984
rect 166809 228926 167427 228928
rect 674880 228984 674972 228986
rect 674880 228928 674930 228984
rect 674880 228926 674972 228928
rect 166809 228923 166875 228926
rect 167361 228923 167427 228926
rect 674925 228924 674972 228926
rect 675036 228924 675042 228988
rect 674925 228923 674991 228924
rect 173157 228850 173223 228853
rect 174813 228850 174879 228853
rect 674046 228850 674052 228852
rect 173157 228848 174879 228850
rect 173157 228792 173162 228848
rect 173218 228792 174818 228848
rect 174874 228792 174879 228848
rect 173157 228790 174879 228792
rect 173157 228787 173223 228790
rect 174813 228787 174879 228790
rect 669270 228790 674052 228850
rect 139301 228714 139367 228717
rect 147305 228714 147371 228717
rect 139301 228712 147371 228714
rect 139301 228656 139306 228712
rect 139362 228656 147310 228712
rect 147366 228656 147371 228712
rect 139301 228654 147371 228656
rect 139301 228651 139367 228654
rect 147305 228651 147371 228654
rect 219617 228714 219683 228717
rect 220537 228714 220603 228717
rect 219617 228712 220603 228714
rect 219617 228656 219622 228712
rect 219678 228656 220542 228712
rect 220598 228656 220603 228712
rect 219617 228654 220603 228656
rect 219617 228651 219683 228654
rect 220537 228651 220603 228654
rect 652569 228578 652635 228581
rect 669270 228578 669330 228790
rect 674046 228788 674052 228790
rect 674116 228788 674122 228852
rect 652569 228576 669330 228578
rect 652569 228520 652574 228576
rect 652630 228520 669330 228576
rect 652569 228518 669330 228520
rect 673729 228578 673795 228581
rect 676673 228578 676739 228581
rect 673729 228576 676739 228578
rect 673729 228520 673734 228576
rect 673790 228520 676678 228576
rect 676734 228520 676739 228576
rect 673729 228518 676739 228520
rect 652569 228515 652635 228518
rect 673729 228515 673795 228518
rect 676673 228515 676739 228518
rect 160001 228170 160067 228173
rect 166809 228170 166875 228173
rect 160001 228168 166875 228170
rect 160001 228112 160006 228168
rect 160062 228112 166814 228168
rect 166870 228112 166875 228168
rect 160001 228110 166875 228112
rect 160001 228107 160067 228110
rect 166809 228107 166875 228110
rect 42425 227626 42491 227629
rect 45553 227626 45619 227629
rect 42425 227624 45619 227626
rect 42425 227568 42430 227624
rect 42486 227568 45558 227624
rect 45614 227568 45619 227624
rect 42425 227566 45619 227568
rect 42425 227563 42491 227566
rect 45553 227563 45619 227566
rect 171225 227626 171291 227629
rect 172145 227626 172211 227629
rect 171225 227624 172211 227626
rect 171225 227568 171230 227624
rect 171286 227568 172150 227624
rect 172206 227568 172211 227624
rect 171225 227566 172211 227568
rect 171225 227563 171291 227566
rect 172145 227563 172211 227566
rect 156689 227490 156755 227493
rect 166533 227490 166599 227493
rect 156689 227488 166599 227490
rect 156689 227432 156694 227488
rect 156750 227432 166538 227488
rect 166594 227432 166599 227488
rect 156689 227430 166599 227432
rect 156689 227427 156755 227430
rect 166533 227427 166599 227430
rect 169477 227354 169543 227357
rect 171685 227354 171751 227357
rect 169477 227352 171751 227354
rect 169477 227296 169482 227352
rect 169538 227296 171690 227352
rect 171746 227296 171751 227352
rect 169477 227294 171751 227296
rect 169477 227291 169543 227294
rect 171685 227291 171751 227294
rect 672257 227082 672323 227085
rect 672574 227082 672580 227084
rect 672257 227080 672580 227082
rect 672257 227024 672262 227080
rect 672318 227024 672580 227080
rect 672257 227022 672580 227024
rect 672257 227019 672323 227022
rect 672574 227020 672580 227022
rect 672644 227020 672650 227084
rect 673729 226538 673795 226541
rect 675201 226538 675267 226541
rect 673729 226536 675267 226538
rect 673729 226480 673734 226536
rect 673790 226480 675206 226536
rect 675262 226480 675267 226536
rect 673729 226478 675267 226480
rect 673729 226475 673795 226478
rect 675201 226475 675267 226478
rect 656157 226402 656223 226405
rect 672717 226402 672783 226405
rect 656157 226400 672783 226402
rect 656157 226344 656162 226400
rect 656218 226344 672722 226400
rect 672778 226344 672783 226400
rect 656157 226342 672783 226344
rect 656157 226339 656223 226342
rect 672717 226339 672783 226342
rect 42609 226266 42675 226269
rect 47209 226266 47275 226269
rect 42609 226264 47275 226266
rect 42609 226208 42614 226264
rect 42670 226208 47214 226264
rect 47270 226208 47275 226264
rect 42609 226206 47275 226208
rect 42609 226203 42675 226206
rect 47209 226203 47275 226206
rect 41965 226132 42031 226133
rect 41965 226128 42012 226132
rect 42076 226130 42082 226132
rect 141141 226130 141207 226133
rect 145189 226130 145255 226133
rect 41965 226072 41970 226128
rect 41965 226068 42012 226072
rect 42076 226070 42122 226130
rect 141141 226128 145255 226130
rect 141141 226072 141146 226128
rect 141202 226072 145194 226128
rect 145250 226072 145255 226128
rect 141141 226070 145255 226072
rect 42076 226068 42082 226070
rect 41965 226067 42031 226068
rect 141141 226067 141207 226070
rect 145189 226067 145255 226070
rect 672597 226130 672663 226133
rect 674833 226130 674899 226133
rect 672597 226128 674899 226130
rect 672597 226072 672602 226128
rect 672658 226072 674838 226128
rect 674894 226072 674899 226128
rect 672597 226070 674899 226072
rect 672597 226067 672663 226070
rect 674833 226067 674899 226070
rect 672257 225858 672323 225861
rect 675017 225858 675083 225861
rect 672257 225856 675083 225858
rect 672257 225800 672262 225856
rect 672318 225800 675022 225856
rect 675078 225800 675083 225856
rect 672257 225798 675083 225800
rect 672257 225795 672323 225798
rect 675017 225795 675083 225798
rect 663057 225722 663123 225725
rect 663057 225720 672090 225722
rect 663057 225664 663062 225720
rect 663118 225664 672090 225720
rect 663057 225662 672090 225664
rect 663057 225659 663123 225662
rect 672030 225453 672090 225662
rect 203885 225450 203951 225453
rect 205081 225450 205147 225453
rect 203885 225448 205147 225450
rect 203885 225392 203890 225448
rect 203946 225392 205086 225448
rect 205142 225392 205147 225448
rect 203885 225390 205147 225392
rect 203885 225387 203951 225390
rect 205081 225387 205147 225390
rect 672027 225448 672093 225453
rect 672027 225392 672032 225448
rect 672088 225392 672093 225448
rect 672027 225387 672093 225392
rect 653397 225314 653463 225317
rect 671245 225314 671311 225317
rect 653397 225312 671311 225314
rect 653397 225256 653402 225312
rect 653458 225256 671250 225312
rect 671306 225256 671311 225312
rect 653397 225254 671311 225256
rect 653397 225251 653463 225254
rect 671245 225251 671311 225254
rect 672149 225314 672215 225317
rect 675661 225314 675727 225317
rect 672149 225312 675727 225314
rect 672149 225256 672154 225312
rect 672210 225256 675666 225312
rect 675722 225256 675727 225312
rect 672149 225254 675727 225256
rect 672149 225251 672215 225254
rect 675661 225251 675727 225254
rect 651465 225042 651531 225045
rect 672257 225042 672323 225045
rect 651465 225040 672323 225042
rect 651465 224984 651470 225040
rect 651526 224984 672262 225040
rect 672318 224984 672323 225040
rect 651465 224982 672323 224984
rect 651465 224979 651531 224982
rect 672257 224979 672323 224982
rect 42425 224906 42491 224909
rect 47025 224906 47091 224909
rect 42425 224904 47091 224906
rect 42425 224848 42430 224904
rect 42486 224848 47030 224904
rect 47086 224848 47091 224904
rect 42425 224846 47091 224848
rect 42425 224843 42491 224846
rect 47025 224843 47091 224846
rect 176285 224906 176351 224909
rect 176837 224906 176903 224909
rect 176285 224904 176903 224906
rect 176285 224848 176290 224904
rect 176346 224848 176842 224904
rect 176898 224848 176903 224904
rect 176285 224846 176903 224848
rect 176285 224843 176351 224846
rect 176837 224843 176903 224846
rect 557257 224770 557323 224773
rect 558545 224770 558611 224773
rect 557257 224768 558611 224770
rect 557257 224712 557262 224768
rect 557318 224712 558550 224768
rect 558606 224712 558611 224768
rect 557257 224710 558611 224712
rect 557257 224707 557323 224710
rect 558545 224707 558611 224710
rect 561397 224770 561463 224773
rect 565169 224770 565235 224773
rect 561397 224768 565235 224770
rect 561397 224712 561402 224768
rect 561458 224712 565174 224768
rect 565230 224712 565235 224768
rect 561397 224710 565235 224712
rect 561397 224707 561463 224710
rect 565169 224707 565235 224710
rect 555785 224498 555851 224501
rect 561673 224498 561739 224501
rect 555785 224496 561739 224498
rect 555785 224440 555790 224496
rect 555846 224440 561678 224496
rect 561734 224440 561739 224496
rect 555785 224438 561739 224440
rect 555785 224435 555851 224438
rect 561673 224435 561739 224438
rect 562593 224498 562659 224501
rect 563145 224498 563211 224501
rect 562593 224496 563211 224498
rect 562593 224440 562598 224496
rect 562654 224440 563150 224496
rect 563206 224440 563211 224496
rect 562593 224438 563211 224440
rect 562593 224435 562659 224438
rect 563145 224435 563211 224438
rect 666829 224362 666895 224365
rect 659610 224360 666895 224362
rect 659610 224304 666834 224360
rect 666890 224304 666895 224360
rect 659610 224302 666895 224304
rect 562685 224090 562751 224093
rect 563421 224090 563487 224093
rect 562685 224088 563487 224090
rect 562685 224032 562690 224088
rect 562746 224032 563426 224088
rect 563482 224032 563487 224088
rect 562685 224030 563487 224032
rect 562685 224027 562751 224030
rect 563421 224027 563487 224030
rect 657537 223682 657603 223685
rect 659610 223682 659670 224302
rect 666829 224299 666895 224302
rect 660205 224090 660271 224093
rect 667013 224090 667079 224093
rect 660205 224088 667079 224090
rect 660205 224032 660210 224088
rect 660266 224032 667018 224088
rect 667074 224032 667079 224088
rect 660205 224030 667079 224032
rect 660205 224027 660271 224030
rect 667013 224027 667079 224030
rect 670785 223954 670851 223957
rect 672073 223954 672139 223957
rect 670785 223952 672139 223954
rect 670785 223896 670790 223952
rect 670846 223896 672078 223952
rect 672134 223896 672139 223952
rect 670785 223894 672139 223896
rect 670785 223891 670851 223894
rect 672073 223891 672139 223894
rect 679249 223818 679315 223821
rect 679206 223816 679315 223818
rect 679206 223760 679254 223816
rect 679310 223760 679315 223816
rect 679206 223755 679315 223760
rect 657537 223680 659670 223682
rect 657537 223624 657542 223680
rect 657598 223624 659670 223680
rect 657537 223622 659670 223624
rect 670785 223682 670851 223685
rect 672257 223682 672323 223685
rect 670785 223680 672323 223682
rect 670785 223624 670790 223680
rect 670846 223624 672262 223680
rect 672318 223624 672323 223680
rect 670785 223622 672323 223624
rect 657537 223619 657603 223622
rect 670785 223619 670851 223622
rect 672257 223619 672323 223622
rect 42149 223546 42215 223549
rect 59997 223546 60063 223549
rect 42149 223544 60063 223546
rect 42149 223488 42154 223544
rect 42210 223488 60002 223544
rect 60058 223488 60063 223544
rect 679206 223516 679266 223755
rect 42149 223486 60063 223488
rect 42149 223483 42215 223486
rect 59997 223483 60063 223486
rect 151905 223274 151971 223277
rect 159817 223274 159883 223277
rect 151905 223272 159883 223274
rect 151905 223216 151910 223272
rect 151966 223216 159822 223272
rect 159878 223216 159883 223272
rect 151905 223214 159883 223216
rect 151905 223211 151971 223214
rect 159817 223211 159883 223214
rect 676029 223138 676095 223141
rect 676029 223136 676292 223138
rect 676029 223080 676034 223136
rect 676090 223080 676292 223136
rect 676029 223078 676292 223080
rect 676029 223075 676095 223078
rect 147305 223002 147371 223005
rect 151445 223002 151511 223005
rect 147305 223000 151511 223002
rect 147305 222944 147310 223000
rect 147366 222944 151450 223000
rect 151506 222944 151511 223000
rect 147305 222942 151511 222944
rect 147305 222939 147371 222942
rect 151445 222939 151511 222942
rect 151629 222730 151695 222733
rect 152089 222730 152155 222733
rect 151629 222728 152155 222730
rect 151629 222672 151634 222728
rect 151690 222672 152094 222728
rect 152150 222672 152155 222728
rect 151629 222670 152155 222672
rect 151629 222667 151695 222670
rect 152089 222667 152155 222670
rect 666001 222730 666067 222733
rect 675201 222730 675267 222733
rect 683665 222730 683731 222733
rect 666001 222728 675267 222730
rect 666001 222672 666006 222728
rect 666062 222672 675206 222728
rect 675262 222672 675267 222728
rect 666001 222670 675267 222672
rect 683652 222728 683731 222730
rect 683652 222672 683670 222728
rect 683726 222672 683731 222728
rect 683652 222670 683731 222672
rect 666001 222667 666067 222670
rect 675201 222667 675267 222670
rect 683665 222667 683731 222670
rect 145925 222322 145991 222325
rect 147121 222322 147187 222325
rect 145925 222320 147187 222322
rect 145925 222264 145930 222320
rect 145986 222264 147126 222320
rect 147182 222264 147187 222320
rect 145925 222262 147187 222264
rect 145925 222259 145991 222262
rect 147121 222259 147187 222262
rect 658181 222322 658247 222325
rect 670785 222322 670851 222325
rect 658181 222320 670851 222322
rect 658181 222264 658186 222320
rect 658242 222264 670790 222320
rect 670846 222264 670851 222320
rect 658181 222262 670851 222264
rect 658181 222259 658247 222262
rect 670785 222259 670851 222262
rect 674649 222322 674715 222325
rect 674649 222320 676292 222322
rect 674649 222264 674654 222320
rect 674710 222264 676292 222320
rect 674649 222262 676292 222264
rect 674649 222259 674715 222262
rect 543687 222210 543753 222213
rect 543584 222208 543753 222210
rect 542261 222186 542327 222189
rect 543584 222186 543692 222208
rect 542261 222184 543692 222186
rect 542261 222128 542266 222184
rect 542322 222152 543692 222184
rect 543748 222152 543753 222208
rect 542322 222147 543753 222152
rect 542322 222128 543750 222147
rect 542261 222126 543750 222128
rect 542261 222123 542327 222126
rect 550633 222050 550699 222053
rect 550817 222050 550883 222053
rect 558729 222050 558795 222053
rect 550633 222048 558795 222050
rect 550633 221992 550638 222048
rect 550694 221992 550822 222048
rect 550878 221992 558734 222048
rect 558790 221992 558795 222048
rect 550633 221990 558795 221992
rect 550633 221987 550699 221990
rect 550817 221987 550883 221990
rect 558729 221987 558795 221990
rect 161427 221914 161493 221917
rect 164509 221914 164575 221917
rect 161427 221912 164575 221914
rect 161427 221856 161432 221912
rect 161488 221856 164514 221912
rect 164570 221856 164575 221912
rect 161427 221854 164575 221856
rect 161427 221851 161493 221854
rect 164509 221851 164575 221854
rect 673729 221914 673795 221917
rect 673729 221912 676292 221914
rect 673729 221856 673734 221912
rect 673790 221856 676292 221912
rect 673729 221854 676292 221856
rect 673729 221851 673795 221854
rect 184657 221778 184723 221781
rect 185761 221778 185827 221781
rect 184657 221776 185827 221778
rect 184657 221720 184662 221776
rect 184718 221720 185766 221776
rect 185822 221720 185827 221776
rect 184657 221718 185827 221720
rect 184657 221715 184723 221718
rect 185761 221715 185827 221718
rect 547137 221778 547203 221781
rect 558545 221778 558611 221781
rect 547137 221776 558611 221778
rect 547137 221720 547142 221776
rect 547198 221720 558550 221776
rect 558606 221720 558611 221776
rect 547137 221718 558611 221720
rect 547137 221715 547203 221718
rect 558545 221715 558611 221718
rect 560937 221778 561003 221781
rect 568941 221778 569007 221781
rect 560937 221776 569007 221778
rect 560937 221720 560942 221776
rect 560998 221720 568946 221776
rect 569002 221720 569007 221776
rect 560937 221718 569007 221720
rect 560937 221715 561003 221718
rect 568941 221715 569007 221718
rect 161657 221642 161723 221645
rect 161614 221640 161723 221642
rect 161614 221584 161662 221640
rect 161718 221584 161723 221640
rect 161614 221579 161723 221584
rect 651925 221642 651991 221645
rect 651925 221640 672090 221642
rect 651925 221584 651930 221640
rect 651986 221584 672090 221640
rect 651925 221582 672090 221584
rect 651925 221579 651991 221582
rect 158253 221506 158319 221509
rect 161614 221506 161674 221579
rect 158253 221504 161674 221506
rect 158253 221448 158258 221504
rect 158314 221448 161674 221504
rect 158253 221446 161674 221448
rect 519629 221506 519695 221509
rect 520181 221506 520247 221509
rect 618253 221506 618319 221509
rect 519629 221504 618319 221506
rect 519629 221448 519634 221504
rect 519690 221448 520186 221504
rect 520242 221448 618258 221504
rect 618314 221448 618319 221504
rect 519629 221446 618319 221448
rect 158253 221443 158319 221446
rect 519629 221443 519695 221446
rect 520181 221443 520247 221446
rect 618253 221443 618319 221446
rect 176469 221370 176535 221373
rect 177297 221370 177363 221373
rect 176469 221368 177363 221370
rect 176469 221312 176474 221368
rect 176530 221312 177302 221368
rect 177358 221312 177363 221368
rect 176469 221310 177363 221312
rect 176469 221307 176535 221310
rect 177297 221307 177363 221310
rect 513557 221234 513623 221237
rect 599485 221234 599551 221237
rect 513557 221232 599551 221234
rect 513557 221176 513562 221232
rect 513618 221176 599490 221232
rect 599546 221176 599551 221232
rect 513557 221174 599551 221176
rect 672030 221234 672090 221582
rect 673085 221506 673151 221509
rect 673085 221504 676292 221506
rect 673085 221448 673090 221504
rect 673146 221448 676292 221504
rect 673085 221446 676292 221448
rect 673085 221443 673151 221446
rect 674833 221234 674899 221237
rect 672030 221232 674899 221234
rect 672030 221176 674838 221232
rect 674894 221176 674899 221232
rect 672030 221174 674899 221176
rect 513557 221171 513623 221174
rect 599485 221171 599551 221174
rect 674833 221171 674899 221174
rect 654317 221098 654383 221101
rect 671337 221098 671403 221101
rect 654317 221096 671403 221098
rect 654317 221040 654322 221096
rect 654378 221040 671342 221096
rect 671398 221040 671403 221096
rect 654317 221038 671403 221040
rect 654317 221035 654383 221038
rect 671337 221035 671403 221038
rect 676029 221098 676095 221101
rect 676029 221096 676292 221098
rect 676029 221040 676034 221096
rect 676090 221040 676292 221096
rect 676029 221038 676292 221040
rect 676029 221035 676095 221038
rect 497733 220962 497799 220965
rect 631317 220962 631383 220965
rect 497733 220960 631383 220962
rect 497733 220904 497738 220960
rect 497794 220904 631322 220960
rect 631378 220904 631383 220960
rect 497733 220902 631383 220904
rect 497733 220899 497799 220902
rect 631317 220899 631383 220902
rect 176469 220826 176535 220829
rect 179781 220826 179847 220829
rect 176469 220824 179847 220826
rect 176469 220768 176474 220824
rect 176530 220768 179786 220824
rect 179842 220768 179847 220824
rect 176469 220766 179847 220768
rect 176469 220763 176535 220766
rect 179781 220763 179847 220766
rect 154021 220690 154087 220693
rect 156965 220690 157031 220693
rect 154021 220688 157031 220690
rect 154021 220632 154026 220688
rect 154082 220632 156970 220688
rect 157026 220632 157031 220688
rect 154021 220630 157031 220632
rect 154021 220627 154087 220630
rect 156965 220627 157031 220630
rect 164141 220690 164207 220693
rect 167085 220690 167151 220693
rect 164141 220688 167151 220690
rect 164141 220632 164146 220688
rect 164202 220632 167090 220688
rect 167146 220632 167151 220688
rect 164141 220630 167151 220632
rect 164141 220627 164207 220630
rect 167085 220627 167151 220630
rect 553577 220690 553643 220693
rect 561489 220690 561555 220693
rect 553577 220688 561555 220690
rect 553577 220632 553582 220688
rect 553638 220632 561494 220688
rect 561550 220632 561555 220688
rect 553577 220630 561555 220632
rect 553577 220627 553643 220630
rect 561489 220627 561555 220630
rect 563053 220690 563119 220693
rect 564801 220690 564867 220693
rect 569953 220690 570019 220693
rect 563053 220688 564867 220690
rect 563053 220632 563058 220688
rect 563114 220632 564806 220688
rect 564862 220632 564867 220688
rect 563053 220630 564867 220632
rect 563053 220627 563119 220630
rect 564801 220627 564867 220630
rect 565310 220688 570019 220690
rect 565310 220632 569958 220688
rect 570014 220632 570019 220688
rect 565310 220630 570019 220632
rect 543549 220554 543615 220557
rect 544745 220554 544811 220557
rect 543549 220552 544811 220554
rect 543549 220496 543554 220552
rect 543610 220496 544750 220552
rect 544806 220496 544811 220552
rect 543549 220494 544811 220496
rect 543549 220491 543615 220494
rect 544745 220491 544811 220494
rect 141969 220418 142035 220421
rect 144177 220418 144243 220421
rect 141969 220416 144243 220418
rect 141969 220360 141974 220416
rect 142030 220360 144182 220416
rect 144238 220360 144243 220416
rect 141969 220358 144243 220360
rect 141969 220355 142035 220358
rect 144177 220355 144243 220358
rect 146753 220418 146819 220421
rect 558361 220418 558427 220421
rect 563237 220418 563303 220421
rect 146753 220416 151830 220418
rect 146753 220360 146758 220416
rect 146814 220387 151830 220416
rect 558361 220416 563303 220418
rect 146814 220382 151833 220387
rect 146814 220360 151772 220382
rect 146753 220358 151772 220360
rect 146753 220355 146819 220358
rect 151767 220326 151772 220358
rect 151828 220326 151833 220382
rect 558361 220360 558366 220416
rect 558422 220360 563242 220416
rect 563298 220360 563303 220416
rect 558361 220358 563303 220360
rect 558361 220355 558427 220358
rect 563237 220355 563303 220358
rect 563421 220418 563487 220421
rect 565310 220418 565370 220630
rect 569953 220627 570019 220630
rect 573357 220690 573423 220693
rect 674097 220690 674163 220693
rect 573357 220688 576870 220690
rect 573357 220632 573362 220688
rect 573418 220632 576870 220688
rect 573357 220630 576870 220632
rect 573357 220627 573423 220630
rect 563421 220416 565370 220418
rect 563421 220360 563426 220416
rect 563482 220360 565370 220416
rect 563421 220358 565370 220360
rect 565629 220418 565695 220421
rect 576577 220418 576643 220421
rect 565629 220416 576643 220418
rect 565629 220360 565634 220416
rect 565690 220360 576582 220416
rect 576638 220360 576643 220416
rect 565629 220358 576643 220360
rect 563421 220355 563487 220358
rect 565629 220355 565695 220358
rect 576577 220355 576643 220358
rect 151767 220321 151833 220326
rect 181529 220282 181595 220285
rect 180750 220280 181595 220282
rect 180750 220224 181534 220280
rect 181590 220224 181595 220280
rect 180750 220222 181595 220224
rect 576810 220282 576870 220630
rect 674097 220688 676292 220690
rect 674097 220632 674102 220688
rect 674158 220632 676292 220688
rect 674097 220630 676292 220632
rect 674097 220627 674163 220630
rect 654133 220418 654199 220421
rect 667013 220418 667079 220421
rect 654133 220416 667079 220418
rect 654133 220360 654138 220416
rect 654194 220360 667018 220416
rect 667074 220360 667079 220416
rect 654133 220358 667079 220360
rect 654133 220355 654199 220358
rect 667013 220355 667079 220358
rect 582465 220282 582531 220285
rect 576810 220280 582531 220282
rect 576810 220224 582470 220280
rect 582526 220224 582531 220280
rect 576810 220222 582531 220224
rect 166947 220146 167013 220149
rect 175549 220146 175615 220149
rect 166947 220144 175615 220146
rect 166947 220088 166952 220144
rect 167008 220088 175554 220144
rect 175610 220088 175615 220144
rect 166947 220086 175615 220088
rect 166947 220083 167013 220086
rect 175549 220083 175615 220086
rect 180517 220146 180583 220149
rect 180750 220146 180810 220222
rect 181529 220219 181595 220222
rect 582465 220219 582531 220222
rect 674649 220282 674715 220285
rect 674649 220280 676292 220282
rect 674649 220224 674654 220280
rect 674710 220224 676292 220280
rect 674649 220222 676292 220224
rect 674649 220219 674715 220222
rect 180517 220144 180810 220146
rect 180517 220088 180522 220144
rect 180578 220088 180810 220144
rect 180517 220086 180810 220088
rect 600129 220146 600195 220149
rect 601141 220146 601207 220149
rect 600129 220144 601207 220146
rect 600129 220088 600134 220144
rect 600190 220088 601146 220144
rect 601202 220088 601207 220144
rect 600129 220086 601207 220088
rect 180517 220083 180583 220086
rect 600129 220083 600195 220086
rect 601141 220083 601207 220086
rect 673545 220146 673611 220149
rect 674097 220146 674163 220149
rect 673545 220144 674163 220146
rect 673545 220088 673550 220144
rect 673606 220088 674102 220144
rect 674158 220088 674163 220144
rect 673545 220086 674163 220088
rect 673545 220083 673611 220086
rect 674097 220083 674163 220086
rect 180885 220010 180951 220013
rect 185117 220010 185183 220013
rect 180885 220008 185183 220010
rect 180885 219952 180890 220008
rect 180946 219952 185122 220008
rect 185178 219952 185183 220008
rect 180885 219950 185183 219952
rect 180885 219947 180951 219950
rect 185117 219947 185183 219950
rect 562869 220010 562935 220013
rect 563053 220010 563119 220013
rect 562869 220008 563119 220010
rect 562869 219952 562874 220008
rect 562930 219952 563058 220008
rect 563114 219952 563119 220008
rect 562869 219950 563119 219952
rect 562869 219947 562935 219950
rect 563053 219947 563119 219950
rect 564801 220010 564867 220013
rect 572529 220010 572595 220013
rect 564801 220008 572595 220010
rect 564801 219952 564806 220008
rect 564862 219952 572534 220008
rect 572590 219952 572595 220008
rect 564801 219950 572595 219952
rect 564801 219947 564867 219950
rect 572529 219947 572595 219950
rect 576577 220010 576643 220013
rect 581821 220010 581887 220013
rect 576577 220008 581887 220010
rect 576577 219952 576582 220008
rect 576638 219952 581826 220008
rect 581882 219952 581887 220008
rect 576577 219950 581887 219952
rect 576577 219947 576643 219950
rect 581821 219947 581887 219950
rect 582649 220010 582715 220013
rect 591941 220010 592007 220013
rect 582649 220008 592007 220010
rect 582649 219952 582654 220008
rect 582710 219952 591946 220008
rect 592002 219952 592007 220008
rect 582649 219950 592007 219952
rect 582649 219947 582715 219950
rect 591941 219947 592007 219950
rect 140773 219874 140839 219877
rect 142153 219874 142219 219877
rect 140773 219872 142219 219874
rect 140773 219816 140778 219872
rect 140834 219816 142158 219872
rect 142214 219816 142219 219872
rect 140773 219814 142219 219816
rect 140773 219811 140839 219814
rect 142153 219811 142219 219814
rect 646037 219874 646103 219877
rect 675017 219874 675083 219877
rect 683297 219874 683363 219877
rect 646037 219872 675083 219874
rect 646037 219816 646042 219872
rect 646098 219816 675022 219872
rect 675078 219816 675083 219872
rect 646037 219814 675083 219816
rect 683284 219872 683363 219874
rect 683284 219816 683302 219872
rect 683358 219816 683363 219872
rect 683284 219814 683363 219816
rect 646037 219811 646103 219814
rect 675017 219811 675083 219814
rect 683297 219811 683363 219814
rect 611445 219738 611511 219741
rect 489870 219736 611511 219738
rect 489870 219680 611450 219736
rect 611506 219680 611511 219736
rect 489870 219678 611511 219680
rect 142153 219602 142219 219605
rect 147765 219602 147831 219605
rect 142153 219600 147831 219602
rect 142153 219544 142158 219600
rect 142214 219544 147770 219600
rect 147826 219544 147831 219600
rect 142153 219542 147831 219544
rect 142153 219539 142219 219542
rect 147765 219539 147831 219542
rect 151629 219602 151695 219605
rect 153653 219602 153719 219605
rect 151629 219600 153719 219602
rect 151629 219544 151634 219600
rect 151690 219544 153658 219600
rect 153714 219544 153719 219600
rect 151629 219542 153719 219544
rect 151629 219539 151695 219542
rect 153653 219539 153719 219542
rect 486969 219466 487035 219469
rect 489870 219466 489930 219678
rect 611445 219675 611511 219678
rect 486969 219464 489930 219466
rect 486969 219408 486974 219464
rect 487030 219408 489930 219464
rect 486969 219406 489930 219408
rect 515213 219466 515279 219469
rect 617241 219466 617307 219469
rect 515213 219464 617307 219466
rect 515213 219408 515218 219464
rect 515274 219408 617246 219464
rect 617302 219408 617307 219464
rect 515213 219406 617307 219408
rect 486969 219403 487035 219406
rect 515213 219403 515279 219406
rect 617241 219403 617307 219406
rect 667013 219466 667079 219469
rect 667013 219464 676292 219466
rect 667013 219408 667018 219464
rect 667074 219408 676292 219464
rect 667013 219406 676292 219408
rect 667013 219403 667079 219406
rect 567285 219194 567351 219197
rect 571517 219194 571583 219197
rect 567285 219192 571583 219194
rect 567285 219136 567290 219192
rect 567346 219136 571522 219192
rect 571578 219136 571583 219192
rect 567285 219134 571583 219136
rect 567285 219131 567351 219134
rect 571517 219131 571583 219134
rect 674925 219058 674991 219061
rect 674925 219056 676292 219058
rect 674925 219000 674930 219056
rect 674986 219000 676292 219056
rect 674925 218998 676292 219000
rect 674925 218995 674991 218998
rect 494697 218922 494763 218925
rect 656801 218922 656867 218925
rect 670785 218922 670851 218925
rect 494697 218920 596190 218922
rect 494697 218864 494702 218920
rect 494758 218864 596190 218920
rect 494697 218862 596190 218864
rect 494697 218859 494763 218862
rect 490373 218650 490439 218653
rect 594793 218650 594859 218653
rect 490373 218648 594859 218650
rect 490373 218592 490378 218648
rect 490434 218592 594798 218648
rect 594854 218592 594859 218648
rect 490373 218590 594859 218592
rect 596130 218650 596190 218862
rect 656801 218920 670851 218922
rect 656801 218864 656806 218920
rect 656862 218864 670790 218920
rect 670846 218864 670851 218920
rect 656801 218862 670851 218864
rect 656801 218859 656867 218862
rect 670785 218859 670851 218862
rect 648613 218650 648679 218653
rect 675385 218650 675451 218653
rect 596130 218590 605850 218650
rect 490373 218587 490439 218590
rect 594793 218587 594859 218590
rect 170949 218514 171015 218517
rect 172881 218514 172947 218517
rect 170949 218512 172947 218514
rect 170949 218456 170954 218512
rect 171010 218456 172886 218512
rect 172942 218456 172947 218512
rect 170949 218454 172947 218456
rect 170949 218451 171015 218454
rect 172881 218451 172947 218454
rect 492673 218378 492739 218381
rect 493777 218378 493843 218381
rect 492673 218376 493843 218378
rect 492673 218320 492678 218376
rect 492734 218320 493782 218376
rect 493838 218320 493843 218376
rect 492673 218318 493843 218320
rect 492673 218315 492739 218318
rect 493777 218315 493843 218318
rect 496905 218378 496971 218381
rect 603349 218378 603415 218381
rect 496905 218376 603415 218378
rect 496905 218320 496910 218376
rect 496966 218320 603354 218376
rect 603410 218320 603415 218376
rect 496905 218318 603415 218320
rect 605790 218378 605850 218590
rect 648613 218648 675451 218650
rect 648613 218592 648618 218648
rect 648674 218592 675390 218648
rect 675446 218592 675451 218648
rect 648613 218590 675451 218592
rect 648613 218587 648679 218590
rect 675385 218587 675451 218590
rect 675702 218588 675708 218652
rect 675772 218650 675778 218652
rect 675772 218590 676292 218650
rect 675772 218588 675778 218590
rect 631133 218378 631199 218381
rect 605790 218376 631199 218378
rect 605790 218320 631138 218376
rect 631194 218320 631199 218376
rect 605790 218318 631199 218320
rect 496905 218315 496971 218318
rect 603349 218315 603415 218318
rect 631133 218315 631199 218318
rect 675293 218242 675359 218245
rect 675293 218240 676292 218242
rect 675293 218184 675298 218240
rect 675354 218184 676292 218240
rect 675293 218182 676292 218184
rect 675293 218179 675359 218182
rect 487797 218106 487863 218109
rect 627453 218106 627519 218109
rect 487797 218104 627519 218106
rect 487797 218048 487802 218104
rect 487858 218048 627458 218104
rect 627514 218048 627519 218104
rect 487797 218046 627519 218048
rect 487797 218043 487863 218046
rect 627453 218043 627519 218046
rect 35801 217970 35867 217973
rect 61285 217970 61351 217973
rect 675661 217970 675727 217973
rect 35801 217968 61351 217970
rect 35801 217912 35806 217968
rect 35862 217912 61290 217968
rect 61346 217912 61351 217968
rect 35801 217910 61351 217912
rect 35801 217907 35867 217910
rect 61285 217907 61351 217910
rect 672950 217968 675727 217970
rect 672950 217912 675666 217968
rect 675722 217912 675727 217968
rect 672950 217910 675727 217912
rect 508497 217834 508563 217837
rect 510153 217836 510219 217837
rect 509182 217834 509188 217836
rect 508497 217832 509188 217834
rect 508497 217776 508502 217832
rect 508558 217776 509188 217832
rect 508497 217774 509188 217776
rect 508497 217771 508563 217774
rect 509182 217772 509188 217774
rect 509252 217772 509258 217836
rect 510102 217834 510108 217836
rect 510062 217774 510108 217834
rect 510172 217832 510219 217836
rect 522573 217836 522639 217837
rect 522573 217834 522620 217836
rect 510214 217776 510219 217832
rect 510102 217772 510108 217774
rect 510172 217772 510219 217776
rect 522528 217832 522620 217834
rect 522528 217776 522578 217832
rect 522528 217774 522620 217776
rect 510153 217771 510219 217772
rect 522573 217772 522620 217774
rect 522684 217772 522690 217836
rect 555693 217834 555759 217837
rect 562685 217834 562751 217837
rect 555693 217832 562751 217834
rect 555693 217776 555698 217832
rect 555754 217776 562690 217832
rect 562746 217776 562751 217832
rect 555693 217774 562751 217776
rect 522573 217771 522639 217772
rect 555693 217771 555759 217774
rect 562685 217771 562751 217774
rect 562869 217834 562935 217837
rect 563605 217834 563671 217837
rect 570965 217836 571031 217837
rect 571333 217836 571399 217837
rect 570965 217834 571012 217836
rect 562869 217832 563671 217834
rect 562869 217776 562874 217832
rect 562930 217776 563610 217832
rect 563666 217776 563671 217832
rect 562869 217774 563671 217776
rect 570920 217832 571012 217834
rect 570920 217776 570970 217832
rect 570920 217774 571012 217776
rect 562869 217771 562935 217774
rect 563605 217771 563671 217774
rect 570965 217772 571012 217774
rect 571076 217772 571082 217836
rect 571333 217834 571380 217836
rect 571288 217832 571380 217834
rect 571288 217776 571338 217832
rect 571288 217774 571380 217776
rect 571333 217772 571380 217774
rect 571444 217772 571450 217836
rect 572437 217834 572503 217837
rect 574093 217834 574159 217837
rect 572437 217832 574159 217834
rect 572437 217776 572442 217832
rect 572498 217776 574098 217832
rect 574154 217776 574159 217832
rect 572437 217774 574159 217776
rect 570965 217771 571031 217772
rect 571333 217771 571399 217772
rect 572437 217771 572503 217774
rect 574093 217771 574159 217774
rect 574318 217772 574324 217836
rect 574388 217834 574394 217836
rect 574553 217834 574619 217837
rect 574388 217832 574619 217834
rect 574388 217776 574558 217832
rect 574614 217776 574619 217832
rect 574388 217774 574619 217776
rect 574388 217772 574394 217774
rect 574553 217771 574619 217774
rect 651097 217834 651163 217837
rect 664253 217834 664319 217837
rect 672073 217834 672139 217837
rect 651097 217832 664319 217834
rect 651097 217776 651102 217832
rect 651158 217776 664258 217832
rect 664314 217776 664319 217832
rect 651097 217774 664319 217776
rect 651097 217771 651163 217774
rect 664253 217771 664319 217774
rect 664486 217832 672139 217834
rect 664486 217776 672078 217832
rect 672134 217776 672139 217832
rect 664486 217774 672139 217776
rect 505645 217562 505711 217565
rect 595161 217562 595227 217565
rect 505645 217560 595227 217562
rect 505645 217504 505650 217560
rect 505706 217504 595166 217560
rect 595222 217504 595227 217560
rect 505645 217502 595227 217504
rect 505645 217499 505711 217502
rect 595161 217499 595227 217502
rect 653765 217562 653831 217565
rect 664486 217562 664546 217774
rect 672073 217771 672139 217774
rect 670601 217562 670667 217565
rect 653765 217560 664546 217562
rect 653765 217504 653770 217560
rect 653826 217504 664546 217560
rect 653765 217502 664546 217504
rect 669270 217560 670667 217562
rect 669270 217504 670606 217560
rect 670662 217504 670667 217560
rect 669270 217502 670667 217504
rect 653765 217499 653831 217502
rect 493777 217292 493843 217293
rect 493726 217228 493732 217292
rect 493796 217290 493843 217292
rect 495341 217290 495407 217293
rect 498469 217290 498535 217293
rect 596357 217290 596423 217293
rect 493796 217288 493888 217290
rect 493838 217232 493888 217288
rect 493796 217230 493888 217232
rect 495341 217288 495450 217290
rect 495341 217232 495346 217288
rect 495402 217232 495450 217288
rect 493796 217228 493843 217230
rect 493777 217227 493843 217228
rect 495341 217227 495450 217232
rect 498469 217288 596423 217290
rect 498469 217232 498474 217288
rect 498530 217232 596362 217288
rect 596418 217232 596423 217288
rect 498469 217230 596423 217232
rect 498469 217227 498535 217230
rect 596357 217227 596423 217230
rect 664253 217290 664319 217293
rect 669270 217290 669330 217502
rect 670601 217499 670667 217502
rect 672073 217562 672139 217565
rect 672950 217562 673010 217910
rect 675661 217907 675727 217910
rect 675886 217908 675892 217972
rect 675956 217970 675962 217972
rect 675956 217910 676230 217970
rect 675956 217908 675962 217910
rect 676170 217834 676230 217910
rect 676170 217774 676292 217834
rect 672073 217560 673010 217562
rect 672073 217504 672078 217560
rect 672134 217504 673010 217560
rect 672073 217502 673010 217504
rect 673177 217562 673243 217565
rect 676029 217562 676095 217565
rect 673177 217560 676095 217562
rect 673177 217504 673182 217560
rect 673238 217504 676034 217560
rect 676090 217504 676095 217560
rect 673177 217502 676095 217504
rect 672073 217499 672139 217502
rect 673177 217499 673243 217502
rect 676029 217499 676095 217502
rect 676170 217366 676292 217426
rect 676170 217290 676230 217366
rect 664253 217288 669330 217290
rect 664253 217232 664258 217288
rect 664314 217232 669330 217288
rect 664253 217230 669330 217232
rect 672766 217230 676230 217290
rect 664253 217227 664319 217230
rect 488671 217154 488737 217157
rect 488671 217152 489930 217154
rect 488671 217096 488676 217152
rect 488732 217096 489930 217152
rect 488671 217094 489930 217096
rect 488671 217091 488737 217094
rect 489870 216746 489930 217094
rect 495390 217018 495450 217227
rect 595713 217018 595779 217021
rect 495390 217016 595779 217018
rect 495390 216960 595718 217016
rect 595774 216960 595779 217016
rect 495390 216958 595779 216960
rect 595713 216955 595779 216958
rect 574093 216746 574159 216749
rect 574369 216748 574435 216749
rect 489870 216744 574159 216746
rect 489870 216688 574098 216744
rect 574154 216688 574159 216744
rect 489870 216686 574159 216688
rect 574093 216683 574159 216686
rect 574318 216684 574324 216748
rect 574388 216746 574435 216748
rect 666829 216746 666895 216749
rect 672766 216746 672826 217230
rect 673361 217018 673427 217021
rect 673361 217016 676292 217018
rect 673361 216960 673366 217016
rect 673422 216960 676292 217016
rect 673361 216958 676292 216960
rect 673361 216955 673427 216958
rect 574388 216744 574480 216746
rect 574430 216688 574480 216744
rect 574388 216686 574480 216688
rect 666829 216744 672826 216746
rect 666829 216688 666834 216744
rect 666890 216688 672826 216744
rect 666829 216686 672826 216688
rect 574388 216684 574435 216686
rect 574369 216683 574435 216684
rect 666829 216683 666895 216686
rect 675886 216548 675892 216612
rect 675956 216610 675962 216612
rect 675956 216550 676292 216610
rect 675956 216548 675962 216550
rect 571006 216412 571012 216476
rect 571076 216474 571082 216476
rect 574921 216474 574987 216477
rect 571076 216472 574987 216474
rect 571076 216416 574926 216472
rect 574982 216416 574987 216472
rect 571076 216414 574987 216416
rect 571076 216412 571082 216414
rect 574921 216411 574987 216414
rect 664713 216474 664779 216477
rect 675661 216474 675727 216477
rect 664713 216472 675727 216474
rect 664713 216416 664718 216472
rect 664774 216416 675666 216472
rect 675722 216416 675727 216472
rect 664713 216414 675727 216416
rect 664713 216411 664779 216414
rect 675661 216411 675727 216414
rect 571374 216140 571380 216204
rect 571444 216202 571450 216204
rect 627913 216202 627979 216205
rect 571444 216200 627979 216202
rect 571444 216144 627918 216200
rect 627974 216144 627979 216200
rect 571444 216142 627979 216144
rect 571444 216140 571450 216142
rect 627913 216139 627979 216142
rect 674741 216202 674807 216205
rect 674741 216200 676292 216202
rect 674741 216144 674746 216200
rect 674802 216144 676292 216200
rect 674741 216142 676292 216144
rect 674741 216139 674807 216142
rect 509182 215868 509188 215932
rect 509252 215930 509258 215932
rect 598473 215930 598539 215933
rect 509252 215928 598539 215930
rect 509252 215872 598478 215928
rect 598534 215872 598539 215928
rect 509252 215870 598539 215872
rect 509252 215868 509258 215870
rect 598473 215867 598539 215870
rect 656525 215930 656591 215933
rect 672257 215930 672323 215933
rect 656525 215928 672323 215930
rect 656525 215872 656530 215928
rect 656586 215872 672262 215928
rect 672318 215872 672323 215928
rect 656525 215870 672323 215872
rect 656525 215867 656591 215870
rect 672257 215867 672323 215870
rect 676170 215734 676292 215794
rect 666645 215658 666711 215661
rect 676170 215658 676230 215734
rect 666645 215656 676230 215658
rect 666645 215600 666650 215656
rect 666706 215600 676230 215656
rect 666645 215598 676230 215600
rect 666645 215595 666711 215598
rect 522614 215324 522620 215388
rect 522684 215386 522690 215388
rect 618897 215386 618963 215389
rect 522684 215384 618963 215386
rect 522684 215328 618902 215384
rect 618958 215328 618963 215384
rect 522684 215326 618963 215328
rect 522684 215324 522690 215326
rect 618897 215323 618963 215326
rect 676029 215386 676095 215389
rect 676029 215384 676292 215386
rect 676029 215328 676034 215384
rect 676090 215328 676292 215384
rect 676029 215326 676292 215328
rect 676029 215323 676095 215326
rect 675661 215250 675727 215253
rect 669270 215248 675727 215250
rect 669270 215192 675666 215248
rect 675722 215192 675727 215248
rect 669270 215190 675727 215192
rect 660389 215114 660455 215117
rect 669270 215114 669330 215190
rect 675661 215187 675727 215190
rect 660389 215112 669330 215114
rect 660389 215056 660394 215112
rect 660450 215056 669330 215112
rect 660389 215054 669330 215056
rect 660389 215051 660455 215054
rect 47945 214978 48011 214981
rect 41492 214976 48011 214978
rect 41492 214920 47950 214976
rect 48006 214920 48011 214976
rect 41492 214918 48011 214920
rect 47945 214915 48011 214918
rect 673545 214978 673611 214981
rect 673545 214976 676292 214978
rect 673545 214920 673550 214976
rect 673606 214920 676292 214976
rect 673545 214918 676292 214920
rect 673545 214915 673611 214918
rect 35801 214706 35867 214709
rect 35758 214704 35867 214706
rect 35758 214648 35806 214704
rect 35862 214648 35867 214704
rect 35758 214643 35867 214648
rect 35758 214540 35818 214643
rect 672993 214570 673059 214573
rect 672993 214568 676292 214570
rect 672993 214512 672998 214568
rect 673054 214512 676292 214568
rect 672993 214510 676292 214512
rect 672993 214507 673059 214510
rect 35801 214298 35867 214301
rect 35758 214296 35867 214298
rect 35758 214240 35806 214296
rect 35862 214240 35867 214296
rect 35758 214235 35867 214240
rect 39665 214298 39731 214301
rect 43805 214298 43871 214301
rect 39665 214296 43871 214298
rect 39665 214240 39670 214296
rect 39726 214240 43810 214296
rect 43866 214240 43871 214296
rect 39665 214238 43871 214240
rect 39665 214235 39731 214238
rect 43805 214235 43871 214238
rect 35758 214132 35818 214235
rect 575982 214026 576042 214404
rect 670785 214162 670851 214165
rect 670785 214160 676292 214162
rect 670785 214104 670790 214160
rect 670846 214104 676292 214160
rect 670785 214102 676292 214104
rect 670785 214099 670851 214102
rect 578877 214026 578943 214029
rect 575982 214024 578943 214026
rect 575982 213968 578882 214024
rect 578938 213968 578943 214024
rect 575982 213966 578943 213968
rect 578877 213963 578943 213966
rect 44357 213754 44423 213757
rect 41492 213752 44423 213754
rect 41492 213696 44362 213752
rect 44418 213696 44423 213752
rect 41492 213694 44423 213696
rect 44357 213691 44423 213694
rect 659377 213754 659443 213757
rect 672073 213754 672139 213757
rect 659377 213752 672139 213754
rect 659377 213696 659382 213752
rect 659438 213696 672078 213752
rect 672134 213696 672139 213752
rect 659377 213694 672139 213696
rect 659377 213691 659443 213694
rect 672073 213691 672139 213694
rect 674281 213754 674347 213757
rect 674281 213752 676292 213754
rect 674281 213696 674286 213752
rect 674342 213696 676292 213752
rect 674281 213694 676292 213696
rect 674281 213691 674347 213694
rect 661493 213482 661559 213485
rect 661493 213480 669330 213482
rect 661493 213424 661498 213480
rect 661554 213424 669330 213480
rect 661493 213422 669330 213424
rect 661493 213419 661559 213422
rect 47761 213346 47827 213349
rect 41492 213344 47827 213346
rect 41492 213288 47766 213344
rect 47822 213288 47827 213344
rect 41492 213286 47827 213288
rect 47761 213283 47827 213286
rect 669270 213074 669330 213422
rect 672073 213346 672139 213349
rect 672073 213344 676292 213346
rect 672073 213288 672078 213344
rect 672134 213288 676292 213344
rect 672073 213286 676292 213288
rect 672073 213283 672139 213286
rect 674465 213074 674531 213077
rect 669270 213072 674531 213074
rect 669270 213016 674470 213072
rect 674526 213016 674531 213072
rect 669270 213014 674531 213016
rect 674465 213011 674531 213014
rect 44817 212938 44883 212941
rect 41492 212936 44883 212938
rect 41492 212880 44822 212936
rect 44878 212880 44883 212936
rect 41492 212878 44883 212880
rect 44817 212875 44883 212878
rect 683070 212533 683130 212908
rect 683070 212528 683179 212533
rect 683070 212500 683118 212528
rect 35758 212261 35818 212500
rect 683100 212472 683118 212500
rect 683174 212472 683179 212528
rect 683100 212470 683179 212472
rect 683113 212467 683179 212470
rect 35758 212256 35867 212261
rect 35758 212200 35806 212256
rect 35862 212200 35867 212256
rect 35758 212198 35867 212200
rect 35801 212195 35867 212198
rect 44173 212122 44239 212125
rect 41492 212120 44239 212122
rect 41492 212064 44178 212120
rect 44234 212064 44239 212120
rect 41492 212062 44239 212064
rect 44173 212059 44239 212062
rect 35617 211850 35683 211853
rect 35574 211848 35683 211850
rect 35574 211792 35622 211848
rect 35678 211792 35683 211848
rect 35574 211787 35683 211792
rect 40125 211850 40191 211853
rect 42793 211850 42859 211853
rect 40125 211848 42859 211850
rect 40125 211792 40130 211848
rect 40186 211792 42798 211848
rect 42854 211792 42859 211848
rect 40125 211790 42859 211792
rect 40125 211787 40191 211790
rect 42793 211787 42859 211790
rect 35574 211684 35634 211787
rect 575982 211714 576042 212228
rect 672257 212122 672323 212125
rect 672257 212120 676292 212122
rect 672257 212064 672262 212120
rect 672318 212064 676292 212120
rect 672257 212062 676292 212064
rect 672257 212059 672323 212062
rect 578325 211714 578391 211717
rect 575982 211712 578391 211714
rect 575982 211656 578330 211712
rect 578386 211656 578391 211712
rect 575982 211654 578391 211656
rect 578325 211651 578391 211654
rect 35801 211442 35867 211445
rect 675477 211444 675543 211445
rect 675477 211442 675524 211444
rect 35758 211440 35867 211442
rect 35758 211384 35806 211440
rect 35862 211384 35867 211440
rect 35758 211379 35867 211384
rect 675396 211440 675524 211442
rect 675588 211442 675594 211444
rect 683113 211442 683179 211445
rect 675588 211440 683179 211442
rect 675396 211384 675482 211440
rect 675588 211384 683118 211440
rect 683174 211384 683179 211440
rect 675396 211382 675524 211384
rect 675477 211380 675524 211382
rect 675588 211382 683179 211384
rect 675588 211380 675594 211382
rect 675477 211379 675543 211380
rect 683113 211379 683179 211382
rect 35758 211276 35818 211379
rect 676581 211172 676647 211173
rect 676581 211168 676628 211172
rect 676692 211170 676698 211172
rect 676581 211112 676586 211168
rect 676581 211108 676628 211112
rect 676692 211110 676738 211170
rect 676692 211108 676698 211110
rect 676581 211107 676647 211108
rect 47945 210898 48011 210901
rect 41492 210896 48011 210898
rect 41492 210840 47950 210896
rect 48006 210840 48011 210896
rect 41492 210838 48011 210840
rect 47945 210835 48011 210838
rect 35574 210221 35634 210460
rect 35525 210216 35634 210221
rect 35801 210218 35867 210221
rect 35525 210160 35530 210216
rect 35586 210160 35634 210216
rect 35525 210158 35634 210160
rect 35758 210216 35867 210218
rect 35758 210160 35806 210216
rect 35862 210160 35867 210216
rect 35525 210155 35591 210158
rect 35758 210155 35867 210160
rect 35758 210052 35818 210155
rect 575982 209810 576042 210052
rect 579521 209810 579587 209813
rect 575982 209808 579587 209810
rect 575982 209752 579526 209808
rect 579582 209752 579587 209808
rect 575982 209750 579587 209752
rect 579521 209747 579587 209750
rect 35758 209405 35818 209644
rect 35758 209400 35867 209405
rect 35758 209344 35806 209400
rect 35862 209344 35867 209400
rect 35758 209342 35867 209344
rect 35801 209339 35867 209342
rect 40769 209402 40835 209405
rect 42977 209402 43043 209405
rect 40769 209400 43043 209402
rect 40769 209344 40774 209400
rect 40830 209344 42982 209400
rect 43038 209344 43043 209400
rect 40769 209342 43043 209344
rect 40769 209339 40835 209342
rect 42977 209339 43043 209342
rect 32998 208997 33058 209236
rect 32998 208992 33107 208997
rect 32998 208936 33046 208992
rect 33102 208936 33107 208992
rect 32998 208934 33107 208936
rect 33041 208931 33107 208934
rect 46933 208858 46999 208861
rect 41492 208856 46999 208858
rect 41492 208800 46938 208856
rect 46994 208800 46999 208856
rect 41492 208798 46999 208800
rect 46933 208795 46999 208798
rect 47117 208450 47183 208453
rect 41492 208448 47183 208450
rect 41492 208392 47122 208448
rect 47178 208392 47183 208448
rect 41492 208390 47183 208392
rect 47117 208387 47183 208390
rect 41505 208178 41571 208181
rect 49601 208178 49667 208181
rect 41505 208176 49667 208178
rect 41505 208120 41510 208176
rect 41566 208120 49606 208176
rect 49662 208120 49667 208176
rect 41505 208118 49667 208120
rect 41505 208115 41571 208118
rect 49601 208115 49667 208118
rect 589457 208042 589523 208045
rect 589457 208040 592572 208042
rect 35758 207773 35818 208012
rect 589457 207984 589462 208040
rect 589518 207984 592572 208040
rect 589457 207982 592572 207984
rect 589457 207979 589523 207982
rect 35758 207768 35867 207773
rect 35758 207712 35806 207768
rect 35862 207712 35867 207768
rect 35758 207710 35867 207712
rect 35801 207707 35867 207710
rect 40902 207708 40908 207772
rect 40972 207708 40978 207772
rect 40910 207604 40970 207708
rect 575982 207498 576042 207876
rect 579521 207498 579587 207501
rect 575982 207496 579587 207498
rect 575982 207440 579526 207496
rect 579582 207440 579587 207496
rect 575982 207438 579587 207440
rect 579521 207435 579587 207438
rect 40125 207362 40191 207365
rect 42006 207362 42012 207364
rect 40125 207360 42012 207362
rect 40125 207304 40130 207360
rect 40186 207304 42012 207360
rect 40125 207302 42012 207304
rect 40125 207299 40191 207302
rect 42006 207300 42012 207302
rect 42076 207300 42082 207364
rect 40542 206956 40602 207196
rect 40534 206892 40540 206956
rect 40604 206892 40610 206956
rect 672441 206954 672507 206957
rect 675477 206954 675543 206957
rect 672441 206952 675543 206954
rect 672441 206896 672446 206952
rect 672502 206896 675482 206952
rect 675538 206896 675543 206952
rect 672441 206894 675543 206896
rect 672441 206891 672507 206894
rect 675477 206891 675543 206894
rect 44357 206818 44423 206821
rect 41492 206816 44423 206818
rect 41492 206760 44362 206816
rect 44418 206760 44423 206816
rect 41492 206758 44423 206760
rect 44357 206755 44423 206758
rect 40953 206546 41019 206549
rect 43161 206546 43227 206549
rect 40953 206544 43227 206546
rect 40953 206488 40958 206544
rect 41014 206488 43166 206544
rect 43222 206488 43227 206544
rect 40953 206486 43227 206488
rect 40953 206483 41019 206486
rect 43161 206483 43227 206486
rect 589457 206410 589523 206413
rect 589457 206408 592572 206410
rect 40726 206140 40786 206380
rect 589457 206352 589462 206408
rect 589518 206352 592572 206408
rect 589457 206350 592572 206352
rect 589457 206347 589523 206350
rect 40718 206076 40724 206140
rect 40788 206076 40794 206140
rect 44173 206002 44239 206005
rect 41492 206000 44239 206002
rect 41492 205944 44178 206000
rect 44234 205944 44239 206000
rect 41492 205942 44239 205944
rect 44173 205939 44239 205942
rect 579521 205866 579587 205869
rect 575798 205864 579587 205866
rect 575798 205808 579526 205864
rect 579582 205808 579587 205864
rect 575798 205806 579587 205808
rect 40769 205730 40835 205733
rect 42793 205730 42859 205733
rect 40769 205728 42859 205730
rect 40769 205672 40774 205728
rect 40830 205672 42798 205728
rect 42854 205672 42859 205728
rect 575798 205700 575858 205806
rect 579521 205803 579587 205806
rect 40769 205670 42859 205672
rect 40769 205667 40835 205670
rect 42793 205667 42859 205670
rect 35574 205325 35634 205564
rect 35574 205320 35683 205325
rect 35574 205264 35622 205320
rect 35678 205264 35683 205320
rect 35574 205262 35683 205264
rect 35617 205259 35683 205262
rect 44541 205186 44607 205189
rect 41492 205184 44607 205186
rect 41492 205128 44546 205184
rect 44602 205128 44607 205184
rect 41492 205126 44607 205128
rect 44541 205123 44607 205126
rect 675753 205050 675819 205053
rect 676254 205050 676260 205052
rect 675753 205048 676260 205050
rect 675753 204992 675758 205048
rect 675814 204992 676260 205048
rect 675753 204990 676260 204992
rect 675753 204987 675819 204990
rect 676254 204988 676260 204990
rect 676324 204988 676330 205052
rect 44817 204778 44883 204781
rect 41492 204776 44883 204778
rect 41492 204720 44822 204776
rect 44878 204720 44883 204776
rect 41492 204718 44883 204720
rect 44817 204715 44883 204718
rect 589457 204778 589523 204781
rect 589457 204776 592572 204778
rect 589457 204720 589462 204776
rect 589518 204720 592572 204776
rect 589457 204718 592572 204720
rect 589457 204715 589523 204718
rect 35801 204506 35867 204509
rect 35758 204504 35867 204506
rect 35758 204448 35806 204504
rect 35862 204448 35867 204504
rect 35758 204443 35867 204448
rect 41689 204506 41755 204509
rect 43805 204506 43871 204509
rect 41689 204504 43871 204506
rect 41689 204448 41694 204504
rect 41750 204448 43810 204504
rect 43866 204448 43871 204504
rect 41689 204446 43871 204448
rect 41689 204443 41755 204446
rect 43805 204443 43871 204446
rect 35758 204340 35818 204443
rect 41689 204098 41755 204101
rect 43989 204098 44055 204101
rect 41689 204096 44055 204098
rect 41689 204040 41694 204096
rect 41750 204040 43994 204096
rect 44050 204040 44055 204096
rect 41689 204038 44055 204040
rect 41689 204035 41755 204038
rect 43989 204035 44055 204038
rect 35758 203693 35818 203932
rect 35758 203688 35867 203693
rect 35758 203632 35806 203688
rect 35862 203632 35867 203688
rect 35758 203630 35867 203632
rect 35801 203627 35867 203630
rect 46197 203554 46263 203557
rect 41492 203552 46263 203554
rect 41492 203496 46202 203552
rect 46258 203496 46263 203552
rect 41492 203494 46263 203496
rect 46197 203491 46263 203494
rect 575982 203282 576042 203524
rect 578325 203282 578391 203285
rect 575982 203280 578391 203282
rect 575982 203224 578330 203280
rect 578386 203224 578391 203280
rect 575982 203222 578391 203224
rect 578325 203219 578391 203222
rect 589457 203146 589523 203149
rect 589457 203144 592572 203146
rect 589457 203088 589462 203144
rect 589518 203088 592572 203144
rect 589457 203086 592572 203088
rect 589457 203083 589523 203086
rect 672533 203012 672599 203013
rect 672533 203010 672580 203012
rect 672488 203008 672580 203010
rect 672488 202952 672538 203008
rect 672488 202950 672580 202952
rect 672533 202948 672580 202950
rect 672644 202948 672650 203012
rect 672533 202947 672599 202948
rect 675753 202738 675819 202741
rect 676438 202738 676444 202740
rect 675753 202736 676444 202738
rect 675753 202680 675758 202736
rect 675814 202680 676444 202736
rect 675753 202678 676444 202680
rect 675753 202675 675819 202678
rect 676438 202676 676444 202678
rect 676508 202676 676514 202740
rect 33041 202194 33107 202197
rect 41638 202194 41644 202196
rect 33041 202192 41644 202194
rect 33041 202136 33046 202192
rect 33102 202136 41644 202192
rect 33041 202134 41644 202136
rect 33041 202131 33107 202134
rect 41638 202132 41644 202134
rect 41708 202132 41714 202196
rect 41873 202194 41939 202197
rect 48589 202194 48655 202197
rect 41873 202192 48655 202194
rect 41873 202136 41878 202192
rect 41934 202136 48594 202192
rect 48650 202136 48655 202192
rect 41873 202134 48655 202136
rect 41873 202131 41939 202134
rect 48589 202131 48655 202134
rect 674741 201922 674807 201925
rect 675385 201922 675451 201925
rect 674741 201920 675451 201922
rect 674741 201864 674746 201920
rect 674802 201864 675390 201920
rect 675446 201864 675451 201920
rect 674741 201862 675451 201864
rect 674741 201859 674807 201862
rect 675385 201859 675451 201862
rect 589457 201514 589523 201517
rect 589457 201512 592572 201514
rect 589457 201456 589462 201512
rect 589518 201456 592572 201512
rect 589457 201454 592572 201456
rect 589457 201451 589523 201454
rect 575982 200834 576042 201348
rect 578785 200834 578851 200837
rect 575982 200832 578851 200834
rect 575982 200776 578790 200832
rect 578846 200776 578851 200832
rect 575982 200774 578851 200776
rect 578785 200771 578851 200774
rect 35801 200698 35867 200701
rect 41822 200698 41828 200700
rect 35801 200696 41828 200698
rect 35801 200640 35806 200696
rect 35862 200640 41828 200696
rect 35801 200638 41828 200640
rect 35801 200635 35867 200638
rect 41822 200636 41828 200638
rect 41892 200636 41898 200700
rect 672993 200562 673059 200565
rect 675477 200562 675543 200565
rect 672993 200560 675543 200562
rect 672993 200504 672998 200560
rect 673054 200504 675482 200560
rect 675538 200504 675543 200560
rect 672993 200502 675543 200504
rect 672993 200499 673059 200502
rect 675477 200499 675543 200502
rect 589457 199882 589523 199885
rect 589457 199880 592572 199882
rect 589457 199824 589462 199880
rect 589518 199824 592572 199880
rect 589457 199822 592572 199824
rect 589457 199819 589523 199822
rect 575982 198930 576042 199172
rect 579521 198930 579587 198933
rect 575982 198928 579587 198930
rect 575982 198872 579526 198928
rect 579582 198872 579587 198928
rect 575982 198870 579587 198872
rect 579521 198867 579587 198870
rect 666645 198658 666711 198661
rect 675109 198658 675175 198661
rect 666645 198656 675175 198658
rect 666645 198600 666650 198656
rect 666706 198600 675114 198656
rect 675170 198600 675175 198656
rect 666645 198598 675175 198600
rect 666645 198595 666711 198598
rect 675109 198595 675175 198598
rect 666829 198386 666895 198389
rect 675385 198386 675451 198389
rect 666829 198384 675451 198386
rect 666829 198328 666834 198384
rect 666890 198328 675390 198384
rect 675446 198328 675451 198384
rect 666829 198326 675451 198328
rect 666829 198323 666895 198326
rect 675385 198323 675451 198326
rect 590377 198250 590443 198253
rect 590377 198248 592572 198250
rect 590377 198192 590382 198248
rect 590438 198192 592572 198248
rect 590377 198190 592572 198192
rect 590377 198187 590443 198190
rect 670785 197570 670851 197573
rect 675477 197570 675543 197573
rect 670785 197568 675543 197570
rect 670785 197512 670790 197568
rect 670846 197512 675482 197568
rect 675538 197512 675543 197568
rect 670785 197510 675543 197512
rect 670785 197507 670851 197510
rect 675477 197507 675543 197510
rect 42425 197298 42491 197301
rect 47117 197298 47183 197301
rect 42425 197296 47183 197298
rect 42425 197240 42430 197296
rect 42486 197240 47122 197296
rect 47178 197240 47183 197296
rect 42425 197238 47183 197240
rect 42425 197235 42491 197238
rect 47117 197235 47183 197238
rect 673545 197162 673611 197165
rect 675385 197162 675451 197165
rect 673545 197160 675451 197162
rect 673545 197104 673550 197160
rect 673606 197104 675390 197160
rect 675446 197104 675451 197160
rect 673545 197102 675451 197104
rect 673545 197099 673611 197102
rect 675385 197099 675451 197102
rect 48589 196482 48655 196485
rect 575982 196482 576042 196996
rect 589457 196618 589523 196621
rect 589457 196616 592572 196618
rect 589457 196560 589462 196616
rect 589518 196560 592572 196616
rect 589457 196558 592572 196560
rect 589457 196555 589523 196558
rect 578509 196482 578575 196485
rect 48589 196480 52164 196482
rect 48589 196424 48594 196480
rect 48650 196424 52164 196480
rect 48589 196422 52164 196424
rect 575982 196480 578575 196482
rect 575982 196424 578514 196480
rect 578570 196424 578575 196480
rect 575982 196422 578575 196424
rect 48589 196419 48655 196422
rect 578509 196419 578575 196422
rect 674281 196074 674347 196077
rect 675109 196074 675175 196077
rect 674281 196072 675175 196074
rect 674281 196016 674286 196072
rect 674342 196016 675114 196072
rect 675170 196016 675175 196072
rect 674281 196014 675175 196016
rect 674281 196011 674347 196014
rect 675109 196011 675175 196014
rect 41781 195804 41847 195805
rect 41781 195800 41828 195804
rect 41892 195802 41898 195804
rect 41781 195744 41786 195800
rect 41781 195740 41828 195744
rect 41892 195742 41938 195802
rect 41892 195740 41898 195742
rect 41781 195739 41847 195740
rect 673177 195258 673243 195261
rect 676806 195258 676812 195260
rect 673177 195256 676812 195258
rect 673177 195200 673182 195256
rect 673238 195200 676812 195256
rect 673177 195198 676812 195200
rect 673177 195195 673243 195198
rect 676806 195196 676812 195198
rect 676876 195196 676882 195260
rect 41965 195124 42031 195125
rect 41965 195120 42012 195124
rect 42076 195122 42082 195124
rect 41965 195064 41970 195120
rect 41965 195060 42012 195064
rect 42076 195062 42122 195122
rect 42076 195060 42082 195062
rect 41965 195059 42031 195060
rect 579521 194986 579587 194989
rect 575798 194984 579587 194986
rect 575798 194928 579526 194984
rect 579582 194928 579587 194984
rect 575798 194926 579587 194928
rect 575798 194820 575858 194926
rect 579521 194923 579587 194926
rect 589273 194986 589339 194989
rect 589273 194984 592572 194986
rect 589273 194928 589278 194984
rect 589334 194928 592572 194984
rect 589273 194926 592572 194928
rect 589273 194923 589339 194926
rect 675753 194578 675819 194581
rect 676622 194578 676628 194580
rect 675753 194576 676628 194578
rect 675753 194520 675758 194576
rect 675814 194520 676628 194576
rect 675753 194518 676628 194520
rect 675753 194515 675819 194518
rect 676622 194516 676628 194518
rect 676692 194516 676698 194580
rect 48313 194442 48379 194445
rect 48313 194440 52164 194442
rect 48313 194384 48318 194440
rect 48374 194384 52164 194440
rect 48313 194382 52164 194384
rect 48313 194379 48379 194382
rect 589457 193354 589523 193357
rect 589457 193352 592572 193354
rect 589457 193296 589462 193352
rect 589518 193296 592572 193352
rect 589457 193294 592572 193296
rect 589457 193291 589523 193294
rect 42425 193218 42491 193221
rect 44357 193218 44423 193221
rect 42425 193216 44423 193218
rect 42425 193160 42430 193216
rect 42486 193160 44362 193216
rect 44418 193160 44423 193216
rect 42425 193158 44423 193160
rect 42425 193155 42491 193158
rect 44357 193155 44423 193158
rect 675753 193218 675819 193221
rect 676070 193218 676076 193220
rect 675753 193216 676076 193218
rect 675753 193160 675758 193216
rect 675814 193160 676076 193216
rect 675753 193158 676076 193160
rect 675753 193155 675819 193158
rect 676070 193156 676076 193158
rect 676140 193156 676146 193220
rect 675661 192810 675727 192813
rect 675886 192810 675892 192812
rect 675661 192808 675892 192810
rect 675661 192752 675666 192808
rect 675722 192752 675892 192808
rect 675661 192750 675892 192752
rect 675661 192747 675727 192750
rect 675886 192748 675892 192750
rect 675956 192748 675962 192812
rect 49601 192402 49667 192405
rect 49601 192400 52164 192402
rect 49601 192344 49606 192400
rect 49662 192344 52164 192400
rect 49601 192342 52164 192344
rect 49601 192339 49667 192342
rect 575982 192266 576042 192644
rect 579521 192266 579587 192269
rect 575982 192264 579587 192266
rect 575982 192208 579526 192264
rect 579582 192208 579587 192264
rect 575982 192206 579587 192208
rect 579521 192203 579587 192206
rect 42333 191722 42399 191725
rect 44541 191722 44607 191725
rect 42333 191720 44607 191722
rect 42333 191664 42338 191720
rect 42394 191664 44546 191720
rect 44602 191664 44607 191720
rect 42333 191662 44607 191664
rect 42333 191659 42399 191662
rect 44541 191659 44607 191662
rect 589457 191722 589523 191725
rect 589457 191720 592572 191722
rect 589457 191664 589462 191720
rect 589518 191664 592572 191720
rect 589457 191662 592572 191664
rect 589457 191659 589523 191662
rect 40718 191524 40724 191588
rect 40788 191586 40794 191588
rect 41781 191586 41847 191589
rect 40788 191584 41847 191586
rect 40788 191528 41786 191584
rect 41842 191528 41847 191584
rect 40788 191526 41847 191528
rect 40788 191524 40794 191526
rect 41781 191523 41847 191526
rect 673361 191178 673427 191181
rect 675109 191178 675175 191181
rect 673361 191176 675175 191178
rect 673361 191120 673366 191176
rect 673422 191120 675114 191176
rect 675170 191120 675175 191176
rect 673361 191118 675175 191120
rect 673361 191115 673427 191118
rect 675109 191115 675175 191118
rect 579521 190770 579587 190773
rect 575798 190768 579587 190770
rect 575798 190712 579526 190768
rect 579582 190712 579587 190768
rect 575798 190710 579587 190712
rect 42425 190498 42491 190501
rect 43989 190498 44055 190501
rect 42425 190496 44055 190498
rect 42425 190440 42430 190496
rect 42486 190440 43994 190496
rect 44050 190440 44055 190496
rect 42425 190438 44055 190440
rect 42425 190435 42491 190438
rect 43989 190435 44055 190438
rect 47761 190498 47827 190501
rect 47761 190496 52164 190498
rect 47761 190440 47766 190496
rect 47822 190440 52164 190496
rect 575798 190468 575858 190710
rect 579521 190707 579587 190710
rect 47761 190438 52164 190440
rect 47761 190435 47827 190438
rect 590561 190090 590627 190093
rect 590561 190088 592572 190090
rect 590561 190032 590566 190088
rect 590622 190032 592572 190088
rect 590561 190030 592572 190032
rect 590561 190027 590627 190030
rect 42425 189954 42491 189957
rect 46933 189954 46999 189957
rect 42425 189952 46999 189954
rect 42425 189896 42430 189952
rect 42486 189896 46938 189952
rect 46994 189896 46999 189952
rect 42425 189894 46999 189896
rect 42425 189891 42491 189894
rect 46933 189891 46999 189894
rect 675334 189076 675340 189140
rect 675404 189138 675410 189140
rect 676121 189138 676187 189141
rect 675404 189136 676187 189138
rect 675404 189080 676126 189136
rect 676182 189080 676187 189136
rect 675404 189078 676187 189080
rect 675404 189076 675410 189078
rect 676121 189075 676187 189078
rect 589641 188458 589707 188461
rect 589641 188456 592572 188458
rect 589641 188400 589646 188456
rect 589702 188400 592572 188456
rect 589641 188398 592572 188400
rect 589641 188395 589707 188398
rect 575982 188050 576042 188292
rect 579521 188050 579587 188053
rect 575982 188048 579587 188050
rect 575982 187992 579526 188048
rect 579582 187992 579587 188048
rect 575982 187990 579587 187992
rect 579521 187987 579587 187990
rect 42425 187642 42491 187645
rect 44173 187642 44239 187645
rect 42425 187640 44239 187642
rect 42425 187584 42430 187640
rect 42486 187584 44178 187640
rect 44234 187584 44239 187640
rect 42425 187582 44239 187584
rect 42425 187579 42491 187582
rect 44173 187579 44239 187582
rect 40534 187172 40540 187236
rect 40604 187234 40610 187236
rect 41781 187234 41847 187237
rect 40604 187232 41847 187234
rect 40604 187176 41786 187232
rect 41842 187176 41847 187232
rect 40604 187174 41847 187176
rect 40604 187172 40610 187174
rect 41781 187171 41847 187174
rect 589457 186826 589523 186829
rect 589457 186824 592572 186826
rect 589457 186768 589462 186824
rect 589518 186768 592572 186824
rect 589457 186766 592572 186768
rect 589457 186763 589523 186766
rect 41454 186356 41460 186420
rect 41524 186418 41530 186420
rect 41781 186418 41847 186421
rect 41524 186416 41847 186418
rect 41524 186360 41786 186416
rect 41842 186360 41847 186416
rect 41524 186358 41847 186360
rect 41524 186356 41530 186358
rect 41781 186355 41847 186358
rect 579521 186282 579587 186285
rect 575798 186280 579587 186282
rect 575798 186224 579526 186280
rect 579582 186224 579587 186280
rect 575798 186222 579587 186224
rect 575798 186116 575858 186222
rect 579521 186219 579587 186222
rect 41781 186012 41847 186013
rect 41781 186008 41828 186012
rect 41892 186010 41898 186012
rect 41781 185952 41786 186008
rect 41781 185948 41828 185952
rect 41892 185950 41938 186010
rect 41892 185948 41898 185950
rect 41781 185947 41847 185948
rect 589457 185194 589523 185197
rect 589457 185192 592572 185194
rect 589457 185136 589462 185192
rect 589518 185136 592572 185192
rect 589457 185134 592572 185136
rect 589457 185131 589523 185134
rect 579521 184378 579587 184381
rect 575798 184376 579587 184378
rect 575798 184320 579526 184376
rect 579582 184320 579587 184376
rect 575798 184318 579587 184320
rect 575798 183940 575858 184318
rect 579521 184315 579587 184318
rect 589457 183562 589523 183565
rect 589457 183560 592572 183562
rect 589457 183504 589462 183560
rect 589518 183504 592572 183560
rect 589457 183502 592572 183504
rect 589457 183499 589523 183502
rect 672533 182066 672599 182069
rect 673126 182066 673132 182068
rect 672533 182064 673132 182066
rect 672533 182008 672538 182064
rect 672594 182008 673132 182064
rect 672533 182006 673132 182008
rect 672533 182003 672599 182006
rect 673126 182004 673132 182006
rect 673196 182004 673202 182068
rect 579521 181930 579587 181933
rect 575798 181928 579587 181930
rect 575798 181872 579526 181928
rect 579582 181872 579587 181928
rect 575798 181870 579587 181872
rect 575798 181764 575858 181870
rect 579521 181867 579587 181870
rect 590561 181930 590627 181933
rect 590561 181928 592572 181930
rect 590561 181872 590566 181928
rect 590622 181872 592572 181928
rect 590561 181870 592572 181872
rect 590561 181867 590627 181870
rect 589641 180298 589707 180301
rect 589641 180296 592572 180298
rect 589641 180240 589646 180296
rect 589702 180240 592572 180296
rect 589641 180238 592572 180240
rect 589641 180235 589707 180238
rect 673310 180236 673316 180300
rect 673380 180298 673386 180300
rect 675937 180298 676003 180301
rect 673380 180296 676003 180298
rect 673380 180240 675942 180296
rect 675998 180240 676003 180296
rect 673380 180238 676003 180240
rect 673380 180236 673386 180238
rect 675937 180235 676003 180238
rect 578785 180162 578851 180165
rect 575798 180160 578851 180162
rect 575798 180104 578790 180160
rect 578846 180104 578851 180160
rect 575798 180102 578851 180104
rect 575798 179588 575858 180102
rect 578785 180099 578851 180102
rect 42057 179346 42123 179349
rect 50705 179346 50771 179349
rect 42057 179344 50771 179346
rect 42057 179288 42062 179344
rect 42118 179288 50710 179344
rect 50766 179288 50771 179344
rect 42057 179286 50771 179288
rect 42057 179283 42123 179286
rect 50705 179283 50771 179286
rect 589457 178666 589523 178669
rect 589457 178664 592572 178666
rect 589457 178608 589462 178664
rect 589518 178608 592572 178664
rect 589457 178606 592572 178608
rect 589457 178603 589523 178606
rect 674097 178530 674163 178533
rect 674097 178528 676292 178530
rect 674097 178472 674102 178528
rect 674158 178472 676292 178528
rect 674097 178470 676292 178472
rect 674097 178467 674163 178470
rect 675937 178122 676003 178125
rect 675937 178120 676292 178122
rect 675937 178064 675942 178120
rect 675998 178064 676292 178120
rect 675937 178062 676292 178064
rect 675937 178059 676003 178062
rect 668025 177986 668091 177989
rect 666694 177984 668091 177986
rect 666694 177928 668030 177984
rect 668086 177928 668091 177984
rect 666694 177926 668091 177928
rect 666694 177918 666754 177926
rect 668025 177923 668091 177926
rect 666356 177858 666754 177918
rect 579521 177714 579587 177717
rect 575798 177712 579587 177714
rect 575798 177656 579526 177712
rect 579582 177656 579587 177712
rect 575798 177654 579587 177656
rect 575798 177412 575858 177654
rect 579521 177651 579587 177654
rect 672717 177714 672783 177717
rect 672717 177712 676292 177714
rect 672717 177656 672722 177712
rect 672778 177656 676292 177712
rect 672717 177654 676292 177656
rect 672717 177651 672783 177654
rect 673637 177306 673703 177309
rect 673637 177304 676292 177306
rect 673637 177248 673642 177304
rect 673698 177248 676292 177304
rect 673637 177246 676292 177248
rect 673637 177243 673703 177246
rect 589641 177034 589707 177037
rect 589641 177032 592572 177034
rect 589641 176976 589646 177032
rect 589702 176976 592572 177032
rect 589641 176974 592572 176976
rect 589641 176971 589707 176974
rect 673637 176898 673703 176901
rect 673637 176896 676292 176898
rect 673637 176840 673642 176896
rect 673698 176840 676292 176896
rect 673637 176838 676292 176840
rect 673637 176835 673703 176838
rect 676806 176608 676812 176672
rect 676876 176608 676882 176672
rect 676814 176460 676874 176608
rect 674649 176082 674715 176085
rect 674649 176080 676292 176082
rect 674649 176024 674654 176080
rect 674710 176024 676292 176080
rect 674649 176022 676292 176024
rect 674649 176019 674715 176022
rect 674465 175674 674531 175677
rect 674465 175672 676292 175674
rect 674465 175616 674470 175672
rect 674526 175616 676292 175672
rect 674465 175614 676292 175616
rect 674465 175611 674531 175614
rect 589457 175402 589523 175405
rect 589457 175400 592572 175402
rect 589457 175344 589462 175400
rect 589518 175344 592572 175400
rect 589457 175342 592572 175344
rect 589457 175339 589523 175342
rect 672533 175266 672599 175269
rect 672533 175264 676292 175266
rect 575982 175130 576042 175236
rect 672533 175208 672538 175264
rect 672594 175208 676292 175264
rect 672533 175206 676292 175208
rect 672533 175203 672599 175206
rect 578785 175130 578851 175133
rect 575982 175128 578851 175130
rect 575982 175072 578790 175128
rect 578846 175072 578851 175128
rect 575982 175070 578851 175072
rect 578785 175067 578851 175070
rect 667013 174994 667079 174997
rect 667013 174992 669330 174994
rect 667013 174936 667018 174992
rect 667074 174936 669330 174992
rect 667013 174934 669330 174936
rect 667013 174931 667079 174934
rect 669270 174858 669330 174934
rect 669270 174798 676292 174858
rect 668025 174722 668091 174725
rect 666694 174720 668091 174722
rect 666694 174664 668030 174720
rect 668086 174664 668091 174720
rect 666694 174662 668091 174664
rect 666694 174654 666754 174662
rect 668025 174659 668091 174662
rect 666356 174594 666754 174654
rect 673361 174450 673427 174453
rect 673361 174448 676292 174450
rect 673361 174392 673366 174448
rect 673422 174392 676292 174448
rect 673361 174390 676292 174392
rect 673361 174387 673427 174390
rect 674833 174042 674899 174045
rect 674833 174040 676292 174042
rect 674833 173984 674838 174040
rect 674894 173984 676292 174040
rect 674833 173982 676292 173984
rect 674833 173979 674899 173982
rect 589457 173770 589523 173773
rect 589457 173768 592572 173770
rect 589457 173712 589462 173768
rect 589518 173712 592572 173768
rect 589457 173710 592572 173712
rect 589457 173707 589523 173710
rect 678237 173634 678303 173637
rect 678237 173632 678316 173634
rect 678237 173576 678242 173632
rect 678298 173576 678316 173632
rect 678237 173574 678316 173576
rect 678237 173571 678303 173574
rect 578417 173498 578483 173501
rect 575798 173496 578483 173498
rect 575798 173440 578422 173496
rect 578478 173440 578483 173496
rect 575798 173438 578483 173440
rect 575798 173060 575858 173438
rect 578417 173435 578483 173438
rect 676029 173226 676095 173229
rect 676029 173224 676292 173226
rect 676029 173168 676034 173224
rect 676090 173168 676292 173224
rect 676029 173166 676292 173168
rect 676029 173163 676095 173166
rect 667933 173090 667999 173093
rect 666694 173088 667999 173090
rect 666694 173032 667938 173088
rect 667994 173032 667999 173088
rect 666694 173030 667999 173032
rect 666694 173022 666754 173030
rect 667933 173027 667999 173030
rect 666356 172962 666754 173022
rect 675886 172756 675892 172820
rect 675956 172818 675962 172820
rect 675956 172758 676292 172818
rect 675956 172756 675962 172758
rect 669589 172410 669655 172413
rect 669589 172408 676292 172410
rect 669589 172352 669594 172408
rect 669650 172352 676292 172408
rect 669589 172350 676292 172352
rect 669589 172347 669655 172350
rect 589457 172138 589523 172141
rect 589457 172136 592572 172138
rect 589457 172080 589462 172136
rect 589518 172080 592572 172136
rect 589457 172078 592572 172080
rect 589457 172075 589523 172078
rect 674557 172002 674623 172005
rect 674557 172000 676292 172002
rect 674557 171944 674562 172000
rect 674618 171944 676292 172000
rect 674557 171942 676292 171944
rect 674557 171939 674623 171942
rect 679617 171594 679683 171597
rect 679604 171592 679683 171594
rect 679604 171536 679622 171592
rect 679678 171536 679683 171592
rect 679604 171534 679683 171536
rect 679617 171531 679683 171534
rect 670969 171186 671035 171189
rect 670969 171184 676292 171186
rect 670969 171128 670974 171184
rect 671030 171128 676292 171184
rect 670969 171126 676292 171128
rect 670969 171123 671035 171126
rect 578233 171050 578299 171053
rect 575798 171048 578299 171050
rect 575798 170992 578238 171048
rect 578294 170992 578299 171048
rect 575798 170990 578299 170992
rect 575798 170884 575858 170990
rect 578233 170987 578299 170990
rect 669446 170988 669452 171052
rect 669516 171050 669522 171052
rect 670601 171050 670667 171053
rect 669516 171048 670667 171050
rect 669516 170992 670606 171048
rect 670662 170992 670667 171048
rect 669516 170990 670667 170992
rect 669516 170988 669522 170990
rect 670601 170987 670667 170990
rect 670325 170778 670391 170781
rect 670325 170776 676292 170778
rect 670325 170720 670330 170776
rect 670386 170720 676292 170776
rect 670325 170718 676292 170720
rect 670325 170715 670391 170718
rect 589641 170506 589707 170509
rect 589641 170504 592572 170506
rect 589641 170448 589646 170504
rect 589702 170448 592572 170504
rect 589641 170446 592572 170448
rect 589641 170443 589707 170446
rect 675886 170308 675892 170372
rect 675956 170370 675962 170372
rect 675956 170310 676292 170370
rect 675956 170308 675962 170310
rect 670417 169962 670483 169965
rect 670417 169960 676292 169962
rect 670417 169904 670422 169960
rect 670478 169904 676292 169960
rect 670417 169902 676292 169904
rect 670417 169899 670483 169902
rect 666356 169698 666754 169758
rect 666694 169690 666754 169698
rect 668209 169690 668275 169693
rect 666694 169688 668275 169690
rect 666694 169632 668214 169688
rect 668270 169632 668275 169688
rect 666694 169630 668275 169632
rect 668209 169627 668275 169630
rect 672993 169554 673059 169557
rect 672993 169552 676292 169554
rect 672993 169496 672998 169552
rect 673054 169496 676292 169552
rect 672993 169494 676292 169496
rect 672993 169491 673059 169494
rect 578693 169282 578759 169285
rect 575798 169280 578759 169282
rect 575798 169224 578698 169280
rect 578754 169224 578759 169280
rect 575798 169222 578759 169224
rect 575798 168708 575858 169222
rect 578693 169219 578759 169222
rect 674373 169146 674439 169149
rect 674373 169144 676292 169146
rect 674373 169088 674378 169144
rect 674434 169088 676292 169144
rect 674373 169086 676292 169088
rect 674373 169083 674439 169086
rect 589457 168874 589523 168877
rect 589457 168872 592572 168874
rect 589457 168816 589462 168872
rect 589518 168816 592572 168872
rect 589457 168814 592572 168816
rect 589457 168811 589523 168814
rect 673177 168738 673243 168741
rect 673177 168736 676292 168738
rect 673177 168680 673182 168736
rect 673238 168680 676292 168736
rect 673177 168678 676292 168680
rect 673177 168675 673243 168678
rect 672717 168330 672783 168333
rect 672717 168328 676292 168330
rect 672717 168272 672722 168328
rect 672778 168272 676292 168328
rect 672717 168270 676292 168272
rect 672717 168267 672783 168270
rect 668209 168194 668275 168197
rect 666694 168192 668275 168194
rect 666694 168136 668214 168192
rect 668270 168136 668275 168192
rect 666694 168134 668275 168136
rect 666694 168126 666754 168134
rect 668209 168131 668275 168134
rect 666356 168066 666754 168126
rect 676029 167922 676095 167925
rect 676029 167920 676292 167922
rect 676029 167864 676034 167920
rect 676090 167864 676292 167920
rect 676029 167862 676292 167864
rect 676029 167859 676095 167862
rect 675334 167452 675340 167516
rect 675404 167514 675410 167516
rect 675661 167514 675727 167517
rect 675404 167512 676292 167514
rect 675404 167456 675666 167512
rect 675722 167456 676292 167512
rect 675404 167454 676292 167456
rect 675404 167452 675410 167454
rect 675661 167451 675727 167454
rect 589457 167242 589523 167245
rect 589457 167240 592572 167242
rect 589457 167184 589462 167240
rect 589518 167184 592572 167240
rect 589457 167182 592572 167184
rect 589457 167179 589523 167182
rect 676170 167046 676292 167106
rect 578233 166970 578299 166973
rect 575798 166968 578299 166970
rect 575798 166912 578238 166968
rect 578294 166912 578299 166968
rect 575798 166910 578299 166912
rect 575798 166532 575858 166910
rect 578233 166907 578299 166910
rect 674097 166970 674163 166973
rect 676170 166970 676230 167046
rect 674097 166968 676230 166970
rect 674097 166912 674102 166968
rect 674158 166912 676230 166968
rect 674097 166910 676230 166912
rect 674097 166907 674163 166910
rect 589457 165610 589523 165613
rect 674281 165610 674347 165613
rect 676029 165610 676095 165613
rect 589457 165608 592572 165610
rect 589457 165552 589462 165608
rect 589518 165552 592572 165608
rect 589457 165550 592572 165552
rect 674281 165608 676095 165610
rect 674281 165552 674286 165608
rect 674342 165552 676034 165608
rect 676090 165552 676095 165608
rect 674281 165550 676095 165552
rect 589457 165547 589523 165550
rect 674281 165547 674347 165550
rect 676029 165547 676095 165550
rect 667933 164930 667999 164933
rect 666694 164928 667999 164930
rect 666694 164872 667938 164928
rect 667994 164872 667999 164928
rect 666694 164870 667999 164872
rect 666694 164862 666754 164870
rect 667933 164867 667999 164870
rect 666356 164802 666754 164862
rect 579521 164522 579587 164525
rect 575798 164520 579587 164522
rect 575798 164464 579526 164520
rect 579582 164464 579587 164520
rect 575798 164462 579587 164464
rect 575798 164356 575858 164462
rect 579521 164459 579587 164462
rect 589457 163978 589523 163981
rect 589457 163976 592572 163978
rect 589457 163920 589462 163976
rect 589518 163920 592572 163976
rect 589457 163918 592572 163920
rect 589457 163915 589523 163918
rect 668393 163298 668459 163301
rect 666694 163296 668459 163298
rect 666694 163240 668398 163296
rect 668454 163240 668459 163296
rect 666694 163238 668459 163240
rect 666694 163230 666754 163238
rect 668393 163235 668459 163238
rect 666356 163170 666754 163230
rect 579337 162754 579403 162757
rect 575798 162752 579403 162754
rect 575798 162696 579342 162752
rect 579398 162696 579403 162752
rect 575798 162694 579403 162696
rect 575798 162180 575858 162694
rect 579337 162691 579403 162694
rect 589457 162346 589523 162349
rect 589457 162344 592572 162346
rect 589457 162288 589462 162344
rect 589518 162288 592572 162344
rect 589457 162286 592572 162288
rect 589457 162283 589523 162286
rect 676070 162148 676076 162212
rect 676140 162210 676146 162212
rect 678237 162210 678303 162213
rect 676140 162208 678303 162210
rect 676140 162152 678242 162208
rect 678298 162152 678303 162208
rect 676140 162150 678303 162152
rect 676140 162148 676146 162150
rect 678237 162147 678303 162150
rect 675937 161396 676003 161397
rect 675886 161394 675892 161396
rect 675846 161334 675892 161394
rect 675956 161392 676003 161396
rect 675998 161336 676003 161392
rect 675886 161332 675892 161334
rect 675956 161332 676003 161336
rect 675937 161331 676003 161332
rect 673126 161060 673132 161124
rect 673196 161122 673202 161124
rect 675385 161122 675451 161125
rect 673196 161120 675451 161122
rect 673196 161064 675390 161120
rect 675446 161064 675451 161120
rect 673196 161062 675451 161064
rect 673196 161060 673202 161062
rect 675385 161059 675451 161062
rect 589457 160714 589523 160717
rect 589457 160712 592572 160714
rect 589457 160656 589462 160712
rect 589518 160656 592572 160712
rect 589457 160654 592572 160656
rect 589457 160651 589523 160654
rect 668393 160442 668459 160445
rect 673821 160442 673887 160445
rect 668393 160440 673887 160442
rect 668393 160384 668398 160440
rect 668454 160384 673826 160440
rect 673882 160384 673887 160440
rect 668393 160382 673887 160384
rect 668393 160379 668459 160382
rect 673821 160379 673887 160382
rect 669313 160034 669379 160037
rect 666694 160032 669379 160034
rect 575982 159898 576042 160004
rect 666694 159976 669318 160032
rect 669374 159976 669379 160032
rect 666694 159974 669379 159976
rect 666694 159966 666754 159974
rect 669313 159971 669379 159974
rect 675661 160034 675727 160037
rect 675886 160034 675892 160036
rect 675661 160032 675892 160034
rect 675661 159976 675666 160032
rect 675722 159976 675892 160032
rect 675661 159974 675892 159976
rect 675661 159971 675727 159974
rect 675886 159972 675892 159974
rect 675956 159972 675962 160036
rect 666356 159906 666754 159966
rect 578233 159898 578299 159901
rect 575982 159896 578299 159898
rect 575982 159840 578238 159896
rect 578294 159840 578299 159896
rect 575982 159838 578299 159840
rect 578233 159835 578299 159838
rect 589457 159082 589523 159085
rect 589457 159080 592572 159082
rect 589457 159024 589462 159080
rect 589518 159024 592572 159080
rect 589457 159022 592572 159024
rect 589457 159019 589523 159022
rect 578417 158402 578483 158405
rect 668393 158402 668459 158405
rect 575798 158400 578483 158402
rect 575798 158344 578422 158400
rect 578478 158344 578483 158400
rect 575798 158342 578483 158344
rect 575798 157828 575858 158342
rect 578417 158339 578483 158342
rect 666694 158400 668459 158402
rect 666694 158344 668398 158400
rect 668454 158344 668459 158400
rect 666694 158342 668459 158344
rect 666694 158334 666754 158342
rect 668393 158339 668459 158342
rect 666356 158274 666754 158334
rect 674373 157588 674439 157589
rect 674373 157584 674420 157588
rect 674484 157586 674490 157588
rect 674741 157586 674807 157589
rect 674373 157528 674378 157584
rect 674373 157524 674420 157528
rect 674484 157526 674530 157586
rect 674741 157584 674850 157586
rect 674741 157528 674746 157584
rect 674802 157528 674850 157584
rect 674484 157524 674490 157526
rect 674373 157523 674439 157524
rect 674741 157523 674850 157528
rect 589273 157450 589339 157453
rect 589273 157448 592572 157450
rect 589273 157392 589278 157448
rect 589334 157392 592572 157448
rect 589273 157390 592572 157392
rect 589273 157387 589339 157390
rect 674790 157181 674850 157523
rect 674741 157176 674850 157181
rect 674741 157120 674746 157176
rect 674802 157120 674850 157176
rect 674741 157118 674850 157120
rect 674741 157115 674807 157118
rect 675753 157042 675819 157045
rect 676438 157042 676444 157044
rect 675753 157040 676444 157042
rect 675753 156984 675758 157040
rect 675814 156984 676444 157040
rect 675753 156982 676444 156984
rect 675753 156979 675819 156982
rect 676438 156980 676444 156982
rect 676508 156980 676514 157044
rect 578877 155954 578943 155957
rect 575798 155952 578943 155954
rect 575798 155896 578882 155952
rect 578938 155896 578943 155952
rect 575798 155894 578943 155896
rect 575798 155652 575858 155894
rect 578877 155891 578943 155894
rect 589457 155818 589523 155821
rect 589457 155816 592572 155818
rect 589457 155760 589462 155816
rect 589518 155760 592572 155816
rect 589457 155758 592572 155760
rect 589457 155755 589523 155758
rect 672993 155546 673059 155549
rect 675109 155546 675175 155549
rect 672993 155544 675175 155546
rect 672993 155488 672998 155544
rect 673054 155488 675114 155544
rect 675170 155488 675175 155544
rect 672993 155486 675175 155488
rect 672993 155483 673059 155486
rect 675109 155483 675175 155486
rect 671153 155410 671219 155413
rect 666878 155408 671219 155410
rect 666878 155352 671158 155408
rect 671214 155352 671219 155408
rect 666878 155350 671219 155352
rect 666878 155070 666938 155350
rect 671153 155347 671219 155350
rect 670417 155138 670483 155141
rect 675017 155138 675083 155141
rect 670417 155136 675083 155138
rect 670417 155080 670422 155136
rect 670478 155080 675022 155136
rect 675078 155080 675083 155136
rect 670417 155078 675083 155080
rect 670417 155075 670483 155078
rect 675017 155075 675083 155078
rect 666356 155010 666938 155070
rect 674465 154868 674531 154869
rect 674414 154804 674420 154868
rect 674484 154866 674531 154868
rect 674484 154864 674576 154866
rect 674526 154808 674576 154864
rect 674484 154806 674576 154808
rect 674484 154804 674531 154806
rect 674465 154803 674531 154804
rect 670785 154458 670851 154461
rect 675017 154458 675083 154461
rect 670785 154456 675083 154458
rect 670785 154400 670790 154456
rect 670846 154400 675022 154456
rect 675078 154400 675083 154456
rect 670785 154398 675083 154400
rect 670785 154395 670851 154398
rect 675017 154395 675083 154398
rect 589457 154186 589523 154189
rect 589457 154184 592572 154186
rect 589457 154128 589462 154184
rect 589518 154128 592572 154184
rect 589457 154126 592572 154128
rect 589457 154123 589523 154126
rect 578325 153642 578391 153645
rect 575798 153640 578391 153642
rect 575798 153584 578330 153640
rect 578386 153584 578391 153640
rect 575798 153582 578391 153584
rect 575798 153476 575858 153582
rect 578325 153579 578391 153582
rect 666356 153378 666938 153438
rect 666878 153370 666938 153378
rect 666878 153310 673470 153370
rect 673410 153234 673470 153310
rect 674230 153234 674236 153236
rect 673410 153174 674236 153234
rect 674230 153172 674236 153174
rect 674300 153172 674306 153236
rect 674465 152690 674531 152693
rect 675109 152690 675175 152693
rect 674465 152688 675175 152690
rect 674465 152632 674470 152688
rect 674526 152632 675114 152688
rect 675170 152632 675175 152688
rect 674465 152630 675175 152632
rect 674465 152627 674531 152630
rect 675109 152627 675175 152630
rect 589457 152554 589523 152557
rect 589457 152552 592572 152554
rect 589457 152496 589462 152552
rect 589518 152496 592572 152552
rect 589457 152494 592572 152496
rect 589457 152491 589523 152494
rect 578233 151738 578299 151741
rect 575798 151736 578299 151738
rect 575798 151680 578238 151736
rect 578294 151680 578299 151736
rect 575798 151678 578299 151680
rect 575798 151300 575858 151678
rect 578233 151675 578299 151678
rect 670601 151738 670667 151741
rect 675109 151738 675175 151741
rect 670601 151736 675175 151738
rect 670601 151680 670606 151736
rect 670662 151680 675114 151736
rect 675170 151680 675175 151736
rect 670601 151678 675175 151680
rect 670601 151675 670667 151678
rect 675109 151675 675175 151678
rect 673177 151058 673243 151061
rect 675109 151058 675175 151061
rect 673177 151056 675175 151058
rect 673177 151000 673182 151056
rect 673238 151000 675114 151056
rect 675170 151000 675175 151056
rect 673177 150998 675175 151000
rect 673177 150995 673243 150998
rect 675109 150995 675175 150998
rect 590009 150922 590075 150925
rect 590009 150920 592572 150922
rect 590009 150864 590014 150920
rect 590070 150864 592572 150920
rect 590009 150862 592572 150864
rect 590009 150859 590075 150862
rect 669589 150378 669655 150381
rect 674925 150378 674991 150381
rect 669589 150376 674991 150378
rect 669589 150320 669594 150376
rect 669650 150320 674930 150376
rect 674986 150320 674991 150376
rect 669589 150318 674991 150320
rect 669589 150315 669655 150318
rect 674925 150315 674991 150318
rect 675753 150378 675819 150381
rect 676254 150378 676260 150380
rect 675753 150376 676260 150378
rect 675753 150320 675758 150376
rect 675814 150320 676260 150376
rect 675753 150318 676260 150320
rect 675753 150315 675819 150318
rect 676254 150316 676260 150318
rect 676324 150316 676330 150380
rect 669129 150242 669195 150245
rect 666694 150240 669195 150242
rect 666694 150184 669134 150240
rect 669190 150184 669195 150240
rect 666694 150182 669195 150184
rect 666694 150174 666754 150182
rect 669129 150179 669195 150182
rect 666356 150114 666754 150174
rect 578877 149698 578943 149701
rect 575798 149696 578943 149698
rect 575798 149640 578882 149696
rect 578938 149640 578943 149696
rect 575798 149638 578943 149640
rect 575798 149124 575858 149638
rect 578877 149635 578943 149638
rect 589457 149290 589523 149293
rect 589457 149288 592572 149290
rect 589457 149232 589462 149288
rect 589518 149232 592572 149288
rect 589457 149230 592572 149232
rect 589457 149227 589523 149230
rect 670785 149154 670851 149157
rect 671521 149154 671587 149157
rect 670785 149152 671587 149154
rect 670785 149096 670790 149152
rect 670846 149096 671526 149152
rect 671582 149096 671587 149152
rect 670785 149094 671587 149096
rect 670785 149091 670851 149094
rect 671521 149091 671587 149094
rect 668945 148610 669011 148613
rect 666694 148608 669011 148610
rect 666694 148552 668950 148608
rect 669006 148552 669011 148608
rect 666694 148550 669011 148552
rect 666694 148542 666754 148550
rect 668945 148547 669011 148550
rect 666356 148482 666754 148542
rect 675753 148474 675819 148477
rect 676070 148474 676076 148476
rect 675753 148472 676076 148474
rect 675753 148416 675758 148472
rect 675814 148416 676076 148472
rect 675753 148414 676076 148416
rect 675753 148411 675819 148414
rect 676070 148412 676076 148414
rect 676140 148412 676146 148476
rect 588537 147658 588603 147661
rect 675385 147660 675451 147661
rect 675334 147658 675340 147660
rect 588537 147656 592572 147658
rect 588537 147600 588542 147656
rect 588598 147600 592572 147656
rect 588537 147598 592572 147600
rect 675294 147598 675340 147658
rect 675404 147656 675451 147660
rect 675446 147600 675451 147656
rect 588537 147595 588603 147598
rect 675334 147596 675340 147598
rect 675404 147596 675451 147600
rect 675385 147595 675451 147596
rect 579521 147522 579587 147525
rect 575798 147520 579587 147522
rect 575798 147464 579526 147520
rect 579582 147464 579587 147520
rect 575798 147462 579587 147464
rect 575798 146948 575858 147462
rect 579521 147459 579587 147462
rect 589457 146026 589523 146029
rect 589457 146024 592572 146026
rect 589457 145968 589462 146024
rect 589518 145968 592572 146024
rect 589457 145966 592572 145968
rect 589457 145963 589523 145966
rect 671889 145346 671955 145349
rect 666694 145344 671955 145346
rect 666694 145288 671894 145344
rect 671950 145288 671955 145344
rect 666694 145286 671955 145288
rect 666694 145278 666754 145286
rect 671889 145283 671955 145286
rect 666356 145218 666754 145278
rect 575982 144666 576042 144772
rect 579245 144666 579311 144669
rect 575982 144664 579311 144666
rect 575982 144608 579250 144664
rect 579306 144608 579311 144664
rect 575982 144606 579311 144608
rect 579245 144603 579311 144606
rect 589457 144394 589523 144397
rect 589457 144392 592572 144394
rect 589457 144336 589462 144392
rect 589518 144336 592572 144392
rect 589457 144334 592572 144336
rect 589457 144331 589523 144334
rect 668577 143714 668643 143717
rect 666694 143712 668643 143714
rect 666694 143656 668582 143712
rect 668638 143656 668643 143712
rect 666694 143654 668643 143656
rect 666694 143646 666754 143654
rect 668577 143651 668643 143654
rect 666356 143586 666754 143646
rect 579521 143034 579587 143037
rect 575798 143032 579587 143034
rect 575798 142976 579526 143032
rect 579582 142976 579587 143032
rect 575798 142974 579587 142976
rect 575798 142596 575858 142974
rect 579521 142971 579587 142974
rect 589825 142762 589891 142765
rect 589825 142760 592572 142762
rect 589825 142704 589830 142760
rect 589886 142704 592572 142760
rect 589825 142702 592572 142704
rect 589825 142699 589891 142702
rect 589457 141130 589523 141133
rect 589457 141128 592572 141130
rect 589457 141072 589462 141128
rect 589518 141072 592572 141128
rect 589457 141070 592572 141072
rect 589457 141067 589523 141070
rect 578601 140586 578667 140589
rect 575798 140584 578667 140586
rect 575798 140528 578606 140584
rect 578662 140528 578667 140584
rect 575798 140526 578667 140528
rect 575798 140420 575858 140526
rect 578601 140523 578667 140526
rect 668209 140450 668275 140453
rect 666694 140448 668275 140450
rect 666694 140392 668214 140448
rect 668270 140392 668275 140448
rect 666694 140390 668275 140392
rect 666694 140382 666754 140390
rect 668209 140387 668275 140390
rect 666356 140322 666754 140382
rect 589457 139498 589523 139501
rect 589457 139496 592572 139498
rect 589457 139440 589462 139496
rect 589518 139440 592572 139496
rect 589457 139438 592572 139440
rect 589457 139435 589523 139438
rect 578601 138818 578667 138821
rect 668393 138818 668459 138821
rect 575798 138816 578667 138818
rect 575798 138760 578606 138816
rect 578662 138760 578667 138816
rect 575798 138758 578667 138760
rect 575798 138244 575858 138758
rect 578601 138755 578667 138758
rect 666694 138816 668459 138818
rect 666694 138760 668398 138816
rect 668454 138760 668459 138816
rect 666694 138758 668459 138760
rect 666694 138750 666754 138758
rect 668393 138755 668459 138758
rect 666356 138690 666754 138750
rect 589457 137866 589523 137869
rect 589457 137864 592572 137866
rect 589457 137808 589462 137864
rect 589518 137808 592572 137864
rect 589457 137806 592572 137808
rect 589457 137803 589523 137806
rect 578877 136642 578943 136645
rect 575798 136640 578943 136642
rect 575798 136584 578882 136640
rect 578938 136584 578943 136640
rect 575798 136582 578943 136584
rect 575798 136068 575858 136582
rect 578877 136579 578943 136582
rect 589457 136234 589523 136237
rect 589457 136232 592572 136234
rect 589457 136176 589462 136232
rect 589518 136176 592572 136232
rect 589457 136174 592572 136176
rect 589457 136171 589523 136174
rect 669446 135554 669452 135556
rect 666694 135494 669452 135554
rect 666694 135486 666754 135494
rect 669446 135492 669452 135494
rect 669516 135492 669522 135556
rect 666356 135426 666754 135486
rect 590377 134602 590443 134605
rect 667749 134602 667815 134605
rect 674833 134602 674899 134605
rect 590377 134600 592572 134602
rect 590377 134544 590382 134600
rect 590438 134544 592572 134600
rect 590377 134542 592572 134544
rect 667749 134600 674899 134602
rect 667749 134544 667754 134600
rect 667810 134544 674838 134600
rect 674894 134544 674899 134600
rect 667749 134542 674899 134544
rect 590377 134539 590443 134542
rect 667749 134539 667815 134542
rect 674833 134539 674899 134542
rect 579521 134466 579587 134469
rect 575798 134464 579587 134466
rect 575798 134408 579526 134464
rect 579582 134408 579587 134464
rect 575798 134406 579587 134408
rect 575798 133892 575858 134406
rect 579521 134403 579587 134406
rect 674833 133922 674899 133925
rect 674833 133920 676322 133922
rect 674833 133864 674838 133920
rect 674894 133864 676322 133920
rect 674833 133862 676322 133864
rect 674833 133859 674899 133862
rect 666356 133794 666754 133854
rect 666694 133786 666754 133794
rect 668761 133786 668827 133789
rect 666694 133784 668827 133786
rect 666694 133728 668766 133784
rect 668822 133728 668827 133784
rect 666694 133726 668827 133728
rect 668761 133723 668827 133726
rect 676262 133348 676322 133862
rect 667565 133106 667631 133109
rect 676489 133106 676555 133109
rect 667565 133104 676555 133106
rect 667565 133048 667570 133104
rect 667626 133048 676494 133104
rect 676550 133048 676555 133104
rect 667565 133046 676555 133048
rect 667565 133043 667631 133046
rect 676489 133043 676555 133046
rect 589457 132970 589523 132973
rect 589457 132968 592572 132970
rect 589457 132912 589462 132968
rect 589518 132912 592572 132968
rect 589457 132910 592572 132912
rect 589457 132907 589523 132910
rect 667381 132698 667447 132701
rect 676262 132698 676322 132940
rect 676489 132698 676555 132701
rect 667381 132696 676322 132698
rect 667381 132640 667386 132696
rect 667442 132640 676322 132696
rect 667381 132638 676322 132640
rect 676446 132696 676555 132698
rect 676446 132640 676494 132696
rect 676550 132640 676555 132696
rect 667381 132635 667447 132638
rect 676446 132635 676555 132640
rect 676446 132532 676506 132635
rect 579061 132290 579127 132293
rect 575798 132288 579127 132290
rect 575798 132232 579066 132288
rect 579122 132232 579127 132288
rect 575798 132230 579127 132232
rect 575798 131716 575858 132230
rect 579061 132227 579127 132230
rect 673637 132154 673703 132157
rect 673637 132152 676292 132154
rect 673637 132096 673642 132152
rect 673698 132096 676292 132152
rect 673637 132094 676292 132096
rect 673637 132091 673703 132094
rect 671337 131746 671403 131749
rect 671337 131744 676292 131746
rect 671337 131688 671342 131744
rect 671398 131688 676292 131744
rect 671337 131686 676292 131688
rect 671337 131683 671403 131686
rect 589457 131338 589523 131341
rect 674649 131338 674715 131341
rect 589457 131336 592572 131338
rect 589457 131280 589462 131336
rect 589518 131280 592572 131336
rect 589457 131278 592572 131280
rect 674649 131336 676292 131338
rect 674649 131280 674654 131336
rect 674710 131280 676292 131336
rect 674649 131278 676292 131280
rect 589457 131275 589523 131278
rect 674649 131275 674715 131278
rect 670141 130930 670207 130933
rect 670141 130928 676292 130930
rect 670141 130872 670146 130928
rect 670202 130872 676292 130928
rect 670141 130870 676292 130872
rect 670141 130867 670207 130870
rect 667933 130658 667999 130661
rect 666694 130656 667999 130658
rect 666694 130600 667938 130656
rect 667994 130600 667999 130656
rect 666694 130598 667999 130600
rect 666694 130590 666754 130598
rect 667933 130595 667999 130598
rect 666356 130530 666754 130590
rect 672533 130522 672599 130525
rect 672533 130520 676292 130522
rect 672533 130464 672538 130520
rect 672594 130464 676292 130520
rect 672533 130462 676292 130464
rect 672533 130459 672599 130462
rect 676213 130250 676279 130253
rect 676213 130248 676322 130250
rect 676213 130192 676218 130248
rect 676274 130192 676322 130248
rect 676213 130187 676322 130192
rect 676262 130084 676322 130187
rect 578877 129706 578943 129709
rect 575798 129704 578943 129706
rect 575798 129648 578882 129704
rect 578938 129648 578943 129704
rect 575798 129646 578943 129648
rect 575798 129540 575858 129646
rect 578877 129643 578943 129646
rect 588721 129706 588787 129709
rect 673361 129706 673427 129709
rect 588721 129704 592572 129706
rect 588721 129648 588726 129704
rect 588782 129648 592572 129704
rect 588721 129646 592572 129648
rect 673361 129704 676292 129706
rect 673361 129648 673366 129704
rect 673422 129648 676292 129704
rect 673361 129646 676292 129648
rect 588721 129643 588787 129646
rect 673361 129643 673427 129646
rect 671521 129298 671587 129301
rect 671521 129296 676292 129298
rect 671521 129240 671526 129296
rect 671582 129240 676292 129296
rect 671521 129238 676292 129240
rect 671521 129235 671587 129238
rect 668577 129026 668643 129029
rect 666694 129024 668643 129026
rect 666694 128968 668582 129024
rect 668638 128968 668643 129024
rect 666694 128966 668643 128968
rect 666694 128958 666754 128966
rect 668577 128963 668643 128966
rect 666356 128898 666754 128958
rect 675845 128890 675911 128893
rect 675845 128888 676292 128890
rect 675845 128832 675850 128888
rect 675906 128832 676292 128888
rect 675845 128830 676292 128832
rect 675845 128827 675911 128830
rect 674974 128422 676292 128482
rect 673913 128346 673979 128349
rect 674974 128346 675034 128422
rect 673913 128344 675034 128346
rect 673913 128288 673918 128344
rect 673974 128288 675034 128344
rect 673913 128286 675034 128288
rect 673913 128283 673979 128286
rect 589457 128074 589523 128077
rect 589457 128072 592572 128074
rect 589457 128016 589462 128072
rect 589518 128016 592572 128072
rect 589457 128014 592572 128016
rect 589457 128011 589523 128014
rect 579521 127938 579587 127941
rect 575798 127936 579587 127938
rect 575798 127880 579526 127936
rect 579582 127880 579587 127936
rect 575798 127878 579587 127880
rect 575798 127364 575858 127878
rect 579521 127875 579587 127878
rect 676446 127805 676506 128044
rect 668577 127802 668643 127805
rect 676213 127802 676279 127805
rect 668577 127800 676279 127802
rect 668577 127744 668582 127800
rect 668638 127744 676218 127800
rect 676274 127744 676279 127800
rect 668577 127742 676279 127744
rect 668577 127739 668643 127742
rect 676213 127739 676279 127742
rect 676397 127800 676506 127805
rect 676397 127744 676402 127800
rect 676458 127744 676506 127800
rect 676397 127742 676506 127744
rect 676397 127739 676463 127742
rect 676262 127396 676322 127636
rect 676254 127332 676260 127396
rect 676324 127332 676330 127396
rect 668945 126986 669011 126989
rect 672257 126986 672323 126989
rect 668945 126984 672323 126986
rect 668945 126928 668950 126984
rect 669006 126928 672262 126984
rect 672318 126928 672323 126984
rect 668945 126926 672323 126928
rect 668945 126923 669011 126926
rect 672257 126923 672323 126926
rect 676070 126924 676076 126988
rect 676140 126986 676146 126988
rect 676262 126986 676322 127228
rect 676140 126926 676322 126986
rect 676140 126924 676146 126926
rect 673361 126578 673427 126581
rect 676262 126578 676322 126820
rect 673361 126576 676322 126578
rect 673361 126520 673366 126576
rect 673422 126520 676322 126576
rect 673361 126518 676322 126520
rect 673361 126515 673427 126518
rect 590101 126442 590167 126445
rect 590101 126440 592572 126442
rect 590101 126384 590106 126440
rect 590162 126384 592572 126440
rect 590101 126382 592572 126384
rect 590101 126379 590167 126382
rect 678286 126173 678346 126412
rect 678237 126168 678346 126173
rect 678237 126112 678242 126168
rect 678298 126112 678346 126168
rect 678237 126110 678346 126112
rect 678237 126107 678303 126110
rect 668761 125762 668827 125765
rect 676630 125764 676690 126004
rect 666694 125760 668827 125762
rect 666694 125704 668766 125760
rect 668822 125704 668827 125760
rect 666694 125702 668827 125704
rect 666694 125694 666754 125702
rect 668761 125699 668827 125702
rect 676622 125700 676628 125764
rect 676692 125700 676698 125764
rect 666356 125634 666754 125694
rect 682334 125357 682394 125596
rect 578325 125354 578391 125357
rect 575798 125352 578391 125354
rect 575798 125296 578330 125352
rect 578386 125296 578391 125352
rect 575798 125294 578391 125296
rect 682334 125352 682443 125357
rect 682334 125296 682382 125352
rect 682438 125296 682443 125352
rect 682334 125294 682443 125296
rect 575798 125188 575858 125294
rect 578325 125291 578391 125294
rect 682377 125291 682443 125294
rect 674649 125218 674715 125221
rect 674649 125216 676292 125218
rect 674649 125160 674654 125216
rect 674710 125160 676292 125216
rect 674649 125158 676292 125160
rect 674649 125155 674715 125158
rect 590561 124810 590627 124813
rect 673177 124810 673243 124813
rect 590561 124808 592572 124810
rect 590561 124752 590566 124808
rect 590622 124752 592572 124808
rect 590561 124750 592572 124752
rect 673177 124808 676292 124810
rect 673177 124752 673182 124808
rect 673238 124752 676292 124808
rect 673177 124750 676292 124752
rect 590561 124747 590627 124750
rect 673177 124747 673243 124750
rect 672073 124130 672139 124133
rect 676446 124132 676506 124372
rect 666694 124128 672139 124130
rect 666694 124072 672078 124128
rect 672134 124072 672139 124128
rect 666694 124070 672139 124072
rect 666694 124062 666754 124070
rect 672073 124067 672139 124070
rect 676438 124068 676444 124132
rect 676508 124068 676514 124132
rect 666356 124002 666754 124062
rect 674465 123994 674531 123997
rect 674465 123992 676292 123994
rect 674465 123936 674470 123992
rect 674526 123936 676292 123992
rect 674465 123934 676292 123936
rect 674465 123931 674531 123934
rect 578693 123586 578759 123589
rect 575798 123584 578759 123586
rect 575798 123528 578698 123584
rect 578754 123528 578759 123584
rect 575798 123526 578759 123528
rect 575798 123012 575858 123526
rect 578693 123523 578759 123526
rect 672993 123586 673059 123589
rect 672993 123584 676292 123586
rect 672993 123528 672998 123584
rect 673054 123528 676292 123584
rect 672993 123526 676292 123528
rect 672993 123523 673059 123526
rect 589457 123178 589523 123181
rect 589457 123176 592572 123178
rect 589457 123120 589462 123176
rect 589518 123120 592572 123176
rect 589457 123118 592572 123120
rect 589457 123115 589523 123118
rect 672533 122906 672599 122909
rect 676262 122906 676322 123148
rect 672533 122904 676322 122906
rect 672533 122848 672538 122904
rect 672594 122848 676322 122904
rect 672533 122846 676322 122848
rect 672533 122843 672599 122846
rect 675017 122498 675083 122501
rect 676262 122498 676322 122740
rect 675017 122496 676322 122498
rect 675017 122440 675022 122496
rect 675078 122440 676322 122496
rect 675017 122438 676322 122440
rect 675017 122435 675083 122438
rect 667197 122090 667263 122093
rect 675334 122090 675340 122092
rect 667197 122088 675340 122090
rect 667197 122032 667202 122088
rect 667258 122032 675340 122088
rect 667197 122030 675340 122032
rect 667197 122027 667263 122030
rect 675334 122028 675340 122030
rect 675404 122090 675410 122092
rect 676262 122090 676322 122332
rect 675404 122030 676322 122090
rect 675404 122028 675410 122030
rect 672073 121682 672139 121685
rect 675017 121682 675083 121685
rect 676262 121682 676322 121924
rect 672073 121680 675083 121682
rect 672073 121624 672078 121680
rect 672134 121624 675022 121680
rect 675078 121624 675083 121680
rect 672073 121622 675083 121624
rect 672073 121619 672139 121622
rect 675017 121619 675083 121622
rect 675894 121622 676322 121682
rect 589273 121546 589339 121549
rect 589273 121544 592572 121546
rect 589273 121488 589278 121544
rect 589334 121488 592572 121544
rect 589273 121486 592572 121488
rect 589273 121483 589339 121486
rect 578877 121410 578943 121413
rect 575798 121408 578943 121410
rect 575798 121352 578882 121408
rect 578938 121352 578943 121408
rect 575798 121350 578943 121352
rect 575798 120836 575858 121350
rect 578877 121347 578943 121350
rect 668945 120866 669011 120869
rect 666694 120864 669011 120866
rect 666694 120808 668950 120864
rect 669006 120808 669011 120864
rect 666694 120806 669011 120808
rect 666694 120798 666754 120806
rect 668945 120803 669011 120806
rect 666356 120738 666754 120798
rect 675894 120730 675954 121622
rect 673410 120670 675954 120730
rect 668761 120594 668827 120597
rect 673410 120594 673470 120670
rect 668761 120592 673470 120594
rect 668761 120536 668766 120592
rect 668822 120536 673470 120592
rect 668761 120534 673470 120536
rect 668761 120531 668827 120534
rect 589641 119914 589707 119917
rect 589641 119912 592572 119914
rect 589641 119856 589646 119912
rect 589702 119856 592572 119912
rect 589641 119854 592572 119856
rect 589641 119851 589707 119854
rect 672717 119234 672783 119237
rect 666694 119232 672783 119234
rect 666694 119176 672722 119232
rect 672778 119176 672783 119232
rect 666694 119174 672783 119176
rect 666694 119166 666754 119174
rect 672717 119171 672783 119174
rect 666356 119106 666754 119166
rect 575982 118418 576042 118660
rect 578509 118418 578575 118421
rect 575982 118416 578575 118418
rect 575982 118360 578514 118416
rect 578570 118360 578575 118416
rect 575982 118358 578575 118360
rect 578509 118355 578575 118358
rect 590101 118282 590167 118285
rect 590101 118280 592572 118282
rect 590101 118224 590106 118280
rect 590162 118224 592572 118280
rect 590101 118222 592572 118224
rect 590101 118219 590167 118222
rect 666356 117474 666938 117534
rect 666878 117466 666938 117474
rect 674281 117466 674347 117469
rect 666878 117464 674347 117466
rect 666878 117408 674286 117464
rect 674342 117408 674347 117464
rect 666878 117406 674347 117408
rect 674281 117403 674347 117406
rect 675702 117268 675708 117332
rect 675772 117330 675778 117332
rect 682377 117330 682443 117333
rect 675772 117328 682443 117330
rect 675772 117272 682382 117328
rect 682438 117272 682443 117328
rect 675772 117270 682443 117272
rect 675772 117268 675778 117270
rect 682377 117267 682443 117270
rect 579521 116922 579587 116925
rect 575798 116920 579587 116922
rect 575798 116864 579526 116920
rect 579582 116864 579587 116920
rect 575798 116862 579587 116864
rect 575798 116484 575858 116862
rect 579521 116859 579587 116862
rect 589457 116650 589523 116653
rect 589457 116648 592572 116650
rect 589457 116592 589462 116648
rect 589518 116592 592572 116648
rect 589457 116590 592572 116592
rect 589457 116587 589523 116590
rect 669037 116514 669103 116517
rect 672533 116514 672599 116517
rect 669037 116512 672599 116514
rect 669037 116456 669042 116512
rect 669098 116456 672538 116512
rect 672594 116456 672599 116512
rect 669037 116454 672599 116456
rect 669037 116451 669103 116454
rect 672533 116451 672599 116454
rect 675109 116378 675175 116381
rect 675845 116378 675911 116381
rect 675109 116376 675911 116378
rect 675109 116320 675114 116376
rect 675170 116320 675850 116376
rect 675906 116320 675911 116376
rect 675109 116318 675911 116320
rect 675109 116315 675175 116318
rect 675845 116315 675911 116318
rect 675109 116106 675175 116109
rect 676029 116106 676095 116109
rect 675109 116104 676095 116106
rect 675109 116048 675114 116104
rect 675170 116048 676034 116104
rect 676090 116048 676095 116104
rect 675109 116046 676095 116048
rect 675109 116043 675175 116046
rect 676029 116043 676095 116046
rect 666356 115842 666754 115902
rect 666694 115834 666754 115842
rect 669221 115834 669287 115837
rect 666694 115832 669287 115834
rect 666694 115776 669226 115832
rect 669282 115776 669287 115832
rect 666694 115774 669287 115776
rect 669221 115771 669287 115774
rect 674046 115772 674052 115836
rect 674116 115834 674122 115836
rect 675477 115834 675543 115837
rect 674116 115832 675543 115834
rect 674116 115776 675482 115832
rect 675538 115776 675543 115832
rect 674116 115774 675543 115776
rect 674116 115772 674122 115774
rect 675477 115771 675543 115774
rect 590285 115018 590351 115021
rect 590285 115016 592572 115018
rect 590285 114960 590290 115016
rect 590346 114960 592572 115016
rect 590285 114958 592572 114960
rect 590285 114955 590351 114958
rect 669221 114610 669287 114613
rect 674097 114610 674163 114613
rect 669221 114608 674163 114610
rect 669221 114552 669226 114608
rect 669282 114552 674102 114608
rect 674158 114552 674163 114608
rect 669221 114550 674163 114552
rect 669221 114547 669287 114550
rect 674097 114547 674163 114550
rect 579245 114474 579311 114477
rect 575798 114472 579311 114474
rect 575798 114416 579250 114472
rect 579306 114416 579311 114472
rect 575798 114414 579311 114416
rect 575798 114308 575858 114414
rect 579245 114411 579311 114414
rect 669037 114338 669103 114341
rect 666694 114336 669103 114338
rect 666694 114280 669042 114336
rect 669098 114280 669103 114336
rect 666694 114278 669103 114280
rect 666694 114270 666754 114278
rect 669037 114275 669103 114278
rect 669221 114338 669287 114341
rect 672073 114338 672139 114341
rect 669221 114336 672139 114338
rect 669221 114280 669226 114336
rect 669282 114280 672078 114336
rect 672134 114280 672139 114336
rect 669221 114278 672139 114280
rect 669221 114275 669287 114278
rect 672073 114275 672139 114278
rect 666356 114210 666754 114270
rect 589457 113386 589523 113389
rect 589457 113384 592572 113386
rect 589457 113328 589462 113384
rect 589518 113328 592572 113384
rect 589457 113326 592572 113328
rect 589457 113323 589523 113326
rect 669221 112706 669287 112709
rect 666694 112704 669287 112706
rect 666694 112648 669226 112704
rect 669282 112648 669287 112704
rect 666694 112646 669287 112648
rect 666694 112638 666754 112646
rect 669221 112643 669287 112646
rect 666356 112578 666754 112638
rect 579521 112570 579587 112573
rect 575798 112568 579587 112570
rect 575798 112512 579526 112568
rect 579582 112512 579587 112568
rect 575798 112510 579587 112512
rect 575798 112132 575858 112510
rect 579521 112507 579587 112510
rect 675753 112434 675819 112437
rect 676254 112434 676260 112436
rect 675753 112432 676260 112434
rect 675753 112376 675758 112432
rect 675814 112376 676260 112432
rect 675753 112374 676260 112376
rect 675753 112371 675819 112374
rect 676254 112372 676260 112374
rect 676324 112372 676330 112436
rect 589457 111754 589523 111757
rect 675753 111754 675819 111757
rect 676622 111754 676628 111756
rect 589457 111752 592572 111754
rect 589457 111696 589462 111752
rect 589518 111696 592572 111752
rect 589457 111694 592572 111696
rect 675753 111752 676628 111754
rect 675753 111696 675758 111752
rect 675814 111696 676628 111752
rect 675753 111694 676628 111696
rect 589457 111691 589523 111694
rect 675753 111691 675819 111694
rect 676622 111692 676628 111694
rect 676692 111692 676698 111756
rect 675753 111348 675819 111349
rect 675702 111284 675708 111348
rect 675772 111346 675819 111348
rect 675772 111344 675864 111346
rect 675814 111288 675864 111344
rect 675772 111286 675864 111288
rect 675772 111284 675819 111286
rect 675753 111283 675819 111284
rect 668761 111074 668827 111077
rect 666694 111072 668827 111074
rect 666694 111016 668766 111072
rect 668822 111016 668827 111072
rect 666694 111014 668827 111016
rect 666694 111006 666754 111014
rect 668761 111011 668827 111014
rect 666356 110946 666754 111006
rect 675753 110394 675819 110397
rect 676438 110394 676444 110396
rect 675753 110392 676444 110394
rect 675753 110336 675758 110392
rect 675814 110336 676444 110392
rect 675753 110334 676444 110336
rect 675753 110331 675819 110334
rect 676438 110332 676444 110334
rect 676508 110332 676514 110396
rect 579337 110122 579403 110125
rect 575798 110120 579403 110122
rect 575798 110064 579342 110120
rect 579398 110064 579403 110120
rect 575798 110062 579403 110064
rect 575798 109956 575858 110062
rect 579337 110059 579403 110062
rect 589457 110122 589523 110125
rect 589457 110120 592572 110122
rect 589457 110064 589462 110120
rect 589518 110064 592572 110120
rect 589457 110062 592572 110064
rect 589457 110059 589523 110062
rect 666645 109374 666711 109377
rect 666356 109372 666711 109374
rect 666356 109316 666650 109372
rect 666706 109316 666711 109372
rect 666356 109314 666711 109316
rect 666645 109311 666711 109314
rect 589457 108490 589523 108493
rect 589457 108488 592572 108490
rect 589457 108432 589462 108488
rect 589518 108432 592572 108488
rect 589457 108430 592572 108432
rect 589457 108427 589523 108430
rect 578325 108354 578391 108357
rect 575798 108352 578391 108354
rect 575798 108296 578330 108352
rect 578386 108296 578391 108352
rect 575798 108294 578391 108296
rect 575798 107780 575858 108294
rect 578325 108291 578391 108294
rect 675753 108218 675819 108221
rect 676070 108218 676076 108220
rect 675753 108216 676076 108218
rect 675753 108160 675758 108216
rect 675814 108160 676076 108216
rect 675753 108158 676076 108160
rect 675753 108155 675819 108158
rect 676070 108156 676076 108158
rect 676140 108156 676146 108220
rect 667933 107810 667999 107813
rect 666694 107808 667999 107810
rect 666694 107752 667938 107808
rect 667994 107752 667999 107808
rect 666694 107750 667999 107752
rect 666694 107742 666754 107750
rect 667933 107747 667999 107750
rect 666356 107682 666754 107742
rect 674465 107538 674531 107541
rect 675385 107538 675451 107541
rect 674465 107536 675451 107538
rect 674465 107480 674470 107536
rect 674526 107480 675390 107536
rect 675446 107480 675451 107536
rect 674465 107478 675451 107480
rect 674465 107475 674531 107478
rect 675385 107475 675451 107478
rect 673177 106994 673243 106997
rect 675385 106994 675451 106997
rect 673177 106992 675451 106994
rect 673177 106936 673182 106992
rect 673238 106936 675390 106992
rect 675446 106936 675451 106992
rect 673177 106934 675451 106936
rect 673177 106931 673243 106934
rect 675385 106931 675451 106934
rect 589457 106858 589523 106861
rect 589457 106856 592572 106858
rect 589457 106800 589462 106856
rect 589518 106800 592572 106856
rect 589457 106798 592572 106800
rect 589457 106795 589523 106798
rect 668117 106178 668183 106181
rect 668393 106178 668459 106181
rect 666694 106176 668459 106178
rect 666694 106120 668122 106176
rect 668178 106120 668398 106176
rect 668454 106120 668459 106176
rect 666694 106118 668459 106120
rect 666694 106110 666754 106118
rect 668117 106115 668183 106118
rect 668393 106115 668459 106118
rect 666356 106050 666754 106110
rect 672993 106042 673059 106045
rect 675385 106042 675451 106045
rect 672993 106040 675451 106042
rect 672993 105984 672998 106040
rect 673054 105984 675390 106040
rect 675446 105984 675451 106040
rect 672993 105982 675451 105984
rect 672993 105979 673059 105982
rect 675385 105979 675451 105982
rect 579061 105906 579127 105909
rect 575798 105904 579127 105906
rect 575798 105848 579066 105904
rect 579122 105848 579127 105904
rect 575798 105846 579127 105848
rect 575798 105604 575858 105846
rect 579061 105843 579127 105846
rect 589825 105226 589891 105229
rect 589825 105224 592572 105226
rect 589825 105168 589830 105224
rect 589886 105168 592572 105224
rect 589825 105166 592572 105168
rect 589825 105163 589891 105166
rect 666356 104418 666754 104478
rect 666694 104410 666754 104418
rect 668301 104410 668367 104413
rect 666694 104408 668367 104410
rect 666694 104352 668306 104408
rect 668362 104352 668367 104408
rect 666694 104350 668367 104352
rect 668301 104347 668367 104350
rect 588537 103594 588603 103597
rect 588537 103592 592572 103594
rect 588537 103536 588542 103592
rect 588598 103536 592572 103592
rect 588537 103534 592572 103536
rect 588537 103531 588603 103534
rect 575982 103186 576042 103428
rect 578509 103186 578575 103189
rect 575982 103184 578575 103186
rect 575982 103128 578514 103184
rect 578570 103128 578575 103184
rect 575982 103126 578575 103128
rect 578509 103123 578575 103126
rect 666356 102786 666754 102846
rect 666694 102778 666754 102786
rect 667933 102778 667999 102781
rect 668577 102778 668643 102781
rect 666694 102776 668643 102778
rect 666694 102720 667938 102776
rect 667994 102720 668582 102776
rect 668638 102720 668643 102776
rect 666694 102718 668643 102720
rect 667933 102715 667999 102718
rect 668577 102715 668643 102718
rect 675385 102644 675451 102645
rect 675334 102642 675340 102644
rect 675294 102582 675340 102642
rect 675404 102640 675451 102644
rect 675446 102584 675451 102640
rect 675334 102580 675340 102582
rect 675404 102580 675451 102584
rect 675385 102579 675451 102580
rect 589457 101962 589523 101965
rect 589457 101960 592572 101962
rect 589457 101904 589462 101960
rect 589518 101904 592572 101960
rect 589457 101902 592572 101904
rect 589457 101899 589523 101902
rect 579153 101690 579219 101693
rect 575798 101688 579219 101690
rect 575798 101632 579158 101688
rect 579214 101632 579219 101688
rect 575798 101630 579219 101632
rect 575798 101252 575858 101630
rect 579153 101627 579219 101630
rect 673361 101010 673427 101013
rect 675109 101010 675175 101013
rect 673361 101008 675175 101010
rect 673361 100952 673366 101008
rect 673422 100952 675114 101008
rect 675170 100952 675175 101008
rect 673361 100950 675175 100952
rect 673361 100947 673427 100950
rect 675109 100947 675175 100950
rect 579521 99242 579587 99245
rect 575798 99240 579587 99242
rect 575798 99184 579526 99240
rect 579582 99184 579587 99240
rect 575798 99182 579587 99184
rect 575798 99076 575858 99182
rect 579521 99179 579587 99182
rect 578601 97474 578667 97477
rect 575798 97472 578667 97474
rect 575798 97416 578606 97472
rect 578662 97416 578667 97472
rect 575798 97414 578667 97416
rect 575798 96900 575858 97414
rect 578601 97411 578667 97414
rect 635549 96930 635615 96933
rect 635774 96930 635780 96932
rect 635549 96928 635780 96930
rect 635549 96872 635554 96928
rect 635610 96872 635780 96928
rect 635549 96870 635780 96872
rect 635549 96867 635615 96870
rect 635774 96868 635780 96870
rect 635844 96868 635850 96932
rect 637021 96930 637087 96933
rect 637246 96930 637252 96932
rect 637021 96928 637252 96930
rect 637021 96872 637026 96928
rect 637082 96872 637252 96928
rect 637021 96870 637252 96872
rect 637021 96867 637087 96870
rect 637246 96868 637252 96870
rect 637316 96868 637322 96932
rect 641989 96522 642055 96525
rect 647182 96522 647188 96524
rect 641989 96520 647188 96522
rect 641989 96464 641994 96520
rect 642050 96464 647188 96520
rect 641989 96462 647188 96464
rect 641989 96459 642055 96462
rect 647182 96460 647188 96462
rect 647252 96460 647258 96524
rect 648061 96522 648127 96525
rect 649257 96522 649323 96525
rect 648061 96520 649323 96522
rect 648061 96464 648066 96520
rect 648122 96464 649262 96520
rect 649318 96464 649323 96520
rect 648061 96462 649323 96464
rect 648061 96459 648127 96462
rect 649257 96459 649323 96462
rect 644933 96114 644999 96117
rect 648613 96114 648679 96117
rect 644933 96112 648679 96114
rect 644933 96056 644938 96112
rect 644994 96056 648618 96112
rect 648674 96056 648679 96112
rect 644933 96054 648679 96056
rect 644933 96051 644999 96054
rect 648613 96051 648679 96054
rect 633934 95916 633940 95980
rect 634004 95978 634010 95980
rect 635733 95978 635799 95981
rect 634004 95976 635799 95978
rect 634004 95920 635738 95976
rect 635794 95920 635799 95976
rect 634004 95918 635799 95920
rect 634004 95916 634010 95918
rect 635733 95915 635799 95918
rect 647877 95842 647943 95845
rect 656341 95842 656407 95845
rect 647877 95840 656407 95842
rect 647877 95784 647882 95840
rect 647938 95784 656346 95840
rect 656402 95784 656407 95840
rect 647877 95782 656407 95784
rect 647877 95779 647943 95782
rect 656341 95779 656407 95782
rect 578325 95026 578391 95029
rect 575798 95024 578391 95026
rect 575798 94968 578330 95024
rect 578386 94968 578391 95024
rect 575798 94966 578391 94968
rect 575798 94724 575858 94966
rect 578325 94963 578391 94966
rect 647325 95026 647391 95029
rect 647325 95024 647434 95026
rect 647325 94968 647330 95024
rect 647386 94968 647434 95024
rect 647325 94963 647434 94968
rect 625429 94482 625495 94485
rect 625429 94480 628268 94482
rect 625429 94424 625434 94480
rect 625490 94424 628268 94480
rect 647374 94452 647434 94963
rect 625429 94422 628268 94424
rect 625429 94419 625495 94422
rect 655237 94210 655303 94213
rect 655237 94208 656788 94210
rect 655237 94152 655242 94208
rect 655298 94152 656788 94208
rect 655237 94150 656788 94152
rect 655237 94147 655303 94150
rect 626441 93666 626507 93669
rect 626441 93664 628268 93666
rect 626441 93608 626446 93664
rect 626502 93608 628268 93664
rect 626441 93606 628268 93608
rect 626441 93603 626507 93606
rect 654685 93394 654751 93397
rect 665357 93394 665423 93397
rect 654685 93392 656788 93394
rect 654685 93336 654690 93392
rect 654746 93336 656788 93392
rect 654685 93334 656788 93336
rect 663596 93392 665423 93394
rect 663596 93336 665362 93392
rect 665418 93336 665423 93392
rect 663596 93334 665423 93336
rect 654685 93331 654751 93334
rect 665357 93331 665423 93334
rect 579245 93122 579311 93125
rect 575798 93120 579311 93122
rect 575798 93064 579250 93120
rect 579306 93064 579311 93120
rect 575798 93062 579311 93064
rect 575798 92548 575858 93062
rect 579245 93059 579311 93062
rect 650310 93060 650316 93124
rect 650380 93122 650386 93124
rect 663793 93122 663859 93125
rect 650380 93062 656818 93122
rect 650380 93060 650386 93062
rect 626257 92850 626323 92853
rect 626257 92848 628268 92850
rect 626257 92792 626262 92848
rect 626318 92792 628268 92848
rect 626257 92790 628268 92792
rect 626257 92787 626323 92790
rect 656758 92548 656818 93062
rect 663566 93120 663859 93122
rect 663566 93064 663798 93120
rect 663854 93064 663859 93120
rect 663566 93062 663859 93064
rect 663566 92548 663626 93062
rect 663793 93059 663859 93062
rect 625797 92034 625863 92037
rect 648797 92034 648863 92037
rect 625797 92032 628268 92034
rect 625797 91976 625802 92032
rect 625858 91976 628268 92032
rect 625797 91974 628268 91976
rect 648140 92032 648863 92034
rect 648140 91976 648802 92032
rect 648858 91976 648863 92032
rect 648140 91974 648863 91976
rect 625797 91971 625863 91974
rect 648797 91971 648863 91974
rect 663977 91762 664043 91765
rect 663596 91760 664043 91762
rect 663596 91704 663982 91760
rect 664038 91704 664043 91760
rect 663596 91702 664043 91704
rect 663977 91699 664043 91702
rect 655421 91490 655487 91493
rect 655421 91488 656788 91490
rect 655421 91432 655426 91488
rect 655482 91432 656788 91488
rect 655421 91430 656788 91432
rect 655421 91427 655487 91430
rect 626441 91218 626507 91221
rect 626441 91216 628268 91218
rect 626441 91160 626446 91216
rect 626502 91160 628268 91216
rect 626441 91158 628268 91160
rect 626441 91155 626507 91158
rect 578601 90946 578667 90949
rect 575798 90944 578667 90946
rect 575798 90888 578606 90944
rect 578662 90888 578667 90944
rect 575798 90886 578667 90888
rect 575798 90372 575858 90886
rect 578601 90883 578667 90886
rect 655421 90674 655487 90677
rect 664345 90674 664411 90677
rect 655421 90672 656788 90674
rect 655421 90616 655426 90672
rect 655482 90616 656788 90672
rect 655421 90614 656788 90616
rect 663596 90672 664411 90674
rect 663596 90616 664350 90672
rect 664406 90616 664411 90672
rect 663596 90614 664411 90616
rect 655421 90611 655487 90614
rect 664345 90611 664411 90614
rect 626441 90402 626507 90405
rect 626441 90400 628268 90402
rect 626441 90344 626446 90400
rect 626502 90344 628268 90400
rect 626441 90342 628268 90344
rect 626441 90339 626507 90342
rect 655789 89858 655855 89861
rect 664529 89858 664595 89861
rect 655789 89856 656788 89858
rect 655789 89800 655794 89856
rect 655850 89800 656788 89856
rect 655789 89798 656788 89800
rect 663596 89856 664595 89858
rect 663596 89800 664534 89856
rect 664590 89800 664595 89856
rect 663596 89798 664595 89800
rect 655789 89795 655855 89798
rect 664529 89795 664595 89798
rect 625245 89586 625311 89589
rect 648245 89586 648311 89589
rect 625245 89584 628268 89586
rect 625245 89528 625250 89584
rect 625306 89528 628268 89584
rect 625245 89526 628268 89528
rect 648140 89584 648311 89586
rect 648140 89528 648250 89584
rect 648306 89528 648311 89584
rect 648140 89526 648311 89528
rect 625245 89523 625311 89526
rect 648245 89523 648311 89526
rect 665173 89042 665239 89045
rect 663596 89040 665239 89042
rect 663596 88984 665178 89040
rect 665234 88984 665239 89040
rect 663596 88982 665239 88984
rect 665173 88979 665239 88982
rect 625429 88770 625495 88773
rect 625429 88768 628268 88770
rect 625429 88712 625434 88768
rect 625490 88712 628268 88768
rect 625429 88710 628268 88712
rect 625429 88707 625495 88710
rect 624969 88634 625035 88637
rect 625245 88634 625311 88637
rect 624969 88632 625311 88634
rect 624969 88576 624974 88632
rect 625030 88576 625250 88632
rect 625306 88576 625311 88632
rect 624969 88574 625311 88576
rect 624969 88571 625035 88574
rect 625245 88571 625311 88574
rect 575982 88090 576042 88196
rect 579245 88090 579311 88093
rect 575982 88088 579311 88090
rect 575982 88032 579250 88088
rect 579306 88032 579311 88088
rect 575982 88030 579311 88032
rect 579245 88027 579311 88030
rect 626441 87954 626507 87957
rect 626441 87952 628268 87954
rect 626441 87896 626446 87952
rect 626502 87896 628268 87952
rect 626441 87894 628268 87896
rect 626441 87891 626507 87894
rect 626257 87138 626323 87141
rect 650545 87138 650611 87141
rect 626257 87136 628268 87138
rect 626257 87080 626262 87136
rect 626318 87080 628268 87136
rect 626257 87078 628268 87080
rect 648140 87136 650611 87138
rect 648140 87080 650550 87136
rect 650606 87080 650611 87136
rect 648140 87078 650611 87080
rect 626257 87075 626323 87078
rect 650545 87075 650611 87078
rect 578325 86458 578391 86461
rect 575798 86456 578391 86458
rect 575798 86400 578330 86456
rect 578386 86400 578391 86456
rect 575798 86398 578391 86400
rect 575798 86020 575858 86398
rect 578325 86395 578391 86398
rect 626441 86322 626507 86325
rect 626441 86320 628268 86322
rect 626441 86264 626446 86320
rect 626502 86264 628268 86320
rect 626441 86262 628268 86264
rect 626441 86259 626507 86262
rect 626441 85506 626507 85509
rect 626441 85504 628268 85506
rect 626441 85448 626446 85504
rect 626502 85448 628268 85504
rect 626441 85446 628268 85448
rect 626441 85443 626507 85446
rect 625245 84690 625311 84693
rect 648613 84690 648679 84693
rect 625245 84688 628268 84690
rect 625245 84632 625250 84688
rect 625306 84632 628268 84688
rect 625245 84630 628268 84632
rect 648140 84688 648679 84690
rect 648140 84632 648618 84688
rect 648674 84632 648679 84688
rect 648140 84630 648679 84632
rect 625245 84627 625311 84630
rect 648613 84627 648679 84630
rect 579245 84010 579311 84013
rect 575798 84008 579311 84010
rect 575798 83952 579250 84008
rect 579306 83952 579311 84008
rect 575798 83950 579311 83952
rect 575798 83844 575858 83950
rect 579245 83947 579311 83950
rect 626441 83874 626507 83877
rect 626441 83872 628268 83874
rect 626441 83816 626446 83872
rect 626502 83816 628268 83872
rect 626441 83814 628268 83816
rect 626441 83811 626507 83814
rect 628741 83330 628807 83333
rect 628741 83328 628850 83330
rect 628741 83272 628746 83328
rect 628802 83272 628850 83328
rect 628741 83267 628850 83272
rect 628790 83028 628850 83267
rect 578877 82242 578943 82245
rect 650269 82242 650335 82245
rect 575798 82240 578943 82242
rect 575798 82184 578882 82240
rect 578938 82184 578943 82240
rect 648140 82240 650335 82242
rect 575798 82182 578943 82184
rect 575798 81668 575858 82182
rect 578877 82179 578943 82182
rect 628790 81698 628850 82212
rect 648140 82184 650274 82240
rect 650330 82184 650335 82240
rect 648140 82182 650335 82184
rect 650269 82179 650335 82182
rect 629201 81698 629267 81701
rect 628790 81696 629267 81698
rect 628790 81640 629206 81696
rect 629262 81640 629267 81696
rect 628790 81638 629267 81640
rect 629201 81635 629267 81638
rect 579429 80066 579495 80069
rect 575798 80064 579495 80066
rect 575798 80008 579434 80064
rect 579490 80008 579495 80064
rect 575798 80006 579495 80008
rect 575798 79492 575858 80006
rect 579429 80003 579495 80006
rect 633893 78572 633959 78573
rect 633893 78570 633940 78572
rect 633848 78568 633940 78570
rect 633848 78512 633898 78568
rect 633848 78510 633940 78512
rect 633893 78508 633940 78510
rect 634004 78508 634010 78572
rect 633893 78507 633959 78508
rect 635774 78100 635780 78164
rect 635844 78162 635850 78164
rect 647509 78162 647575 78165
rect 635844 78160 647575 78162
rect 635844 78104 647514 78160
rect 647570 78104 647575 78160
rect 635844 78102 647575 78104
rect 635844 78100 635850 78102
rect 647509 78099 647575 78102
rect 578233 77890 578299 77893
rect 575798 77888 578299 77890
rect 575798 77832 578238 77888
rect 578294 77832 578299 77888
rect 575798 77830 578299 77832
rect 575798 77316 575858 77830
rect 578233 77827 578299 77830
rect 580441 77890 580507 77893
rect 580441 77888 625170 77890
rect 580441 77832 580446 77888
rect 580502 77832 625170 77888
rect 580441 77830 625170 77832
rect 580441 77827 580507 77830
rect 625110 77618 625170 77830
rect 637062 77618 637068 77620
rect 625110 77558 637068 77618
rect 637062 77556 637068 77558
rect 637132 77618 637138 77620
rect 639597 77618 639663 77621
rect 637132 77616 639663 77618
rect 637132 77560 639602 77616
rect 639658 77560 639663 77616
rect 637132 77558 639663 77560
rect 637132 77556 637138 77558
rect 639597 77555 639663 77558
rect 623037 77346 623103 77349
rect 633893 77346 633959 77349
rect 623037 77344 633959 77346
rect 623037 77288 623042 77344
rect 623098 77288 633898 77344
rect 633954 77288 633959 77344
rect 623037 77286 633959 77288
rect 623037 77283 623103 77286
rect 633893 77283 633959 77286
rect 579245 75714 579311 75717
rect 575798 75712 579311 75714
rect 575798 75656 579250 75712
rect 579306 75656 579311 75712
rect 575798 75654 579311 75656
rect 575798 75140 575858 75654
rect 579245 75651 579311 75654
rect 646497 74218 646563 74221
rect 646454 74216 646563 74218
rect 646454 74160 646502 74216
rect 646558 74160 646563 74216
rect 646454 74155 646563 74160
rect 646454 73848 646514 74155
rect 579521 73130 579587 73133
rect 575798 73128 579587 73130
rect 575798 73072 579526 73128
rect 579582 73072 579587 73128
rect 575798 73070 579587 73072
rect 575798 72964 575858 73070
rect 579521 73067 579587 73070
rect 646681 71770 646747 71773
rect 646638 71768 646747 71770
rect 646638 71712 646686 71768
rect 646742 71712 646747 71768
rect 646638 71707 646747 71712
rect 646638 71400 646698 71707
rect 578509 71226 578575 71229
rect 575798 71224 578575 71226
rect 575798 71168 578514 71224
rect 578570 71168 578575 71224
rect 575798 71166 578575 71168
rect 575798 70788 575858 71166
rect 578509 71163 578575 71166
rect 646313 69186 646379 69189
rect 646270 69184 646379 69186
rect 646270 69128 646318 69184
rect 646374 69128 646379 69184
rect 646270 69123 646379 69128
rect 646270 68952 646330 69123
rect 575798 66874 575858 68612
rect 646129 67146 646195 67149
rect 646086 67144 646195 67146
rect 646086 67088 646134 67144
rect 646190 67088 646195 67144
rect 646086 67083 646195 67088
rect 579521 66874 579587 66877
rect 575798 66872 579587 66874
rect 575798 66816 579526 66872
rect 579582 66816 579587 66872
rect 575798 66814 579587 66816
rect 575798 66436 575858 66814
rect 579521 66811 579587 66814
rect 646086 66504 646146 67083
rect 579521 64562 579587 64565
rect 575798 64560 579587 64562
rect 575798 64504 579526 64560
rect 579582 64504 579587 64560
rect 575798 64502 579587 64504
rect 575798 64260 575858 64502
rect 579521 64499 579587 64502
rect 647325 64426 647391 64429
rect 646638 64424 647391 64426
rect 646638 64368 647330 64424
rect 647386 64368 647391 64424
rect 646638 64366 647391 64368
rect 646638 64056 646698 64366
rect 647325 64363 647391 64366
rect 648981 62114 649047 62117
rect 646638 62112 649047 62114
rect 575982 61842 576042 62084
rect 646638 62056 648986 62112
rect 649042 62056 649047 62112
rect 646638 62054 649047 62056
rect 579521 61842 579587 61845
rect 575982 61840 579587 61842
rect 575982 61784 579526 61840
rect 579582 61784 579587 61840
rect 575982 61782 579587 61784
rect 579521 61779 579587 61782
rect 646638 61608 646698 62054
rect 648981 62051 649047 62054
rect 578877 60482 578943 60485
rect 575798 60480 578943 60482
rect 575798 60424 578882 60480
rect 578938 60424 578943 60480
rect 575798 60422 578943 60424
rect 575798 59908 575858 60422
rect 578877 60419 578943 60422
rect 648613 59258 648679 59261
rect 646638 59256 648679 59258
rect 646638 59200 648618 59256
rect 648674 59200 648679 59256
rect 646638 59198 648679 59200
rect 646638 59160 646698 59198
rect 648613 59195 648679 59198
rect 579521 57898 579587 57901
rect 575798 57896 579587 57898
rect 575798 57840 579526 57896
rect 579582 57840 579587 57896
rect 575798 57838 579587 57840
rect 575798 57732 575858 57838
rect 579521 57835 579587 57838
rect 647509 57354 647575 57357
rect 646638 57352 647575 57354
rect 646638 57296 647514 57352
rect 647570 57296 647575 57352
rect 646638 57294 647575 57296
rect 646638 56712 646698 57294
rect 647509 57291 647575 57294
rect 578325 56130 578391 56133
rect 575798 56128 578391 56130
rect 575798 56072 578330 56128
rect 578386 56072 578391 56128
rect 575798 56070 578391 56072
rect 575798 55556 575858 56070
rect 578325 56067 578391 56070
rect 462630 54980 462636 55044
rect 462700 55042 462706 55044
rect 577497 55042 577563 55045
rect 462700 55040 577563 55042
rect 462700 54984 577502 55040
rect 577558 54984 577563 55040
rect 462700 54982 577563 54984
rect 462700 54980 462706 54982
rect 577497 54979 577563 54982
rect 574461 54770 574527 54773
rect 459878 54768 574527 54770
rect 459878 54712 574466 54768
rect 574522 54712 574527 54768
rect 459878 54710 574527 54712
rect 459878 53685 459938 54710
rect 574461 54707 574527 54710
rect 591297 54498 591363 54501
rect 466410 54496 591363 54498
rect 466410 54440 591302 54496
rect 591358 54440 591363 54496
rect 466410 54438 591363 54440
rect 466410 54226 466470 54438
rect 591297 54435 591363 54438
rect 576117 54226 576183 54229
rect 460798 54166 466470 54226
rect 476070 54224 576183 54226
rect 476070 54168 576122 54224
rect 576178 54168 576183 54224
rect 476070 54166 576183 54168
rect 460798 53685 460858 54166
rect 476070 53954 476130 54166
rect 576117 54163 576183 54166
rect 461718 53894 476130 53954
rect 461718 53685 461778 53894
rect 459829 53680 459938 53685
rect 459829 53624 459834 53680
rect 459890 53624 459938 53680
rect 459829 53622 459938 53624
rect 460749 53680 460858 53685
rect 460749 53624 460754 53680
rect 460810 53624 460858 53680
rect 460749 53622 460858 53624
rect 461669 53680 461778 53685
rect 462589 53684 462655 53685
rect 462589 53682 462636 53684
rect 461669 53624 461674 53680
rect 461730 53624 461778 53680
rect 461669 53622 461778 53624
rect 462544 53680 462636 53682
rect 462544 53624 462594 53680
rect 462544 53622 462636 53624
rect 459829 53619 459895 53622
rect 460749 53619 460815 53622
rect 461669 53619 461735 53622
rect 462589 53620 462636 53622
rect 462700 53620 462706 53684
rect 462589 53619 462655 53620
rect 468293 53274 468359 53277
rect 475193 53274 475259 53277
rect 468293 53272 475259 53274
rect 468293 53216 468298 53272
rect 468354 53216 475198 53272
rect 475254 53216 475259 53272
rect 468293 53214 475259 53216
rect 468293 53211 468359 53214
rect 475193 53211 475259 53214
rect 194358 50220 194364 50284
rect 194428 50282 194434 50284
rect 308029 50282 308095 50285
rect 194428 50280 308095 50282
rect 194428 50224 308034 50280
rect 308090 50224 308095 50280
rect 194428 50222 308095 50224
rect 194428 50220 194434 50222
rect 308029 50219 308095 50222
rect 518750 48860 518756 48924
rect 518820 48922 518826 48924
rect 549989 48922 550055 48925
rect 518820 48920 550055 48922
rect 518820 48864 549994 48920
rect 550050 48864 550055 48920
rect 518820 48862 550055 48864
rect 518820 48860 518826 48862
rect 549989 48859 550055 48862
rect 661585 48512 661651 48515
rect 661480 48510 661651 48512
rect 661480 48454 661590 48510
rect 661646 48454 661651 48510
rect 661480 48452 661651 48454
rect 661585 48449 661651 48452
rect 529606 48044 529612 48108
rect 529676 48106 529682 48108
rect 553669 48106 553735 48109
rect 529676 48104 553735 48106
rect 529676 48048 553674 48104
rect 553730 48048 553735 48104
rect 529676 48046 553735 48048
rect 529676 48044 529682 48046
rect 553669 48043 553735 48046
rect 515438 47772 515444 47836
rect 515508 47834 515514 47836
rect 522941 47834 523007 47837
rect 515508 47832 523007 47834
rect 515508 47776 522946 47832
rect 523002 47776 523007 47832
rect 515508 47774 523007 47776
rect 515508 47772 515514 47774
rect 522941 47771 523007 47774
rect 526478 47772 526484 47836
rect 526548 47834 526554 47836
rect 552013 47834 552079 47837
rect 526548 47832 552079 47834
rect 526548 47776 552018 47832
rect 552074 47776 552079 47832
rect 661769 47791 661835 47794
rect 526548 47774 552079 47776
rect 526548 47772 526554 47774
rect 552013 47771 552079 47774
rect 661388 47789 661835 47791
rect 661388 47733 661774 47789
rect 661830 47733 661835 47789
rect 661388 47731 661835 47733
rect 661769 47728 661835 47731
rect 520958 47500 520964 47564
rect 521028 47562 521034 47564
rect 547873 47562 547939 47565
rect 521028 47560 547939 47562
rect 521028 47504 547878 47560
rect 547934 47504 547939 47560
rect 521028 47502 547939 47504
rect 521028 47500 521034 47502
rect 547873 47499 547939 47502
rect 662413 47426 662479 47429
rect 661388 47424 662479 47426
rect 661388 47368 662418 47424
rect 662474 47368 662479 47424
rect 661388 47366 662479 47368
rect 662413 47363 662479 47366
rect 522062 47228 522068 47292
rect 522132 47290 522138 47292
rect 545665 47290 545731 47293
rect 522132 47288 545731 47290
rect 522132 47232 545670 47288
rect 545726 47232 545731 47288
rect 522132 47230 545731 47232
rect 522132 47228 522138 47230
rect 545665 47227 545731 47230
rect 458173 47018 458239 47021
rect 465257 47018 465323 47021
rect 458173 47016 465323 47018
rect 458173 46960 458178 47016
rect 458234 46960 465262 47016
rect 465318 46960 465323 47016
rect 458173 46958 465323 46960
rect 458173 46955 458239 46958
rect 465257 46955 465323 46958
rect 458357 46746 458423 46749
rect 465073 46746 465139 46749
rect 458357 46744 465139 46746
rect 458357 46688 458362 46744
rect 458418 46688 465078 46744
rect 465134 46688 465139 46744
rect 458357 46686 465139 46688
rect 458357 46683 458423 46686
rect 465073 46683 465139 46686
rect 130561 44434 130627 44437
rect 132585 44434 132651 44437
rect 130561 44432 132651 44434
rect 130561 44376 130566 44432
rect 130622 44376 132590 44432
rect 132646 44376 132651 44432
rect 130561 44374 132651 44376
rect 130561 44371 130627 44374
rect 132585 44371 132651 44374
rect 458214 44372 458220 44436
rect 458284 44434 458290 44436
rect 459185 44434 459251 44437
rect 458284 44432 459251 44434
rect 458284 44376 459190 44432
rect 459246 44376 459251 44432
rect 458284 44374 459251 44376
rect 458284 44372 458290 44374
rect 459185 44371 459251 44374
rect 461342 44372 461348 44436
rect 461412 44434 461418 44436
rect 461945 44434 462011 44437
rect 461412 44432 462011 44434
rect 461412 44376 461950 44432
rect 462006 44376 462011 44432
rect 461412 44374 462011 44376
rect 461412 44372 461418 44374
rect 461945 44371 462011 44374
rect 462262 44372 462268 44436
rect 462332 44434 462338 44436
rect 462497 44434 462563 44437
rect 462332 44432 462563 44434
rect 462332 44376 462502 44432
rect 462558 44376 462563 44432
rect 462332 44374 462563 44376
rect 462332 44372 462338 44374
rect 462497 44371 462563 44374
rect 142613 44298 142679 44301
rect 142110 44296 142679 44298
rect 142110 44240 142618 44296
rect 142674 44240 142679 44296
rect 142110 44238 142679 44240
rect 141734 43964 141740 44028
rect 141804 44026 141810 44028
rect 142110 44026 142170 44238
rect 142613 44235 142679 44238
rect 255865 44162 255931 44165
rect 460105 44162 460171 44165
rect 463877 44162 463943 44165
rect 255865 44160 460171 44162
rect 255865 44104 255870 44160
rect 255926 44104 460110 44160
rect 460166 44104 460171 44160
rect 255865 44102 460171 44104
rect 255865 44099 255931 44102
rect 460105 44099 460171 44102
rect 460890 44160 463943 44162
rect 460890 44104 463882 44160
rect 463938 44104 463943 44160
rect 460890 44102 463943 44104
rect 141804 43966 142170 44026
rect 141804 43964 141810 43966
rect 307293 43890 307359 43893
rect 440233 43890 440299 43893
rect 307293 43888 440299 43890
rect 307293 43832 307298 43888
rect 307354 43832 440238 43888
rect 440294 43832 440299 43888
rect 307293 43830 440299 43832
rect 307293 43827 307359 43830
rect 440233 43827 440299 43830
rect 441061 43890 441127 43893
rect 460890 43890 460950 44102
rect 463877 44099 463943 44102
rect 441061 43888 460950 43890
rect 441061 43832 441066 43888
rect 441122 43832 460950 43888
rect 441061 43830 460950 43832
rect 441061 43827 441127 43830
rect 460841 43482 460907 43485
rect 471053 43482 471119 43485
rect 460841 43480 471119 43482
rect 460841 43424 460846 43480
rect 460902 43424 471058 43480
rect 471114 43424 471119 43480
rect 460841 43422 471119 43424
rect 460841 43419 460907 43422
rect 471053 43419 471119 43422
rect 462313 43210 462379 43213
rect 465809 43210 465875 43213
rect 462313 43208 465875 43210
rect 462313 43152 462318 43208
rect 462374 43152 465814 43208
rect 465870 43152 465875 43208
rect 462313 43150 465875 43152
rect 462313 43147 462379 43150
rect 465809 43147 465875 43150
rect 461761 42938 461827 42941
rect 463969 42938 464035 42941
rect 461761 42936 464035 42938
rect 461761 42880 461766 42936
rect 461822 42880 463974 42936
rect 464030 42880 464035 42936
rect 461761 42878 464035 42880
rect 461761 42875 461827 42878
rect 463969 42875 464035 42878
rect 518801 42804 518867 42805
rect 518750 42802 518756 42804
rect 518710 42742 518756 42802
rect 518820 42800 518867 42804
rect 518862 42744 518867 42800
rect 518750 42740 518756 42742
rect 518820 42740 518867 42744
rect 518801 42739 518867 42740
rect 416589 42394 416655 42397
rect 416589 42392 422310 42394
rect 416589 42336 416594 42392
rect 416650 42336 422310 42392
rect 416589 42334 422310 42336
rect 416589 42331 416655 42334
rect 422250 42258 422310 42334
rect 446213 42258 446279 42261
rect 461117 42258 461183 42261
rect 422250 42198 427830 42258
rect 194317 42124 194383 42125
rect 194317 42122 194364 42124
rect 194272 42120 194364 42122
rect 194272 42064 194322 42120
rect 194272 42062 194364 42064
rect 194317 42060 194364 42062
rect 194428 42060 194434 42124
rect 415761 42122 415827 42125
rect 421966 42122 421972 42124
rect 415761 42120 421972 42122
rect 415761 42064 415766 42120
rect 415822 42064 421972 42120
rect 415761 42062 421972 42064
rect 194317 42059 194383 42060
rect 415761 42059 415827 42062
rect 421966 42060 421972 42062
rect 422036 42060 422042 42124
rect 405641 41852 405707 41853
rect 405590 41850 405596 41852
rect 405550 41790 405596 41850
rect 405660 41848 405707 41852
rect 405702 41792 405707 41848
rect 405590 41788 405596 41790
rect 405660 41788 405707 41792
rect 405641 41787 405707 41788
rect 419901 41852 419967 41853
rect 419901 41848 419948 41852
rect 420012 41850 420018 41852
rect 419901 41792 419906 41848
rect 419901 41788 419948 41792
rect 420012 41790 420058 41850
rect 420012 41788 420018 41790
rect 419901 41787 419967 41788
rect 427770 41578 427830 42198
rect 446213 42256 461183 42258
rect 446213 42200 446218 42256
rect 446274 42200 461122 42256
rect 461178 42200 461183 42256
rect 446213 42198 461183 42200
rect 446213 42195 446279 42198
rect 461117 42195 461183 42198
rect 515397 42124 515463 42125
rect 520917 42124 520983 42125
rect 522021 42124 522087 42125
rect 526437 42124 526503 42125
rect 529565 42124 529631 42125
rect 515397 42122 515444 42124
rect 515352 42120 515444 42122
rect 515352 42064 515402 42120
rect 515352 42062 515444 42064
rect 515397 42060 515444 42062
rect 515508 42060 515514 42124
rect 520917 42122 520964 42124
rect 520872 42120 520964 42122
rect 520872 42064 520922 42120
rect 520872 42062 520964 42064
rect 520917 42060 520964 42062
rect 521028 42060 521034 42124
rect 522021 42122 522068 42124
rect 521976 42120 522068 42122
rect 521976 42064 522026 42120
rect 521976 42062 522068 42064
rect 522021 42060 522068 42062
rect 522132 42060 522138 42124
rect 526437 42122 526484 42124
rect 526392 42120 526484 42122
rect 526392 42064 526442 42120
rect 526392 42062 526484 42064
rect 526437 42060 526484 42062
rect 526548 42060 526554 42124
rect 529565 42122 529612 42124
rect 529520 42120 529612 42122
rect 529520 42064 529570 42120
rect 529520 42062 529612 42064
rect 529565 42060 529612 42062
rect 529676 42060 529682 42124
rect 515397 42059 515463 42060
rect 520917 42059 520983 42060
rect 522021 42059 522087 42060
rect 526437 42059 526503 42060
rect 529565 42059 529631 42060
rect 441838 41788 441844 41852
rect 441908 41850 441914 41852
rect 460606 41850 460612 41852
rect 441908 41790 460612 41850
rect 441908 41788 441914 41790
rect 460606 41788 460612 41790
rect 460676 41788 460682 41852
rect 446213 41578 446279 41581
rect 427770 41576 446279 41578
rect 427770 41520 446218 41576
rect 446274 41520 446279 41576
rect 427770 41518 446279 41520
rect 446213 41515 446279 41518
rect 141693 40356 141759 40357
rect 141693 40352 141740 40356
rect 141804 40354 141810 40356
rect 141693 40296 141698 40352
rect 141693 40292 141740 40296
rect 141804 40294 141850 40354
rect 141804 40292 141810 40294
rect 141693 40291 141759 40292
<< via3 >>
rect 675708 892196 675772 892260
rect 675524 887436 675588 887500
rect 676444 883416 676508 883420
rect 676444 883360 676494 883416
rect 676494 883360 676508 883416
rect 676444 883356 676508 883360
rect 676260 883280 676324 883284
rect 676260 883224 676310 883280
rect 676310 883224 676324 883280
rect 676260 883220 676324 883224
rect 675708 881860 675772 881924
rect 675156 876556 675220 876620
rect 675156 874108 675220 874172
rect 675524 873564 675588 873628
rect 676444 873564 676508 873628
rect 676260 872340 676324 872404
rect 675524 869816 675588 869820
rect 675524 869760 675574 869816
rect 675574 869760 675588 869816
rect 675524 869756 675588 869760
rect 675708 867172 675772 867236
rect 675892 865676 675956 865740
rect 676076 865404 676140 865468
rect 42012 813180 42076 813244
rect 42196 811276 42260 811340
rect 40540 805564 40604 805628
rect 40908 804748 40972 804812
rect 40724 804476 40788 804540
rect 41828 802436 41892 802500
rect 41092 800668 41156 800732
rect 40356 800532 40420 800596
rect 40908 794820 40972 794884
rect 40356 793052 40420 793116
rect 41092 792644 41156 792708
rect 41828 791556 41892 791620
rect 40724 791284 40788 791348
rect 41644 788156 41708 788220
rect 676076 788020 676140 788084
rect 41460 786796 41524 786860
rect 674420 786660 674484 786724
rect 40540 786116 40604 786180
rect 674604 784620 674668 784684
rect 675156 780540 675220 780604
rect 676812 776052 676876 776116
rect 675156 775568 675220 775572
rect 675156 775512 675170 775568
rect 675170 775512 675220 775568
rect 675156 775508 675220 775512
rect 41460 769796 41524 769860
rect 41644 766940 41708 767004
rect 40724 766532 40788 766596
rect 40540 765308 40604 765372
rect 40908 764900 40972 764964
rect 41828 757692 41892 757756
rect 40356 757284 40420 757348
rect 42012 757208 42076 757212
rect 42012 757152 42026 757208
rect 42026 757152 42076 757208
rect 42012 757148 42076 757152
rect 40908 754020 40972 754084
rect 40356 753612 40420 753676
rect 42196 753400 42260 753404
rect 42196 753344 42210 753400
rect 42210 753344 42260 753400
rect 42196 753340 42260 753344
rect 42196 750484 42260 750548
rect 42012 749728 42076 749732
rect 42012 749672 42026 749728
rect 42026 749672 42076 749728
rect 42012 749668 42076 749672
rect 40540 749396 40604 749460
rect 40724 746812 40788 746876
rect 41828 745316 41892 745380
rect 41644 744364 41708 744428
rect 41460 743684 41524 743748
rect 675340 742248 675404 742252
rect 675340 742192 675390 742248
rect 675390 742192 675404 742248
rect 675340 742188 675404 742192
rect 674236 738108 674300 738172
rect 675340 727228 675404 727292
rect 676076 726548 676140 726612
rect 41828 725792 41892 725796
rect 41828 725736 41842 725792
rect 41842 725736 41892 725792
rect 41828 725732 41892 725736
rect 673868 722392 673932 722396
rect 673868 722336 673882 722392
rect 673882 722336 673932 722392
rect 673868 722332 673932 722336
rect 41828 721924 41892 721988
rect 674052 721848 674116 721852
rect 674052 721792 674102 721848
rect 674102 721792 674116 721848
rect 674052 721788 674116 721792
rect 675340 721516 675404 721580
rect 673868 720020 673932 720084
rect 40540 718524 40604 718588
rect 40724 718252 40788 718316
rect 41828 718252 41892 718316
rect 41644 717572 41708 717636
rect 674052 717088 674116 717092
rect 674052 717032 674066 717088
rect 674066 717032 674116 717088
rect 674052 717028 674116 717032
rect 41828 716756 41892 716820
rect 42012 714640 42076 714644
rect 42012 714584 42062 714640
rect 42062 714584 42076 714640
rect 42012 714580 42076 714584
rect 40356 714172 40420 714236
rect 674420 711996 674484 712060
rect 40356 709820 40420 709884
rect 674604 709140 674668 709204
rect 675892 707508 675956 707572
rect 40724 707372 40788 707436
rect 42012 706420 42076 706484
rect 40540 704244 40604 704308
rect 41460 703564 41524 703628
rect 41828 701796 41892 701860
rect 41644 701524 41708 701588
rect 676812 701388 676876 701452
rect 675524 696824 675588 696828
rect 675524 696768 675538 696824
rect 675538 696768 675588 696824
rect 675524 696764 675588 696768
rect 673868 693228 673932 693292
rect 673868 688060 673932 688124
rect 42012 683572 42076 683636
rect 42196 682756 42260 682820
rect 674236 682348 674300 682412
rect 675524 681396 675588 681460
rect 675340 681048 675404 681052
rect 675340 680992 675390 681048
rect 675390 680992 675404 681048
rect 675340 680988 675404 680992
rect 40540 678928 40604 678992
rect 40724 678928 40788 678992
rect 41828 678268 41892 678332
rect 675156 676364 675220 676428
rect 676076 676364 676140 676428
rect 41828 672692 41892 672756
rect 42012 671604 42076 671668
rect 42012 668536 42076 668540
rect 42012 668480 42062 668536
rect 42062 668480 42076 668536
rect 42012 668476 42076 668480
rect 676812 666572 676876 666636
rect 40908 665076 40972 665140
rect 40724 663988 40788 664052
rect 40540 662764 40604 662828
rect 41644 658548 41708 658612
rect 41828 658336 41892 658340
rect 41828 658280 41842 658336
rect 41842 658280 41892 658336
rect 41828 658276 41892 658280
rect 41460 657188 41524 657252
rect 674420 652836 674484 652900
rect 675156 650176 675220 650180
rect 675156 650120 675206 650176
rect 675206 650120 675220 650176
rect 675156 650116 675220 650120
rect 677180 648620 677244 648684
rect 676812 644676 676876 644740
rect 44220 642228 44284 642292
rect 41460 640596 41524 640660
rect 40908 636516 40972 636580
rect 676076 636108 676140 636172
rect 40540 635292 40604 635356
rect 40724 634884 40788 634948
rect 676076 631348 676140 631412
rect 41644 629852 41708 629916
rect 41828 629172 41892 629236
rect 40908 623324 40972 623388
rect 40724 621964 40788 622028
rect 40540 620740 40604 620804
rect 673868 616116 673932 616180
rect 41460 615980 41524 616044
rect 41828 615436 41892 615500
rect 41828 613456 41892 613460
rect 41828 613400 41878 613456
rect 41878 613400 41892 613456
rect 41828 613396 41892 613400
rect 675892 607004 675956 607068
rect 674236 602788 674300 602852
rect 44220 599660 44284 599724
rect 43116 599252 43180 599316
rect 675892 599116 675956 599180
rect 676996 598844 677060 598908
rect 41092 596974 41156 597038
rect 43116 597000 43180 597004
rect 43116 596944 43130 597000
rect 43130 596944 43180 597000
rect 43116 596940 43180 596944
rect 41828 596396 41892 596460
rect 40540 594118 40604 594182
rect 677180 592860 677244 592924
rect 676076 592588 676140 592652
rect 674420 591228 674484 591292
rect 40724 589596 40788 589660
rect 40908 589052 40972 589116
rect 674972 586528 675036 586532
rect 674972 586472 674986 586528
rect 674986 586472 675036 586528
rect 674972 586468 675036 586472
rect 676076 586196 676140 586260
rect 40356 586060 40420 586124
rect 41828 585108 41892 585172
rect 40356 580212 40420 580276
rect 40908 577764 40972 577828
rect 676996 576404 677060 576468
rect 40724 574636 40788 574700
rect 40540 573820 40604 573884
rect 676812 572732 676876 572796
rect 41828 572188 41892 572252
rect 41644 571916 41708 571980
rect 41460 570828 41524 570892
rect 675340 561912 675404 561916
rect 675340 561856 675390 561912
rect 675390 561856 675404 561912
rect 675340 561852 675404 561856
rect 675156 559404 675220 559468
rect 41092 558724 41156 558788
rect 41092 557488 41156 557552
rect 674972 555520 675036 555524
rect 674972 555464 674986 555520
rect 674986 555464 675036 555520
rect 674972 555460 675036 555464
rect 42196 553964 42260 554028
rect 676444 553964 676508 554028
rect 41368 553348 41432 553412
rect 676996 552060 677060 552124
rect 42380 551788 42444 551852
rect 675156 550428 675220 550492
rect 674972 549476 675036 549540
rect 675340 548388 675404 548452
rect 676812 548252 676876 548316
rect 676444 547572 676508 547636
rect 674236 547300 674300 547364
rect 675892 547028 675956 547092
rect 676076 546756 676140 546820
rect 41644 546348 41708 546412
rect 42380 546348 42444 546412
rect 40908 545668 40972 545732
rect 40724 545396 40788 545460
rect 41460 542268 41524 542332
rect 675156 541240 675220 541244
rect 675156 541184 675206 541240
rect 675206 541184 675220 541240
rect 675156 541180 675220 541184
rect 675156 539608 675220 539612
rect 675156 539552 675170 539608
rect 675170 539552 675220 539608
rect 675156 539548 675220 539552
rect 40724 537236 40788 537300
rect 40908 536964 40972 537028
rect 41460 533700 41524 533764
rect 40540 532884 40604 532948
rect 41828 529892 41892 529956
rect 41828 529408 41892 529412
rect 41828 529352 41878 529408
rect 41878 529352 41892 529408
rect 41828 529348 41892 529352
rect 676812 503644 676876 503708
rect 675708 488004 675772 488068
rect 675892 483924 675956 483988
rect 677180 482522 677244 482526
rect 677180 482466 677194 482522
rect 677194 482466 677244 482522
rect 677180 482462 677244 482466
rect 673868 455228 673932 455292
rect 41828 422316 41892 422380
rect 40540 418644 40604 418708
rect 41460 415244 41524 415308
rect 41828 414836 41892 414900
rect 41644 414564 41708 414628
rect 40724 406948 40788 407012
rect 40540 403820 40604 403884
rect 41828 401976 41892 401980
rect 41828 401920 41842 401976
rect 41842 401920 41892 401976
rect 41828 401916 41892 401920
rect 677180 401236 677244 401300
rect 676812 400420 676876 400484
rect 41828 399392 41892 399396
rect 41828 399336 41842 399392
rect 41842 399336 41892 399392
rect 41828 399332 41892 399336
rect 41460 398788 41524 398852
rect 676076 398788 676140 398852
rect 676628 396748 676692 396812
rect 676444 396340 676508 396404
rect 676260 395116 676324 395180
rect 675892 392804 675956 392868
rect 675708 387636 675772 387700
rect 676628 384916 676692 384980
rect 41460 383012 41524 383076
rect 676444 382196 676508 382260
rect 40724 379340 40788 379404
rect 41644 378932 41708 378996
rect 675708 378720 675772 378724
rect 675708 378664 675758 378720
rect 675758 378664 675772 378720
rect 675708 378660 675772 378664
rect 40540 378116 40604 378180
rect 40908 377708 40972 377772
rect 676260 377300 676324 377364
rect 41828 376892 41892 376956
rect 676076 373628 676140 373692
rect 675708 373008 675772 373012
rect 675708 372952 675722 373008
rect 675722 372952 675772 373008
rect 675708 372948 675772 372952
rect 40724 365604 40788 365668
rect 40908 364244 40972 364308
rect 40540 363700 40604 363764
rect 41828 358728 41892 358732
rect 41828 358672 41878 358728
rect 41878 358672 41892 358728
rect 41828 358668 41892 358672
rect 41460 356900 41524 356964
rect 41828 355600 41892 355604
rect 41828 355544 41878 355600
rect 41878 355544 41892 355600
rect 41828 355540 41892 355544
rect 675524 354180 675588 354244
rect 675892 353908 675956 353972
rect 675708 352956 675772 353020
rect 675892 351596 675956 351660
rect 675340 347652 675404 347716
rect 676444 346564 676508 346628
rect 44220 342892 44284 342956
rect 44588 340988 44652 341052
rect 42748 340444 42812 340508
rect 676260 340308 676324 340372
rect 44404 340172 44468 340236
rect 675524 339416 675588 339420
rect 675524 339360 675538 339416
rect 675538 339360 675588 339416
rect 675524 339356 675588 339360
rect 676076 337860 676140 337924
rect 42932 337588 42996 337652
rect 40540 336908 40604 336972
rect 40724 336500 40788 336564
rect 40908 336092 40972 336156
rect 41828 335684 41892 335748
rect 676444 335276 676508 335340
rect 41460 331196 41524 331260
rect 41644 330380 41708 330444
rect 675340 327992 675404 327996
rect 675340 327936 675390 327992
rect 675390 327936 675404 327992
rect 675340 327932 675404 327936
rect 676628 325620 676692 325684
rect 41828 324864 41892 324868
rect 41828 324808 41842 324864
rect 41842 324808 41892 324864
rect 41828 324804 41892 324808
rect 40908 322764 40972 322828
rect 40724 316780 40788 316844
rect 40540 315964 40604 316028
rect 41828 315616 41892 315620
rect 41828 315560 41842 315616
rect 41842 315560 41892 315616
rect 41828 315556 41892 315560
rect 41460 313652 41524 313716
rect 42932 312700 42996 312764
rect 675892 308756 675956 308820
rect 676076 304540 676140 304604
rect 675892 302636 675956 302700
rect 676444 301608 676508 301612
rect 676444 301552 676458 301608
rect 676458 301552 676508 301608
rect 676444 301548 676508 301552
rect 676628 301472 676692 301476
rect 676628 301416 676678 301472
rect 676678 301416 676692 301472
rect 676628 301412 676692 301416
rect 44220 300052 44284 300116
rect 44404 299236 44468 299300
rect 44588 298420 44652 298484
rect 42748 297604 42812 297668
rect 674788 297392 674852 297396
rect 674788 297336 674838 297392
rect 674838 297336 674852 297392
rect 674788 297332 674852 297336
rect 675708 297332 675772 297396
rect 42012 296788 42076 296852
rect 675524 296516 675588 296580
rect 676628 295700 676692 295764
rect 41828 293116 41892 293180
rect 674788 292844 674852 292908
rect 40540 292528 40604 292592
rect 40724 292588 40788 292592
rect 40724 292532 40774 292588
rect 40774 292532 40788 292588
rect 40724 292528 40788 292532
rect 41828 292496 41892 292500
rect 41828 292440 41842 292496
rect 41842 292440 41892 292496
rect 41828 292436 41892 292440
rect 675524 292224 675588 292228
rect 675524 292168 675574 292224
rect 675574 292168 675588 292224
rect 675524 292164 675588 292168
rect 676444 290940 676508 291004
rect 676260 286996 676324 287060
rect 42012 284276 42076 284340
rect 676076 283596 676140 283660
rect 675892 282644 675956 282708
rect 675708 281616 675772 281620
rect 675708 281560 675722 281616
rect 675722 281560 675772 281616
rect 675708 281556 675772 281560
rect 40908 279788 40972 279852
rect 40724 277068 40788 277132
rect 40540 274212 40604 274276
rect 41828 272368 41892 272372
rect 41828 272312 41842 272368
rect 41842 272312 41892 272368
rect 41828 272308 41892 272312
rect 41460 270404 41524 270468
rect 42012 269104 42076 269108
rect 42012 269048 42062 269104
rect 42062 269048 42076 269104
rect 42012 269044 42076 269048
rect 675340 264148 675404 264212
rect 676996 261564 677060 261628
rect 675892 261156 675956 261220
rect 676812 260748 676876 260812
rect 675340 258028 675404 258092
rect 40540 250548 40604 250612
rect 676996 250140 677060 250204
rect 676076 249868 676140 249932
rect 40724 249732 40788 249796
rect 675340 249596 675404 249660
rect 676812 246604 676876 246668
rect 673316 246196 673380 246260
rect 42012 238036 42076 238100
rect 674236 236676 674300 236740
rect 40724 236540 40788 236604
rect 40540 229604 40604 229668
rect 674972 228984 675036 228988
rect 674972 228928 674986 228984
rect 674986 228928 675036 228984
rect 674972 228924 675036 228928
rect 674052 228788 674116 228852
rect 672580 227020 672644 227084
rect 42012 226128 42076 226132
rect 42012 226072 42026 226128
rect 42026 226072 42076 226128
rect 42012 226068 42076 226072
rect 675708 218588 675772 218652
rect 509188 217772 509252 217836
rect 510108 217832 510172 217836
rect 510108 217776 510158 217832
rect 510158 217776 510172 217832
rect 510108 217772 510172 217776
rect 522620 217832 522684 217836
rect 522620 217776 522634 217832
rect 522634 217776 522684 217832
rect 522620 217772 522684 217776
rect 571012 217832 571076 217836
rect 571012 217776 571026 217832
rect 571026 217776 571076 217832
rect 571012 217772 571076 217776
rect 571380 217832 571444 217836
rect 571380 217776 571394 217832
rect 571394 217776 571444 217832
rect 571380 217772 571444 217776
rect 574324 217772 574388 217836
rect 493732 217288 493796 217292
rect 493732 217232 493782 217288
rect 493782 217232 493796 217288
rect 493732 217228 493796 217232
rect 675892 217908 675956 217972
rect 574324 216744 574388 216748
rect 574324 216688 574374 216744
rect 574374 216688 574388 216744
rect 574324 216684 574388 216688
rect 675892 216548 675956 216612
rect 571012 216412 571076 216476
rect 571380 216140 571444 216204
rect 509188 215868 509252 215932
rect 522620 215324 522684 215388
rect 675524 211440 675588 211444
rect 675524 211384 675538 211440
rect 675538 211384 675588 211440
rect 675524 211380 675588 211384
rect 676628 211168 676692 211172
rect 676628 211112 676642 211168
rect 676642 211112 676692 211168
rect 676628 211108 676692 211112
rect 40908 207708 40972 207772
rect 42012 207300 42076 207364
rect 40540 206892 40604 206956
rect 40724 206076 40788 206140
rect 676260 204988 676324 205052
rect 672580 203008 672644 203012
rect 672580 202952 672594 203008
rect 672594 202952 672644 203008
rect 672580 202948 672644 202952
rect 676444 202676 676508 202740
rect 41644 202132 41708 202196
rect 41828 200636 41892 200700
rect 41828 195800 41892 195804
rect 41828 195744 41842 195800
rect 41842 195744 41892 195800
rect 41828 195740 41892 195744
rect 676812 195196 676876 195260
rect 42012 195120 42076 195124
rect 42012 195064 42026 195120
rect 42026 195064 42076 195120
rect 42012 195060 42076 195064
rect 676628 194516 676692 194580
rect 676076 193156 676140 193220
rect 675892 192748 675956 192812
rect 40724 191524 40788 191588
rect 675340 189076 675404 189140
rect 40540 187172 40604 187236
rect 41460 186356 41524 186420
rect 41828 186008 41892 186012
rect 41828 185952 41842 186008
rect 41842 185952 41892 186008
rect 41828 185948 41892 185952
rect 673132 182004 673196 182068
rect 673316 180236 673380 180300
rect 676812 176608 676876 176672
rect 675892 172756 675956 172820
rect 669452 170988 669516 171052
rect 675892 170308 675956 170372
rect 675340 167452 675404 167516
rect 676076 162148 676140 162212
rect 675892 161392 675956 161396
rect 675892 161336 675942 161392
rect 675942 161336 675956 161392
rect 675892 161332 675956 161336
rect 673132 161060 673196 161124
rect 675892 159972 675956 160036
rect 674420 157584 674484 157588
rect 674420 157528 674434 157584
rect 674434 157528 674484 157584
rect 674420 157524 674484 157528
rect 676444 156980 676508 157044
rect 674420 154864 674484 154868
rect 674420 154808 674470 154864
rect 674470 154808 674484 154864
rect 674420 154804 674484 154808
rect 674236 153172 674300 153236
rect 676260 150316 676324 150380
rect 676076 148412 676140 148476
rect 675340 147656 675404 147660
rect 675340 147600 675390 147656
rect 675390 147600 675404 147656
rect 675340 147596 675404 147600
rect 669452 135492 669516 135556
rect 676260 127332 676324 127396
rect 676076 126924 676140 126988
rect 676628 125700 676692 125764
rect 676444 124068 676508 124132
rect 675340 122028 675404 122092
rect 675708 117268 675772 117332
rect 674052 115772 674116 115836
rect 676260 112372 676324 112436
rect 676628 111692 676692 111756
rect 675708 111344 675772 111348
rect 675708 111288 675758 111344
rect 675758 111288 675772 111344
rect 675708 111284 675772 111288
rect 676444 110332 676508 110396
rect 676076 108156 676140 108220
rect 675340 102640 675404 102644
rect 675340 102584 675390 102640
rect 675390 102584 675404 102640
rect 675340 102580 675404 102584
rect 635780 96868 635844 96932
rect 637252 96868 637316 96932
rect 647188 96460 647252 96524
rect 633940 95916 634004 95980
rect 650316 93060 650380 93124
rect 633940 78568 634004 78572
rect 633940 78512 633954 78568
rect 633954 78512 634004 78568
rect 633940 78508 634004 78512
rect 635780 78100 635844 78164
rect 637068 77556 637132 77620
rect 462636 54980 462700 55044
rect 462636 53680 462700 53684
rect 462636 53624 462650 53680
rect 462650 53624 462700 53680
rect 462636 53620 462700 53624
rect 194364 50220 194428 50284
rect 518756 48860 518820 48924
rect 529612 48044 529676 48108
rect 515444 47772 515508 47836
rect 526484 47772 526548 47836
rect 520964 47500 521028 47564
rect 522068 47228 522132 47292
rect 458220 44372 458284 44436
rect 461348 44372 461412 44436
rect 462268 44372 462332 44436
rect 141740 43964 141804 44028
rect 518756 42800 518820 42804
rect 518756 42744 518806 42800
rect 518806 42744 518820 42800
rect 518756 42740 518820 42744
rect 194364 42120 194428 42124
rect 194364 42064 194378 42120
rect 194378 42064 194428 42120
rect 194364 42060 194428 42064
rect 421972 42060 422036 42124
rect 405596 41848 405660 41852
rect 405596 41792 405646 41848
rect 405646 41792 405660 41848
rect 405596 41788 405660 41792
rect 419948 41848 420012 41852
rect 419948 41792 419962 41848
rect 419962 41792 420012 41848
rect 419948 41788 420012 41792
rect 515444 42120 515508 42124
rect 515444 42064 515458 42120
rect 515458 42064 515508 42120
rect 515444 42060 515508 42064
rect 520964 42120 521028 42124
rect 520964 42064 520978 42120
rect 520978 42064 521028 42120
rect 520964 42060 521028 42064
rect 522068 42120 522132 42124
rect 522068 42064 522082 42120
rect 522082 42064 522132 42120
rect 522068 42060 522132 42064
rect 526484 42120 526548 42124
rect 526484 42064 526498 42120
rect 526498 42064 526548 42120
rect 526484 42060 526548 42064
rect 529612 42120 529676 42124
rect 529612 42064 529626 42120
rect 529626 42064 529676 42120
rect 529612 42060 529676 42064
rect 441844 41788 441908 41852
rect 460612 41788 460676 41852
rect 141740 40352 141804 40356
rect 141740 40296 141754 40352
rect 141754 40296 141804 40352
rect 141740 40292 141804 40296
<< metal4 >>
rect 675707 892260 675773 892261
rect 675707 892196 675708 892260
rect 675772 892196 675773 892260
rect 675707 892195 675773 892196
rect 675523 887500 675589 887501
rect 675523 887436 675524 887500
rect 675588 887436 675589 887500
rect 675523 887435 675589 887436
rect 675526 885730 675586 887435
rect 675710 886410 675770 892195
rect 675710 886350 676138 886410
rect 675526 885670 675954 885730
rect 675707 881924 675773 881925
rect 675707 881860 675708 881924
rect 675772 881860 675773 881924
rect 675707 881859 675773 881860
rect 675155 876620 675221 876621
rect 675155 876556 675156 876620
rect 675220 876556 675221 876620
rect 675155 876555 675221 876556
rect 675158 874173 675218 876555
rect 675155 874172 675221 874173
rect 675155 874108 675156 874172
rect 675220 874108 675221 874172
rect 675155 874107 675221 874108
rect 675523 873628 675589 873629
rect 675523 873564 675524 873628
rect 675588 873564 675589 873628
rect 675523 873563 675589 873564
rect 675526 869821 675586 873563
rect 675523 869820 675589 869821
rect 675523 869756 675524 869820
rect 675588 869756 675589 869820
rect 675523 869755 675589 869756
rect 675710 867237 675770 881859
rect 675707 867236 675773 867237
rect 675707 867172 675708 867236
rect 675772 867172 675773 867236
rect 675707 867171 675773 867172
rect 675894 865741 675954 885670
rect 675891 865740 675957 865741
rect 675891 865676 675892 865740
rect 675956 865676 675957 865740
rect 675891 865675 675957 865676
rect 676078 865469 676138 886350
rect 676443 883420 676509 883421
rect 676443 883356 676444 883420
rect 676508 883356 676509 883420
rect 676443 883355 676509 883356
rect 676259 883284 676325 883285
rect 676259 883220 676260 883284
rect 676324 883220 676325 883284
rect 676259 883219 676325 883220
rect 676262 872405 676322 883219
rect 676446 873629 676506 883355
rect 676443 873628 676509 873629
rect 676443 873564 676444 873628
rect 676508 873564 676509 873628
rect 676443 873563 676509 873564
rect 676259 872404 676325 872405
rect 676259 872340 676260 872404
rect 676324 872340 676325 872404
rect 676259 872339 676325 872340
rect 676075 865468 676141 865469
rect 676075 865404 676076 865468
rect 676140 865404 676141 865468
rect 676075 865403 676141 865404
rect 42011 813244 42077 813245
rect 42011 813180 42012 813244
rect 42076 813180 42077 813244
rect 42011 813179 42077 813180
rect 42014 809570 42074 813179
rect 42195 811340 42261 811341
rect 42195 811276 42196 811340
rect 42260 811276 42261 811340
rect 42195 811275 42261 811276
rect 41462 809510 42074 809570
rect 40539 805628 40605 805629
rect 40539 805564 40540 805628
rect 40604 805564 40605 805628
rect 40539 805563 40605 805564
rect 40355 800596 40421 800597
rect 40355 800532 40356 800596
rect 40420 800532 40421 800596
rect 40355 800531 40421 800532
rect 40358 793117 40418 800531
rect 40355 793116 40421 793117
rect 40355 793052 40356 793116
rect 40420 793052 40421 793116
rect 40355 793051 40421 793052
rect 40542 786181 40602 805563
rect 40907 804812 40973 804813
rect 40907 804748 40908 804812
rect 40972 804748 40973 804812
rect 40907 804747 40973 804748
rect 40723 804540 40789 804541
rect 40723 804476 40724 804540
rect 40788 804476 40789 804540
rect 40723 804475 40789 804476
rect 40726 791349 40786 804475
rect 40910 794885 40970 804747
rect 41091 800732 41157 800733
rect 41091 800668 41092 800732
rect 41156 800668 41157 800732
rect 41091 800667 41157 800668
rect 40907 794884 40973 794885
rect 40907 794820 40908 794884
rect 40972 794820 40973 794884
rect 40907 794819 40973 794820
rect 41094 792709 41154 800667
rect 41091 792708 41157 792709
rect 41091 792644 41092 792708
rect 41156 792644 41157 792708
rect 41091 792643 41157 792644
rect 40723 791348 40789 791349
rect 40723 791284 40724 791348
rect 40788 791284 40789 791348
rect 40723 791283 40789 791284
rect 41462 786861 41522 809510
rect 42198 808710 42258 811275
rect 41646 808650 42258 808710
rect 41646 788221 41706 808650
rect 41827 802500 41893 802501
rect 41827 802436 41828 802500
rect 41892 802436 41893 802500
rect 41827 802435 41893 802436
rect 41830 791621 41890 802435
rect 41827 791620 41893 791621
rect 41827 791556 41828 791620
rect 41892 791556 41893 791620
rect 41827 791555 41893 791556
rect 41643 788220 41709 788221
rect 41643 788156 41644 788220
rect 41708 788156 41709 788220
rect 41643 788155 41709 788156
rect 676075 788084 676141 788085
rect 676075 788020 676076 788084
rect 676140 788020 676141 788084
rect 676075 788019 676141 788020
rect 41459 786860 41525 786861
rect 41459 786796 41460 786860
rect 41524 786796 41525 786860
rect 41459 786795 41525 786796
rect 674419 786724 674485 786725
rect 674419 786660 674420 786724
rect 674484 786660 674485 786724
rect 674419 786659 674485 786660
rect 40539 786180 40605 786181
rect 40539 786116 40540 786180
rect 40604 786116 40605 786180
rect 40539 786115 40605 786116
rect 41459 769860 41525 769861
rect 41459 769796 41460 769860
rect 41524 769796 41525 769860
rect 41459 769795 41525 769796
rect 40723 766596 40789 766597
rect 40723 766532 40724 766596
rect 40788 766532 40789 766596
rect 40723 766531 40789 766532
rect 40539 765372 40605 765373
rect 40539 765308 40540 765372
rect 40604 765308 40605 765372
rect 40539 765307 40605 765308
rect 40355 757348 40421 757349
rect 40355 757284 40356 757348
rect 40420 757284 40421 757348
rect 40355 757283 40421 757284
rect 40358 753677 40418 757283
rect 40355 753676 40421 753677
rect 40355 753612 40356 753676
rect 40420 753612 40421 753676
rect 40355 753611 40421 753612
rect 40542 749461 40602 765307
rect 40539 749460 40605 749461
rect 40539 749396 40540 749460
rect 40604 749396 40605 749460
rect 40539 749395 40605 749396
rect 40726 746877 40786 766531
rect 40907 764964 40973 764965
rect 40907 764900 40908 764964
rect 40972 764900 40973 764964
rect 40907 764899 40973 764900
rect 40910 754085 40970 764899
rect 40907 754084 40973 754085
rect 40907 754020 40908 754084
rect 40972 754020 40973 754084
rect 40907 754019 40973 754020
rect 40723 746876 40789 746877
rect 40723 746812 40724 746876
rect 40788 746812 40789 746876
rect 40723 746811 40789 746812
rect 41462 743749 41522 769795
rect 41643 767004 41709 767005
rect 41643 766940 41644 767004
rect 41708 766940 41709 767004
rect 41643 766939 41709 766940
rect 41646 744429 41706 766939
rect 41827 757756 41893 757757
rect 41827 757692 41828 757756
rect 41892 757692 41893 757756
rect 41827 757691 41893 757692
rect 41830 745381 41890 757691
rect 42011 757212 42077 757213
rect 42011 757148 42012 757212
rect 42076 757148 42077 757212
rect 42011 757147 42077 757148
rect 42014 749733 42074 757147
rect 42195 753404 42261 753405
rect 42195 753340 42196 753404
rect 42260 753340 42261 753404
rect 42195 753339 42261 753340
rect 42198 750549 42258 753339
rect 42195 750548 42261 750549
rect 42195 750484 42196 750548
rect 42260 750484 42261 750548
rect 42195 750483 42261 750484
rect 42011 749732 42077 749733
rect 42011 749668 42012 749732
rect 42076 749668 42077 749732
rect 42011 749667 42077 749668
rect 41827 745380 41893 745381
rect 41827 745316 41828 745380
rect 41892 745316 41893 745380
rect 41827 745315 41893 745316
rect 41643 744428 41709 744429
rect 41643 744364 41644 744428
rect 41708 744364 41709 744428
rect 41643 744363 41709 744364
rect 41459 743748 41525 743749
rect 41459 743684 41460 743748
rect 41524 743684 41525 743748
rect 41459 743683 41525 743684
rect 674235 738172 674301 738173
rect 674235 738108 674236 738172
rect 674300 738108 674301 738172
rect 674235 738107 674301 738108
rect 41827 725796 41893 725797
rect 41827 725732 41828 725796
rect 41892 725732 41893 725796
rect 41827 725731 41893 725732
rect 41830 725250 41890 725731
rect 41462 725190 41890 725250
rect 40539 718588 40605 718589
rect 40539 718524 40540 718588
rect 40604 718524 40605 718588
rect 40539 718523 40605 718524
rect 40355 714236 40421 714237
rect 40355 714172 40356 714236
rect 40420 714172 40421 714236
rect 40355 714171 40421 714172
rect 40358 709885 40418 714171
rect 40355 709884 40421 709885
rect 40355 709820 40356 709884
rect 40420 709820 40421 709884
rect 40355 709819 40421 709820
rect 40542 704309 40602 718523
rect 40723 718316 40789 718317
rect 40723 718252 40724 718316
rect 40788 718252 40789 718316
rect 40723 718251 40789 718252
rect 40726 707437 40786 718251
rect 40723 707436 40789 707437
rect 40723 707372 40724 707436
rect 40788 707372 40789 707436
rect 40723 707371 40789 707372
rect 40539 704308 40605 704309
rect 40539 704244 40540 704308
rect 40604 704244 40605 704308
rect 40539 704243 40605 704244
rect 41462 703629 41522 725190
rect 673867 722396 673933 722397
rect 673867 722332 673868 722396
rect 673932 722332 673933 722396
rect 673867 722331 673933 722332
rect 41827 721988 41893 721989
rect 41827 721924 41828 721988
rect 41892 721924 41893 721988
rect 41827 721923 41893 721924
rect 41830 718317 41890 721923
rect 673870 720085 673930 722331
rect 674051 721852 674117 721853
rect 674051 721788 674052 721852
rect 674116 721788 674117 721852
rect 674051 721787 674117 721788
rect 673867 720084 673933 720085
rect 673867 720020 673868 720084
rect 673932 720020 673933 720084
rect 673867 720019 673933 720020
rect 41827 718316 41893 718317
rect 41827 718252 41828 718316
rect 41892 718252 41893 718316
rect 41827 718251 41893 718252
rect 41643 717636 41709 717637
rect 41643 717572 41644 717636
rect 41708 717572 41709 717636
rect 41643 717571 41709 717572
rect 41459 703628 41525 703629
rect 41459 703564 41460 703628
rect 41524 703564 41525 703628
rect 41459 703563 41525 703564
rect 41646 701589 41706 717571
rect 674054 717093 674114 721787
rect 674051 717092 674117 717093
rect 674051 717028 674052 717092
rect 674116 717028 674117 717092
rect 674051 717027 674117 717028
rect 41827 716820 41893 716821
rect 41827 716756 41828 716820
rect 41892 716756 41893 716820
rect 41827 716755 41893 716756
rect 41830 701861 41890 716755
rect 42011 714644 42077 714645
rect 42011 714580 42012 714644
rect 42076 714580 42077 714644
rect 42011 714579 42077 714580
rect 42014 706485 42074 714579
rect 42011 706484 42077 706485
rect 42011 706420 42012 706484
rect 42076 706420 42077 706484
rect 42011 706419 42077 706420
rect 41827 701860 41893 701861
rect 41827 701796 41828 701860
rect 41892 701796 41893 701860
rect 41827 701795 41893 701796
rect 41643 701588 41709 701589
rect 41643 701524 41644 701588
rect 41708 701524 41709 701588
rect 41643 701523 41709 701524
rect 673867 693292 673933 693293
rect 673867 693228 673868 693292
rect 673932 693228 673933 693292
rect 673867 693227 673933 693228
rect 673870 688125 673930 693227
rect 673867 688124 673933 688125
rect 673867 688060 673868 688124
rect 673932 688060 673933 688124
rect 673867 688059 673933 688060
rect 42011 683636 42077 683637
rect 42011 683572 42012 683636
rect 42076 683572 42077 683636
rect 42011 683571 42077 683572
rect 40539 678992 40605 678993
rect 40539 678928 40540 678992
rect 40604 678928 40605 678992
rect 40539 678927 40605 678928
rect 40723 678992 40789 678993
rect 40723 678928 40724 678992
rect 40788 678928 40789 678992
rect 40723 678927 40789 678928
rect 40542 662829 40602 678927
rect 40726 664053 40786 678927
rect 41827 678332 41893 678333
rect 41827 678330 41828 678332
rect 40910 678270 41828 678330
rect 40910 665141 40970 678270
rect 41827 678268 41828 678270
rect 41892 678268 41893 678332
rect 41827 678267 41893 678268
rect 42014 674930 42074 683571
rect 42195 682820 42261 682821
rect 42195 682756 42196 682820
rect 42260 682756 42261 682820
rect 42195 682755 42261 682756
rect 41462 674870 42074 674930
rect 40907 665140 40973 665141
rect 40907 665076 40908 665140
rect 40972 665076 40973 665140
rect 40907 665075 40973 665076
rect 40723 664052 40789 664053
rect 40723 663988 40724 664052
rect 40788 663988 40789 664052
rect 40723 663987 40789 663988
rect 40539 662828 40605 662829
rect 40539 662764 40540 662828
rect 40604 662764 40605 662828
rect 40539 662763 40605 662764
rect 41462 657253 41522 674870
rect 42198 674250 42258 682755
rect 674238 682413 674298 738107
rect 674422 712061 674482 786659
rect 674603 784684 674669 784685
rect 674603 784620 674604 784684
rect 674668 784620 674669 784684
rect 674603 784619 674669 784620
rect 674419 712060 674485 712061
rect 674419 711996 674420 712060
rect 674484 711996 674485 712060
rect 674419 711995 674485 711996
rect 674606 709205 674666 784619
rect 675155 780604 675221 780605
rect 675155 780540 675156 780604
rect 675220 780540 675221 780604
rect 675155 780539 675221 780540
rect 675158 775573 675218 780539
rect 675155 775572 675221 775573
rect 675155 775508 675156 775572
rect 675220 775508 675221 775572
rect 675155 775507 675221 775508
rect 675339 742252 675405 742253
rect 675339 742188 675340 742252
rect 675404 742188 675405 742252
rect 675339 742187 675405 742188
rect 675342 727293 675402 742187
rect 675339 727292 675405 727293
rect 675339 727228 675340 727292
rect 675404 727228 675405 727292
rect 675339 727227 675405 727228
rect 676078 726613 676138 788019
rect 676811 776116 676877 776117
rect 676811 776052 676812 776116
rect 676876 776052 676877 776116
rect 676811 776051 676877 776052
rect 676075 726612 676141 726613
rect 676075 726548 676076 726612
rect 676140 726548 676141 726612
rect 676075 726547 676141 726548
rect 675339 721580 675405 721581
rect 675339 721516 675340 721580
rect 675404 721516 675405 721580
rect 675339 721515 675405 721516
rect 674603 709204 674669 709205
rect 674603 709140 674604 709204
rect 674668 709140 674669 709204
rect 674603 709139 674669 709140
rect 674235 682412 674301 682413
rect 674235 682348 674236 682412
rect 674300 682348 674301 682412
rect 674235 682347 674301 682348
rect 675342 681053 675402 721515
rect 675891 707572 675957 707573
rect 675891 707508 675892 707572
rect 675956 707570 675957 707572
rect 676814 707570 676874 776051
rect 675956 707510 676874 707570
rect 675956 707508 675957 707510
rect 675891 707507 675957 707508
rect 676811 701452 676877 701453
rect 676811 701388 676812 701452
rect 676876 701388 676877 701452
rect 676811 701387 676877 701388
rect 675523 696828 675589 696829
rect 675523 696764 675524 696828
rect 675588 696764 675589 696828
rect 675523 696763 675589 696764
rect 675526 681461 675586 696763
rect 675523 681460 675589 681461
rect 675523 681396 675524 681460
rect 675588 681396 675589 681460
rect 675523 681395 675589 681396
rect 675339 681052 675405 681053
rect 675339 680988 675340 681052
rect 675404 680988 675405 681052
rect 675339 680987 675405 680988
rect 675155 676428 675221 676429
rect 675155 676364 675156 676428
rect 675220 676364 675221 676428
rect 675155 676363 675221 676364
rect 676075 676428 676141 676429
rect 676075 676364 676076 676428
rect 676140 676364 676141 676428
rect 676075 676363 676141 676364
rect 41646 674190 42258 674250
rect 41646 658613 41706 674190
rect 41827 672756 41893 672757
rect 41827 672692 41828 672756
rect 41892 672692 41893 672756
rect 41827 672691 41893 672692
rect 41643 658612 41709 658613
rect 41643 658548 41644 658612
rect 41708 658548 41709 658612
rect 41643 658547 41709 658548
rect 41830 658341 41890 672691
rect 42011 671668 42077 671669
rect 42011 671604 42012 671668
rect 42076 671604 42077 671668
rect 42011 671603 42077 671604
rect 42014 668541 42074 671603
rect 42011 668540 42077 668541
rect 42011 668476 42012 668540
rect 42076 668476 42077 668540
rect 42011 668475 42077 668476
rect 41827 658340 41893 658341
rect 41827 658276 41828 658340
rect 41892 658276 41893 658340
rect 41827 658275 41893 658276
rect 41459 657252 41525 657253
rect 41459 657188 41460 657252
rect 41524 657188 41525 657252
rect 41459 657187 41525 657188
rect 674419 652900 674485 652901
rect 674419 652836 674420 652900
rect 674484 652836 674485 652900
rect 674419 652835 674485 652836
rect 44219 642292 44285 642293
rect 44219 642228 44220 642292
rect 44284 642228 44285 642292
rect 44219 642227 44285 642228
rect 41459 640660 41525 640661
rect 41459 640596 41460 640660
rect 41524 640596 41525 640660
rect 41459 640595 41525 640596
rect 40907 636580 40973 636581
rect 40907 636516 40908 636580
rect 40972 636516 40973 636580
rect 40907 636515 40973 636516
rect 40539 635356 40605 635357
rect 40539 635292 40540 635356
rect 40604 635292 40605 635356
rect 40539 635291 40605 635292
rect 40542 620805 40602 635291
rect 40723 634948 40789 634949
rect 40723 634884 40724 634948
rect 40788 634884 40789 634948
rect 40723 634883 40789 634884
rect 40726 622029 40786 634883
rect 40910 623389 40970 636515
rect 40907 623388 40973 623389
rect 40907 623324 40908 623388
rect 40972 623324 40973 623388
rect 40907 623323 40973 623324
rect 40723 622028 40789 622029
rect 40723 621964 40724 622028
rect 40788 621964 40789 622028
rect 40723 621963 40789 621964
rect 40539 620804 40605 620805
rect 40539 620740 40540 620804
rect 40604 620740 40605 620804
rect 40539 620739 40605 620740
rect 41462 616045 41522 640595
rect 41643 629916 41709 629917
rect 41643 629852 41644 629916
rect 41708 629852 41709 629916
rect 41643 629851 41709 629852
rect 41459 616044 41525 616045
rect 41459 615980 41460 616044
rect 41524 615980 41525 616044
rect 41459 615979 41525 615980
rect 41646 615090 41706 629851
rect 41827 629236 41893 629237
rect 41827 629172 41828 629236
rect 41892 629172 41893 629236
rect 41827 629171 41893 629172
rect 41830 615501 41890 629171
rect 41827 615500 41893 615501
rect 41827 615436 41828 615500
rect 41892 615436 41893 615500
rect 41827 615435 41893 615436
rect 41646 615030 41890 615090
rect 41830 613461 41890 615030
rect 41827 613460 41893 613461
rect 41827 613396 41828 613460
rect 41892 613396 41893 613460
rect 41827 613395 41893 613396
rect 44222 599725 44282 642227
rect 673867 616180 673933 616181
rect 673867 616116 673868 616180
rect 673932 616116 673933 616180
rect 673867 616115 673933 616116
rect 44219 599724 44285 599725
rect 44219 599660 44220 599724
rect 44284 599660 44285 599724
rect 44219 599659 44285 599660
rect 43115 599316 43181 599317
rect 43115 599252 43116 599316
rect 43180 599252 43181 599316
rect 43115 599251 43181 599252
rect 41091 597038 41157 597039
rect 41091 596974 41092 597038
rect 41156 596974 41157 597038
rect 43118 597005 43178 599251
rect 41091 596973 41157 596974
rect 43115 597004 43181 597005
rect 40539 594182 40605 594183
rect 40539 594118 40540 594182
rect 40604 594118 40605 594182
rect 40539 594117 40605 594118
rect 40355 586124 40421 586125
rect 40355 586060 40356 586124
rect 40420 586060 40421 586124
rect 40355 586059 40421 586060
rect 40358 580277 40418 586059
rect 40355 580276 40421 580277
rect 40355 580212 40356 580276
rect 40420 580212 40421 580276
rect 40355 580211 40421 580212
rect 40542 573885 40602 594117
rect 41094 592514 41154 596973
rect 43115 596940 43116 597004
rect 43180 596940 43181 597004
rect 43115 596939 43181 596940
rect 41827 596460 41893 596461
rect 41827 596396 41828 596460
rect 41892 596396 41893 596460
rect 41827 596395 41893 596396
rect 41094 592454 41338 592514
rect 40723 589660 40789 589661
rect 40723 589596 40724 589660
rect 40788 589596 40789 589660
rect 40723 589595 40789 589596
rect 40726 574701 40786 589595
rect 41278 589290 41338 592454
rect 41278 589230 41522 589290
rect 40907 589116 40973 589117
rect 40907 589052 40908 589116
rect 40972 589052 40973 589116
rect 40907 589051 40973 589052
rect 40910 577829 40970 589051
rect 40907 577828 40973 577829
rect 40907 577764 40908 577828
rect 40972 577764 40973 577828
rect 40907 577763 40973 577764
rect 40723 574700 40789 574701
rect 40723 574636 40724 574700
rect 40788 574636 40789 574700
rect 40723 574635 40789 574636
rect 40539 573884 40605 573885
rect 40539 573820 40540 573884
rect 40604 573820 40605 573884
rect 40539 573819 40605 573820
rect 41462 570893 41522 589230
rect 41830 587210 41890 596395
rect 41646 587150 41890 587210
rect 41646 571981 41706 587150
rect 41827 585172 41893 585173
rect 41827 585108 41828 585172
rect 41892 585108 41893 585172
rect 41827 585107 41893 585108
rect 41830 572253 41890 585107
rect 41827 572252 41893 572253
rect 41827 572188 41828 572252
rect 41892 572188 41893 572252
rect 41827 572187 41893 572188
rect 41643 571980 41709 571981
rect 41643 571916 41644 571980
rect 41708 571916 41709 571980
rect 41643 571915 41709 571916
rect 41459 570892 41525 570893
rect 41459 570828 41460 570892
rect 41524 570828 41525 570892
rect 41459 570827 41525 570828
rect 41091 558788 41157 558789
rect 41091 558724 41092 558788
rect 41156 558724 41157 558788
rect 41091 558723 41157 558724
rect 41094 557553 41154 558723
rect 41091 557552 41157 557553
rect 41091 557488 41092 557552
rect 41156 557488 41157 557552
rect 41091 557487 41157 557488
rect 42195 554028 42261 554029
rect 42195 553964 42196 554028
rect 42260 553964 42261 554028
rect 42195 553963 42261 553964
rect 41367 553412 41433 553413
rect 41367 553348 41368 553412
rect 41432 553348 41433 553412
rect 41367 553347 41433 553348
rect 41370 553210 41430 553347
rect 40542 553150 41430 553210
rect 40542 532949 40602 553150
rect 41643 546412 41709 546413
rect 41643 546348 41644 546412
rect 41708 546348 41709 546412
rect 41643 546347 41709 546348
rect 40907 545732 40973 545733
rect 40907 545668 40908 545732
rect 40972 545668 40973 545732
rect 40907 545667 40973 545668
rect 40723 545460 40789 545461
rect 40723 545396 40724 545460
rect 40788 545396 40789 545460
rect 40723 545395 40789 545396
rect 40726 537301 40786 545395
rect 40723 537300 40789 537301
rect 40723 537236 40724 537300
rect 40788 537236 40789 537300
rect 40723 537235 40789 537236
rect 40910 537029 40970 545667
rect 41459 542332 41525 542333
rect 41459 542268 41460 542332
rect 41524 542268 41525 542332
rect 41459 542267 41525 542268
rect 40907 537028 40973 537029
rect 40907 536964 40908 537028
rect 40972 536964 40973 537028
rect 40907 536963 40973 536964
rect 41462 533765 41522 542267
rect 41459 533764 41525 533765
rect 41459 533700 41460 533764
rect 41524 533700 41525 533764
rect 41459 533699 41525 533700
rect 40539 532948 40605 532949
rect 40539 532884 40540 532948
rect 40604 532884 40605 532948
rect 40539 532883 40605 532884
rect 41646 529410 41706 546347
rect 42198 543750 42258 553963
rect 42379 551852 42445 551853
rect 42379 551788 42380 551852
rect 42444 551788 42445 551852
rect 42379 551787 42445 551788
rect 42382 546413 42442 551787
rect 42379 546412 42445 546413
rect 42379 546348 42380 546412
rect 42444 546348 42445 546412
rect 42379 546347 42445 546348
rect 41830 543690 42258 543750
rect 41830 529957 41890 543690
rect 41827 529956 41893 529957
rect 41827 529892 41828 529956
rect 41892 529892 41893 529956
rect 41827 529891 41893 529892
rect 41827 529412 41893 529413
rect 41827 529410 41828 529412
rect 41646 529350 41828 529410
rect 41827 529348 41828 529350
rect 41892 529348 41893 529412
rect 41827 529347 41893 529348
rect 673870 455293 673930 616115
rect 674235 602852 674301 602853
rect 674235 602788 674236 602852
rect 674300 602788 674301 602852
rect 674235 602787 674301 602788
rect 674238 547365 674298 602787
rect 674422 591293 674482 652835
rect 675158 650181 675218 676363
rect 675155 650180 675221 650181
rect 675155 650116 675156 650180
rect 675220 650116 675221 650180
rect 675155 650115 675221 650116
rect 676078 636173 676138 676363
rect 676814 666637 676874 701387
rect 676811 666636 676877 666637
rect 676811 666572 676812 666636
rect 676876 666572 676877 666636
rect 676811 666571 676877 666572
rect 677179 648684 677245 648685
rect 677179 648620 677180 648684
rect 677244 648620 677245 648684
rect 677179 648619 677245 648620
rect 676811 644740 676877 644741
rect 676811 644676 676812 644740
rect 676876 644676 676877 644740
rect 676811 644675 676877 644676
rect 676075 636172 676141 636173
rect 676075 636108 676076 636172
rect 676140 636108 676141 636172
rect 676075 636107 676141 636108
rect 676075 631412 676141 631413
rect 676075 631348 676076 631412
rect 676140 631348 676141 631412
rect 676075 631347 676141 631348
rect 675891 607068 675957 607069
rect 675891 607004 675892 607068
rect 675956 607004 675957 607068
rect 675891 607003 675957 607004
rect 675894 599181 675954 607003
rect 675891 599180 675957 599181
rect 675891 599116 675892 599180
rect 675956 599116 675957 599180
rect 675891 599115 675957 599116
rect 676078 592653 676138 631347
rect 676075 592652 676141 592653
rect 676075 592588 676076 592652
rect 676140 592588 676141 592652
rect 676075 592587 676141 592588
rect 674419 591292 674485 591293
rect 674419 591228 674420 591292
rect 674484 591228 674485 591292
rect 674419 591227 674485 591228
rect 674971 586532 675037 586533
rect 674971 586468 674972 586532
rect 675036 586468 675037 586532
rect 674971 586467 675037 586468
rect 674974 582390 675034 586467
rect 676075 586260 676141 586261
rect 676075 586196 676076 586260
rect 676140 586196 676141 586260
rect 676075 586195 676141 586196
rect 674974 582330 675954 582390
rect 675339 561916 675405 561917
rect 675339 561852 675340 561916
rect 675404 561852 675405 561916
rect 675339 561851 675405 561852
rect 675155 559468 675221 559469
rect 675155 559404 675156 559468
rect 675220 559404 675221 559468
rect 675155 559403 675221 559404
rect 674971 555524 675037 555525
rect 674971 555460 674972 555524
rect 675036 555460 675037 555524
rect 674971 555459 675037 555460
rect 674974 549541 675034 555459
rect 675158 550493 675218 559403
rect 675155 550492 675221 550493
rect 675155 550428 675156 550492
rect 675220 550428 675221 550492
rect 675155 550427 675221 550428
rect 674971 549540 675037 549541
rect 674971 549476 674972 549540
rect 675036 549476 675037 549540
rect 674971 549475 675037 549476
rect 675342 548453 675402 561851
rect 675339 548452 675405 548453
rect 675339 548388 675340 548452
rect 675404 548388 675405 548452
rect 675339 548387 675405 548388
rect 674235 547364 674301 547365
rect 674235 547300 674236 547364
rect 674300 547300 674301 547364
rect 674235 547299 674301 547300
rect 675894 547093 675954 582330
rect 675891 547092 675957 547093
rect 675891 547028 675892 547092
rect 675956 547028 675957 547092
rect 675891 547027 675957 547028
rect 676078 546821 676138 586195
rect 676814 572797 676874 644675
rect 676995 598908 677061 598909
rect 676995 598844 676996 598908
rect 677060 598844 677061 598908
rect 676995 598843 677061 598844
rect 676998 576469 677058 598843
rect 677182 592925 677242 648619
rect 677179 592924 677245 592925
rect 677179 592860 677180 592924
rect 677244 592860 677245 592924
rect 677179 592859 677245 592860
rect 676995 576468 677061 576469
rect 676995 576404 676996 576468
rect 677060 576404 677061 576468
rect 676995 576403 677061 576404
rect 676811 572796 676877 572797
rect 676811 572732 676812 572796
rect 676876 572732 676877 572796
rect 676811 572731 676877 572732
rect 676443 554028 676509 554029
rect 676443 553964 676444 554028
rect 676508 553964 676509 554028
rect 676443 553963 676509 553964
rect 676446 547637 676506 553963
rect 676995 552124 677061 552125
rect 676995 552060 676996 552124
rect 677060 552060 677061 552124
rect 676995 552059 677061 552060
rect 676811 548316 676877 548317
rect 676811 548252 676812 548316
rect 676876 548252 676877 548316
rect 676811 548251 676877 548252
rect 676443 547636 676509 547637
rect 676443 547572 676444 547636
rect 676508 547572 676509 547636
rect 676443 547571 676509 547572
rect 676075 546820 676141 546821
rect 676075 546756 676076 546820
rect 676140 546756 676141 546820
rect 676075 546755 676141 546756
rect 675155 541244 675221 541245
rect 675155 541180 675156 541244
rect 675220 541180 675221 541244
rect 675155 541179 675221 541180
rect 675158 539613 675218 541179
rect 675155 539612 675221 539613
rect 675155 539548 675156 539612
rect 675220 539548 675221 539612
rect 675155 539547 675221 539548
rect 676814 503709 676874 548251
rect 676811 503708 676877 503709
rect 676811 503644 676812 503708
rect 676876 503644 676877 503708
rect 676811 503643 676877 503644
rect 676998 492690 677058 552059
rect 676998 492630 677426 492690
rect 677366 491310 677426 492630
rect 675894 491250 677426 491310
rect 675707 488068 675773 488069
rect 675707 488004 675708 488068
rect 675772 488004 675773 488068
rect 675707 488003 675773 488004
rect 675710 481650 675770 488003
rect 675894 483989 675954 491250
rect 675891 483988 675957 483989
rect 675891 483924 675892 483988
rect 675956 483924 675957 483988
rect 675891 483923 675957 483924
rect 677179 482526 677245 482527
rect 677179 482462 677180 482526
rect 677244 482462 677245 482526
rect 677179 482461 677245 482462
rect 675710 481590 676690 481650
rect 676630 476130 676690 481590
rect 676630 476070 676874 476130
rect 673867 455292 673933 455293
rect 673867 455228 673868 455292
rect 673932 455228 673933 455292
rect 673867 455227 673933 455228
rect 41827 422380 41893 422381
rect 41827 422316 41828 422380
rect 41892 422316 41893 422380
rect 41827 422315 41893 422316
rect 41830 421970 41890 422315
rect 40726 421910 41890 421970
rect 40539 418708 40605 418709
rect 40539 418644 40540 418708
rect 40604 418644 40605 418708
rect 40539 418643 40605 418644
rect 40542 403885 40602 418643
rect 40726 407013 40786 421910
rect 41459 415308 41525 415309
rect 41459 415244 41460 415308
rect 41524 415244 41525 415308
rect 41459 415243 41525 415244
rect 40723 407012 40789 407013
rect 40723 406948 40724 407012
rect 40788 406948 40789 407012
rect 40723 406947 40789 406948
rect 40539 403884 40605 403885
rect 40539 403820 40540 403884
rect 40604 403820 40605 403884
rect 40539 403819 40605 403820
rect 41462 398853 41522 415243
rect 41827 414900 41893 414901
rect 41827 414836 41828 414900
rect 41892 414836 41893 414900
rect 41827 414835 41893 414836
rect 41643 414628 41709 414629
rect 41643 414564 41644 414628
rect 41708 414564 41709 414628
rect 41643 414563 41709 414564
rect 41646 400890 41706 414563
rect 41830 401981 41890 414835
rect 41827 401980 41893 401981
rect 41827 401916 41828 401980
rect 41892 401916 41893 401980
rect 41827 401915 41893 401916
rect 41646 400830 41890 400890
rect 41830 399397 41890 400830
rect 676814 400485 676874 476070
rect 677182 401301 677242 482461
rect 677179 401300 677245 401301
rect 677179 401236 677180 401300
rect 677244 401236 677245 401300
rect 677179 401235 677245 401236
rect 676811 400484 676877 400485
rect 676811 400420 676812 400484
rect 676876 400420 676877 400484
rect 676811 400419 676877 400420
rect 41827 399396 41893 399397
rect 41827 399332 41828 399396
rect 41892 399332 41893 399396
rect 41827 399331 41893 399332
rect 41459 398852 41525 398853
rect 41459 398788 41460 398852
rect 41524 398788 41525 398852
rect 41459 398787 41525 398788
rect 676075 398852 676141 398853
rect 676075 398788 676076 398852
rect 676140 398788 676141 398852
rect 676075 398787 676141 398788
rect 675891 392868 675957 392869
rect 675891 392804 675892 392868
rect 675956 392804 675957 392868
rect 675891 392803 675957 392804
rect 675707 387700 675773 387701
rect 675707 387636 675708 387700
rect 675772 387636 675773 387700
rect 675707 387635 675773 387636
rect 41459 383076 41525 383077
rect 41459 383012 41460 383076
rect 41524 383012 41525 383076
rect 41459 383011 41525 383012
rect 40723 379404 40789 379405
rect 40723 379340 40724 379404
rect 40788 379340 40789 379404
rect 40723 379339 40789 379340
rect 40539 378180 40605 378181
rect 40539 378116 40540 378180
rect 40604 378116 40605 378180
rect 40539 378115 40605 378116
rect 40542 363765 40602 378115
rect 40726 365669 40786 379339
rect 40907 377772 40973 377773
rect 40907 377708 40908 377772
rect 40972 377708 40973 377772
rect 40907 377707 40973 377708
rect 40723 365668 40789 365669
rect 40723 365604 40724 365668
rect 40788 365604 40789 365668
rect 40723 365603 40789 365604
rect 40910 364309 40970 377707
rect 40907 364308 40973 364309
rect 40907 364244 40908 364308
rect 40972 364244 40973 364308
rect 40907 364243 40973 364244
rect 40539 363764 40605 363765
rect 40539 363700 40540 363764
rect 40604 363700 40605 363764
rect 40539 363699 40605 363700
rect 41462 356965 41522 383011
rect 41643 378996 41709 378997
rect 41643 378932 41644 378996
rect 41708 378932 41709 378996
rect 41643 378931 41709 378932
rect 41646 358050 41706 378931
rect 675710 378725 675770 387635
rect 675707 378724 675773 378725
rect 675707 378660 675708 378724
rect 675772 378660 675773 378724
rect 675707 378659 675773 378660
rect 41827 376956 41893 376957
rect 41827 376892 41828 376956
rect 41892 376892 41893 376956
rect 41827 376891 41893 376892
rect 41830 358733 41890 376891
rect 675894 374010 675954 392803
rect 675710 373950 675954 374010
rect 675710 373013 675770 373950
rect 676078 373693 676138 398787
rect 676627 396812 676693 396813
rect 676627 396748 676628 396812
rect 676692 396748 676693 396812
rect 676627 396747 676693 396748
rect 676443 396404 676509 396405
rect 676443 396340 676444 396404
rect 676508 396340 676509 396404
rect 676443 396339 676509 396340
rect 676259 395180 676325 395181
rect 676259 395116 676260 395180
rect 676324 395116 676325 395180
rect 676259 395115 676325 395116
rect 676262 377365 676322 395115
rect 676446 382261 676506 396339
rect 676630 384981 676690 396747
rect 676627 384980 676693 384981
rect 676627 384916 676628 384980
rect 676692 384916 676693 384980
rect 676627 384915 676693 384916
rect 676443 382260 676509 382261
rect 676443 382196 676444 382260
rect 676508 382196 676509 382260
rect 676443 382195 676509 382196
rect 676259 377364 676325 377365
rect 676259 377300 676260 377364
rect 676324 377300 676325 377364
rect 676259 377299 676325 377300
rect 676075 373692 676141 373693
rect 676075 373628 676076 373692
rect 676140 373628 676141 373692
rect 676075 373627 676141 373628
rect 675707 373012 675773 373013
rect 675707 372948 675708 373012
rect 675772 372948 675773 373012
rect 675707 372947 675773 372948
rect 41827 358732 41893 358733
rect 41827 358668 41828 358732
rect 41892 358668 41893 358732
rect 41827 358667 41893 358668
rect 41646 357990 41890 358050
rect 41459 356964 41525 356965
rect 41459 356900 41460 356964
rect 41524 356900 41525 356964
rect 41459 356899 41525 356900
rect 41830 355605 41890 357990
rect 41827 355604 41893 355605
rect 41827 355540 41828 355604
rect 41892 355540 41893 355604
rect 41827 355539 41893 355540
rect 675523 354244 675589 354245
rect 675523 354180 675524 354244
rect 675588 354180 675589 354244
rect 675523 354179 675589 354180
rect 675339 347716 675405 347717
rect 675339 347652 675340 347716
rect 675404 347652 675405 347716
rect 675339 347651 675405 347652
rect 44219 342956 44285 342957
rect 44219 342892 44220 342956
rect 44284 342892 44285 342956
rect 44219 342891 44285 342892
rect 42747 340508 42813 340509
rect 42747 340444 42748 340508
rect 42812 340444 42813 340508
rect 42747 340443 42813 340444
rect 40539 336972 40605 336973
rect 40539 336908 40540 336972
rect 40604 336908 40605 336972
rect 40539 336907 40605 336908
rect 40542 316029 40602 336907
rect 40723 336564 40789 336565
rect 40723 336500 40724 336564
rect 40788 336500 40789 336564
rect 40723 336499 40789 336500
rect 40726 316845 40786 336499
rect 40907 336156 40973 336157
rect 40907 336092 40908 336156
rect 40972 336092 40973 336156
rect 40907 336091 40973 336092
rect 40910 322829 40970 336091
rect 41827 335748 41893 335749
rect 41827 335684 41828 335748
rect 41892 335684 41893 335748
rect 41827 335683 41893 335684
rect 41459 331260 41525 331261
rect 41459 331196 41460 331260
rect 41524 331196 41525 331260
rect 41459 331195 41525 331196
rect 40907 322828 40973 322829
rect 40907 322764 40908 322828
rect 40972 322764 40973 322828
rect 40907 322763 40973 322764
rect 40723 316844 40789 316845
rect 40723 316780 40724 316844
rect 40788 316780 40789 316844
rect 40723 316779 40789 316780
rect 40539 316028 40605 316029
rect 40539 315964 40540 316028
rect 40604 315964 40605 316028
rect 40539 315963 40605 315964
rect 41462 313717 41522 331195
rect 41643 330444 41709 330445
rect 41643 330380 41644 330444
rect 41708 330380 41709 330444
rect 41643 330379 41709 330380
rect 41646 316050 41706 330379
rect 41830 324869 41890 335683
rect 41827 324868 41893 324869
rect 41827 324804 41828 324868
rect 41892 324804 41893 324868
rect 41827 324803 41893 324804
rect 41646 315990 41890 316050
rect 41830 315621 41890 315990
rect 41827 315620 41893 315621
rect 41827 315556 41828 315620
rect 41892 315556 41893 315620
rect 41827 315555 41893 315556
rect 41459 313716 41525 313717
rect 41459 313652 41460 313716
rect 41524 313652 41525 313716
rect 41459 313651 41525 313652
rect 42750 297669 42810 340443
rect 42931 337652 42997 337653
rect 42931 337588 42932 337652
rect 42996 337588 42997 337652
rect 42931 337587 42997 337588
rect 42934 312765 42994 337587
rect 42931 312764 42997 312765
rect 42931 312700 42932 312764
rect 42996 312700 42997 312764
rect 42931 312699 42997 312700
rect 44222 300117 44282 342891
rect 44587 341052 44653 341053
rect 44587 340988 44588 341052
rect 44652 340988 44653 341052
rect 44587 340987 44653 340988
rect 44403 340236 44469 340237
rect 44403 340172 44404 340236
rect 44468 340172 44469 340236
rect 44403 340171 44469 340172
rect 44219 300116 44285 300117
rect 44219 300052 44220 300116
rect 44284 300052 44285 300116
rect 44219 300051 44285 300052
rect 44406 299301 44466 340171
rect 44403 299300 44469 299301
rect 44403 299236 44404 299300
rect 44468 299236 44469 299300
rect 44403 299235 44469 299236
rect 44590 298485 44650 340987
rect 675342 327997 675402 347651
rect 675526 339421 675586 354179
rect 675891 353972 675957 353973
rect 675891 353908 675892 353972
rect 675956 353970 675957 353972
rect 675956 353910 676506 353970
rect 675956 353908 675957 353910
rect 675891 353907 675957 353908
rect 675707 353020 675773 353021
rect 675707 352956 675708 353020
rect 675772 352956 675773 353020
rect 675707 352955 675773 352956
rect 675710 350550 675770 352955
rect 675891 351660 675957 351661
rect 675891 351596 675892 351660
rect 675956 351596 675957 351660
rect 675891 351595 675957 351596
rect 675894 351250 675954 351595
rect 675894 351190 676322 351250
rect 675710 350490 676138 350550
rect 675523 339420 675589 339421
rect 675523 339356 675524 339420
rect 675588 339356 675589 339420
rect 675523 339355 675589 339356
rect 676078 337925 676138 350490
rect 676262 340373 676322 351190
rect 676446 347790 676506 353910
rect 676446 347730 676690 347790
rect 676443 346628 676509 346629
rect 676443 346564 676444 346628
rect 676508 346564 676509 346628
rect 676443 346563 676509 346564
rect 676259 340372 676325 340373
rect 676259 340308 676260 340372
rect 676324 340308 676325 340372
rect 676259 340307 676325 340308
rect 676075 337924 676141 337925
rect 676075 337860 676076 337924
rect 676140 337860 676141 337924
rect 676075 337859 676141 337860
rect 676446 335341 676506 346563
rect 676443 335340 676509 335341
rect 676443 335276 676444 335340
rect 676508 335276 676509 335340
rect 676443 335275 676509 335276
rect 675339 327996 675405 327997
rect 675339 327932 675340 327996
rect 675404 327932 675405 327996
rect 675339 327931 675405 327932
rect 676630 325685 676690 347730
rect 676627 325684 676693 325685
rect 676627 325620 676628 325684
rect 676692 325620 676693 325684
rect 676627 325619 676693 325620
rect 675891 308820 675957 308821
rect 675891 308756 675892 308820
rect 675956 308756 675957 308820
rect 675891 308755 675957 308756
rect 675894 303650 675954 308755
rect 676075 304604 676141 304605
rect 676075 304540 676076 304604
rect 676140 304540 676141 304604
rect 676075 304539 676141 304540
rect 676078 304330 676138 304539
rect 676078 304270 676322 304330
rect 675894 303590 676138 303650
rect 675891 302700 675957 302701
rect 675891 302636 675892 302700
rect 675956 302636 675957 302700
rect 675891 302635 675957 302636
rect 44587 298484 44653 298485
rect 44587 298420 44588 298484
rect 44652 298420 44653 298484
rect 44587 298419 44653 298420
rect 42747 297668 42813 297669
rect 42747 297604 42748 297668
rect 42812 297604 42813 297668
rect 42747 297603 42813 297604
rect 674787 297396 674853 297397
rect 674787 297332 674788 297396
rect 674852 297332 674853 297396
rect 674787 297331 674853 297332
rect 675707 297396 675773 297397
rect 675707 297332 675708 297396
rect 675772 297332 675773 297396
rect 675707 297331 675773 297332
rect 42011 296852 42077 296853
rect 42011 296788 42012 296852
rect 42076 296788 42077 296852
rect 42011 296787 42077 296788
rect 40910 293390 41890 293450
rect 40539 292592 40605 292593
rect 40539 292528 40540 292592
rect 40604 292528 40605 292592
rect 40539 292527 40605 292528
rect 40723 292592 40789 292593
rect 40723 292528 40724 292592
rect 40788 292528 40789 292592
rect 40723 292527 40789 292528
rect 40542 274277 40602 292527
rect 40726 277133 40786 292527
rect 40910 279853 40970 293390
rect 41830 293181 41890 293390
rect 41827 293180 41893 293181
rect 41827 293116 41828 293180
rect 41892 293116 41893 293180
rect 41827 293115 41893 293116
rect 42014 292770 42074 296787
rect 674790 292909 674850 297331
rect 675523 296580 675589 296581
rect 675523 296516 675524 296580
rect 675588 296516 675589 296580
rect 675523 296515 675589 296516
rect 674787 292908 674853 292909
rect 674787 292844 674788 292908
rect 674852 292844 674853 292908
rect 674787 292843 674853 292844
rect 41646 292710 42074 292770
rect 41646 292590 41706 292710
rect 41462 292530 41706 292590
rect 40907 279852 40973 279853
rect 40907 279788 40908 279852
rect 40972 279788 40973 279852
rect 40907 279787 40973 279788
rect 40723 277132 40789 277133
rect 40723 277068 40724 277132
rect 40788 277068 40789 277132
rect 40723 277067 40789 277068
rect 40539 274276 40605 274277
rect 40539 274212 40540 274276
rect 40604 274212 40605 274276
rect 40539 274211 40605 274212
rect 41462 270469 41522 292530
rect 41827 292500 41893 292501
rect 41827 292436 41828 292500
rect 41892 292436 41893 292500
rect 41827 292435 41893 292436
rect 41830 272373 41890 292435
rect 675526 292229 675586 296515
rect 675523 292228 675589 292229
rect 675523 292164 675524 292228
rect 675588 292164 675589 292228
rect 675523 292163 675589 292164
rect 42011 284340 42077 284341
rect 42011 284276 42012 284340
rect 42076 284276 42077 284340
rect 42011 284275 42077 284276
rect 41827 272372 41893 272373
rect 41827 272308 41828 272372
rect 41892 272308 41893 272372
rect 41827 272307 41893 272308
rect 41459 270468 41525 270469
rect 41459 270404 41460 270468
rect 41524 270404 41525 270468
rect 41459 270403 41525 270404
rect 42014 269109 42074 284275
rect 675710 281621 675770 297331
rect 675894 282709 675954 302635
rect 676078 283661 676138 303590
rect 676262 287061 676322 304270
rect 676443 301612 676509 301613
rect 676443 301548 676444 301612
rect 676508 301548 676509 301612
rect 676443 301547 676509 301548
rect 676446 291005 676506 301547
rect 676627 301476 676693 301477
rect 676627 301412 676628 301476
rect 676692 301412 676693 301476
rect 676627 301411 676693 301412
rect 676630 295765 676690 301411
rect 676627 295764 676693 295765
rect 676627 295700 676628 295764
rect 676692 295700 676693 295764
rect 676627 295699 676693 295700
rect 676443 291004 676509 291005
rect 676443 290940 676444 291004
rect 676508 290940 676509 291004
rect 676443 290939 676509 290940
rect 676259 287060 676325 287061
rect 676259 286996 676260 287060
rect 676324 286996 676325 287060
rect 676259 286995 676325 286996
rect 676075 283660 676141 283661
rect 676075 283596 676076 283660
rect 676140 283596 676141 283660
rect 676075 283595 676141 283596
rect 675891 282708 675957 282709
rect 675891 282644 675892 282708
rect 675956 282644 675957 282708
rect 675891 282643 675957 282644
rect 675707 281620 675773 281621
rect 675707 281556 675708 281620
rect 675772 281556 675773 281620
rect 675707 281555 675773 281556
rect 42011 269108 42077 269109
rect 42011 269044 42012 269108
rect 42076 269044 42077 269108
rect 42011 269043 42077 269044
rect 675339 264212 675405 264213
rect 675339 264148 675340 264212
rect 675404 264148 675405 264212
rect 675339 264147 675405 264148
rect 675342 258093 675402 264147
rect 676995 261628 677061 261629
rect 676995 261564 676996 261628
rect 677060 261564 677061 261628
rect 676995 261563 677061 261564
rect 675891 261220 675957 261221
rect 675891 261156 675892 261220
rect 675956 261156 675957 261220
rect 675891 261155 675957 261156
rect 675339 258092 675405 258093
rect 675339 258028 675340 258092
rect 675404 258028 675405 258092
rect 675339 258027 675405 258028
rect 40539 250612 40605 250613
rect 40539 250548 40540 250612
rect 40604 250548 40605 250612
rect 40539 250547 40605 250548
rect 40542 229669 40602 250547
rect 40723 249796 40789 249797
rect 40723 249732 40724 249796
rect 40788 249732 40789 249796
rect 40723 249731 40789 249732
rect 40726 236605 40786 249731
rect 675342 249661 675402 258027
rect 675894 253950 675954 261155
rect 676811 260812 676877 260813
rect 676811 260748 676812 260812
rect 676876 260748 676877 260812
rect 676811 260747 676877 260748
rect 675894 253890 676138 253950
rect 676078 249933 676138 253890
rect 676075 249932 676141 249933
rect 676075 249868 676076 249932
rect 676140 249868 676141 249932
rect 676075 249867 676141 249868
rect 675339 249660 675405 249661
rect 675339 249596 675340 249660
rect 675404 249596 675405 249660
rect 675339 249595 675405 249596
rect 676814 246669 676874 260747
rect 676998 250205 677058 261563
rect 676995 250204 677061 250205
rect 676995 250140 676996 250204
rect 677060 250140 677061 250204
rect 676995 250139 677061 250140
rect 676811 246668 676877 246669
rect 676811 246604 676812 246668
rect 676876 246604 676877 246668
rect 676811 246603 676877 246604
rect 673315 246260 673381 246261
rect 673315 246196 673316 246260
rect 673380 246196 673381 246260
rect 673315 246195 673381 246196
rect 42011 238100 42077 238101
rect 42011 238036 42012 238100
rect 42076 238036 42077 238100
rect 42011 238035 42077 238036
rect 40723 236604 40789 236605
rect 40723 236540 40724 236604
rect 40788 236540 40789 236604
rect 40723 236539 40789 236540
rect 40539 229668 40605 229669
rect 40539 229604 40540 229668
rect 40604 229604 40605 229668
rect 40539 229603 40605 229604
rect 42014 226133 42074 238035
rect 672579 227084 672645 227085
rect 672579 227020 672580 227084
rect 672644 227020 672645 227084
rect 672579 227019 672645 227020
rect 42011 226132 42077 226133
rect 42011 226068 42012 226132
rect 42076 226068 42077 226132
rect 42011 226067 42077 226068
rect 509187 217836 509253 217837
rect 509187 217772 509188 217836
rect 509252 217772 509253 217836
rect 522619 217836 522685 217837
rect 509187 217771 509253 217772
rect 510107 217772 510108 217822
rect 510172 217772 510173 217822
rect 510107 217771 510173 217772
rect 522619 217772 522620 217836
rect 522684 217772 522685 217836
rect 522619 217771 522685 217772
rect 571011 217836 571077 217837
rect 571011 217772 571012 217836
rect 571076 217772 571077 217836
rect 571011 217771 571077 217772
rect 571379 217836 571445 217837
rect 571379 217772 571380 217836
rect 571444 217772 571445 217836
rect 571379 217771 571445 217772
rect 574323 217772 574324 217822
rect 574388 217772 574389 217822
rect 574323 217771 574389 217772
rect 509190 215933 509250 217771
rect 509187 215932 509253 215933
rect 509187 215868 509188 215932
rect 509252 215868 509253 215932
rect 509187 215867 509253 215868
rect 522622 215389 522682 217771
rect 571014 216477 571074 217771
rect 571011 216476 571077 216477
rect 571011 216412 571012 216476
rect 571076 216412 571077 216476
rect 571011 216411 571077 216412
rect 571382 216205 571442 217771
rect 574326 216749 574386 217142
rect 574323 216748 574389 216749
rect 574323 216684 574324 216748
rect 574388 216684 574389 216748
rect 574323 216683 574389 216684
rect 571379 216204 571445 216205
rect 571379 216140 571380 216204
rect 571444 216140 571445 216204
rect 571379 216139 571445 216140
rect 522619 215388 522685 215389
rect 522619 215324 522620 215388
rect 522684 215324 522685 215388
rect 522619 215323 522685 215324
rect 40907 207772 40973 207773
rect 40907 207708 40908 207772
rect 40972 207708 40973 207772
rect 40907 207707 40973 207708
rect 40539 206956 40605 206957
rect 40539 206892 40540 206956
rect 40604 206892 40605 206956
rect 40539 206891 40605 206892
rect 40542 187237 40602 206891
rect 40723 206140 40789 206141
rect 40723 206076 40724 206140
rect 40788 206076 40789 206140
rect 40723 206075 40789 206076
rect 40726 191589 40786 206075
rect 40910 195530 40970 207707
rect 42011 207364 42077 207365
rect 42011 207300 42012 207364
rect 42076 207300 42077 207364
rect 42011 207299 42077 207300
rect 41643 202196 41709 202197
rect 41643 202132 41644 202196
rect 41708 202132 41709 202196
rect 41643 202131 41709 202132
rect 40910 195470 41522 195530
rect 40723 191588 40789 191589
rect 40723 191524 40724 191588
rect 40788 191524 40789 191588
rect 40723 191523 40789 191524
rect 40539 187236 40605 187237
rect 40539 187172 40540 187236
rect 40604 187172 40605 187236
rect 40539 187171 40605 187172
rect 41462 186421 41522 195470
rect 41646 190470 41706 202131
rect 41827 200700 41893 200701
rect 41827 200636 41828 200700
rect 41892 200636 41893 200700
rect 41827 200635 41893 200636
rect 41830 195805 41890 200635
rect 41827 195804 41893 195805
rect 41827 195740 41828 195804
rect 41892 195740 41893 195804
rect 41827 195739 41893 195740
rect 42014 195125 42074 207299
rect 672582 203013 672642 227019
rect 672579 203012 672645 203013
rect 672579 202948 672580 203012
rect 672644 202948 672645 203012
rect 672579 202947 672645 202948
rect 42011 195124 42077 195125
rect 42011 195060 42012 195124
rect 42076 195060 42077 195124
rect 42011 195059 42077 195060
rect 41646 190410 41890 190470
rect 41459 186420 41525 186421
rect 41459 186356 41460 186420
rect 41524 186356 41525 186420
rect 41459 186355 41525 186356
rect 41830 186013 41890 190410
rect 41827 186012 41893 186013
rect 41827 185948 41828 186012
rect 41892 185948 41893 186012
rect 41827 185947 41893 185948
rect 673131 182068 673197 182069
rect 673131 182004 673132 182068
rect 673196 182004 673197 182068
rect 673131 182003 673197 182004
rect 669451 171052 669517 171053
rect 669451 170988 669452 171052
rect 669516 170988 669517 171052
rect 669451 170987 669517 170988
rect 669454 157350 669514 170987
rect 673134 161125 673194 182003
rect 673318 180301 673378 246195
rect 674235 236740 674301 236741
rect 674235 236676 674236 236740
rect 674300 236676 674301 236740
rect 674235 236675 674301 236676
rect 674051 228852 674117 228853
rect 674051 228788 674052 228852
rect 674116 228788 674117 228852
rect 674051 228787 674117 228788
rect 673315 180300 673381 180301
rect 673315 180236 673316 180300
rect 673380 180236 673381 180300
rect 673315 180235 673381 180236
rect 673131 161124 673197 161125
rect 673131 161060 673132 161124
rect 673196 161060 673197 161124
rect 673131 161059 673197 161060
rect 669270 157290 669514 157350
rect 669270 138030 669330 157290
rect 669270 137970 669514 138030
rect 669454 135557 669514 137970
rect 669451 135556 669517 135557
rect 669451 135492 669452 135556
rect 669516 135492 669517 135556
rect 669451 135491 669517 135492
rect 674054 115837 674114 228787
rect 674238 153237 674298 236675
rect 674971 228988 675037 228989
rect 674971 228924 674972 228988
rect 675036 228924 675037 228988
rect 674971 228923 675037 228924
rect 674974 224970 675034 228923
rect 674974 224910 675402 224970
rect 675342 189141 675402 224910
rect 675707 218652 675773 218653
rect 675707 218588 675708 218652
rect 675772 218588 675773 218652
rect 675707 218587 675773 218588
rect 675523 211444 675589 211445
rect 675523 211380 675524 211444
rect 675588 211380 675589 211444
rect 675523 211379 675589 211380
rect 675526 205650 675586 211379
rect 675710 210490 675770 218587
rect 675891 217972 675957 217973
rect 675891 217908 675892 217972
rect 675956 217970 675957 217972
rect 675956 217910 676322 217970
rect 675956 217908 675957 217910
rect 675891 217907 675957 217908
rect 676262 217290 676322 217910
rect 676262 217230 676506 217290
rect 675891 216612 675957 216613
rect 675891 216548 675892 216612
rect 675956 216610 675957 216612
rect 675956 216550 676322 216610
rect 675956 216548 675957 216550
rect 675891 216547 675957 216548
rect 675710 210430 676138 210490
rect 675526 205590 675954 205650
rect 675894 192813 675954 205590
rect 676078 193221 676138 210430
rect 676262 205053 676322 216550
rect 676259 205052 676325 205053
rect 676259 204988 676260 205052
rect 676324 204988 676325 205052
rect 676259 204987 676325 204988
rect 676446 202741 676506 217230
rect 676627 211172 676693 211173
rect 676627 211108 676628 211172
rect 676692 211108 676693 211172
rect 676627 211107 676693 211108
rect 676443 202740 676509 202741
rect 676443 202676 676444 202740
rect 676508 202676 676509 202740
rect 676443 202675 676509 202676
rect 676630 194581 676690 211107
rect 676811 195260 676877 195261
rect 676811 195196 676812 195260
rect 676876 195196 676877 195260
rect 676811 195195 676877 195196
rect 676627 194580 676693 194581
rect 676627 194516 676628 194580
rect 676692 194516 676693 194580
rect 676627 194515 676693 194516
rect 676075 193220 676141 193221
rect 676075 193156 676076 193220
rect 676140 193156 676141 193220
rect 676075 193155 676141 193156
rect 675891 192812 675957 192813
rect 675891 192748 675892 192812
rect 675956 192748 675957 192812
rect 675891 192747 675957 192748
rect 675339 189140 675405 189141
rect 675339 189076 675340 189140
rect 675404 189076 675405 189140
rect 675339 189075 675405 189076
rect 676814 176673 676874 195195
rect 676811 176672 676877 176673
rect 676811 176608 676812 176672
rect 676876 176608 676877 176672
rect 676811 176607 676877 176608
rect 675891 172820 675957 172821
rect 675891 172756 675892 172820
rect 675956 172756 675957 172820
rect 675891 172755 675957 172756
rect 675894 172410 675954 172755
rect 675894 172350 676506 172410
rect 675891 170372 675957 170373
rect 675891 170308 675892 170372
rect 675956 170370 675957 170372
rect 675956 170310 676322 170370
rect 675956 170308 675957 170310
rect 675891 170307 675957 170308
rect 675339 167516 675405 167517
rect 675339 167452 675340 167516
rect 675404 167452 675405 167516
rect 675339 167451 675405 167452
rect 674419 157588 674485 157589
rect 674419 157524 674420 157588
rect 674484 157524 674485 157588
rect 674419 157523 674485 157524
rect 674422 154869 674482 157523
rect 674419 154868 674485 154869
rect 674419 154804 674420 154868
rect 674484 154804 674485 154868
rect 674419 154803 674485 154804
rect 674235 153236 674301 153237
rect 674235 153172 674236 153236
rect 674300 153172 674301 153236
rect 674235 153171 674301 153172
rect 675342 147661 675402 167451
rect 676075 162212 676141 162213
rect 676075 162148 676076 162212
rect 676140 162148 676141 162212
rect 676075 162147 676141 162148
rect 675891 161396 675957 161397
rect 675891 161332 675892 161396
rect 675956 161332 675957 161396
rect 675891 161331 675957 161332
rect 675894 160037 675954 161331
rect 675891 160036 675957 160037
rect 675891 159972 675892 160036
rect 675956 159972 675957 160036
rect 675891 159971 675957 159972
rect 676078 148477 676138 162147
rect 676262 150381 676322 170310
rect 676446 157045 676506 172350
rect 676443 157044 676509 157045
rect 676443 156980 676444 157044
rect 676508 156980 676509 157044
rect 676443 156979 676509 156980
rect 676259 150380 676325 150381
rect 676259 150316 676260 150380
rect 676324 150316 676325 150380
rect 676259 150315 676325 150316
rect 676075 148476 676141 148477
rect 676075 148412 676076 148476
rect 676140 148412 676141 148476
rect 676075 148411 676141 148412
rect 675339 147660 675405 147661
rect 675339 147596 675340 147660
rect 675404 147596 675405 147660
rect 675339 147595 675405 147596
rect 676259 127396 676325 127397
rect 676259 127332 676260 127396
rect 676324 127332 676325 127396
rect 676259 127331 676325 127332
rect 676075 126988 676141 126989
rect 676075 126924 676076 126988
rect 676140 126924 676141 126988
rect 676075 126923 676141 126924
rect 675339 122092 675405 122093
rect 675339 122028 675340 122092
rect 675404 122028 675405 122092
rect 675339 122027 675405 122028
rect 674051 115836 674117 115837
rect 674051 115772 674052 115836
rect 674116 115772 674117 115836
rect 674051 115771 674117 115772
rect 675342 102645 675402 122027
rect 675707 117332 675773 117333
rect 675707 117268 675708 117332
rect 675772 117268 675773 117332
rect 675707 117267 675773 117268
rect 675710 111349 675770 117267
rect 675707 111348 675773 111349
rect 675707 111284 675708 111348
rect 675772 111284 675773 111348
rect 675707 111283 675773 111284
rect 676078 108221 676138 126923
rect 676262 112437 676322 127331
rect 676627 125764 676693 125765
rect 676627 125700 676628 125764
rect 676692 125700 676693 125764
rect 676627 125699 676693 125700
rect 676443 124132 676509 124133
rect 676443 124068 676444 124132
rect 676508 124068 676509 124132
rect 676443 124067 676509 124068
rect 676259 112436 676325 112437
rect 676259 112372 676260 112436
rect 676324 112372 676325 112436
rect 676259 112371 676325 112372
rect 676446 110397 676506 124067
rect 676630 111757 676690 125699
rect 676627 111756 676693 111757
rect 676627 111692 676628 111756
rect 676692 111692 676693 111756
rect 676627 111691 676693 111692
rect 676443 110396 676509 110397
rect 676443 110332 676444 110396
rect 676508 110332 676509 110396
rect 676443 110331 676509 110332
rect 676075 108220 676141 108221
rect 676075 108156 676076 108220
rect 676140 108156 676141 108220
rect 676075 108155 676141 108156
rect 675339 102644 675405 102645
rect 675339 102580 675340 102644
rect 675404 102580 675405 102644
rect 675339 102579 675405 102580
rect 635779 96932 635845 96933
rect 635779 96868 635780 96932
rect 635844 96868 635845 96932
rect 635779 96867 635845 96868
rect 637251 96932 637317 96933
rect 637251 96868 637252 96932
rect 637316 96868 637317 96932
rect 637251 96867 637317 96868
rect 633939 95980 634005 95981
rect 633939 95916 633940 95980
rect 634004 95916 634005 95980
rect 633939 95915 634005 95916
rect 633942 78573 634002 95915
rect 633939 78572 634005 78573
rect 633939 78508 633940 78572
rect 634004 78508 634005 78572
rect 633939 78507 634005 78508
rect 635782 78165 635842 96867
rect 637254 84210 637314 96867
rect 647187 96524 647253 96525
rect 647187 96460 647188 96524
rect 647252 96460 647253 96524
rect 647187 96459 647253 96460
rect 647190 94298 647250 96459
rect 650318 93125 650378 93382
rect 650315 93124 650381 93125
rect 650315 93060 650316 93124
rect 650380 93060 650381 93124
rect 650315 93059 650381 93060
rect 637070 84150 637314 84210
rect 635779 78164 635845 78165
rect 635779 78100 635780 78164
rect 635844 78100 635845 78164
rect 635779 78099 635845 78100
rect 637070 77621 637130 84150
rect 637067 77620 637133 77621
rect 637067 77556 637068 77620
rect 637132 77556 637133 77620
rect 637067 77555 637133 77556
rect 462635 55044 462701 55045
rect 462635 54980 462636 55044
rect 462700 54980 462701 55044
rect 462635 54979 462701 54980
rect 462638 53685 462698 54979
rect 462635 53684 462701 53685
rect 462635 53620 462636 53684
rect 462700 53620 462701 53684
rect 462635 53619 462701 53620
rect 194363 50284 194429 50285
rect 194363 50220 194364 50284
rect 194428 50220 194429 50284
rect 194363 50219 194429 50220
rect 141739 44028 141805 44029
rect 141739 43964 141740 44028
rect 141804 43964 141805 44028
rect 141739 43963 141805 43964
rect 141742 40357 141802 43963
rect 194366 42125 194426 50219
rect 518755 48924 518821 48925
rect 518755 48860 518756 48924
rect 518820 48860 518821 48924
rect 518755 48859 518821 48860
rect 515443 47836 515509 47837
rect 515443 47772 515444 47836
rect 515508 47772 515509 47836
rect 515443 47771 515509 47772
rect 458219 44436 458285 44437
rect 458219 44372 458220 44436
rect 458284 44372 458285 44436
rect 458219 44371 458285 44372
rect 461347 44436 461413 44437
rect 461347 44372 461348 44436
rect 461412 44372 461413 44436
rect 461347 44371 461413 44372
rect 462267 44436 462333 44437
rect 462267 44372 462268 44436
rect 462332 44372 462333 44436
rect 462267 44371 462333 44372
rect 194363 42124 194429 42125
rect 194363 42060 194364 42124
rect 194428 42060 194429 42124
rect 194363 42059 194429 42060
rect 421971 42124 422037 42125
rect 421971 42060 421972 42124
rect 422036 42060 422037 42124
rect 421971 42059 422037 42060
rect 405595 41852 405661 41853
rect 405595 41788 405596 41852
rect 405660 41788 405661 41852
rect 405595 41787 405661 41788
rect 421974 41850 422034 42059
rect 421974 41790 422162 41850
rect 405598 40578 405658 41787
rect 441843 41852 441909 41853
rect 441843 41850 441844 41852
rect 441626 41790 441844 41850
rect 441843 41788 441844 41790
rect 441908 41788 441909 41852
rect 441843 41787 441909 41788
rect 458222 40578 458282 44371
rect 461350 41938 461410 44371
rect 462270 41938 462330 44371
rect 515446 42125 515506 47771
rect 518758 42805 518818 48859
rect 529611 48108 529677 48109
rect 529611 48044 529612 48108
rect 529676 48044 529677 48108
rect 529611 48043 529677 48044
rect 526483 47836 526549 47837
rect 526483 47772 526484 47836
rect 526548 47772 526549 47836
rect 526483 47771 526549 47772
rect 520963 47564 521029 47565
rect 520963 47500 520964 47564
rect 521028 47500 521029 47564
rect 520963 47499 521029 47500
rect 518755 42804 518821 42805
rect 518755 42740 518756 42804
rect 518820 42740 518821 42804
rect 518755 42739 518821 42740
rect 520966 42125 521026 47499
rect 522067 47292 522133 47293
rect 522067 47228 522068 47292
rect 522132 47228 522133 47292
rect 522067 47227 522133 47228
rect 522070 42125 522130 47227
rect 526486 42125 526546 47771
rect 529614 42125 529674 48043
rect 515443 42124 515509 42125
rect 515443 42060 515444 42124
rect 515508 42060 515509 42124
rect 515443 42059 515509 42060
rect 520963 42124 521029 42125
rect 520963 42060 520964 42124
rect 521028 42060 521029 42124
rect 520963 42059 521029 42060
rect 522067 42124 522133 42125
rect 522067 42060 522068 42124
rect 522132 42060 522133 42124
rect 522067 42059 522133 42060
rect 526483 42124 526549 42125
rect 526483 42060 526484 42124
rect 526548 42060 526549 42124
rect 526483 42059 526549 42060
rect 529611 42124 529677 42125
rect 529611 42060 529612 42124
rect 529676 42060 529677 42124
rect 529611 42059 529677 42060
rect 460611 41852 460677 41853
rect 460611 41788 460612 41852
rect 460676 41850 460677 41852
rect 460676 41790 460802 41850
rect 460676 41788 460677 41790
rect 460611 41787 460677 41788
rect 141739 40356 141805 40357
rect 141739 40292 141740 40356
rect 141804 40292 141805 40356
rect 141739 40291 141805 40292
<< via4 >>
rect 510022 217836 510258 218058
rect 510022 217822 510108 217836
rect 510108 217822 510172 217836
rect 510172 217822 510258 217836
rect 574238 217836 574474 218058
rect 574238 217822 574324 217836
rect 574324 217822 574388 217836
rect 574388 217822 574474 217836
rect 493646 217292 493882 217378
rect 493646 217228 493732 217292
rect 493732 217228 493796 217292
rect 493796 217228 493882 217292
rect 493646 217142 493882 217228
rect 574238 217142 574474 217378
rect 647102 94062 647338 94298
rect 650230 93382 650466 93618
rect 419862 41852 420098 41938
rect 419862 41788 419948 41852
rect 419948 41788 420012 41852
rect 420012 41788 420098 41852
rect 419862 41702 420098 41788
rect 422162 41702 422398 41938
rect 441390 41702 441626 41938
rect 460802 41702 461038 41938
rect 461262 41702 461498 41938
rect 462182 41702 462418 41938
rect 405510 40342 405746 40578
rect 458134 40342 458370 40578
<< metal5 >>
rect 78610 1018624 90778 1030789
rect 130010 1018624 142178 1030789
rect 181410 1018624 193578 1030789
rect 231810 1018624 243978 1030789
rect 284410 1018624 296578 1030789
rect 334810 1018624 346978 1030789
rect 386210 1018624 398378 1030789
rect 475210 1018624 487378 1030789
rect 526610 1018624 538778 1030789
rect 577010 1018624 589178 1030789
rect 628410 1018624 640578 1030789
rect 6811 956610 18976 968778
rect 698624 953022 710789 965190
rect 6167 914054 19620 924934
rect 697980 909666 711433 920546
rect 6811 871210 18976 883378
rect 698512 863640 711002 876160
rect 6811 829010 18976 841178
rect 698624 819822 710789 831990
rect 6598 786640 19088 799160
rect 698512 774440 711002 786960
rect 6598 743440 19088 755960
rect 698512 729440 711002 741960
rect 6598 700240 19088 712760
rect 698512 684440 711002 696960
rect 6598 657040 19088 669560
rect 698512 639240 711002 651760
rect 6598 613840 19088 626360
rect 698512 594240 711002 606760
rect 6598 570640 19088 583160
rect 698512 549040 711002 561560
rect 6598 527440 19088 539960
rect 698624 505222 710789 517390
rect 6811 484410 18976 496578
rect 697980 461866 711433 472746
rect 6167 442854 19620 453734
rect 698624 417022 710789 429190
rect 6598 399840 19088 412360
rect 698512 371840 711002 384360
rect 6598 356640 19088 369160
rect 698512 326640 711002 339160
rect 6598 313440 19088 325960
rect 6598 270240 19088 282760
rect 698512 281640 711002 294160
rect 6598 227040 19088 239560
rect 698512 236640 711002 249160
rect 509980 218058 574516 218100
rect 509980 217822 510022 218058
rect 510258 217822 574238 218058
rect 574474 217822 574516 218058
rect 509980 217780 574516 217822
rect 493604 217378 574516 217420
rect 493604 217142 493646 217378
rect 493882 217142 574238 217378
rect 574474 217142 574516 217378
rect 493604 217100 574516 217142
rect 6598 183840 19088 196360
rect 698512 191440 711002 203960
rect 698512 146440 711002 158960
rect 6811 111610 18976 123778
rect 698512 101240 711002 113760
rect 647060 94298 647748 94340
rect 647060 94062 647102 94298
rect 647338 94062 647748 94298
rect 647060 94020 647748 94062
rect 647428 93660 647748 94020
rect 647428 93618 650508 93660
rect 647428 93382 650230 93618
rect 650466 93382 650508 93618
rect 647428 93340 650508 93382
rect 6167 70054 19620 80934
rect 419820 41938 421796 41980
rect 419820 41702 419862 41938
rect 420098 41702 421796 41938
rect 419820 41660 421796 41702
rect 422120 41938 441668 41980
rect 422120 41702 422162 41938
rect 422398 41702 441390 41938
rect 441626 41702 441668 41938
rect 422120 41660 441668 41702
rect 442084 41660 450684 41980
rect 421476 41300 421796 41660
rect 442084 41300 442404 41660
rect 421476 40980 442404 41300
rect 450364 41300 450684 41660
rect 451100 41660 460436 41980
rect 460760 41938 461540 41980
rect 460760 41702 460802 41938
rect 461038 41702 461262 41938
rect 461498 41702 461540 41938
rect 460760 41660 461540 41702
rect 461956 41938 462460 41980
rect 461956 41702 462182 41938
rect 462418 41702 462460 41938
rect 461956 41660 462460 41702
rect 451100 41300 451420 41660
rect 450364 40980 451420 41300
rect 460116 41300 460436 41660
rect 461956 41300 462276 41660
rect 460116 40980 462276 41300
rect 405468 40578 458412 40620
rect 405468 40342 405510 40578
rect 405746 40342 458134 40578
rect 458370 40342 458412 40578
rect 405468 40300 458412 40342
rect 80222 6811 92390 18976
rect 136713 7143 144150 18309
rect 187640 6598 200160 19088
rect 243266 6167 254146 19620
rect 296240 6598 308760 19088
rect 351040 6598 363560 19088
rect 405840 6598 418360 19088
rect 460640 6598 473160 19088
rect 515440 6598 527960 19088
rect 570422 6811 582590 18976
rect 624222 6811 636390 18976
use caravan_logo  caravan_logo
timestamp 1636751500
transform 1 0 255300 0 1 6032
box 2240 2560 37000 11520
use caravan_motto  caravan_motto
timestamp 1637698689
transform 1 0 -54560 0 1 -52
box 367960 10204 399802 14768
use caravan_power_routing  caravan_power_routing
timestamp 1666269678
transform 1 0 0 0 1 0
box 6022 30806 711814 997678
use caravan_signal_routing  caravan_signal_routing
timestamp 1666277172
transform 1 0 0 0 1 0
box 39764 415548 677806 997846
use caravel_clocking  clock_ctrl
timestamp 1666097791
transform 1 0 626764 0 1 55284
box 136 496 20000 20000
use copyright_block_a  copyright_block_a
timestamp 1665519472
transform 1 0 149582 0 1 16298
box -262 -10162 35048 2764
use buff_flash_clkrst  flash_clkrst_buffers
timestamp 1665682149
transform 1 0 458400 0 1 47600
box 330 0 7699 5000
use gpio_control_block  gpio_control_bidir_1\[0\]
timestamp 1666126335
transform -1 0 710203 0 1 121000
box 872 416 34000 13000
use gpio_control_block  gpio_control_bidir_1\[1\]
timestamp 1666126335
transform -1 0 710203 0 1 166200
box 872 416 34000 13000
use gpio_control_block  gpio_control_bidir_2\[0\]
timestamp 1666126335
transform 1 0 7631 0 1 289000
box 872 416 34000 13000
use gpio_control_block  gpio_control_bidir_2\[1\]
timestamp 1666126335
transform 1 0 7631 0 1 245800
box 872 416 34000 13000
use gpio_control_block  gpio_control_bidir_2\[2\]
timestamp 1666126335
transform 1 0 7631 0 1 202600
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[0\]
timestamp 1666126335
transform -1 0 710203 0 1 523800
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[1\]
timestamp 1666126335
transform -1 0 710203 0 1 568800
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[2\]
timestamp 1666126335
transform -1 0 710203 0 1 614000
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[3\]
timestamp 1666126335
transform -1 0 710203 0 1 659000
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[4\]
timestamp 1666126335
transform -1 0 710203 0 1 704200
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[5\]
timestamp 1666126335
transform -1 0 710203 0 1 884800
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[0\]
timestamp 1666126335
transform -1 0 710203 0 1 211200
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[1\]
timestamp 1666126335
transform -1 0 710203 0 1 256400
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[2\]
timestamp 1666126335
transform -1 0 710203 0 1 301400
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[3\]
timestamp 1666126335
transform -1 0 710203 0 1 346400
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[4\]
timestamp 1666126335
transform -1 0 710203 0 1 391600
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[5\]
timestamp 1666126335
transform -1 0 710203 0 1 479800
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[0\]
timestamp 1666126335
transform 1 0 7631 0 1 805400
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[1\]
timestamp 1666126335
transform 1 0 7631 0 1 762200
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[2\]
timestamp 1666126335
transform 1 0 7631 0 1 719000
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[3\]
timestamp 1666126335
transform 1 0 7631 0 1 675800
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[4\]
timestamp 1666126335
transform 1 0 7631 0 1 632600
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[5\]
timestamp 1666126335
transform 1 0 7631 0 1 589400
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[6\]
timestamp 1666126335
transform 1 0 7631 0 1 546200
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[7\]
timestamp 1666126335
transform 1 0 7631 0 1 418600
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[8\]
timestamp 1666126335
transform 1 0 7631 0 1 375400
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[9\]
timestamp 1666126335
transform 1 0 7631 0 1 332200
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_0
timestamp 1638587925
transform -1 0 709467 0 1 134000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_1
timestamp 1638587925
transform -1 0 709467 0 1 179200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_2
timestamp 1638587925
transform -1 0 709467 0 1 224200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_3
timestamp 1638587925
transform -1 0 709467 0 1 269400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_4
timestamp 1638587925
transform -1 0 709467 0 1 314400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_5
timestamp 1638587925
transform -1 0 709467 0 1 359400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_6
timestamp 1638587925
transform -1 0 709467 0 1 404600
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_7
timestamp 1638587925
transform -1 0 709467 0 1 492800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_8
timestamp 1638587925
transform -1 0 709467 0 1 536800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_9
timestamp 1638587925
transform -1 0 709467 0 1 581800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_10
timestamp 1638587925
transform -1 0 709467 0 1 627000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_11
timestamp 1638587925
transform -1 0 709467 0 1 672000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_12
timestamp 1638587925
transform -1 0 709467 0 1 717200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_13
timestamp 1638587925
transform -1 0 709467 0 1 897800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_25
timestamp 1638587925
transform 1 0 8367 0 1 818400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_26
timestamp 1638587925
transform 1 0 8367 0 1 775200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_27
timestamp 1638587925
transform 1 0 8367 0 1 732000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_28
timestamp 1638587925
transform 1 0 8367 0 1 688800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_29
timestamp 1638587925
transform 1 0 8367 0 1 645600
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_30
timestamp 1638587925
transform 1 0 8367 0 1 602400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_31
timestamp 1638587925
transform 1 0 8367 0 1 559200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_32
timestamp 1638587925
transform 1 0 8367 0 1 431600
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_33
timestamp 1638587925
transform 1 0 8367 0 1 388400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_34
timestamp 1638587925
transform 1 0 8367 0 1 345200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_35
timestamp 1638587925
transform 1 0 8367 0 1 302000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_36
timestamp 1638587925
transform 1 0 8367 0 1 258800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_37
timestamp 1638587925
transform 1 0 8367 0 1 215600
box -38 0 6018 2224
use housekeeping  housekeeping
timestamp 1666084955
transform 1 0 592434 0 1 100002
box 0 0 74046 110190
use mgmt_protect  mgmt_buffers
timestamp 1666114774
transform 1 0 128180 0 1 232036
box 1066 -400 424400 32400
use user_analog_project_wrapper  mprj
timestamp 1632839657
transform 1 0 65308 0 1 278718
box -800 -800 584800 704800
use open_source  open_source
timestamp 1666123577
transform 1 0 206074 0 1 2336
box 752 5164 29030 16242
use chip_io_alt  padframe
timestamp 1666101961
transform 1 0 0 0 1 0
box 0 0 717600 1037600
use digital_pll  pll
timestamp 1666101174
transform 1 0 628146 0 1 80944
box 0 0 20000 15000
use simple_por  por
timestamp 1650914729
transform 1 0 650146 0 -1 55282
box -52 -62 11344 8684
use xres_buf  rstb_level
timestamp 1649268499
transform -1 0 145710 0 -1 50488
box 374 -400 3540 3800
use gpio_signal_buffering_alt  sigbuf
timestamp 1666028682
transform 1 0 0 0 1 0
box 40023 41960 677583 728321
use mgmt_core_wrapper  soc
timestamp 1665963385
transform 1 0 52034 0 1 53002
box -156 0 524096 164000
use spare_logic_block  spare_logic\[0\]
timestamp 1638030917
transform 1 0 88632 0 1 232528
box 0 0 9000 9000
use spare_logic_block  spare_logic\[1\]
timestamp 1638030917
transform 1 0 108632 0 1 232528
box 0 0 9000 9000
use spare_logic_block  spare_logic\[2\]
timestamp 1638030917
transform 1 0 640874 0 1 220592
box 0 0 9000 9000
use spare_logic_block  spare_logic\[3\]
timestamp 1638030917
transform 1 0 578632 0 1 232528
box 0 0 9000 9000
use user_id_textblock  user_id_textblock
timestamp 1608324878
transform 1 0 96272 0 1 6890
box -656 1508 33720 10344
use user_id_programming  user_id_value
timestamp 1650371074
transform 1 0 656624 0 1 88126
box 0 0 7109 7077
<< labels >>
flabel metal5 s 187640 6598 200160 19088 0 FreeSans 16000 0 0 0 clock
port 0 nsew signal input
flabel metal5 s 351040 6598 363560 19088 0 FreeSans 16000 0 0 0 flash_clk
port 1 nsew signal tristate
flabel metal5 s 296240 6598 308760 19088 0 FreeSans 16000 0 0 0 flash_csb
port 2 nsew signal tristate
flabel metal5 s 405840 6598 418360 19088 0 FreeSans 16000 0 0 0 flash_io0
port 3 nsew signal tristate
flabel metal5 s 460640 6598 473160 19088 0 FreeSans 16000 0 0 0 flash_io1
port 4 nsew signal tristate
flabel metal5 s 515440 6598 527960 19088 0 FreeSans 16000 0 0 0 gpio
port 5 nsew signal bidirectional
flabel metal5 s 698512 101240 711002 113760 0 FreeSans 16000 0 0 0 mprj_io[0]
port 6 nsew signal bidirectional
flabel metal5 s 698512 684440 711002 696960 0 FreeSans 16000 0 0 0 mprj_io[10]
port 7 nsew signal bidirectional
flabel metal5 s 698512 729440 711002 741960 0 FreeSans 16000 0 0 0 mprj_io[11]
port 8 nsew signal bidirectional
flabel metal5 s 698512 774440 711002 786960 0 FreeSans 16000 0 0 0 mprj_io[12]
port 9 nsew signal bidirectional
flabel metal5 s 698512 863640 711002 876160 0 FreeSans 16000 0 0 0 mprj_io[13]
port 10 nsew signal bidirectional
flabel metal5 s 698624 953022 710789 965190 0 FreeSans 16000 0 0 0 mprj_io[14]
port 11 nsew signal bidirectional
flabel metal5 s 628410 1018624 640578 1030789 0 FreeSans 16000 0 0 0 mprj_io[15]
port 12 nsew signal bidirectional
flabel metal5 s 526610 1018624 538778 1030789 0 FreeSans 16000 0 0 0 mprj_io[16]
port 13 nsew signal bidirectional
flabel metal5 s 475210 1018624 487378 1030789 0 FreeSans 16000 0 0 0 mprj_io[17]
port 14 nsew signal bidirectional
flabel metal5 s 386210 1018624 398378 1030789 0 FreeSans 16000 0 0 0 mprj_io[18]
port 15 nsew signal bidirectional
flabel metal5 s 284410 1018624 296578 1030789 0 FreeSans 16000 0 0 0 mprj_io[19]
port 16 nsew signal bidirectional
flabel metal5 s 698512 146440 711002 158960 0 FreeSans 16000 0 0 0 mprj_io[1]
port 17 nsew signal bidirectional
flabel metal5 s 231810 1018624 243978 1030789 0 FreeSans 16000 0 0 0 mprj_io[20]
port 18 nsew signal bidirectional
flabel metal5 s 181410 1018624 193578 1030789 0 FreeSans 16000 0 0 0 mprj_io[21]
port 19 nsew signal bidirectional
flabel metal5 s 130010 1018624 142178 1030789 0 FreeSans 16000 0 0 0 mprj_io[22]
port 20 nsew signal bidirectional
flabel metal5 s 78610 1018624 90778 1030789 0 FreeSans 16000 0 0 0 mprj_io[23]
port 21 nsew signal bidirectional
flabel metal5 s 6811 956610 18976 968778 0 FreeSans 16000 0 0 0 mprj_io[24]
port 22 nsew signal bidirectional
flabel metal5 s 6598 786640 19088 799160 0 FreeSans 16000 0 0 0 mprj_io[25]
port 23 nsew signal bidirectional
flabel metal5 s 6598 743440 19088 755960 0 FreeSans 16000 0 0 0 mprj_io[26]
port 24 nsew signal bidirectional
flabel metal5 s 6598 700240 19088 712760 0 FreeSans 16000 0 0 0 mprj_io[27]
port 25 nsew signal bidirectional
flabel metal5 s 6598 657040 19088 669560 0 FreeSans 16000 0 0 0 mprj_io[28]
port 26 nsew signal bidirectional
flabel metal5 s 6598 613840 19088 626360 0 FreeSans 16000 0 0 0 mprj_io[29]
port 27 nsew signal bidirectional
flabel metal5 s 698512 191440 711002 203960 0 FreeSans 16000 0 0 0 mprj_io[2]
port 28 nsew signal bidirectional
flabel metal5 s 6598 570640 19088 583160 0 FreeSans 16000 0 0 0 mprj_io[30]
port 29 nsew signal bidirectional
flabel metal5 s 6598 527440 19088 539960 0 FreeSans 16000 0 0 0 mprj_io[31]
port 30 nsew signal bidirectional
flabel metal5 s 6598 399840 19088 412360 0 FreeSans 16000 0 0 0 mprj_io[32]
port 31 nsew signal bidirectional
flabel metal5 s 6598 356640 19088 369160 0 FreeSans 16000 0 0 0 mprj_io[33]
port 32 nsew signal bidirectional
flabel metal5 s 6598 313440 19088 325960 0 FreeSans 16000 0 0 0 mprj_io[34]
port 33 nsew signal bidirectional
flabel metal5 s 6598 270240 19088 282760 0 FreeSans 16000 0 0 0 mprj_io[35]
port 34 nsew signal bidirectional
flabel metal5 s 6598 227040 19088 239560 0 FreeSans 16000 0 0 0 mprj_io[36]
port 35 nsew signal bidirectional
flabel metal5 s 6598 183840 19088 196360 0 FreeSans 16000 0 0 0 mprj_io[37]
port 36 nsew signal bidirectional
flabel metal5 s 698512 236640 711002 249160 0 FreeSans 16000 0 0 0 mprj_io[3]
port 37 nsew signal bidirectional
flabel metal5 s 698512 281640 711002 294160 0 FreeSans 16000 0 0 0 mprj_io[4]
port 38 nsew signal bidirectional
flabel metal5 s 698512 326640 711002 339160 0 FreeSans 16000 0 0 0 mprj_io[5]
port 39 nsew signal bidirectional
flabel metal5 s 698512 371840 711002 384360 0 FreeSans 16000 0 0 0 mprj_io[6]
port 40 nsew signal bidirectional
flabel metal5 s 698512 549040 711002 561560 0 FreeSans 16000 0 0 0 mprj_io[7]
port 41 nsew signal bidirectional
flabel metal5 s 698512 594240 711002 606760 0 FreeSans 16000 0 0 0 mprj_io[8]
port 42 nsew signal bidirectional
flabel metal5 s 698512 639240 711002 651760 0 FreeSans 16000 0 0 0 mprj_io[9]
port 43 nsew signal bidirectional
flabel metal5 s 136713 7143 144150 18309 0 FreeSans 16000 0 0 0 resetb
port 44 nsew signal input
flabel metal5 s 6167 70054 19620 80934 0 FreeSans 16000 0 0 0 vccd
port 45 nsew signal bidirectional
flabel metal5 s 697980 909666 711433 920546 0 FreeSans 16000 0 0 0 vccd1
port 46 nsew signal bidirectional
flabel metal5 s 6167 914054 19620 924934 0 FreeSans 16000 0 0 0 vccd2
port 47 nsew signal bidirectional
flabel metal5 s 624222 6811 636390 18976 0 FreeSans 16000 0 0 0 vdda
port 48 nsew signal bidirectional
flabel metal5 s 698624 819822 710789 831990 0 FreeSans 16000 0 0 0 vdda1
port 49 nsew signal bidirectional
flabel metal5 s 698624 505222 710789 517390 0 FreeSans 16000 0 0 0 vdda1_2
port 50 nsew signal bidirectional
flabel metal5 s 6811 484410 18976 496578 0 FreeSans 16000 0 0 0 vdda2
port 51 nsew signal bidirectional
flabel metal5 s 6811 111610 18976 123778 0 FreeSans 16000 0 0 0 vddio
port 52 nsew signal bidirectional
flabel metal5 s 6811 871210 18976 883378 0 FreeSans 16000 0 0 0 vddio_2
port 53 nsew signal bidirectional
flabel metal5 s 80222 6811 92390 18976 0 FreeSans 16000 0 0 0 vssa
port 54 nsew signal bidirectional
flabel metal5 s 577010 1018624 589178 1030789 0 FreeSans 16000 0 0 0 vssa1
port 55 nsew signal bidirectional
flabel metal5 s 698624 417022 710789 429190 0 FreeSans 16000 0 0 0 vssa1_2
port 56 nsew signal bidirectional
flabel metal5 s 6811 829010 18976 841178 0 FreeSans 16000 0 0 0 vssa2
port 57 nsew signal bidirectional
flabel metal5 s 243266 6167 254146 19620 0 FreeSans 16000 0 0 0 vssd
port 58 nsew signal bidirectional
flabel metal5 s 697980 461866 711433 472746 0 FreeSans 16000 0 0 0 vssd1
port 59 nsew signal bidirectional
flabel metal5 s 6167 442854 19620 453734 0 FreeSans 16000 0 0 0 vssd2
port 60 nsew signal bidirectional
flabel metal5 s 570422 6811 582590 18976 0 FreeSans 16000 0 0 0 vssio
port 61 nsew signal bidirectional
flabel metal5 s 334810 1018624 346978 1030789 0 FreeSans 16000 0 0 0 vssio_2
port 62 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 717600 1037600
<< end >>
