* NGSPICE file created from gpio_control_block.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfbbn_2 abstract view
.subckt sky130_fd_sc_hd__dfbbn_2 CLK_N D RESET_B SET_B VGND VNB VPB VPWR Q Q_N
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__einvp_8 abstract view
.subckt sky130_fd_sc_hd__einvp_8 A TE VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_2 abstract view
.subckt sky130_fd_sc_hd__ebufn_2 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for gpio_logic_high abstract view
.subckt gpio_logic_high gpio_logic1 vccd1 vssd1
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd2_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd2_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s50_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s50_1 A VGND VNB VPB VPWR X
.ends

.subckt gpio_control_block gpio_defaults[0] gpio_defaults[10] gpio_defaults[11] gpio_defaults[12]
+ gpio_defaults[1] gpio_defaults[2] gpio_defaults[3] gpio_defaults[4] gpio_defaults[5]
+ gpio_defaults[6] gpio_defaults[7] gpio_defaults[8] gpio_defaults[9] mgmt_gpio_in
+ mgmt_gpio_oeb mgmt_gpio_out one pad_gpio_ana_en pad_gpio_ana_pol pad_gpio_ana_sel
+ pad_gpio_dm[0] pad_gpio_dm[1] pad_gpio_dm[2] pad_gpio_holdover pad_gpio_ib_mode_sel
+ pad_gpio_in pad_gpio_inenb pad_gpio_out pad_gpio_outenb pad_gpio_slow_sel pad_gpio_vtrip_sel
+ resetn resetn_out serial_clock serial_clock_out serial_data_in serial_data_out serial_load
+ serial_load_out user_gpio_in user_gpio_oeb user_gpio_out vccd vccd1 vssd vssd1 zero
X_200_ _207_/CLK _200_/D resetn vssd vssd vccd vccd _201_/D sky130_fd_sc_hd__dfrtp_2
XFILLER_18_31 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__127__B_N gpio_defaults[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_114_ resetn vssd vssd vccd vccd _177_/A sky130_fd_sc_hd__buf_1
XFILLER_13_3 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_57 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_130_ _130_/A vssd vssd vccd vccd _130_/X sky130_fd_sc_hd__buf_1
XANTENNA__124__B gpio_defaults[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__160__B_N gpio_defaults[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xhold20 hold20/A vssd vssd vccd vccd _190_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_179__3 _179__3/A vssd vssd vccd vccd _179__3/Y sky130_fd_sc_hd__inv_2
X_189_ _154__11/Y _189_/D _153_/X _156_/X vssd vssd vccd vccd pad_gpio_dm[0] _104_/A2
+ sky130_fd_sc_hd__dfbbn_2
XANTENNA__200__RESET_B resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xclkbuf_1_1_0__077_ clkbuf_0__077_/X vssd vssd vccd vccd _131__7/A sky130_fd_sc_hd__clkbuf_2
X_112_ _210_/A vssd vssd vccd vccd _112_/X sky130_fd_sc_hd__buf_1
Xhold10 _207_/D vssd vssd vccd vccd hold20/A sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold21 _203_/D vssd vssd vccd vccd _194_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_3_26 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_111_ _111_/A vssd vssd vccd vccd _111_/X sky130_fd_sc_hd__buf_1
XANTENNA__146__B gpio_defaults[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_188_ _148__10/Y _188_/D _147_/X _150_/X vssd vssd vccd vccd _188_/Q _188_/Q_N sky130_fd_sc_hd__dfbbn_2
XFILLER_15_24 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xhold22 _202_/D vssd vssd vccd vccd _193_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_6_26 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xhold11 hold1/X vssd vssd vccd vccd _187_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_187_ _142__9/Y _187_/D _140_/X _145_/X vssd vssd vccd vccd pad_gpio_ib_mode_sel
+ _187_/Q_N sky130_fd_sc_hd__dfbbn_2
X_110_ _180_/A gpio_defaults[0] vssd vssd vccd vccd _111_/A sky130_fd_sc_hd__or2_2
Xhold12 _200_/D vssd vssd vccd vccd hold1/A sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold23 _201_/D vssd vssd vccd vccd _192_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_1_82 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__162__B gpio_defaults[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_93 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__157__B gpio_defaults[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_186_ _136__8/Y _186_/D _135_/X _138_/X vssd vssd vccd vccd pad_gpio_inenb _186_/Q_N
+ sky130_fd_sc_hd__dfbbn_2
Xhold13 hold2/X vssd vssd vccd vccd _191_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XPHY_0 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__203__RESET_B resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_185_ _131__7/Y _185_/D _130_/X _133_/X vssd vssd vccd vccd pad_gpio_vtrip_sel _185_/Q_N
+ sky130_fd_sc_hd__dfbbn_2
XANTENNA__196__RESET_B resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_099_ _188_/Q mgmt_gpio_oeb _182_/Q _098_/X vssd vssd vccd vccd pad_gpio_outenb sky130_fd_sc_hd__a31o_2
Xhold14 hold4/X vssd vssd vccd vccd _188_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_168_ _168_/A vssd vssd vccd vccd _168_/X sky130_fd_sc_hd__buf_1
XPHY_1 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_164__13 _164__13/A vssd vssd vccd vccd _164__13/Y sky130_fd_sc_hd__inv_2
X_184_ _126__6/Y hold8/X _125_/X _128_/X vssd vssd vccd vccd pad_gpio_slow_sel _184_/Q_N
+ sky130_fd_sc_hd__dfbbn_2
XFILLER_18_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xconst_source vssd vssd vccd vccd one zero sky130_fd_sc_hd__conb_1
X_098_ _182_/Q user_gpio_oeb vssd vssd vccd vccd _098_/X sky130_fd_sc_hd__and2b_2
Xhold15 hold5/X vssd vssd vccd vccd _183_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_167_ _172_/A gpio_defaults[5] vssd vssd vccd vccd _168_/A sky130_fd_sc_hd__or2_2
XFILLER_16_93 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_2 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_183_ _120__5/Y _183_/D _119_/X _122_/X vssd vssd vccd vccd pad_gpio_holdover _183_/Q_N
+ sky130_fd_sc_hd__dfbbn_2
X_166_ _166_/A vssd vssd vccd vccd _166_/X sky130_fd_sc_hd__buf_1
X_097_ _097_/A vssd vssd vccd vccd _097_/X sky130_fd_sc_hd__buf_1
Xhold16 hold6/X vssd vssd vccd vccd _182_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_149_ _165_/A gpio_defaults[1] vssd vssd vccd vccd _150_/A sky130_fd_sc_hd__or2b_2
XPHY_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__100__A user_gpio_out vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_182_ _113__4/Y _182_/D _111_/X _117_/X vssd vssd vccd vccd _182_/Q _182_/Q_N sky130_fd_sc_hd__dfbbn_2
Xhold17 hold3/X vssd vssd vccd vccd _189_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_096_ pad_gpio_inenb _188_/Q vssd vssd vccd vccd _097_/A sky130_fd_sc_hd__or2b_2
X_165_ _165_/A gpio_defaults[12] vssd vssd vccd vccd _166_/A sky130_fd_sc_hd__or2b_2
XANTENNA__206__RESET_B resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_4 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__199__RESET_B resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xclkbuf_1_1_0_serial_load clkbuf_0_serial_load/X vssd vssd vccd vccd _210_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__195__D serial_data_in vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_181_ _181_/A vssd vssd vccd vccd _181_/X sky130_fd_sc_hd__buf_1
XFILLER_18_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_147_ _147_/A vssd vssd vccd vccd _147_/X sky130_fd_sc_hd__buf_1
Xhold18 hold7/X vssd vssd vccd vccd _186_/D sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA__106__A pad_gpio_in vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_5 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__114__A resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_180_ _180_/A gpio_defaults[7] vssd vssd vccd vccd _181_/A sky130_fd_sc_hd__or2b_2
X_169__1 _179__3/A vssd vssd vccd vccd _169__1/Y sky130_fd_sc_hd__inv_2
XANTENNA__109__A resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xhold19 hold9/X vssd vssd vccd vccd _185_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_163_ _163_/A vssd vssd vccd vccd _163_/X sky130_fd_sc_hd__buf_1
XANTENNA__149__B_N gpio_defaults[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_34 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_78 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_129_ _146_/A gpio_defaults[9] vssd vssd vccd vccd _130_/A sky130_fd_sc_hd__or2_2
Xclkbuf_0__077_ _112_/X vssd vssd vccd vccd clkbuf_0__077_/X sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_0_0__077_ clkbuf_0__077_/X vssd vssd vccd vccd _136__8/A sky130_fd_sc_hd__clkbuf_2
X_146_ _146_/A gpio_defaults[1] vssd vssd vccd vccd _147_/A sky130_fd_sc_hd__or2_2
XPHY_6 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_174__2 _179__3/A vssd vssd vccd vccd _174__2/Y sky130_fd_sc_hd__inv_2
X_162_ _172_/A gpio_defaults[12] vssd vssd vccd vccd _163_/A sky130_fd_sc_hd__or2_2
X_145_ _145_/A vssd vssd vccd vccd _145_/X sky130_fd_sc_hd__buf_1
XANTENNA__116__B_N gpio_defaults[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_128_ _128_/A vssd vssd vccd vccd _128_/X sky130_fd_sc_hd__buf_1
XFILLER_7_78 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_7 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_161_ _161_/A vssd vssd vccd vccd _161_/X sky130_fd_sc_hd__buf_1
Xgpio_in_buf _106_/Y gpio_in_buf/TE vssd vssd vccd vccd user_gpio_in sky130_fd_sc_hd__einvp_8
XANTENNA_clkbuf_0_serial_load_A serial_load vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_127_ _137_/A gpio_defaults[8] vssd vssd vccd vccd _128_/A sky130_fd_sc_hd__or2b_2
XFILLER_16_3 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_144_ _165_/A gpio_defaults[4] vssd vssd vccd vccd _145_/A sky130_fd_sc_hd__or2b_2
XPHY_8 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_143_ _177_/A vssd vssd vccd vccd _165_/A sky130_fd_sc_hd__buf_1
X_136__8 _136__8/A vssd vssd vccd vccd _136__8/Y sky130_fd_sc_hd__inv_2
X_160_ _165_/A gpio_defaults[11] vssd vssd vccd vccd _161_/A sky130_fd_sc_hd__or2b_2
XFILLER_1_26 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_9 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__139__B gpio_defaults[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_109_ resetn vssd vssd vccd vccd _180_/A sky130_fd_sc_hd__buf_1
XTAP_60 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__152__B gpio_defaults[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_125_ _125_/A vssd vssd vccd vccd _125_/X sky130_fd_sc_hd__buf_1
X_211_ pad_gpio_in _097_/X vssd vssd vccd vccd mgmt_gpio_in sky130_fd_sc_hd__ebufn_2
X_108_ _108_/A vssd vssd vccd vccd serial_data_out sky130_fd_sc_hd__buf_1
X_154__11 _142__9/A vssd vssd vccd vccd _154__11/Y sky130_fd_sc_hd__inv_2
XFILLER_13_69 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__175__B_N gpio_defaults[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_210_ _210_/A vssd vssd vccd vccd serial_load_out sky130_fd_sc_hd__buf_2
XTAP_61 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_50 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_141_ _210_/A vssd vssd vccd vccd _141_/X sky130_fd_sc_hd__buf_1
X_124_ _146_/A gpio_defaults[8] vssd vssd vccd vccd _125_/A sky130_fd_sc_hd__or2_2
Xclkbuf_1_1_0_serial_clock clkbuf_0_serial_clock/X vssd vssd vccd vccd _209_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__202__RESET_B resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__195__RESET_B resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_3 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_107_ one _107_/B vssd vssd vccd vccd _108_/A sky130_fd_sc_hd__and2_2
XANTENNA__165__B_N gpio_defaults[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_62 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_140_ _140_/A vssd vssd vccd vccd _140_/X sky130_fd_sc_hd__buf_1
XFILLER_10_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_51 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_40 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_123_ _177_/A vssd vssd vccd vccd _146_/A sky130_fd_sc_hd__buf_1
X_106_ pad_gpio_in vssd vssd vccd vccd _106_/Y sky130_fd_sc_hd__inv_2
X_148__10 _142__9/A vssd vssd vccd vccd _148__10/Y sky130_fd_sc_hd__inv_2
XANTENNA__177__B gpio_defaults[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__132__B_N gpio_defaults[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_63 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_52 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_41 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__155__B_N gpio_defaults[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_60 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_122_ _122_/A vssd vssd vccd vccd _122_/X sky130_fd_sc_hd__buf_1
X_199_ _207_/CLK hold7/A resetn vssd vssd vccd vccd _200_/D sky130_fd_sc_hd__dfrtp_2
X_105_ _182_/Q _100_/Y _103_/X _104_/Y vssd vssd vccd vccd pad_gpio_out sky130_fd_sc_hd__o22ai_2
XTAP_64 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_93 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_53 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_198_ _209_/A hold5/A resetn vssd vssd vccd vccd hold7/A sky130_fd_sc_hd__dfrtp_2
XTAP_42 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__098__B user_gpio_oeb vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_121_ _137_/A gpio_defaults[2] vssd vssd vccd vccd _122_/A sky130_fd_sc_hd__or2b_2
X_104_ pad_gpio_dm[2] _104_/A2 _101_/Y _182_/Q vssd vssd vccd vccd _104_/Y sky130_fd_sc_hd__o31ai_2
XFILLER_12_3 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_65 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__205__RESET_B resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_54 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_43 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_197_ _209_/A hold4/A resetn vssd vssd vccd vccd hold5/A sky130_fd_sc_hd__dfrtp_2
XANTENNA__198__RESET_B resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_103_ pad_gpio_dm[2] _101_/Y _102_/Y vssd vssd vccd vccd _103_/X sky130_fd_sc_hd__o21a_2
X_120__5 _136__8/A vssd vssd vccd vccd _120__5/Y sky130_fd_sc_hd__inv_2
Xhold1 hold1/A vssd vssd vccd vccd hold1/X sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_55 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_196_ _209_/A hold6/A resetn vssd vssd vccd vccd hold4/A sky130_fd_sc_hd__dfrtp_2
XANTENNA__101__A mgmt_gpio_oeb vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_44 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_102_ mgmt_gpio_out vssd vssd vccd vccd _102_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_0_serial_load serial_load vssd vssd vccd vccd clkbuf_0_serial_load/X sky130_fd_sc_hd__clkbuf_16
Xhold2 hold2/A vssd vssd vccd vccd hold2/X sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_56 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_45 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xgpio_logic_high gpio_in_buf/TE vccd1 vssd1 gpio_logic_high
X_195_ _209_/A serial_data_in resetn vssd vssd vccd vccd hold6/A sky130_fd_sc_hd__dfrtp_2
X_101_ mgmt_gpio_oeb pad_gpio_dm[1] vssd vssd vccd vccd _101_/Y sky130_fd_sc_hd__nand2_2
X_178_ _178_/A vssd vssd vccd vccd _178_/X sky130_fd_sc_hd__buf_1
Xhold3 hold3/A vssd vssd vccd vccd hold3/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xclkbuf_1_1_0__049_ clkbuf_0__049_/X vssd vssd vccd vccd _142__9/A sky130_fd_sc_hd__clkbuf_2
Xclkbuf_1_0_0_serial_load clkbuf_0_serial_load/X vssd vssd vccd vccd _179__3/A sky130_fd_sc_hd__clkbuf_2
XFILLER_10_3 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_126__6 _131__7/A vssd vssd vccd vccd _126__6/Y sky130_fd_sc_hd__inv_2
XFILLER_14_42 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_57 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_46 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_194_ _179__3/Y _194_/D _178_/X _181_/X vssd vssd vccd vccd pad_gpio_ana_pol _194_/Q_N
+ sky130_fd_sc_hd__dfbbn_2
X_100_ user_gpio_out vssd vssd vccd vccd _100_/Y sky130_fd_sc_hd__inv_2
XANTENNA__208__A resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_177_ _177_/A gpio_defaults[7] vssd vssd vccd vccd _178_/A sky130_fd_sc_hd__or2_2
Xhold4 hold4/A vssd vssd vccd vccd hold4/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_131__7 _131__7/A vssd vssd vccd vccd _131__7/Y sky130_fd_sc_hd__inv_2
XTAP_58 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_47 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_20 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_193_ _174__2/Y _193_/D _173_/X _176_/X vssd vssd vccd vccd pad_gpio_ana_sel _193_/Q_N
+ sky130_fd_sc_hd__dfbbn_2
XANTENNA__118__B gpio_defaults[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_176_ _176_/A vssd vssd vccd vccd _176_/X sky130_fd_sc_hd__buf_1
Xhold5 hold5/A vssd vssd vccd vccd hold5/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xdata_delay_1 hold2/A vssd vssd vccd vccd data_delay_2/A sky130_fd_sc_hd__dlygate4sd2_1
XPHY_32 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_59 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_48 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_192_ _169__1/Y _192_/D _168_/X _171_/X vssd vssd vccd vccd pad_gpio_ana_en _192_/Q_N
+ sky130_fd_sc_hd__dfbbn_2
X_175_ _180_/A gpio_defaults[6] vssd vssd vccd vccd _176_/A sky130_fd_sc_hd__or2b_2
XFILLER_2_47 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__129__B gpio_defaults[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__134__B gpio_defaults[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xhold6 hold6/A vssd vssd vccd vccd hold6/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_158_ _158_/A vssd vssd vccd vccd _158_/X sky130_fd_sc_hd__buf_1
XTAP_49 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_38 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0_0_serial_clock clkbuf_0_serial_clock/X vssd vssd vccd vccd _207_/CLK sky130_fd_sc_hd__clkbuf_2
Xdata_delay_2 data_delay_2/A vssd vssd vccd vccd _107_/B sky130_fd_sc_hd__dlygate4sd2_1
XPHY_33 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_24 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_22 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xclkbuf_0_serial_clock serial_clock vssd vssd vccd vccd clkbuf_0_serial_clock/X sky130_fd_sc_hd__clkbuf_16
X_191_ _164__13/Y _191_/D _163_/X _166_/X vssd vssd vccd vccd pad_gpio_dm[2] _191_/Q_N
+ sky130_fd_sc_hd__dfbbn_2
XPHY_11 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_157_ _172_/A gpio_defaults[11] vssd vssd vccd vccd _158_/A sky130_fd_sc_hd__or2_2
X_209_ _209_/A vssd vssd vccd vccd serial_clock_out sky130_fd_sc_hd__buf_2
Xhold7 hold7/A vssd vssd vccd vccd hold7/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_5_26 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_142__9 _142__9/A vssd vssd vccd vccd _142__9/Y sky130_fd_sc_hd__inv_2
XANTENNA__201__RESET_B resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_39 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_34 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_23 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_190_ _159__12/Y _190_/D _158_/X _161_/X vssd vssd vccd vccd pad_gpio_dm[1] _190_/Q_N
+ sky130_fd_sc_hd__dfbbn_2
X_173_ _173_/A vssd vssd vccd vccd _173_/X sky130_fd_sc_hd__buf_1
X_156_ _156_/A vssd vssd vccd vccd _156_/X sky130_fd_sc_hd__buf_1
XFILLER_8_37 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xhold8 hold8/A vssd vssd vccd vccd hold8/X sky130_fd_sc_hd__clkdlybuf4s50_1
X_208_ resetn vssd vssd vccd vccd resetn_out sky130_fd_sc_hd__buf_2
X_139_ _146_/A gpio_defaults[4] vssd vssd vccd vccd _140_/A sky130_fd_sc_hd__or2_2
XPHY_35 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_24 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_13 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_3 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_155_ _165_/A gpio_defaults[10] vssd vssd vccd vccd _156_/A sky130_fd_sc_hd__or2b_2
X_172_ _172_/A gpio_defaults[6] vssd vssd vccd vccd _173_/A sky130_fd_sc_hd__or2_2
XFILLER_3_93 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_138_ _138_/A vssd vssd vccd vccd _138_/X sky130_fd_sc_hd__buf_1
Xhold9 hold9/A vssd vssd vccd vccd hold9/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_72 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_207_ _207_/CLK _207_/D resetn vssd vssd vccd vccd hold2/A sky130_fd_sc_hd__dfrtp_2
XANTENNA__172__B gpio_defaults[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__167__B gpio_defaults[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_36 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_25 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_171_ _171_/A vssd vssd vccd vccd _171_/X sky130_fd_sc_hd__buf_1
XPHY_14 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_80 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_137_ _137_/A gpio_defaults[3] vssd vssd vccd vccd _138_/A sky130_fd_sc_hd__or2b_2
XFILLER_17_3 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__096__A pad_gpio_inenb vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_206_ _209_/A hold3/A resetn vssd vssd vccd vccd _207_/D sky130_fd_sc_hd__dfrtp_2
XPHY_37 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_26 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__121__B_N gpio_defaults[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_170_ _180_/A gpio_defaults[5] vssd vssd vccd vccd _171_/A sky130_fd_sc_hd__or2b_2
XANTENNA__204__RESET_B resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_93 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_205_ _209_/A hold9/A resetn vssd vssd vccd vccd hold3/A sky130_fd_sc_hd__dfrtp_2
X_153_ _153_/A vssd vssd vccd vccd _153_/X sky130_fd_sc_hd__buf_1
XANTENNA__144__B_N gpio_defaults[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_119_ _119_/A vssd vssd vccd vccd _119_/X sky130_fd_sc_hd__buf_1
XANTENNA__197__RESET_B resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_93 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_16 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_113__4 _136__8/A vssd vssd vccd vccd _113__4/Y sky130_fd_sc_hd__inv_2
X_152_ _172_/A gpio_defaults[10] vssd vssd vccd vccd _153_/A sky130_fd_sc_hd__or2_2
X_135_ _135_/A vssd vssd vccd vccd _135_/X sky130_fd_sc_hd__buf_1
X_204_ _209_/A hold8/A resetn vssd vssd vccd vccd hold9/A sky130_fd_sc_hd__dfrtp_2
X_118_ _180_/A gpio_defaults[2] vssd vssd vccd vccd _119_/A sky130_fd_sc_hd__or2_2
XPHY_28 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_17 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xclkbuf_0__049_ _141_/X vssd vssd vccd vccd clkbuf_0__049_/X sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_0_0__049_ clkbuf_0__049_/X vssd vssd vccd vccd _164__13/A sky130_fd_sc_hd__clkbuf_2
X_134_ _146_/A gpio_defaults[3] vssd vssd vccd vccd _135_/A sky130_fd_sc_hd__or2_2
X_203_ _207_/CLK _203_/D resetn vssd vssd vccd vccd hold8/A sky130_fd_sc_hd__dfrtp_2
X_151_ _177_/A vssd vssd vccd vccd _172_/A sky130_fd_sc_hd__buf_1
XFILLER_18_61 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_117_ _117_/A vssd vssd vccd vccd _117_/X sky130_fd_sc_hd__buf_1
XPHY_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_18 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__102__A mgmt_gpio_out vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_150_ _150_/A vssd vssd vccd vccd _150_/X sky130_fd_sc_hd__buf_1
X_159__12 _164__13/A vssd vssd vccd vccd _159__12/Y sky130_fd_sc_hd__inv_2
X_133_ _133_/A vssd vssd vccd vccd _133_/X sky130_fd_sc_hd__buf_1
X_202_ _207_/CLK _202_/D resetn vssd vssd vccd vccd _203_/D sky130_fd_sc_hd__dfrtp_2
X_116_ _137_/A gpio_defaults[0] vssd vssd vccd vccd _117_/A sky130_fd_sc_hd__or2b_2
XPHY_19 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__180__B_N gpio_defaults[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__207__RESET_B resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_0_serial_clock_A serial_clock vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__137__B_N gpio_defaults[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_132_ _137_/A gpio_defaults[9] vssd vssd vccd vccd _133_/A sky130_fd_sc_hd__or2b_2
XANTENNA__099__A2 mgmt_gpio_oeb vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_201_ _207_/CLK _201_/D resetn vssd vssd vccd vccd _202_/D sky130_fd_sc_hd__dfrtp_2
XANTENNA__110__B gpio_defaults[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_115_ _177_/A vssd vssd vccd vccd _137_/A sky130_fd_sc_hd__buf_1
XANTENNA__211__A pad_gpio_in vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__170__B_N gpio_defaults[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
.ends

