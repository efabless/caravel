VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO padframe_power_connections
  CLASS BLOCK ;
  FOREIGN padframe_power_connections ;
  ORIGIN 0.000 0.000 ;
  SIZE 0 BY 0 ;
END padframe_power_connections
END LIBRARY

