magic
tech sky130A
magscale 1 2
timestamp 1636038210
<< locali >>
rect 4537 10455 4571 10693
rect 3617 10047 3651 10149
rect 10517 9775 10551 10489
rect 5181 8279 5215 8585
rect 5181 8245 5273 8279
rect 2789 6783 2823 6953
rect 3985 6647 4019 6817
rect 1593 5695 1627 6409
rect 10367 6409 10517 6443
rect 2237 5559 2271 6409
rect 2697 4879 2731 5865
rect 2881 5355 2915 5661
rect 2973 5559 3007 5865
rect 8125 5559 8159 5865
rect 3341 3043 3375 3145
<< viali >>
rect 1317 11305 1351 11339
rect 1869 11305 1903 11339
rect 2973 11305 3007 11339
rect 7021 11305 7055 11339
rect 2329 11237 2363 11271
rect 3249 11237 3283 11271
rect 5457 11237 5491 11271
rect 5917 11237 5951 11271
rect 6285 11237 6319 11271
rect 6653 11237 6687 11271
rect 7941 11169 7975 11203
rect 1501 11101 1535 11135
rect 2053 11101 2087 11135
rect 2513 11101 2547 11135
rect 2881 11101 2915 11135
rect 3157 11101 3191 11135
rect 3433 11101 3467 11135
rect 3617 11101 3651 11135
rect 5641 11101 5675 11135
rect 5733 11101 5767 11135
rect 6193 11101 6227 11135
rect 6469 11101 6503 11135
rect 6837 11101 6871 11135
rect 7389 11101 7423 11135
rect 8861 11101 8895 11135
rect 9229 11101 9263 11135
rect 3893 11033 3927 11067
rect 5365 10965 5399 10999
rect 9045 10965 9079 10999
rect 9413 10965 9447 10999
rect 9045 10761 9079 10795
rect 4537 10693 4571 10727
rect 1685 10625 1719 10659
rect 2053 10625 2087 10659
rect 2329 10625 2363 10659
rect 2605 10625 2639 10659
rect 2697 10557 2731 10591
rect 2973 10557 3007 10591
rect 4445 10557 4479 10591
rect 1501 10489 1535 10523
rect 2421 10489 2455 10523
rect 4813 10625 4847 10659
rect 5089 10625 5123 10659
rect 5365 10625 5399 10659
rect 5641 10625 5675 10659
rect 5733 10625 5767 10659
rect 6193 10625 6227 10659
rect 6561 10625 6595 10659
rect 8493 10625 8527 10659
rect 8861 10625 8895 10659
rect 9229 10625 9263 10659
rect 6837 10557 6871 10591
rect 4905 10489 4939 10523
rect 5917 10489 5951 10523
rect 6377 10489 6411 10523
rect 10517 10489 10551 10523
rect 2145 10421 2179 10455
rect 4537 10421 4571 10455
rect 4629 10421 4663 10455
rect 5181 10421 5215 10455
rect 5457 10421 5491 10455
rect 8309 10421 8343 10455
rect 8677 10421 8711 10455
rect 9413 10421 9447 10455
rect 2697 10217 2731 10251
rect 8585 10217 8619 10251
rect 8769 10217 8803 10251
rect 2973 10149 3007 10183
rect 3617 10149 3651 10183
rect 3709 10149 3743 10183
rect 6285 10149 6319 10183
rect 8125 10149 8159 10183
rect 3985 10081 4019 10115
rect 4353 10081 4387 10115
rect 9321 10081 9355 10115
rect 2605 10013 2639 10047
rect 2881 10013 2915 10047
rect 3157 10013 3191 10047
rect 3433 10013 3467 10047
rect 3617 10013 3651 10047
rect 3893 10013 3927 10047
rect 5825 10013 5859 10047
rect 6377 10013 6411 10047
rect 8401 10013 8435 10047
rect 9137 10013 9171 10047
rect 6653 9945 6687 9979
rect 8217 9945 8251 9979
rect 2421 9877 2455 9911
rect 3249 9877 3283 9911
rect 9229 9877 9263 9911
rect 10517 9741 10551 9775
rect 4629 9673 4663 9707
rect 5365 9673 5399 9707
rect 9321 9673 9355 9707
rect 3065 9605 3099 9639
rect 1501 9537 1535 9571
rect 1777 9537 1811 9571
rect 2421 9537 2455 9571
rect 2697 9537 2731 9571
rect 4813 9537 4847 9571
rect 4905 9537 4939 9571
rect 5641 9537 5675 9571
rect 5825 9537 5859 9571
rect 6009 9537 6043 9571
rect 6377 9537 6411 9571
rect 7389 9537 7423 9571
rect 8861 9537 8895 9571
rect 2789 9469 2823 9503
rect 6837 9469 6871 9503
rect 7021 9469 7055 9503
rect 2237 9401 2271 9435
rect 2513 9401 2547 9435
rect 1317 9333 1351 9367
rect 1593 9333 1627 9367
rect 2053 9333 2087 9367
rect 4537 9333 4571 9367
rect 4997 9333 5031 9367
rect 6469 9333 6503 9367
rect 1501 9129 1535 9163
rect 2697 9129 2731 9163
rect 3617 9129 3651 9163
rect 7481 9129 7515 9163
rect 8217 9129 8251 9163
rect 8769 9129 8803 9163
rect 1869 9061 1903 9095
rect 2053 9061 2087 9095
rect 3249 9061 3283 9095
rect 7941 9061 7975 9095
rect 2605 8993 2639 9027
rect 5187 8993 5221 9027
rect 5549 8993 5583 9027
rect 9321 8993 9355 9027
rect 1409 8925 1443 8959
rect 1685 8925 1719 8959
rect 1777 8925 1811 8959
rect 2237 8925 2271 8959
rect 2881 8925 2915 8959
rect 3157 8925 3191 8959
rect 3433 8925 3467 8959
rect 3801 8925 3835 8959
rect 4077 8925 4111 8959
rect 4353 8925 4387 8959
rect 4629 8925 4663 8959
rect 5089 8925 5123 8959
rect 7021 8925 7055 8959
rect 7757 8925 7791 8959
rect 8125 8925 8159 8959
rect 9137 8925 9171 8959
rect 9229 8857 9263 8891
rect 2973 8789 3007 8823
rect 3893 8789 3927 8823
rect 4169 8789 4203 8823
rect 4445 8789 4479 8823
rect 4905 8789 4939 8823
rect 8585 8789 8619 8823
rect 1501 8585 1535 8619
rect 2329 8585 2363 8619
rect 2421 8585 2455 8619
rect 5181 8585 5215 8619
rect 5917 8585 5951 8619
rect 6929 8585 6963 8619
rect 1409 8449 1443 8483
rect 1685 8449 1719 8483
rect 1961 8449 1995 8483
rect 2605 8449 2639 8483
rect 2973 8449 3007 8483
rect 5089 8433 5123 8467
rect 3065 8381 3099 8415
rect 3341 8381 3375 8415
rect 1777 8313 1811 8347
rect 4905 8313 4939 8347
rect 5457 8517 5491 8551
rect 5641 8517 5675 8551
rect 6285 8517 6319 8551
rect 5273 8449 5307 8483
rect 5825 8449 5859 8483
rect 6469 8449 6503 8483
rect 6745 8449 6779 8483
rect 7665 8449 7699 8483
rect 7757 8449 7791 8483
rect 8401 8449 8435 8483
rect 8585 8449 8619 8483
rect 8677 8449 8711 8483
rect 8861 8449 8895 8483
rect 6653 8381 6687 8415
rect 7113 8381 7147 8415
rect 8217 8381 8251 8415
rect 9321 8381 9355 8415
rect 7573 8313 7607 8347
rect 7941 8313 7975 8347
rect 1225 8245 1259 8279
rect 2789 8245 2823 8279
rect 4813 8245 4847 8279
rect 5273 8245 5307 8279
rect 1593 8041 1627 8075
rect 7113 8041 7147 8075
rect 8033 8041 8067 8075
rect 8769 8041 8803 8075
rect 1501 7973 1535 8007
rect 2237 7973 2271 8007
rect 2513 7973 2547 8007
rect 3801 7973 3835 8007
rect 7573 7973 7607 8007
rect 8493 7973 8527 8007
rect 4813 7905 4847 7939
rect 9321 7905 9355 7939
rect 1777 7837 1811 7871
rect 2053 7837 2087 7871
rect 2421 7837 2455 7871
rect 2697 7837 2731 7871
rect 3157 7837 3191 7871
rect 3985 7837 4019 7871
rect 4261 7837 4295 7871
rect 4721 7837 4755 7871
rect 5181 7837 5215 7871
rect 6653 7837 6687 7871
rect 7389 7837 7423 7871
rect 7757 7837 7791 7871
rect 8309 7837 8343 7871
rect 1225 7701 1259 7735
rect 1869 7701 1903 7735
rect 2973 7701 3007 7735
rect 3433 7701 3467 7735
rect 4077 7701 4111 7735
rect 4537 7701 4571 7735
rect 8217 7701 8251 7735
rect 9137 7701 9171 7735
rect 9229 7701 9263 7735
rect 2881 7497 2915 7531
rect 3157 7497 3191 7531
rect 6009 7497 6043 7531
rect 9137 7497 9171 7531
rect 1593 7361 1627 7395
rect 2513 7361 2547 7395
rect 2789 7361 2823 7395
rect 3065 7361 3099 7395
rect 3341 7361 3375 7395
rect 3617 7361 3651 7395
rect 4077 7361 4111 7395
rect 5549 7361 5583 7395
rect 6193 7361 6227 7395
rect 8677 7361 8711 7395
rect 9229 7361 9263 7395
rect 2145 7293 2179 7327
rect 3709 7293 3743 7327
rect 6837 7293 6871 7327
rect 7205 7293 7239 7327
rect 1961 7225 1995 7259
rect 2605 7225 2639 7259
rect 8861 7225 8895 7259
rect 1409 7157 1443 7191
rect 2329 7157 2363 7191
rect 3433 7157 3467 7191
rect 6469 7157 6503 7191
rect 6653 7157 6687 7191
rect 9413 7157 9447 7191
rect 2789 6953 2823 6987
rect 3065 6953 3099 6987
rect 5549 6953 5583 6987
rect 7481 6953 7515 6987
rect 8769 6953 8803 6987
rect 3249 6817 3283 6851
rect 3985 6817 4019 6851
rect 5733 6817 5767 6851
rect 9321 6817 9355 6851
rect 1501 6749 1535 6783
rect 1777 6749 1811 6783
rect 2145 6749 2179 6783
rect 2421 6749 2455 6783
rect 2697 6749 2731 6783
rect 2789 6749 2823 6783
rect 4169 6749 4203 6783
rect 4445 6749 4479 6783
rect 5273 6749 5307 6783
rect 6009 6749 6043 6783
rect 6193 6749 6227 6783
rect 8217 6749 8251 6783
rect 8309 6749 8343 6783
rect 9137 6749 9171 6783
rect 9229 6749 9263 6783
rect 1317 6613 1351 6647
rect 1593 6613 1627 6647
rect 1961 6613 1995 6647
rect 2237 6613 2271 6647
rect 2513 6613 2547 6647
rect 3341 6613 3375 6647
rect 3617 6613 3651 6647
rect 3801 6613 3835 6647
rect 3985 6613 4019 6647
rect 5825 6613 5859 6647
rect 8033 6613 8067 6647
rect 8493 6613 8527 6647
rect 1593 6409 1627 6443
rect 1593 5661 1627 5695
rect 2237 6409 2271 6443
rect 10333 6409 10367 6443
rect 10517 6409 10551 6443
rect 3617 6341 3651 6375
rect 5457 6341 5491 6375
rect 7389 6341 7423 6375
rect 7757 6341 7791 6375
rect 3341 6273 3375 6307
rect 7021 6273 7055 6307
rect 7205 6273 7239 6307
rect 7665 6273 7699 6307
rect 7941 6273 7975 6307
rect 8309 6273 8343 6307
rect 8861 6273 8895 6307
rect 5181 6205 5215 6239
rect 8769 6137 8803 6171
rect 5089 6069 5123 6103
rect 6929 6069 6963 6103
rect 7481 6069 7515 6103
rect 8125 6069 8159 6103
rect 8401 6069 8435 6103
rect 8953 6069 8987 6103
rect 9321 6069 9355 6103
rect 2237 5525 2271 5559
rect 2697 5865 2731 5899
rect 2973 5865 3007 5899
rect 8033 5865 8067 5899
rect 8125 5865 8159 5899
rect 2881 5661 2915 5695
rect 6101 5729 6135 5763
rect 3341 5661 3375 5695
rect 5549 5661 5583 5695
rect 5733 5661 5767 5695
rect 7573 5661 7607 5695
rect 3617 5593 3651 5627
rect 8861 5797 8895 5831
rect 9413 5797 9447 5831
rect 8401 5729 8435 5763
rect 8493 5729 8527 5763
rect 8677 5661 8711 5695
rect 9137 5661 9171 5695
rect 9229 5661 9263 5695
rect 2973 5525 3007 5559
rect 5089 5525 5123 5559
rect 5365 5525 5399 5559
rect 8125 5525 8159 5559
rect 8953 5525 8987 5559
rect 2881 5321 2915 5355
rect 7665 5321 7699 5355
rect 9137 5321 9171 5355
rect 9229 5321 9263 5355
rect 6193 5253 6227 5287
rect 7941 5253 7975 5287
rect 3433 5185 3467 5219
rect 3801 5185 3835 5219
rect 5273 5185 5307 5219
rect 7757 5185 7791 5219
rect 8677 5185 8711 5219
rect 8787 5185 8821 5219
rect 8953 5185 8987 5219
rect 9413 5185 9447 5219
rect 5917 5117 5951 5151
rect 5733 4981 5767 5015
rect 8125 4981 8159 5015
rect 8493 4981 8527 5015
rect 2697 4845 2731 4879
rect 3341 4777 3375 4811
rect 4445 4777 4479 4811
rect 4629 4777 4663 4811
rect 6101 4777 6135 4811
rect 6745 4777 6779 4811
rect 7113 4777 7147 4811
rect 9505 4777 9539 4811
rect 3617 4709 3651 4743
rect 7205 4641 7239 4675
rect 7573 4641 7607 4675
rect 3525 4573 3559 4607
rect 3801 4573 3835 4607
rect 4077 4573 4111 4607
rect 4169 4573 4203 4607
rect 4721 4573 4755 4607
rect 4997 4573 5031 4607
rect 6469 4573 6503 4607
rect 6653 4573 6687 4607
rect 9045 4573 9079 4607
rect 5733 4505 5767 4539
rect 5917 4505 5951 4539
rect 6285 4505 6319 4539
rect 3893 4437 3927 4471
rect 8309 4233 8343 4267
rect 9045 4233 9079 4267
rect 3433 4097 3467 4131
rect 3801 4097 3835 4131
rect 5273 4097 5307 4131
rect 6193 4097 6227 4131
rect 7665 4097 7699 4131
rect 8493 4097 8527 4131
rect 8585 4097 8619 4131
rect 9321 4097 9355 4131
rect 5825 4029 5859 4063
rect 9137 3961 9171 3995
rect 5733 3893 5767 3927
rect 8125 3893 8159 3927
rect 8861 3893 8895 3927
rect 6009 3689 6043 3723
rect 8585 3689 8619 3723
rect 9229 3689 9263 3723
rect 8953 3621 8987 3655
rect 3341 3553 3375 3587
rect 3617 3553 3651 3587
rect 6285 3553 6319 3587
rect 5733 3485 5767 3519
rect 6653 3485 6687 3519
rect 8125 3485 8159 3519
rect 8861 3485 8895 3519
rect 9137 3485 9171 3519
rect 9413 3485 9447 3519
rect 5181 3417 5215 3451
rect 5365 3417 5399 3451
rect 5089 3349 5123 3383
rect 5549 3349 5583 3383
rect 6193 3349 6227 3383
rect 8677 3349 8711 3383
rect 3341 3145 3375 3179
rect 4629 3145 4663 3179
rect 7205 3145 7239 3179
rect 8769 3145 8803 3179
rect 9137 3145 9171 3179
rect 9229 3145 9263 3179
rect 3709 3077 3743 3111
rect 3341 3009 3375 3043
rect 3617 3009 3651 3043
rect 3893 3009 3927 3043
rect 4169 3009 4203 3043
rect 5089 3009 5123 3043
rect 6561 3009 6595 3043
rect 7389 3009 7423 3043
rect 7481 3009 7515 3043
rect 8309 3009 8343 3043
rect 4721 2941 4755 2975
rect 7021 2941 7055 2975
rect 3433 2873 3467 2907
rect 4077 2805 4111 2839
rect 4261 2805 4295 2839
rect 7573 2805 7607 2839
rect 7941 2805 7975 2839
rect 8401 2805 8435 2839
rect 9413 2805 9447 2839
rect 3525 2601 3559 2635
rect 7573 2601 7607 2635
rect 7941 2601 7975 2635
rect 9229 2601 9263 2635
rect 9321 2601 9355 2635
rect 5549 2533 5583 2567
rect 8677 2533 8711 2567
rect 3801 2465 3835 2499
rect 5733 2465 5767 2499
rect 6009 2465 6043 2499
rect 3709 2397 3743 2431
rect 7757 2397 7791 2431
rect 8125 2397 8159 2431
rect 8309 2397 8343 2431
rect 8861 2397 8895 2431
rect 9505 2397 9539 2431
rect 4077 2329 4111 2363
rect 8493 2329 8527 2363
rect 9045 2329 9079 2363
rect 7481 2261 7515 2295
<< metal1 >>
rect 1210 11772 1216 11824
rect 1268 11812 1274 11824
rect 4982 11812 4988 11824
rect 1268 11784 4988 11812
rect 1268 11772 1274 11784
rect 4982 11772 4988 11784
rect 5040 11772 5046 11824
rect 3418 11704 3424 11756
rect 3476 11744 3482 11756
rect 7650 11744 7656 11756
rect 3476 11716 7656 11744
rect 3476 11704 3482 11716
rect 7650 11704 7656 11716
rect 7708 11704 7714 11756
rect 3234 11636 3240 11688
rect 3292 11676 3298 11688
rect 5074 11676 5080 11688
rect 3292 11648 5080 11676
rect 3292 11636 3298 11648
rect 5074 11636 5080 11648
rect 5132 11676 5138 11688
rect 6270 11676 6276 11688
rect 5132 11648 6276 11676
rect 5132 11636 5138 11648
rect 6270 11636 6276 11648
rect 6328 11636 6334 11688
rect 1854 11568 1860 11620
rect 1912 11608 1918 11620
rect 16574 11608 16580 11620
rect 1912 11580 16580 11608
rect 1912 11568 1918 11580
rect 16574 11568 16580 11580
rect 16632 11568 16638 11620
rect 1302 11500 1308 11552
rect 1360 11540 1366 11552
rect 8570 11540 8576 11552
rect 1360 11512 8576 11540
rect 1360 11500 1366 11512
rect 8570 11500 8576 11512
rect 8628 11500 8634 11552
rect 920 11450 9844 11472
rect 920 11398 2566 11450
rect 2618 11398 2630 11450
rect 2682 11398 2694 11450
rect 2746 11398 2758 11450
rect 2810 11398 2822 11450
rect 2874 11398 5666 11450
rect 5718 11398 5730 11450
rect 5782 11398 5794 11450
rect 5846 11398 5858 11450
rect 5910 11398 5922 11450
rect 5974 11398 8766 11450
rect 8818 11398 8830 11450
rect 8882 11398 8894 11450
rect 8946 11398 8958 11450
rect 9010 11398 9022 11450
rect 9074 11398 9844 11450
rect 920 11376 9844 11398
rect 1302 11336 1308 11348
rect 1263 11308 1308 11336
rect 1302 11296 1308 11308
rect 1360 11296 1366 11348
rect 1854 11336 1860 11348
rect 1815 11308 1860 11336
rect 1854 11296 1860 11308
rect 1912 11296 1918 11348
rect 2961 11339 3019 11345
rect 2961 11305 2973 11339
rect 3007 11336 3019 11339
rect 6454 11336 6460 11348
rect 3007 11308 6460 11336
rect 3007 11305 3019 11308
rect 2961 11299 3019 11305
rect 6454 11296 6460 11308
rect 6512 11296 6518 11348
rect 7009 11339 7067 11345
rect 7009 11305 7021 11339
rect 7055 11336 7067 11339
rect 9674 11336 9680 11348
rect 7055 11308 9680 11336
rect 7055 11305 7067 11308
rect 7009 11299 7067 11305
rect 9674 11296 9680 11308
rect 9732 11296 9738 11348
rect 2317 11271 2375 11277
rect 2317 11237 2329 11271
rect 2363 11268 2375 11271
rect 3050 11268 3056 11280
rect 2363 11240 3056 11268
rect 2363 11237 2375 11240
rect 2317 11231 2375 11237
rect 3050 11228 3056 11240
rect 3108 11228 3114 11280
rect 3237 11271 3295 11277
rect 3237 11237 3249 11271
rect 3283 11237 3295 11271
rect 3237 11231 3295 11237
rect 5445 11271 5503 11277
rect 5445 11237 5457 11271
rect 5491 11268 5503 11271
rect 5905 11271 5963 11277
rect 5491 11240 5856 11268
rect 5491 11237 5503 11240
rect 5445 11231 5503 11237
rect 3252 11200 3280 11231
rect 5828 11200 5856 11240
rect 5905 11237 5917 11271
rect 5951 11268 5963 11271
rect 5994 11268 6000 11280
rect 5951 11240 6000 11268
rect 5951 11237 5963 11240
rect 5905 11231 5963 11237
rect 5994 11228 6000 11240
rect 6052 11228 6058 11280
rect 6270 11268 6276 11280
rect 6231 11240 6276 11268
rect 6270 11228 6276 11240
rect 6328 11228 6334 11280
rect 6641 11271 6699 11277
rect 6641 11237 6653 11271
rect 6687 11268 6699 11271
rect 9490 11268 9496 11280
rect 6687 11240 9496 11268
rect 6687 11237 6699 11240
rect 6641 11231 6699 11237
rect 9490 11228 9496 11240
rect 9548 11228 9554 11280
rect 7098 11200 7104 11212
rect 3252 11172 5764 11200
rect 5828 11172 7104 11200
rect 1489 11135 1547 11141
rect 1489 11101 1501 11135
rect 1535 11132 1547 11135
rect 1854 11132 1860 11144
rect 1535 11104 1860 11132
rect 1535 11101 1547 11104
rect 1489 11095 1547 11101
rect 1854 11092 1860 11104
rect 1912 11092 1918 11144
rect 2041 11135 2099 11141
rect 2041 11101 2053 11135
rect 2087 11132 2099 11135
rect 2406 11132 2412 11144
rect 2087 11104 2412 11132
rect 2087 11101 2099 11104
rect 2041 11095 2099 11101
rect 2406 11092 2412 11104
rect 2464 11132 2470 11144
rect 2501 11135 2559 11141
rect 2501 11132 2513 11135
rect 2464 11104 2513 11132
rect 2464 11092 2470 11104
rect 2501 11101 2513 11104
rect 2547 11101 2559 11135
rect 2501 11095 2559 11101
rect 2869 11135 2927 11141
rect 2869 11101 2881 11135
rect 2915 11132 2927 11135
rect 3142 11132 3148 11144
rect 2915 11104 3148 11132
rect 2915 11101 2927 11104
rect 2869 11095 2927 11101
rect 3142 11092 3148 11104
rect 3200 11092 3206 11144
rect 3418 11132 3424 11144
rect 3379 11104 3424 11132
rect 3418 11092 3424 11104
rect 3476 11092 3482 11144
rect 3602 11132 3608 11144
rect 3563 11104 3608 11132
rect 3602 11092 3608 11104
rect 3660 11092 3666 11144
rect 5258 11092 5264 11144
rect 5316 11132 5322 11144
rect 5736 11141 5764 11172
rect 7098 11160 7104 11172
rect 7156 11160 7162 11212
rect 7926 11200 7932 11212
rect 7887 11172 7932 11200
rect 7926 11160 7932 11172
rect 7984 11160 7990 11212
rect 5629 11135 5687 11141
rect 5629 11132 5641 11135
rect 5316 11104 5641 11132
rect 5316 11092 5322 11104
rect 5629 11101 5641 11104
rect 5675 11101 5687 11135
rect 5629 11095 5687 11101
rect 5721 11135 5779 11141
rect 5721 11101 5733 11135
rect 5767 11101 5779 11135
rect 6178 11132 6184 11144
rect 6139 11104 6184 11132
rect 5721 11095 5779 11101
rect 6178 11092 6184 11104
rect 6236 11092 6242 11144
rect 6457 11135 6515 11141
rect 6457 11101 6469 11135
rect 6503 11101 6515 11135
rect 6822 11132 6828 11144
rect 6783 11104 6828 11132
rect 6457 11095 6515 11101
rect 3881 11067 3939 11073
rect 2746 11036 3096 11064
rect 2406 10956 2412 11008
rect 2464 10996 2470 11008
rect 2746 10996 2774 11036
rect 2464 10968 2774 10996
rect 3068 10996 3096 11036
rect 3881 11033 3893 11067
rect 3927 11064 3939 11067
rect 3970 11064 3976 11076
rect 3927 11036 3976 11064
rect 3927 11033 3939 11036
rect 3881 11027 3939 11033
rect 3970 11024 3976 11036
rect 4028 11024 4034 11076
rect 4338 11024 4344 11076
rect 4396 11024 4402 11076
rect 6472 11064 6500 11095
rect 6822 11092 6828 11104
rect 6880 11092 6886 11144
rect 7377 11135 7435 11141
rect 7377 11101 7389 11135
rect 7423 11132 7435 11135
rect 8294 11132 8300 11144
rect 7423 11104 8300 11132
rect 7423 11101 7435 11104
rect 7377 11095 7435 11101
rect 8294 11092 8300 11104
rect 8352 11092 8358 11144
rect 8849 11135 8907 11141
rect 8849 11101 8861 11135
rect 8895 11101 8907 11135
rect 9214 11132 9220 11144
rect 9175 11104 9220 11132
rect 8849 11095 8907 11101
rect 8864 11064 8892 11095
rect 9214 11092 9220 11104
rect 9272 11092 9278 11144
rect 13814 11064 13820 11076
rect 5276 11036 6500 11064
rect 6932 11036 8892 11064
rect 9048 11036 13820 11064
rect 5276 10996 5304 11036
rect 3068 10968 5304 10996
rect 5353 10999 5411 11005
rect 2464 10956 2470 10968
rect 5353 10965 5365 10999
rect 5399 10996 5411 10999
rect 6178 10996 6184 11008
rect 5399 10968 6184 10996
rect 5399 10965 5411 10968
rect 5353 10959 5411 10965
rect 6178 10956 6184 10968
rect 6236 10956 6242 11008
rect 6362 10956 6368 11008
rect 6420 10996 6426 11008
rect 6932 10996 6960 11036
rect 9048 11005 9076 11036
rect 13814 11024 13820 11036
rect 13872 11024 13878 11076
rect 6420 10968 6960 10996
rect 9033 10999 9091 11005
rect 6420 10956 6426 10968
rect 9033 10965 9045 10999
rect 9079 10965 9091 10999
rect 9398 10996 9404 11008
rect 9359 10968 9404 10996
rect 9033 10959 9091 10965
rect 9398 10956 9404 10968
rect 9456 10956 9462 11008
rect 920 10906 9844 10928
rect 920 10854 4116 10906
rect 4168 10854 4180 10906
rect 4232 10854 4244 10906
rect 4296 10854 4308 10906
rect 4360 10854 4372 10906
rect 4424 10854 7216 10906
rect 7268 10854 7280 10906
rect 7332 10854 7344 10906
rect 7396 10854 7408 10906
rect 7460 10854 7472 10906
rect 7524 10854 9844 10906
rect 920 10832 9844 10854
rect 9033 10795 9091 10801
rect 9033 10792 9045 10795
rect 1688 10764 9045 10792
rect 1688 10665 1716 10764
rect 9033 10761 9045 10764
rect 9079 10761 9091 10795
rect 9033 10755 9091 10761
rect 3418 10724 3424 10736
rect 2608 10696 3424 10724
rect 1673 10659 1731 10665
rect 1673 10625 1685 10659
rect 1719 10625 1731 10659
rect 1673 10619 1731 10625
rect 2041 10659 2099 10665
rect 2041 10625 2053 10659
rect 2087 10656 2099 10659
rect 2314 10656 2320 10668
rect 2087 10628 2320 10656
rect 2087 10625 2099 10628
rect 2041 10619 2099 10625
rect 2314 10616 2320 10628
rect 2372 10616 2378 10668
rect 2608 10665 2636 10696
rect 3418 10684 3424 10696
rect 3476 10684 3482 10736
rect 4525 10727 4583 10733
rect 4525 10693 4537 10727
rect 4571 10724 4583 10727
rect 6914 10724 6920 10736
rect 4571 10696 6224 10724
rect 4571 10693 4583 10696
rect 4525 10687 4583 10693
rect 2593 10659 2651 10665
rect 2593 10625 2605 10659
rect 2639 10625 2651 10659
rect 4798 10656 4804 10668
rect 4759 10628 4804 10656
rect 2593 10619 2651 10625
rect 4798 10616 4804 10628
rect 4856 10616 4862 10668
rect 5074 10656 5080 10668
rect 5035 10628 5080 10656
rect 5074 10616 5080 10628
rect 5132 10616 5138 10668
rect 5353 10659 5411 10665
rect 5353 10625 5365 10659
rect 5399 10656 5411 10659
rect 5534 10656 5540 10668
rect 5399 10628 5540 10656
rect 5399 10625 5411 10628
rect 5353 10619 5411 10625
rect 5534 10616 5540 10628
rect 5592 10616 5598 10668
rect 6196 10665 6224 10696
rect 6380 10696 6920 10724
rect 5629 10659 5687 10665
rect 5629 10625 5641 10659
rect 5675 10625 5687 10659
rect 5629 10619 5687 10625
rect 5721 10659 5779 10665
rect 5721 10625 5733 10659
rect 5767 10656 5779 10659
rect 6181 10659 6239 10665
rect 5767 10628 6132 10656
rect 5767 10625 5779 10628
rect 5721 10619 5779 10625
rect 2685 10591 2743 10597
rect 2685 10557 2697 10591
rect 2731 10557 2743 10591
rect 2685 10551 2743 10557
rect 2961 10591 3019 10597
rect 2961 10557 2973 10591
rect 3007 10588 3019 10591
rect 3510 10588 3516 10600
rect 3007 10560 3516 10588
rect 3007 10557 3019 10560
rect 2961 10551 3019 10557
rect 1486 10520 1492 10532
rect 1447 10492 1492 10520
rect 1486 10480 1492 10492
rect 1544 10480 1550 10532
rect 2406 10520 2412 10532
rect 2367 10492 2412 10520
rect 2406 10480 2412 10492
rect 2464 10480 2470 10532
rect 2130 10452 2136 10464
rect 2091 10424 2136 10452
rect 2130 10412 2136 10424
rect 2188 10412 2194 10464
rect 2700 10452 2728 10551
rect 3510 10548 3516 10560
rect 3568 10548 3574 10600
rect 3970 10548 3976 10600
rect 4028 10588 4034 10600
rect 4338 10588 4344 10600
rect 4028 10560 4344 10588
rect 4028 10548 4034 10560
rect 4338 10548 4344 10560
rect 4396 10588 4402 10600
rect 4433 10591 4491 10597
rect 4433 10588 4445 10591
rect 4396 10560 4445 10588
rect 4396 10548 4402 10560
rect 4433 10557 4445 10560
rect 4479 10557 4491 10591
rect 5644 10588 5672 10619
rect 5994 10588 6000 10600
rect 5644 10560 6000 10588
rect 4433 10551 4491 10557
rect 5994 10548 6000 10560
rect 6052 10548 6058 10600
rect 6104 10588 6132 10628
rect 6181 10625 6193 10659
rect 6227 10625 6239 10659
rect 6181 10619 6239 10625
rect 6270 10588 6276 10600
rect 6104 10560 6276 10588
rect 6270 10548 6276 10560
rect 6328 10548 6334 10600
rect 4893 10523 4951 10529
rect 4893 10489 4905 10523
rect 4939 10520 4951 10523
rect 5258 10520 5264 10532
rect 4939 10492 5264 10520
rect 4939 10489 4951 10492
rect 4893 10483 4951 10489
rect 5258 10480 5264 10492
rect 5316 10480 5322 10532
rect 5905 10523 5963 10529
rect 5905 10489 5917 10523
rect 5951 10520 5963 10523
rect 6086 10520 6092 10532
rect 5951 10492 6092 10520
rect 5951 10489 5963 10492
rect 5905 10483 5963 10489
rect 6086 10480 6092 10492
rect 6144 10480 6150 10532
rect 6380 10529 6408 10696
rect 6914 10684 6920 10696
rect 6972 10684 6978 10736
rect 8772 10696 12434 10724
rect 6546 10656 6552 10668
rect 6507 10628 6552 10656
rect 6546 10616 6552 10628
rect 6604 10616 6610 10668
rect 7926 10616 7932 10668
rect 7984 10656 7990 10668
rect 8202 10656 8208 10668
rect 7984 10628 8208 10656
rect 7984 10616 7990 10628
rect 8202 10616 8208 10628
rect 8260 10616 8266 10668
rect 8478 10656 8484 10668
rect 8439 10628 8484 10656
rect 8478 10616 8484 10628
rect 8536 10616 8542 10668
rect 6454 10548 6460 10600
rect 6512 10588 6518 10600
rect 6825 10591 6883 10597
rect 6825 10588 6837 10591
rect 6512 10560 6837 10588
rect 6512 10548 6518 10560
rect 6825 10557 6837 10560
rect 6871 10557 6883 10591
rect 6825 10551 6883 10557
rect 6914 10548 6920 10600
rect 6972 10588 6978 10600
rect 8772 10588 8800 10696
rect 8849 10659 8907 10665
rect 8849 10625 8861 10659
rect 8895 10625 8907 10659
rect 8849 10619 8907 10625
rect 6972 10560 8800 10588
rect 6972 10548 6978 10560
rect 6365 10523 6423 10529
rect 6365 10489 6377 10523
rect 6411 10489 6423 10523
rect 8864 10520 8892 10619
rect 9122 10616 9128 10668
rect 9180 10656 9186 10668
rect 9217 10659 9275 10665
rect 9217 10656 9229 10659
rect 9180 10628 9229 10656
rect 9180 10616 9186 10628
rect 9217 10625 9229 10628
rect 9263 10625 9275 10659
rect 9217 10619 9275 10625
rect 12406 10588 12434 10696
rect 16758 10588 16764 10600
rect 12406 10560 16764 10588
rect 16758 10548 16764 10560
rect 16816 10548 16822 10600
rect 10505 10523 10563 10529
rect 10505 10520 10517 10523
rect 6365 10483 6423 10489
rect 7852 10492 8892 10520
rect 9324 10492 10517 10520
rect 3050 10452 3056 10464
rect 2700 10424 3056 10452
rect 3050 10412 3056 10424
rect 3108 10452 3114 10464
rect 3602 10452 3608 10464
rect 3108 10424 3608 10452
rect 3108 10412 3114 10424
rect 3602 10412 3608 10424
rect 3660 10412 3666 10464
rect 3694 10412 3700 10464
rect 3752 10452 3758 10464
rect 4525 10455 4583 10461
rect 4525 10452 4537 10455
rect 3752 10424 4537 10452
rect 3752 10412 3758 10424
rect 4525 10421 4537 10424
rect 4571 10421 4583 10455
rect 4525 10415 4583 10421
rect 4617 10455 4675 10461
rect 4617 10421 4629 10455
rect 4663 10452 4675 10455
rect 5074 10452 5080 10464
rect 4663 10424 5080 10452
rect 4663 10421 4675 10424
rect 4617 10415 4675 10421
rect 5074 10412 5080 10424
rect 5132 10412 5138 10464
rect 5169 10455 5227 10461
rect 5169 10421 5181 10455
rect 5215 10452 5227 10455
rect 5350 10452 5356 10464
rect 5215 10424 5356 10452
rect 5215 10421 5227 10424
rect 5169 10415 5227 10421
rect 5350 10412 5356 10424
rect 5408 10412 5414 10464
rect 5445 10455 5503 10461
rect 5445 10421 5457 10455
rect 5491 10452 5503 10455
rect 6454 10452 6460 10464
rect 5491 10424 6460 10452
rect 5491 10421 5503 10424
rect 5445 10415 5503 10421
rect 6454 10412 6460 10424
rect 6512 10412 6518 10464
rect 6546 10412 6552 10464
rect 6604 10452 6610 10464
rect 7852 10452 7880 10492
rect 8294 10452 8300 10464
rect 6604 10424 7880 10452
rect 8255 10424 8300 10452
rect 6604 10412 6610 10424
rect 8294 10412 8300 10424
rect 8352 10412 8358 10464
rect 8665 10455 8723 10461
rect 8665 10421 8677 10455
rect 8711 10452 8723 10455
rect 9324 10452 9352 10492
rect 10505 10489 10517 10492
rect 10551 10489 10563 10523
rect 10505 10483 10563 10489
rect 8711 10424 9352 10452
rect 9401 10455 9459 10461
rect 8711 10421 8723 10424
rect 8665 10415 8723 10421
rect 9401 10421 9413 10455
rect 9447 10452 9459 10455
rect 13538 10452 13544 10464
rect 9447 10424 13544 10452
rect 9447 10421 9459 10424
rect 9401 10415 9459 10421
rect 13538 10412 13544 10424
rect 13596 10412 13602 10464
rect 920 10362 9844 10384
rect 920 10310 2566 10362
rect 2618 10310 2630 10362
rect 2682 10310 2694 10362
rect 2746 10310 2758 10362
rect 2810 10310 2822 10362
rect 2874 10310 5666 10362
rect 5718 10310 5730 10362
rect 5782 10310 5794 10362
rect 5846 10310 5858 10362
rect 5910 10310 5922 10362
rect 5974 10310 8766 10362
rect 8818 10310 8830 10362
rect 8882 10310 8894 10362
rect 8946 10310 8958 10362
rect 9010 10310 9022 10362
rect 9074 10310 9844 10362
rect 920 10288 9844 10310
rect 2685 10251 2743 10257
rect 2685 10217 2697 10251
rect 2731 10248 2743 10251
rect 3786 10248 3792 10260
rect 2731 10220 3792 10248
rect 2731 10217 2743 10220
rect 2685 10211 2743 10217
rect 3786 10208 3792 10220
rect 3844 10208 3850 10260
rect 4062 10208 4068 10260
rect 4120 10248 4126 10260
rect 8573 10251 8631 10257
rect 8573 10248 8585 10251
rect 4120 10220 8585 10248
rect 4120 10208 4126 10220
rect 8573 10217 8585 10220
rect 8619 10217 8631 10251
rect 8573 10211 8631 10217
rect 8757 10251 8815 10257
rect 8757 10217 8769 10251
rect 8803 10248 8815 10251
rect 9214 10248 9220 10260
rect 8803 10220 9220 10248
rect 8803 10217 8815 10220
rect 8757 10211 8815 10217
rect 9214 10208 9220 10220
rect 9272 10208 9278 10260
rect 2406 10140 2412 10192
rect 2464 10180 2470 10192
rect 2961 10183 3019 10189
rect 2961 10180 2973 10183
rect 2464 10152 2973 10180
rect 2464 10140 2470 10152
rect 2961 10149 2973 10152
rect 3007 10149 3019 10183
rect 3602 10180 3608 10192
rect 3563 10152 3608 10180
rect 2961 10143 3019 10149
rect 3602 10140 3608 10152
rect 3660 10140 3666 10192
rect 3697 10183 3755 10189
rect 3697 10149 3709 10183
rect 3743 10149 3755 10183
rect 3697 10143 3755 10149
rect 2130 10072 2136 10124
rect 2188 10112 2194 10124
rect 3712 10112 3740 10143
rect 5258 10140 5264 10192
rect 5316 10180 5322 10192
rect 6086 10180 6092 10192
rect 5316 10152 6092 10180
rect 5316 10140 5322 10152
rect 6086 10140 6092 10152
rect 6144 10140 6150 10192
rect 6273 10183 6331 10189
rect 6273 10149 6285 10183
rect 6319 10180 6331 10183
rect 6362 10180 6368 10192
rect 6319 10152 6368 10180
rect 6319 10149 6331 10152
rect 6273 10143 6331 10149
rect 6362 10140 6368 10152
rect 6420 10140 6426 10192
rect 7834 10140 7840 10192
rect 7892 10180 7898 10192
rect 8113 10183 8171 10189
rect 8113 10180 8125 10183
rect 7892 10152 8125 10180
rect 7892 10140 7898 10152
rect 8113 10149 8125 10152
rect 8159 10149 8171 10183
rect 8113 10143 8171 10149
rect 8386 10140 8392 10192
rect 8444 10140 8450 10192
rect 3973 10115 4031 10121
rect 3973 10112 3985 10115
rect 2188 10084 2912 10112
rect 3712 10084 3985 10112
rect 2188 10072 2194 10084
rect 2884 10053 2912 10084
rect 3973 10081 3985 10084
rect 4019 10081 4031 10115
rect 4338 10112 4344 10124
rect 4299 10084 4344 10112
rect 3973 10075 4031 10081
rect 4338 10072 4344 10084
rect 4396 10072 4402 10124
rect 6730 10072 6736 10124
rect 6788 10112 6794 10124
rect 8404 10112 8432 10140
rect 9306 10112 9312 10124
rect 6788 10084 8432 10112
rect 9267 10084 9312 10112
rect 6788 10072 6794 10084
rect 9306 10072 9312 10084
rect 9364 10072 9370 10124
rect 2593 10047 2651 10053
rect 2593 10044 2605 10047
rect 2148 10016 2605 10044
rect 2148 9988 2176 10016
rect 2593 10013 2605 10016
rect 2639 10013 2651 10047
rect 2593 10007 2651 10013
rect 2869 10047 2927 10053
rect 2869 10013 2881 10047
rect 2915 10044 2927 10047
rect 2958 10044 2964 10056
rect 2915 10016 2964 10044
rect 2915 10013 2927 10016
rect 2869 10007 2927 10013
rect 2958 10004 2964 10016
rect 3016 10004 3022 10056
rect 3145 10047 3203 10053
rect 3145 10013 3157 10047
rect 3191 10044 3203 10047
rect 3234 10044 3240 10056
rect 3191 10016 3240 10044
rect 3191 10013 3203 10016
rect 3145 10007 3203 10013
rect 3234 10004 3240 10016
rect 3292 10004 3298 10056
rect 3421 10047 3479 10053
rect 3421 10013 3433 10047
rect 3467 10044 3479 10047
rect 3605 10047 3663 10053
rect 3605 10044 3617 10047
rect 3467 10016 3617 10044
rect 3467 10013 3479 10016
rect 3421 10007 3479 10013
rect 3605 10013 3617 10016
rect 3651 10013 3663 10047
rect 3878 10044 3884 10056
rect 3839 10016 3884 10044
rect 3605 10007 3663 10013
rect 3878 10004 3884 10016
rect 3936 10004 3942 10056
rect 5350 10004 5356 10056
rect 5408 10044 5414 10056
rect 5813 10047 5871 10053
rect 5813 10044 5825 10047
rect 5408 10016 5825 10044
rect 5408 10004 5414 10016
rect 5813 10013 5825 10016
rect 5859 10013 5871 10047
rect 6362 10044 6368 10056
rect 6323 10016 6368 10044
rect 5813 10007 5871 10013
rect 6362 10004 6368 10016
rect 6420 10004 6426 10056
rect 7926 10004 7932 10056
rect 7984 10044 7990 10056
rect 8389 10047 8447 10053
rect 8389 10044 8401 10047
rect 7984 10016 8401 10044
rect 7984 10004 7990 10016
rect 8389 10013 8401 10016
rect 8435 10013 8447 10047
rect 8389 10007 8447 10013
rect 8570 10004 8576 10056
rect 8628 10044 8634 10056
rect 9125 10047 9183 10053
rect 9125 10044 9137 10047
rect 8628 10016 9137 10044
rect 8628 10004 8634 10016
rect 9125 10013 9137 10016
rect 9171 10013 9183 10047
rect 9125 10007 9183 10013
rect 2130 9936 2136 9988
rect 2188 9936 2194 9988
rect 3252 9948 4016 9976
rect 2409 9911 2467 9917
rect 2409 9877 2421 9911
rect 2455 9908 2467 9911
rect 2958 9908 2964 9920
rect 2455 9880 2964 9908
rect 2455 9877 2467 9880
rect 2409 9871 2467 9877
rect 2958 9868 2964 9880
rect 3016 9868 3022 9920
rect 3252 9917 3280 9948
rect 3237 9911 3295 9917
rect 3237 9877 3249 9911
rect 3283 9877 3295 9911
rect 3237 9871 3295 9877
rect 3418 9868 3424 9920
rect 3476 9908 3482 9920
rect 3694 9908 3700 9920
rect 3476 9880 3700 9908
rect 3476 9868 3482 9880
rect 3694 9868 3700 9880
rect 3752 9868 3758 9920
rect 3988 9908 4016 9948
rect 4614 9936 4620 9988
rect 4672 9976 4678 9988
rect 4672 9948 4738 9976
rect 4672 9936 4678 9948
rect 6178 9936 6184 9988
rect 6236 9976 6242 9988
rect 6641 9979 6699 9985
rect 6641 9976 6653 9979
rect 6236 9948 6653 9976
rect 6236 9936 6242 9948
rect 6641 9945 6653 9948
rect 6687 9945 6699 9979
rect 6641 9939 6699 9945
rect 6730 9936 6736 9988
rect 6788 9976 6794 9988
rect 8202 9976 8208 9988
rect 6788 9962 7130 9976
rect 7866 9962 8208 9976
rect 6788 9948 7144 9962
rect 6788 9936 6794 9948
rect 5626 9908 5632 9920
rect 3988 9880 5632 9908
rect 5626 9868 5632 9880
rect 5684 9868 5690 9920
rect 6454 9868 6460 9920
rect 6512 9908 6518 9920
rect 7006 9908 7012 9920
rect 6512 9880 7012 9908
rect 6512 9868 6518 9880
rect 7006 9868 7012 9880
rect 7064 9868 7070 9920
rect 7116 9908 7144 9948
rect 7852 9948 8208 9962
rect 7852 9908 7880 9948
rect 8202 9936 8208 9948
rect 8260 9936 8266 9988
rect 7116 9880 7880 9908
rect 9214 9868 9220 9920
rect 9272 9908 9278 9920
rect 9272 9880 9317 9908
rect 9272 9868 9278 9880
rect 920 9818 9844 9840
rect 920 9766 4116 9818
rect 4168 9766 4180 9818
rect 4232 9766 4244 9818
rect 4296 9766 4308 9818
rect 4360 9766 4372 9818
rect 4424 9766 7216 9818
rect 7268 9766 7280 9818
rect 7332 9766 7344 9818
rect 7396 9766 7408 9818
rect 7460 9766 7472 9818
rect 7524 9766 9844 9818
rect 920 9744 9844 9766
rect 10505 9775 10563 9781
rect 10505 9741 10517 9775
rect 10551 9772 10563 9775
rect 13814 9772 13820 9784
rect 10551 9744 13820 9772
rect 10551 9741 10563 9744
rect 10505 9735 10563 9741
rect 13814 9732 13820 9744
rect 13872 9732 13878 9784
rect 2958 9664 2964 9716
rect 3016 9704 3022 9716
rect 3234 9704 3240 9716
rect 3016 9676 3240 9704
rect 3016 9664 3022 9676
rect 3234 9664 3240 9676
rect 3292 9664 3298 9716
rect 4522 9704 4528 9716
rect 3436 9676 4528 9704
rect 2774 9636 2780 9648
rect 2700 9608 2780 9636
rect 1026 9528 1032 9580
rect 1084 9568 1090 9580
rect 1489 9571 1547 9577
rect 1489 9568 1501 9571
rect 1084 9540 1501 9568
rect 1084 9528 1090 9540
rect 1489 9537 1501 9540
rect 1535 9537 1547 9571
rect 1489 9531 1547 9537
rect 1765 9571 1823 9577
rect 1765 9537 1777 9571
rect 1811 9537 1823 9571
rect 2406 9568 2412 9580
rect 2367 9540 2412 9568
rect 1765 9531 1823 9537
rect 1118 9460 1124 9512
rect 1176 9500 1182 9512
rect 1780 9500 1808 9531
rect 2406 9528 2412 9540
rect 2464 9528 2470 9580
rect 2700 9577 2728 9608
rect 2774 9596 2780 9608
rect 2832 9596 2838 9648
rect 3053 9639 3111 9645
rect 3053 9605 3065 9639
rect 3099 9636 3111 9639
rect 3436 9636 3464 9676
rect 4522 9664 4528 9676
rect 4580 9664 4586 9716
rect 4617 9707 4675 9713
rect 4617 9673 4629 9707
rect 4663 9704 4675 9707
rect 4798 9704 4804 9716
rect 4663 9676 4804 9704
rect 4663 9673 4675 9676
rect 4617 9667 4675 9673
rect 4798 9664 4804 9676
rect 4856 9664 4862 9716
rect 5353 9707 5411 9713
rect 5353 9673 5365 9707
rect 5399 9673 5411 9707
rect 5353 9667 5411 9673
rect 3099 9608 3464 9636
rect 3099 9605 3111 9608
rect 3053 9599 3111 9605
rect 3694 9596 3700 9648
rect 3752 9596 3758 9648
rect 4430 9596 4436 9648
rect 4488 9636 4494 9648
rect 5368 9636 5396 9667
rect 5626 9664 5632 9716
rect 5684 9704 5690 9716
rect 5684 9676 7788 9704
rect 5684 9664 5690 9676
rect 4488 9608 5396 9636
rect 5644 9608 6408 9636
rect 7760 9622 7788 9676
rect 7926 9664 7932 9716
rect 7984 9704 7990 9716
rect 9122 9704 9128 9716
rect 7984 9676 9128 9704
rect 7984 9664 7990 9676
rect 9122 9664 9128 9676
rect 9180 9664 9186 9716
rect 9306 9704 9312 9716
rect 9267 9676 9312 9704
rect 9306 9664 9312 9676
rect 9364 9664 9370 9716
rect 4488 9596 4494 9608
rect 2685 9571 2743 9577
rect 2685 9537 2697 9571
rect 2731 9537 2743 9571
rect 2685 9531 2743 9537
rect 4338 9528 4344 9580
rect 4396 9568 4402 9580
rect 4801 9571 4859 9577
rect 4801 9568 4813 9571
rect 4396 9540 4813 9568
rect 4396 9528 4402 9540
rect 4801 9537 4813 9540
rect 4847 9537 4859 9571
rect 4801 9531 4859 9537
rect 4893 9571 4951 9577
rect 4893 9537 4905 9571
rect 4939 9568 4951 9571
rect 5074 9568 5080 9580
rect 4939 9540 5080 9568
rect 4939 9537 4951 9540
rect 4893 9531 4951 9537
rect 5074 9528 5080 9540
rect 5132 9528 5138 9580
rect 5644 9577 5672 9608
rect 5629 9571 5687 9577
rect 5629 9568 5641 9571
rect 5184 9540 5641 9568
rect 1176 9472 1808 9500
rect 2777 9503 2835 9509
rect 1176 9460 1182 9472
rect 2777 9469 2789 9503
rect 2823 9500 2835 9503
rect 3050 9500 3056 9512
rect 2823 9472 3056 9500
rect 2823 9469 2835 9472
rect 2777 9463 2835 9469
rect 3050 9460 3056 9472
rect 3108 9460 3114 9512
rect 4062 9460 4068 9512
rect 4120 9500 4126 9512
rect 5184 9500 5212 9540
rect 5629 9537 5641 9540
rect 5675 9537 5687 9571
rect 5810 9568 5816 9580
rect 5771 9540 5816 9568
rect 5629 9531 5687 9537
rect 5810 9528 5816 9540
rect 5868 9528 5874 9580
rect 5994 9568 6000 9580
rect 5955 9540 6000 9568
rect 5994 9528 6000 9540
rect 6052 9528 6058 9580
rect 6380 9577 6408 9608
rect 6365 9571 6423 9577
rect 6365 9537 6377 9571
rect 6411 9537 6423 9571
rect 6365 9531 6423 9537
rect 6914 9528 6920 9580
rect 6972 9568 6978 9580
rect 7374 9568 7380 9580
rect 6972 9540 7380 9568
rect 6972 9528 6978 9540
rect 7374 9528 7380 9540
rect 7432 9528 7438 9580
rect 8849 9571 8907 9577
rect 8849 9537 8861 9571
rect 8895 9537 8907 9571
rect 8849 9531 8907 9537
rect 6825 9503 6883 9509
rect 6825 9500 6837 9503
rect 4120 9472 5212 9500
rect 5276 9472 6837 9500
rect 4120 9460 4126 9472
rect 1946 9392 1952 9444
rect 2004 9432 2010 9444
rect 2225 9435 2283 9441
rect 2225 9432 2237 9435
rect 2004 9404 2237 9432
rect 2004 9392 2010 9404
rect 2225 9401 2237 9404
rect 2271 9401 2283 9435
rect 2225 9395 2283 9401
rect 2501 9435 2559 9441
rect 2501 9401 2513 9435
rect 2547 9432 2559 9435
rect 2682 9432 2688 9444
rect 2547 9404 2688 9432
rect 2547 9401 2559 9404
rect 2501 9395 2559 9401
rect 2682 9392 2688 9404
rect 2740 9392 2746 9444
rect 4154 9392 4160 9444
rect 4212 9432 4218 9444
rect 5276 9432 5304 9472
rect 6825 9469 6837 9472
rect 6871 9469 6883 9503
rect 6825 9463 6883 9469
rect 7009 9503 7067 9509
rect 7009 9469 7021 9503
rect 7055 9500 7067 9503
rect 7098 9500 7104 9512
rect 7055 9472 7104 9500
rect 7055 9469 7067 9472
rect 7009 9463 7067 9469
rect 7098 9460 7104 9472
rect 7156 9460 7162 9512
rect 4212 9404 5304 9432
rect 4212 9392 4218 9404
rect 5810 9392 5816 9444
rect 5868 9392 5874 9444
rect 1305 9367 1363 9373
rect 1305 9333 1317 9367
rect 1351 9364 1363 9367
rect 1394 9364 1400 9376
rect 1351 9336 1400 9364
rect 1351 9333 1363 9336
rect 1305 9327 1363 9333
rect 1394 9324 1400 9336
rect 1452 9324 1458 9376
rect 1578 9364 1584 9376
rect 1539 9336 1584 9364
rect 1578 9324 1584 9336
rect 1636 9324 1642 9376
rect 1762 9324 1768 9376
rect 1820 9364 1826 9376
rect 2041 9367 2099 9373
rect 2041 9364 2053 9367
rect 1820 9336 2053 9364
rect 1820 9324 1826 9336
rect 2041 9333 2053 9336
rect 2087 9333 2099 9367
rect 2041 9327 2099 9333
rect 3602 9324 3608 9376
rect 3660 9364 3666 9376
rect 4338 9364 4344 9376
rect 3660 9336 4344 9364
rect 3660 9324 3666 9336
rect 4338 9324 4344 9336
rect 4396 9324 4402 9376
rect 4522 9364 4528 9376
rect 4483 9336 4528 9364
rect 4522 9324 4528 9336
rect 4580 9324 4586 9376
rect 4706 9324 4712 9376
rect 4764 9364 4770 9376
rect 4985 9367 5043 9373
rect 4985 9364 4997 9367
rect 4764 9336 4997 9364
rect 4764 9324 4770 9336
rect 4985 9333 4997 9336
rect 5031 9364 5043 9367
rect 5828 9364 5856 9392
rect 6454 9364 6460 9376
rect 5031 9336 6460 9364
rect 5031 9333 5043 9336
rect 4985 9327 5043 9333
rect 6454 9324 6460 9336
rect 6512 9324 6518 9376
rect 6730 9324 6736 9376
rect 6788 9364 6794 9376
rect 8864 9364 8892 9531
rect 6788 9336 8892 9364
rect 6788 9324 6794 9336
rect 920 9274 9844 9296
rect 920 9222 2566 9274
rect 2618 9222 2630 9274
rect 2682 9222 2694 9274
rect 2746 9222 2758 9274
rect 2810 9222 2822 9274
rect 2874 9222 5666 9274
rect 5718 9222 5730 9274
rect 5782 9222 5794 9274
rect 5846 9222 5858 9274
rect 5910 9222 5922 9274
rect 5974 9222 8766 9274
rect 8818 9222 8830 9274
rect 8882 9222 8894 9274
rect 8946 9222 8958 9274
rect 9010 9222 9022 9274
rect 9074 9222 9844 9274
rect 920 9200 9844 9222
rect 1489 9163 1547 9169
rect 1489 9129 1501 9163
rect 1535 9160 1547 9163
rect 1535 9132 2176 9160
rect 1535 9129 1547 9132
rect 1489 9123 1547 9129
rect 1854 9092 1860 9104
rect 1815 9064 1860 9092
rect 1854 9052 1860 9064
rect 1912 9052 1918 9104
rect 2038 9092 2044 9104
rect 1999 9064 2044 9092
rect 2038 9052 2044 9064
rect 2096 9052 2102 9104
rect 2148 9092 2176 9132
rect 2314 9120 2320 9172
rect 2372 9160 2378 9172
rect 2685 9163 2743 9169
rect 2685 9160 2697 9163
rect 2372 9132 2697 9160
rect 2372 9120 2378 9132
rect 2685 9129 2697 9132
rect 2731 9129 2743 9163
rect 3510 9160 3516 9172
rect 2685 9123 2743 9129
rect 3160 9132 3516 9160
rect 3160 9092 3188 9132
rect 3510 9120 3516 9132
rect 3568 9120 3574 9172
rect 3605 9163 3663 9169
rect 3605 9129 3617 9163
rect 3651 9160 3663 9163
rect 3786 9160 3792 9172
rect 3651 9132 3792 9160
rect 3651 9129 3663 9132
rect 3605 9123 3663 9129
rect 3786 9120 3792 9132
rect 3844 9120 3850 9172
rect 4614 9160 4620 9172
rect 3896 9132 4620 9160
rect 2148 9064 3188 9092
rect 3237 9095 3295 9101
rect 3237 9061 3249 9095
rect 3283 9092 3295 9095
rect 3896 9092 3924 9132
rect 4614 9120 4620 9132
rect 4672 9120 4678 9172
rect 4798 9120 4804 9172
rect 4856 9160 4862 9172
rect 4856 9132 6500 9160
rect 4856 9120 4862 9132
rect 6472 9092 6500 9132
rect 6822 9120 6828 9172
rect 6880 9160 6886 9172
rect 7469 9163 7527 9169
rect 7469 9160 7481 9163
rect 6880 9132 7481 9160
rect 6880 9120 6886 9132
rect 7469 9129 7481 9132
rect 7515 9129 7527 9163
rect 8202 9160 8208 9172
rect 8163 9132 8208 9160
rect 7469 9123 7527 9129
rect 8202 9120 8208 9132
rect 8260 9120 8266 9172
rect 8478 9120 8484 9172
rect 8536 9160 8542 9172
rect 8757 9163 8815 9169
rect 8757 9160 8769 9163
rect 8536 9132 8769 9160
rect 8536 9120 8542 9132
rect 8757 9129 8769 9132
rect 8803 9129 8815 9163
rect 8757 9123 8815 9129
rect 7929 9095 7987 9101
rect 3283 9064 3924 9092
rect 5000 9064 5304 9092
rect 6472 9064 7052 9092
rect 3283 9061 3295 9064
rect 3237 9055 3295 9061
rect 2314 9024 2320 9036
rect 1780 8996 2320 9024
rect 1397 8959 1455 8965
rect 1397 8925 1409 8959
rect 1443 8956 1455 8959
rect 1670 8956 1676 8968
rect 1443 8928 1676 8956
rect 1443 8925 1455 8928
rect 1397 8919 1455 8925
rect 1670 8916 1676 8928
rect 1728 8916 1734 8968
rect 1780 8965 1808 8996
rect 2314 8984 2320 8996
rect 2372 8984 2378 9036
rect 2593 9027 2651 9033
rect 2593 8993 2605 9027
rect 2639 9024 2651 9027
rect 3326 9024 3332 9036
rect 2639 8996 3332 9024
rect 2639 8993 2651 8996
rect 2593 8987 2651 8993
rect 1765 8959 1823 8965
rect 1765 8925 1777 8959
rect 1811 8925 1823 8959
rect 2222 8956 2228 8968
rect 2183 8928 2228 8956
rect 1765 8919 1823 8925
rect 2222 8916 2228 8928
rect 2280 8916 2286 8968
rect 2884 8965 2912 8996
rect 3326 8984 3332 8996
rect 3384 8984 3390 9036
rect 2869 8959 2927 8965
rect 2869 8925 2881 8959
rect 2915 8956 2927 8959
rect 3142 8956 3148 8968
rect 2915 8928 2949 8956
rect 3103 8928 3148 8956
rect 2915 8925 2927 8928
rect 2869 8919 2927 8925
rect 3142 8916 3148 8928
rect 3200 8916 3206 8968
rect 3421 8959 3479 8965
rect 3421 8925 3433 8959
rect 3467 8956 3479 8959
rect 3602 8956 3608 8968
rect 3467 8928 3608 8956
rect 3467 8925 3479 8928
rect 3421 8919 3479 8925
rect 3602 8916 3608 8928
rect 3660 8916 3666 8968
rect 3789 8959 3847 8965
rect 3789 8925 3801 8959
rect 3835 8925 3847 8959
rect 3789 8919 3847 8925
rect 3050 8848 3056 8900
rect 3108 8888 3114 8900
rect 3326 8888 3332 8900
rect 3108 8860 3332 8888
rect 3108 8848 3114 8860
rect 3326 8848 3332 8860
rect 3384 8848 3390 8900
rect 3804 8888 3832 8919
rect 4062 8916 4068 8968
rect 4120 8956 4126 8968
rect 4341 8959 4399 8965
rect 4120 8928 4165 8956
rect 4120 8916 4126 8928
rect 4341 8925 4353 8959
rect 4387 8925 4399 8959
rect 4341 8919 4399 8925
rect 4617 8959 4675 8965
rect 4617 8925 4629 8959
rect 4663 8956 4675 8959
rect 4890 8956 4896 8968
rect 4663 8928 4896 8956
rect 4663 8925 4675 8928
rect 4617 8919 4675 8925
rect 4246 8888 4252 8900
rect 3712 8860 4252 8888
rect 3712 8832 3740 8860
rect 4246 8848 4252 8860
rect 4304 8848 4310 8900
rect 4356 8888 4384 8919
rect 4890 8916 4896 8928
rect 4948 8916 4954 8968
rect 5000 8888 5028 9064
rect 5166 9024 5172 9036
rect 5224 9033 5230 9036
rect 5133 8996 5172 9024
rect 5166 8984 5172 8996
rect 5224 8987 5233 9033
rect 5224 8984 5230 8987
rect 5077 8959 5135 8965
rect 5077 8925 5089 8959
rect 5123 8956 5135 8959
rect 5276 8956 5304 9064
rect 5537 9027 5595 9033
rect 5537 8993 5549 9027
rect 5583 9024 5595 9027
rect 6178 9024 6184 9036
rect 5583 8996 6184 9024
rect 5583 8993 5595 8996
rect 5537 8987 5595 8993
rect 6178 8984 6184 8996
rect 6236 8984 6242 9036
rect 7024 9024 7052 9064
rect 7929 9061 7941 9095
rect 7975 9092 7987 9095
rect 10134 9092 10140 9104
rect 7975 9064 10140 9092
rect 7975 9061 7987 9064
rect 7929 9055 7987 9061
rect 10134 9052 10140 9064
rect 10192 9052 10198 9104
rect 8662 9024 8668 9036
rect 7024 8996 8668 9024
rect 8662 8984 8668 8996
rect 8720 8984 8726 9036
rect 9306 9024 9312 9036
rect 9267 8996 9312 9024
rect 9306 8984 9312 8996
rect 9364 8984 9370 9036
rect 5626 8956 5632 8968
rect 5123 8928 5212 8956
rect 5276 8928 5632 8956
rect 5123 8925 5135 8928
rect 5077 8919 5135 8925
rect 5184 8900 5212 8928
rect 5626 8916 5632 8928
rect 5684 8916 5690 8968
rect 7006 8956 7012 8968
rect 6967 8928 7012 8956
rect 7006 8916 7012 8928
rect 7064 8916 7070 8968
rect 7742 8956 7748 8968
rect 7703 8928 7748 8956
rect 7742 8916 7748 8928
rect 7800 8916 7806 8968
rect 7834 8916 7840 8968
rect 7892 8956 7898 8968
rect 8113 8959 8171 8965
rect 8113 8956 8125 8959
rect 7892 8928 8125 8956
rect 7892 8916 7898 8928
rect 8113 8925 8125 8928
rect 8159 8925 8171 8959
rect 8113 8919 8171 8925
rect 8202 8916 8208 8968
rect 8260 8956 8266 8968
rect 9125 8959 9183 8965
rect 9125 8956 9137 8959
rect 8260 8928 9137 8956
rect 8260 8916 8266 8928
rect 9125 8925 9137 8928
rect 9171 8925 9183 8959
rect 9125 8919 9183 8925
rect 4356 8860 5028 8888
rect 5166 8848 5172 8900
rect 5224 8848 5230 8900
rect 5902 8848 5908 8900
rect 5960 8848 5966 8900
rect 6914 8848 6920 8900
rect 6972 8888 6978 8900
rect 9217 8891 9275 8897
rect 9217 8888 9229 8891
rect 6972 8860 9229 8888
rect 6972 8848 6978 8860
rect 9217 8857 9229 8860
rect 9263 8857 9275 8891
rect 9217 8851 9275 8857
rect 13446 8848 13452 8900
rect 13504 8888 13510 8900
rect 22370 8888 22376 8900
rect 13504 8860 22376 8888
rect 13504 8848 13510 8860
rect 22370 8848 22376 8860
rect 22428 8848 22434 8900
rect 2958 8780 2964 8832
rect 3016 8820 3022 8832
rect 3016 8792 3061 8820
rect 3016 8780 3022 8792
rect 3694 8780 3700 8832
rect 3752 8780 3758 8832
rect 3878 8820 3884 8832
rect 3839 8792 3884 8820
rect 3878 8780 3884 8792
rect 3936 8780 3942 8832
rect 3970 8780 3976 8832
rect 4028 8820 4034 8832
rect 4157 8823 4215 8829
rect 4157 8820 4169 8823
rect 4028 8792 4169 8820
rect 4028 8780 4034 8792
rect 4157 8789 4169 8792
rect 4203 8789 4215 8823
rect 4157 8783 4215 8789
rect 4433 8823 4491 8829
rect 4433 8789 4445 8823
rect 4479 8820 4491 8823
rect 4706 8820 4712 8832
rect 4479 8792 4712 8820
rect 4479 8789 4491 8792
rect 4433 8783 4491 8789
rect 4706 8780 4712 8792
rect 4764 8780 4770 8832
rect 4893 8823 4951 8829
rect 4893 8789 4905 8823
rect 4939 8820 4951 8823
rect 5810 8820 5816 8832
rect 4939 8792 5816 8820
rect 4939 8789 4951 8792
rect 4893 8783 4951 8789
rect 5810 8780 5816 8792
rect 5868 8780 5874 8832
rect 6270 8780 6276 8832
rect 6328 8820 6334 8832
rect 6546 8820 6552 8832
rect 6328 8792 6552 8820
rect 6328 8780 6334 8792
rect 6546 8780 6552 8792
rect 6604 8780 6610 8832
rect 8386 8780 8392 8832
rect 8444 8820 8450 8832
rect 8573 8823 8631 8829
rect 8573 8820 8585 8823
rect 8444 8792 8585 8820
rect 8444 8780 8450 8792
rect 8573 8789 8585 8792
rect 8619 8789 8631 8823
rect 8573 8783 8631 8789
rect 920 8730 9844 8752
rect 920 8678 4116 8730
rect 4168 8678 4180 8730
rect 4232 8678 4244 8730
rect 4296 8678 4308 8730
rect 4360 8678 4372 8730
rect 4424 8678 7216 8730
rect 7268 8678 7280 8730
rect 7332 8678 7344 8730
rect 7396 8678 7408 8730
rect 7460 8678 7472 8730
rect 7524 8678 9844 8730
rect 920 8656 9844 8678
rect 1486 8616 1492 8628
rect 1447 8588 1492 8616
rect 1486 8576 1492 8588
rect 1544 8576 1550 8628
rect 1854 8576 1860 8628
rect 1912 8616 1918 8628
rect 2038 8616 2044 8628
rect 1912 8588 2044 8616
rect 1912 8576 1918 8588
rect 2038 8576 2044 8588
rect 2096 8616 2102 8628
rect 2317 8619 2375 8625
rect 2317 8616 2329 8619
rect 2096 8588 2329 8616
rect 2096 8576 2102 8588
rect 2317 8585 2329 8588
rect 2363 8585 2375 8619
rect 2317 8579 2375 8585
rect 2409 8619 2467 8625
rect 2409 8585 2421 8619
rect 2455 8616 2467 8619
rect 2866 8616 2872 8628
rect 2455 8588 2872 8616
rect 2455 8585 2467 8588
rect 2409 8579 2467 8585
rect 2866 8576 2872 8588
rect 2924 8576 2930 8628
rect 4890 8576 4896 8628
rect 4948 8616 4954 8628
rect 5074 8616 5080 8628
rect 4948 8588 5080 8616
rect 4948 8576 4954 8588
rect 5074 8576 5080 8588
rect 5132 8616 5138 8628
rect 5169 8619 5227 8625
rect 5169 8616 5181 8619
rect 5132 8588 5181 8616
rect 5132 8576 5138 8588
rect 5169 8585 5181 8588
rect 5215 8585 5227 8619
rect 5169 8579 5227 8585
rect 5350 8576 5356 8628
rect 5408 8616 5414 8628
rect 5905 8619 5963 8625
rect 5905 8616 5917 8619
rect 5408 8588 5917 8616
rect 5408 8576 5414 8588
rect 5905 8585 5917 8588
rect 5951 8616 5963 8619
rect 6362 8616 6368 8628
rect 5951 8588 6368 8616
rect 5951 8585 5963 8588
rect 5905 8579 5963 8585
rect 6362 8576 6368 8588
rect 6420 8576 6426 8628
rect 6917 8619 6975 8625
rect 6917 8585 6929 8619
rect 6963 8616 6975 8619
rect 9582 8616 9588 8628
rect 6963 8588 9588 8616
rect 6963 8585 6975 8588
rect 6917 8579 6975 8585
rect 9582 8576 9588 8588
rect 9640 8576 9646 8628
rect 1210 8508 1216 8560
rect 1268 8548 1274 8560
rect 1268 8520 1716 8548
rect 1268 8508 1274 8520
rect 1688 8489 1716 8520
rect 2222 8508 2228 8560
rect 2280 8548 2286 8560
rect 2280 8520 2636 8548
rect 2280 8508 2286 8520
rect 1397 8483 1455 8489
rect 1397 8449 1409 8483
rect 1443 8449 1455 8483
rect 1397 8443 1455 8449
rect 1673 8483 1731 8489
rect 1673 8449 1685 8483
rect 1719 8449 1731 8483
rect 1673 8443 1731 8449
rect 1949 8483 2007 8489
rect 1949 8449 1961 8483
rect 1995 8480 2007 8483
rect 2314 8480 2320 8492
rect 1995 8452 2320 8480
rect 1995 8449 2007 8452
rect 1949 8443 2007 8449
rect 1412 8412 1440 8443
rect 2314 8440 2320 8452
rect 2372 8440 2378 8492
rect 2608 8489 2636 8520
rect 3050 8508 3056 8560
rect 3108 8508 3114 8560
rect 4798 8548 4804 8560
rect 4554 8520 4804 8548
rect 4798 8508 4804 8520
rect 4856 8548 4862 8560
rect 5445 8551 5503 8557
rect 5445 8548 5457 8551
rect 4856 8520 5457 8548
rect 4856 8508 4862 8520
rect 5445 8517 5457 8520
rect 5491 8517 5503 8551
rect 5445 8511 5503 8517
rect 5629 8551 5687 8557
rect 5629 8517 5641 8551
rect 5675 8548 5687 8551
rect 5994 8548 6000 8560
rect 5675 8520 6000 8548
rect 5675 8517 5687 8520
rect 5629 8511 5687 8517
rect 5994 8508 6000 8520
rect 6052 8508 6058 8560
rect 6178 8508 6184 8560
rect 6236 8548 6242 8560
rect 6273 8551 6331 8557
rect 6273 8548 6285 8551
rect 6236 8520 6285 8548
rect 6236 8508 6242 8520
rect 6273 8517 6285 8520
rect 6319 8517 6331 8551
rect 7098 8548 7104 8560
rect 6273 8511 6331 8517
rect 6380 8520 7104 8548
rect 2593 8483 2651 8489
rect 2593 8449 2605 8483
rect 2639 8449 2651 8483
rect 2958 8480 2964 8492
rect 2919 8452 2964 8480
rect 2593 8443 2651 8449
rect 2958 8440 2964 8452
rect 3016 8440 3022 8492
rect 2682 8412 2688 8424
rect 1412 8384 2688 8412
rect 2682 8372 2688 8384
rect 2740 8372 2746 8424
rect 3068 8421 3096 8508
rect 5261 8484 5319 8489
rect 5261 8483 5396 8484
rect 5074 8424 5080 8476
rect 5132 8464 5138 8476
rect 5132 8436 5177 8464
rect 5261 8449 5273 8483
rect 5307 8456 5396 8483
rect 5307 8449 5319 8456
rect 5261 8443 5319 8449
rect 5132 8424 5138 8436
rect 3053 8415 3111 8421
rect 3053 8381 3065 8415
rect 3099 8381 3111 8415
rect 3053 8375 3111 8381
rect 3329 8415 3387 8421
rect 3329 8381 3341 8415
rect 3375 8412 3387 8415
rect 3878 8412 3884 8424
rect 3375 8384 3884 8412
rect 3375 8381 3387 8384
rect 3329 8375 3387 8381
rect 3878 8372 3884 8384
rect 3936 8412 3942 8424
rect 4522 8412 4528 8424
rect 3936 8384 4528 8412
rect 3936 8372 3942 8384
rect 4522 8372 4528 8384
rect 4580 8372 4586 8424
rect 1762 8344 1768 8356
rect 1723 8316 1768 8344
rect 1762 8304 1768 8316
rect 1820 8304 1826 8356
rect 4430 8304 4436 8356
rect 4488 8344 4494 8356
rect 4893 8347 4951 8353
rect 4893 8344 4905 8347
rect 4488 8316 4905 8344
rect 4488 8304 4494 8316
rect 4893 8313 4905 8316
rect 4939 8313 4951 8347
rect 4893 8307 4951 8313
rect 1210 8276 1216 8288
rect 1171 8248 1216 8276
rect 1210 8236 1216 8248
rect 1268 8236 1274 8288
rect 2777 8279 2835 8285
rect 2777 8245 2789 8279
rect 2823 8276 2835 8279
rect 4522 8276 4528 8288
rect 2823 8248 4528 8276
rect 2823 8245 2835 8248
rect 2777 8239 2835 8245
rect 4522 8236 4528 8248
rect 4580 8236 4586 8288
rect 4801 8279 4859 8285
rect 4801 8245 4813 8279
rect 4847 8276 4859 8279
rect 5166 8276 5172 8288
rect 4847 8248 5172 8276
rect 4847 8245 4859 8248
rect 4801 8239 4859 8245
rect 5166 8236 5172 8248
rect 5224 8236 5230 8288
rect 5261 8279 5319 8285
rect 5261 8245 5273 8279
rect 5307 8276 5319 8279
rect 5368 8276 5396 8456
rect 5813 8483 5871 8489
rect 5813 8449 5825 8483
rect 5859 8480 5871 8483
rect 6380 8480 6408 8520
rect 7098 8508 7104 8520
rect 7156 8508 7162 8560
rect 8202 8508 8208 8560
rect 8260 8548 8266 8560
rect 13814 8548 13820 8560
rect 8260 8520 8892 8548
rect 8260 8508 8266 8520
rect 5859 8452 6408 8480
rect 5859 8449 5871 8452
rect 5813 8443 5871 8449
rect 6454 8440 6460 8492
rect 6512 8480 6518 8492
rect 6730 8480 6736 8492
rect 6512 8452 6557 8480
rect 6691 8452 6736 8480
rect 6512 8440 6518 8452
rect 6730 8440 6736 8452
rect 6788 8440 6794 8492
rect 6822 8440 6828 8492
rect 6880 8480 6886 8492
rect 7653 8483 7711 8489
rect 7653 8480 7665 8483
rect 6880 8452 7665 8480
rect 6880 8440 6886 8452
rect 7653 8449 7665 8452
rect 7699 8449 7711 8483
rect 7653 8443 7711 8449
rect 7745 8483 7803 8489
rect 7745 8449 7757 8483
rect 7791 8480 7803 8483
rect 8294 8480 8300 8492
rect 7791 8452 8300 8480
rect 7791 8449 7803 8452
rect 7745 8443 7803 8449
rect 8294 8440 8300 8452
rect 8352 8440 8358 8492
rect 8386 8440 8392 8492
rect 8444 8480 8450 8492
rect 8570 8480 8576 8492
rect 8444 8452 8489 8480
rect 8531 8452 8576 8480
rect 8444 8440 8450 8452
rect 8570 8440 8576 8452
rect 8628 8440 8634 8492
rect 8662 8440 8668 8492
rect 8720 8480 8726 8492
rect 8864 8489 8892 8520
rect 12406 8520 13820 8548
rect 8849 8483 8907 8489
rect 8720 8452 8765 8480
rect 8720 8440 8726 8452
rect 8849 8449 8861 8483
rect 8895 8449 8907 8483
rect 8849 8443 8907 8449
rect 6270 8372 6276 8424
rect 6328 8412 6334 8424
rect 6641 8415 6699 8421
rect 6641 8412 6653 8415
rect 6328 8384 6653 8412
rect 6328 8372 6334 8384
rect 6641 8381 6653 8384
rect 6687 8381 6699 8415
rect 6641 8375 6699 8381
rect 7006 8372 7012 8424
rect 7064 8412 7070 8424
rect 7101 8415 7159 8421
rect 7101 8412 7113 8415
rect 7064 8384 7113 8412
rect 7064 8372 7070 8384
rect 7101 8381 7113 8384
rect 7147 8381 7159 8415
rect 7101 8375 7159 8381
rect 7834 8372 7840 8424
rect 7892 8412 7898 8424
rect 8205 8415 8263 8421
rect 8205 8412 8217 8415
rect 7892 8384 8217 8412
rect 7892 8372 7898 8384
rect 8205 8381 8217 8384
rect 8251 8381 8263 8415
rect 8205 8375 8263 8381
rect 9309 8415 9367 8421
rect 9309 8381 9321 8415
rect 9355 8412 9367 8415
rect 10870 8412 10876 8424
rect 9355 8384 10876 8412
rect 9355 8381 9367 8384
rect 9309 8375 9367 8381
rect 10870 8372 10876 8384
rect 10928 8372 10934 8424
rect 5718 8304 5724 8356
rect 5776 8344 5782 8356
rect 6362 8344 6368 8356
rect 5776 8316 6368 8344
rect 5776 8304 5782 8316
rect 6362 8304 6368 8316
rect 6420 8304 6426 8356
rect 6546 8304 6552 8356
rect 6604 8344 6610 8356
rect 7561 8347 7619 8353
rect 7561 8344 7573 8347
rect 6604 8316 7573 8344
rect 6604 8304 6610 8316
rect 7561 8313 7573 8316
rect 7607 8313 7619 8347
rect 7561 8307 7619 8313
rect 7929 8347 7987 8353
rect 7929 8313 7941 8347
rect 7975 8344 7987 8347
rect 12406 8344 12434 8520
rect 13814 8508 13820 8520
rect 13872 8508 13878 8560
rect 7975 8316 12434 8344
rect 7975 8313 7987 8316
rect 7929 8307 7987 8313
rect 5307 8248 5396 8276
rect 5307 8245 5319 8248
rect 5261 8239 5319 8245
rect 5442 8236 5448 8288
rect 5500 8276 5506 8288
rect 8478 8276 8484 8288
rect 5500 8248 8484 8276
rect 5500 8236 5506 8248
rect 8478 8236 8484 8248
rect 8536 8236 8542 8288
rect 920 8186 9844 8208
rect 920 8134 2566 8186
rect 2618 8134 2630 8186
rect 2682 8134 2694 8186
rect 2746 8134 2758 8186
rect 2810 8134 2822 8186
rect 2874 8134 5666 8186
rect 5718 8134 5730 8186
rect 5782 8134 5794 8186
rect 5846 8134 5858 8186
rect 5910 8134 5922 8186
rect 5974 8134 8766 8186
rect 8818 8134 8830 8186
rect 8882 8134 8894 8186
rect 8946 8134 8958 8186
rect 9010 8134 9022 8186
rect 9074 8134 9844 8186
rect 920 8112 9844 8134
rect 1581 8075 1639 8081
rect 1581 8041 1593 8075
rect 1627 8072 1639 8075
rect 3050 8072 3056 8084
rect 1627 8044 3056 8072
rect 1627 8041 1639 8044
rect 1581 8035 1639 8041
rect 3050 8032 3056 8044
rect 3108 8032 3114 8084
rect 3142 8032 3148 8084
rect 3200 8072 3206 8084
rect 6178 8072 6184 8084
rect 3200 8044 6184 8072
rect 3200 8032 3206 8044
rect 6178 8032 6184 8044
rect 6236 8032 6242 8084
rect 7101 8075 7159 8081
rect 7101 8041 7113 8075
rect 7147 8072 7159 8075
rect 7742 8072 7748 8084
rect 7147 8044 7748 8072
rect 7147 8041 7159 8044
rect 7101 8035 7159 8041
rect 7742 8032 7748 8044
rect 7800 8032 7806 8084
rect 8018 8072 8024 8084
rect 7979 8044 8024 8072
rect 8018 8032 8024 8044
rect 8076 8032 8082 8084
rect 8757 8075 8815 8081
rect 8404 8044 8708 8072
rect 1489 8007 1547 8013
rect 1489 7973 1501 8007
rect 1535 8004 1547 8007
rect 2130 8004 2136 8016
rect 1535 7976 2136 8004
rect 1535 7973 1547 7976
rect 1489 7967 1547 7973
rect 2130 7964 2136 7976
rect 2188 7964 2194 8016
rect 2225 8007 2283 8013
rect 2225 7973 2237 8007
rect 2271 8004 2283 8007
rect 2406 8004 2412 8016
rect 2271 7976 2412 8004
rect 2271 7973 2283 7976
rect 2225 7967 2283 7973
rect 2406 7964 2412 7976
rect 2464 7964 2470 8016
rect 2501 8007 2559 8013
rect 2501 7973 2513 8007
rect 2547 8004 2559 8007
rect 3694 8004 3700 8016
rect 2547 7976 3700 8004
rect 2547 7973 2559 7976
rect 2501 7967 2559 7973
rect 3694 7964 3700 7976
rect 3752 7964 3758 8016
rect 3789 8007 3847 8013
rect 3789 7973 3801 8007
rect 3835 7973 3847 8007
rect 3789 7967 3847 7973
rect 2958 7896 2964 7948
rect 3016 7936 3022 7948
rect 3804 7936 3832 7967
rect 4430 7964 4436 8016
rect 4488 8004 4494 8016
rect 4890 8004 4896 8016
rect 4488 7976 4896 8004
rect 4488 7964 4494 7976
rect 4890 7964 4896 7976
rect 4948 7964 4954 8016
rect 7561 8007 7619 8013
rect 7561 7973 7573 8007
rect 7607 8004 7619 8007
rect 8404 8004 8432 8044
rect 7607 7976 8432 8004
rect 8481 8007 8539 8013
rect 7607 7973 7619 7976
rect 7561 7967 7619 7973
rect 8481 7973 8493 8007
rect 8527 7973 8539 8007
rect 8680 8004 8708 8044
rect 8757 8041 8769 8075
rect 8803 8072 8815 8075
rect 9214 8072 9220 8084
rect 8803 8044 9220 8072
rect 8803 8041 8815 8044
rect 8757 8035 8815 8041
rect 9214 8032 9220 8044
rect 9272 8032 9278 8084
rect 13538 8004 13544 8016
rect 8680 7976 13544 8004
rect 8481 7967 8539 7973
rect 3016 7908 3648 7936
rect 3804 7908 4292 7936
rect 3016 7896 3022 7908
rect 1762 7868 1768 7880
rect 1723 7840 1768 7868
rect 1762 7828 1768 7840
rect 1820 7828 1826 7880
rect 2038 7868 2044 7880
rect 1999 7840 2044 7868
rect 2038 7828 2044 7840
rect 2096 7828 2102 7880
rect 2409 7871 2467 7877
rect 2409 7837 2421 7871
rect 2455 7837 2467 7871
rect 2682 7868 2688 7880
rect 2643 7840 2688 7868
rect 2409 7831 2467 7837
rect 1026 7760 1032 7812
rect 1084 7800 1090 7812
rect 2424 7800 2452 7831
rect 2682 7828 2688 7840
rect 2740 7868 2746 7880
rect 3145 7871 3203 7877
rect 3145 7868 3157 7871
rect 2740 7840 3157 7868
rect 2740 7828 2746 7840
rect 3145 7837 3157 7840
rect 3191 7837 3203 7871
rect 3145 7831 3203 7837
rect 3620 7800 3648 7908
rect 3786 7828 3792 7880
rect 3844 7868 3850 7880
rect 4264 7877 4292 7908
rect 4522 7896 4528 7948
rect 4580 7936 4586 7948
rect 4801 7939 4859 7945
rect 4801 7936 4813 7939
rect 4580 7908 4813 7936
rect 4580 7896 4586 7908
rect 4801 7905 4813 7908
rect 4847 7905 4859 7939
rect 5442 7936 5448 7948
rect 4801 7899 4859 7905
rect 5000 7908 5448 7936
rect 3973 7871 4031 7877
rect 3973 7868 3985 7871
rect 3844 7840 3985 7868
rect 3844 7828 3850 7840
rect 3973 7837 3985 7840
rect 4019 7837 4031 7871
rect 3973 7831 4031 7837
rect 4249 7871 4307 7877
rect 4249 7837 4261 7871
rect 4295 7837 4307 7871
rect 4249 7831 4307 7837
rect 4709 7871 4767 7877
rect 4709 7837 4721 7871
rect 4755 7868 4767 7871
rect 5000 7868 5028 7908
rect 5442 7896 5448 7908
rect 5500 7896 5506 7948
rect 7926 7936 7932 7948
rect 7392 7908 7932 7936
rect 5166 7868 5172 7880
rect 4755 7840 5028 7868
rect 5127 7840 5172 7868
rect 4755 7837 4767 7840
rect 4709 7831 4767 7837
rect 5166 7828 5172 7840
rect 5224 7828 5230 7880
rect 6638 7868 6644 7880
rect 6599 7840 6644 7868
rect 6638 7828 6644 7840
rect 6696 7828 6702 7880
rect 7392 7877 7420 7908
rect 7926 7896 7932 7908
rect 7984 7896 7990 7948
rect 7377 7871 7435 7877
rect 7377 7837 7389 7871
rect 7423 7837 7435 7871
rect 7742 7868 7748 7880
rect 7703 7840 7748 7868
rect 7377 7831 7435 7837
rect 7742 7828 7748 7840
rect 7800 7828 7806 7880
rect 8297 7871 8355 7877
rect 8297 7837 8309 7871
rect 8343 7868 8355 7871
rect 8386 7868 8392 7880
rect 8343 7840 8392 7868
rect 8343 7837 8355 7840
rect 8297 7831 8355 7837
rect 8386 7828 8392 7840
rect 8444 7828 8450 7880
rect 8496 7868 8524 7967
rect 13538 7964 13544 7976
rect 13596 7964 13602 8016
rect 9306 7936 9312 7948
rect 9267 7908 9312 7936
rect 9306 7896 9312 7908
rect 9364 7896 9370 7948
rect 13630 7868 13636 7880
rect 8496 7840 13636 7868
rect 13630 7828 13636 7840
rect 13688 7828 13694 7880
rect 1084 7772 2360 7800
rect 2424 7772 3464 7800
rect 3620 7772 4844 7800
rect 1084 7760 1090 7772
rect 1118 7692 1124 7744
rect 1176 7732 1182 7744
rect 1213 7735 1271 7741
rect 1213 7732 1225 7735
rect 1176 7704 1225 7732
rect 1176 7692 1182 7704
rect 1213 7701 1225 7704
rect 1259 7701 1271 7735
rect 1213 7695 1271 7701
rect 1857 7735 1915 7741
rect 1857 7701 1869 7735
rect 1903 7732 1915 7735
rect 2222 7732 2228 7744
rect 1903 7704 2228 7732
rect 1903 7701 1915 7704
rect 1857 7695 1915 7701
rect 2222 7692 2228 7704
rect 2280 7692 2286 7744
rect 2332 7732 2360 7772
rect 3436 7744 3464 7772
rect 2961 7735 3019 7741
rect 2961 7732 2973 7735
rect 2332 7704 2973 7732
rect 2961 7701 2973 7704
rect 3007 7732 3019 7735
rect 3142 7732 3148 7744
rect 3007 7704 3148 7732
rect 3007 7701 3019 7704
rect 2961 7695 3019 7701
rect 3142 7692 3148 7704
rect 3200 7692 3206 7744
rect 3418 7732 3424 7744
rect 3379 7704 3424 7732
rect 3418 7692 3424 7704
rect 3476 7692 3482 7744
rect 3510 7692 3516 7744
rect 3568 7732 3574 7744
rect 4065 7735 4123 7741
rect 4065 7732 4077 7735
rect 3568 7704 4077 7732
rect 3568 7692 3574 7704
rect 4065 7701 4077 7704
rect 4111 7701 4123 7735
rect 4522 7732 4528 7744
rect 4483 7704 4528 7732
rect 4065 7695 4123 7701
rect 4522 7692 4528 7704
rect 4580 7692 4586 7744
rect 4816 7732 4844 7772
rect 5534 7760 5540 7812
rect 5592 7760 5598 7812
rect 6822 7760 6828 7812
rect 6880 7800 6886 7812
rect 6880 7772 12434 7800
rect 6880 7760 6886 7772
rect 8205 7735 8263 7741
rect 8205 7732 8217 7735
rect 4816 7704 8217 7732
rect 8205 7701 8217 7704
rect 8251 7701 8263 7735
rect 8205 7695 8263 7701
rect 8478 7692 8484 7744
rect 8536 7732 8542 7744
rect 9122 7732 9128 7744
rect 8536 7704 9128 7732
rect 8536 7692 8542 7704
rect 9122 7692 9128 7704
rect 9180 7692 9186 7744
rect 9214 7692 9220 7744
rect 9272 7732 9278 7744
rect 12406 7732 12434 7772
rect 13722 7732 13728 7744
rect 9272 7704 9317 7732
rect 12406 7704 13728 7732
rect 9272 7692 9278 7704
rect 13722 7692 13728 7704
rect 13780 7692 13786 7744
rect 920 7642 9844 7664
rect 920 7590 4116 7642
rect 4168 7590 4180 7642
rect 4232 7590 4244 7642
rect 4296 7590 4308 7642
rect 4360 7590 4372 7642
rect 4424 7590 7216 7642
rect 7268 7590 7280 7642
rect 7332 7590 7344 7642
rect 7396 7590 7408 7642
rect 7460 7590 7472 7642
rect 7524 7590 9844 7642
rect 13446 7624 13452 7676
rect 13504 7664 13510 7676
rect 22278 7664 22284 7676
rect 13504 7636 22284 7664
rect 13504 7624 13510 7636
rect 22278 7624 22284 7636
rect 22336 7624 22342 7676
rect 920 7568 9844 7590
rect 2130 7488 2136 7540
rect 2188 7528 2194 7540
rect 2869 7531 2927 7537
rect 2869 7528 2881 7531
rect 2188 7500 2881 7528
rect 2188 7488 2194 7500
rect 2869 7497 2881 7500
rect 2915 7497 2927 7531
rect 2869 7491 2927 7497
rect 3050 7488 3056 7540
rect 3108 7528 3114 7540
rect 3145 7531 3203 7537
rect 3145 7528 3157 7531
rect 3108 7500 3157 7528
rect 3108 7488 3114 7500
rect 3145 7497 3157 7500
rect 3191 7497 3203 7531
rect 3145 7491 3203 7497
rect 3234 7488 3240 7540
rect 3292 7528 3298 7540
rect 3292 7500 4384 7528
rect 3292 7488 3298 7500
rect 4356 7472 4384 7500
rect 4890 7488 4896 7540
rect 4948 7488 4954 7540
rect 4982 7488 4988 7540
rect 5040 7528 5046 7540
rect 5902 7528 5908 7540
rect 5040 7500 5908 7528
rect 5040 7488 5046 7500
rect 5902 7488 5908 7500
rect 5960 7488 5966 7540
rect 5997 7531 6055 7537
rect 5997 7497 6009 7531
rect 6043 7528 6055 7531
rect 7742 7528 7748 7540
rect 6043 7500 7748 7528
rect 6043 7497 6055 7500
rect 5997 7491 6055 7497
rect 7742 7488 7748 7500
rect 7800 7488 7806 7540
rect 7834 7488 7840 7540
rect 7892 7528 7898 7540
rect 8018 7528 8024 7540
rect 7892 7500 8024 7528
rect 7892 7488 7898 7500
rect 8018 7488 8024 7500
rect 8076 7488 8082 7540
rect 8478 7488 8484 7540
rect 8536 7528 8542 7540
rect 9125 7531 9183 7537
rect 9125 7528 9137 7531
rect 8536 7500 9137 7528
rect 8536 7488 8542 7500
rect 9125 7497 9137 7500
rect 9171 7497 9183 7531
rect 9125 7491 9183 7497
rect 1762 7420 1768 7472
rect 1820 7460 1826 7472
rect 1820 7432 2176 7460
rect 1820 7420 1826 7432
rect 1581 7395 1639 7401
rect 1581 7361 1593 7395
rect 1627 7392 1639 7395
rect 1627 7364 1992 7392
rect 1627 7361 1639 7364
rect 1581 7355 1639 7361
rect 1964 7265 1992 7364
rect 2148 7333 2176 7432
rect 4338 7420 4344 7472
rect 4396 7420 4402 7472
rect 4908 7446 4936 7488
rect 8110 7420 8116 7472
rect 8168 7420 8174 7472
rect 8570 7420 8576 7472
rect 8628 7460 8634 7472
rect 8628 7432 9260 7460
rect 8628 7420 8634 7432
rect 2501 7395 2559 7401
rect 2501 7361 2513 7395
rect 2547 7392 2559 7395
rect 2774 7392 2780 7404
rect 2547 7364 2636 7392
rect 2735 7364 2780 7392
rect 2547 7361 2559 7364
rect 2501 7355 2559 7361
rect 2133 7327 2191 7333
rect 2133 7293 2145 7327
rect 2179 7324 2191 7327
rect 2314 7324 2320 7336
rect 2179 7296 2320 7324
rect 2179 7293 2191 7296
rect 2133 7287 2191 7293
rect 2314 7284 2320 7296
rect 2372 7284 2378 7336
rect 1949 7259 2007 7265
rect 1949 7225 1961 7259
rect 1995 7256 2007 7259
rect 2406 7256 2412 7268
rect 1995 7228 2412 7256
rect 1995 7225 2007 7228
rect 1949 7219 2007 7225
rect 2406 7216 2412 7228
rect 2464 7216 2470 7268
rect 2608 7265 2636 7364
rect 2774 7352 2780 7364
rect 2832 7352 2838 7404
rect 3050 7392 3056 7404
rect 3011 7364 3056 7392
rect 3050 7352 3056 7364
rect 3108 7352 3114 7404
rect 3329 7395 3387 7401
rect 3329 7361 3341 7395
rect 3375 7361 3387 7395
rect 3329 7355 3387 7361
rect 3605 7395 3663 7401
rect 3605 7361 3617 7395
rect 3651 7392 3663 7395
rect 4062 7392 4068 7404
rect 3651 7364 3832 7392
rect 4023 7364 4068 7392
rect 3651 7361 3663 7364
rect 3605 7355 3663 7361
rect 2593 7259 2651 7265
rect 2593 7225 2605 7259
rect 2639 7225 2651 7259
rect 3344 7256 3372 7355
rect 3510 7284 3516 7336
rect 3568 7324 3574 7336
rect 3697 7327 3755 7333
rect 3697 7324 3709 7327
rect 3568 7296 3709 7324
rect 3568 7284 3574 7296
rect 3697 7293 3709 7296
rect 3743 7293 3755 7327
rect 3804 7324 3832 7364
rect 4062 7352 4068 7364
rect 4120 7352 4126 7404
rect 5537 7395 5595 7401
rect 5537 7361 5549 7395
rect 5583 7392 5595 7395
rect 5994 7392 6000 7404
rect 5583 7364 6000 7392
rect 5583 7361 5595 7364
rect 5537 7355 5595 7361
rect 5994 7352 6000 7364
rect 6052 7352 6058 7404
rect 6178 7392 6184 7404
rect 6139 7364 6184 7392
rect 6178 7352 6184 7364
rect 6236 7352 6242 7404
rect 8662 7392 8668 7404
rect 8623 7364 8668 7392
rect 8662 7352 8668 7364
rect 8720 7352 8726 7404
rect 9232 7401 9260 7432
rect 9217 7395 9275 7401
rect 9217 7361 9229 7395
rect 9263 7361 9275 7395
rect 9217 7355 9275 7361
rect 4522 7324 4528 7336
rect 3804 7296 4528 7324
rect 3697 7287 3755 7293
rect 4522 7284 4528 7296
rect 4580 7284 4586 7336
rect 6825 7327 6883 7333
rect 6825 7324 6837 7327
rect 5552 7296 6837 7324
rect 3602 7256 3608 7268
rect 2593 7219 2651 7225
rect 2746 7228 3004 7256
rect 3344 7228 3608 7256
rect 1394 7188 1400 7200
rect 1355 7160 1400 7188
rect 1394 7148 1400 7160
rect 1452 7148 1458 7200
rect 2317 7191 2375 7197
rect 2317 7157 2329 7191
rect 2363 7188 2375 7191
rect 2746 7188 2774 7228
rect 2363 7160 2774 7188
rect 2976 7188 3004 7228
rect 3602 7216 3608 7228
rect 3660 7216 3666 7268
rect 5074 7216 5080 7268
rect 5132 7256 5138 7268
rect 5350 7256 5356 7268
rect 5132 7228 5356 7256
rect 5132 7216 5138 7228
rect 5350 7216 5356 7228
rect 5408 7216 5414 7268
rect 3234 7188 3240 7200
rect 2976 7160 3240 7188
rect 2363 7157 2375 7160
rect 2317 7151 2375 7157
rect 3234 7148 3240 7160
rect 3292 7148 3298 7200
rect 3421 7191 3479 7197
rect 3421 7157 3433 7191
rect 3467 7188 3479 7191
rect 5552 7188 5580 7296
rect 6825 7293 6837 7296
rect 6871 7293 6883 7327
rect 7193 7327 7251 7333
rect 7193 7324 7205 7327
rect 6825 7287 6883 7293
rect 6932 7296 7205 7324
rect 5626 7216 5632 7268
rect 5684 7256 5690 7268
rect 6932 7256 6960 7296
rect 7193 7293 7205 7296
rect 7239 7324 7251 7327
rect 7558 7324 7564 7336
rect 7239 7296 7564 7324
rect 7239 7293 7251 7296
rect 7193 7287 7251 7293
rect 7558 7284 7564 7296
rect 7616 7284 7622 7336
rect 13814 7284 13820 7336
rect 13872 7324 13878 7336
rect 19426 7324 19432 7336
rect 13872 7296 19432 7324
rect 13872 7284 13878 7296
rect 19426 7284 19432 7296
rect 19484 7284 19490 7336
rect 5684 7228 6960 7256
rect 8849 7259 8907 7265
rect 5684 7216 5690 7228
rect 8849 7225 8861 7259
rect 8895 7256 8907 7259
rect 9030 7256 9036 7268
rect 8895 7228 9036 7256
rect 8895 7225 8907 7228
rect 8849 7219 8907 7225
rect 9030 7216 9036 7228
rect 9088 7216 9094 7268
rect 6454 7188 6460 7200
rect 3467 7160 5580 7188
rect 6415 7160 6460 7188
rect 3467 7157 3479 7160
rect 3421 7151 3479 7157
rect 6454 7148 6460 7160
rect 6512 7148 6518 7200
rect 6638 7188 6644 7200
rect 6599 7160 6644 7188
rect 6638 7148 6644 7160
rect 6696 7148 6702 7200
rect 9401 7191 9459 7197
rect 9401 7157 9413 7191
rect 9447 7188 9459 7191
rect 13722 7188 13728 7200
rect 9447 7160 13728 7188
rect 9447 7157 9459 7160
rect 9401 7151 9459 7157
rect 13722 7148 13728 7160
rect 13780 7148 13786 7200
rect 920 7098 9844 7120
rect 920 7046 2566 7098
rect 2618 7046 2630 7098
rect 2682 7046 2694 7098
rect 2746 7046 2758 7098
rect 2810 7046 2822 7098
rect 2874 7046 5666 7098
rect 5718 7046 5730 7098
rect 5782 7046 5794 7098
rect 5846 7046 5858 7098
rect 5910 7046 5922 7098
rect 5974 7046 8766 7098
rect 8818 7046 8830 7098
rect 8882 7046 8894 7098
rect 8946 7046 8958 7098
rect 9010 7046 9022 7098
rect 9074 7046 9844 7098
rect 920 7024 9844 7046
rect 2038 6944 2044 6996
rect 2096 6944 2102 6996
rect 2777 6987 2835 6993
rect 2777 6953 2789 6987
rect 2823 6984 2835 6987
rect 3053 6987 3111 6993
rect 3053 6984 3065 6987
rect 2823 6956 3065 6984
rect 2823 6953 2835 6956
rect 2777 6947 2835 6953
rect 3053 6953 3065 6956
rect 3099 6984 3111 6987
rect 4246 6984 4252 6996
rect 3099 6956 4252 6984
rect 3099 6953 3111 6956
rect 3053 6947 3111 6953
rect 4246 6944 4252 6956
rect 4304 6944 4310 6996
rect 5074 6944 5080 6996
rect 5132 6984 5138 6996
rect 5537 6987 5595 6993
rect 5537 6984 5549 6987
rect 5132 6956 5549 6984
rect 5132 6944 5138 6956
rect 5537 6953 5549 6956
rect 5583 6984 5595 6987
rect 6454 6984 6460 6996
rect 5583 6956 6460 6984
rect 5583 6953 5595 6956
rect 5537 6947 5595 6953
rect 6454 6944 6460 6956
rect 6512 6944 6518 6996
rect 7098 6944 7104 6996
rect 7156 6984 7162 6996
rect 7469 6987 7527 6993
rect 7469 6984 7481 6987
rect 7156 6956 7481 6984
rect 7156 6944 7162 6956
rect 7469 6953 7481 6956
rect 7515 6953 7527 6987
rect 7469 6947 7527 6953
rect 8757 6987 8815 6993
rect 8757 6953 8769 6987
rect 8803 6984 8815 6987
rect 9214 6984 9220 6996
rect 8803 6956 9220 6984
rect 8803 6953 8815 6956
rect 8757 6947 8815 6953
rect 9214 6944 9220 6956
rect 9272 6944 9278 6996
rect 2056 6916 2084 6944
rect 3510 6916 3516 6928
rect 2056 6888 3516 6916
rect 3510 6876 3516 6888
rect 3568 6876 3574 6928
rect 3694 6876 3700 6928
rect 3752 6916 3758 6928
rect 6638 6916 6644 6928
rect 3752 6888 6644 6916
rect 3752 6876 3758 6888
rect 6638 6876 6644 6888
rect 6696 6876 6702 6928
rect 8202 6876 8208 6928
rect 8260 6876 8266 6928
rect 1670 6848 1676 6860
rect 1504 6820 1676 6848
rect 1504 6789 1532 6820
rect 1670 6808 1676 6820
rect 1728 6808 1734 6860
rect 3237 6851 3295 6857
rect 3237 6848 3249 6851
rect 2424 6820 3249 6848
rect 1489 6783 1547 6789
rect 1489 6749 1501 6783
rect 1535 6749 1547 6783
rect 1762 6780 1768 6792
rect 1723 6752 1768 6780
rect 1489 6743 1547 6749
rect 1762 6740 1768 6752
rect 1820 6740 1826 6792
rect 2130 6780 2136 6792
rect 2091 6752 2136 6780
rect 2130 6740 2136 6752
rect 2188 6740 2194 6792
rect 2222 6740 2228 6792
rect 2280 6740 2286 6792
rect 2424 6789 2452 6820
rect 3237 6817 3249 6820
rect 3283 6848 3295 6851
rect 3973 6851 4031 6857
rect 3973 6848 3985 6851
rect 3283 6820 3985 6848
rect 3283 6817 3295 6820
rect 3237 6811 3295 6817
rect 3973 6817 3985 6820
rect 4019 6817 4031 6851
rect 3973 6811 4031 6817
rect 4246 6808 4252 6860
rect 4304 6848 4310 6860
rect 4982 6848 4988 6860
rect 4304 6820 4988 6848
rect 4304 6808 4310 6820
rect 4982 6808 4988 6820
rect 5040 6808 5046 6860
rect 5350 6808 5356 6860
rect 5408 6848 5414 6860
rect 5721 6851 5779 6857
rect 5721 6848 5733 6851
rect 5408 6820 5733 6848
rect 5408 6808 5414 6820
rect 5721 6817 5733 6820
rect 5767 6817 5779 6851
rect 5721 6811 5779 6817
rect 5810 6808 5816 6860
rect 5868 6848 5874 6860
rect 8220 6848 8248 6876
rect 9306 6848 9312 6860
rect 5868 6820 8248 6848
rect 9267 6820 9312 6848
rect 5868 6808 5874 6820
rect 9306 6808 9312 6820
rect 9364 6808 9370 6860
rect 2409 6783 2467 6789
rect 2409 6749 2421 6783
rect 2455 6749 2467 6783
rect 2409 6743 2467 6749
rect 2685 6783 2743 6789
rect 2685 6749 2697 6783
rect 2731 6780 2743 6783
rect 2777 6783 2835 6789
rect 2777 6780 2789 6783
rect 2731 6752 2789 6780
rect 2731 6749 2743 6752
rect 2685 6743 2743 6749
rect 2777 6749 2789 6752
rect 2823 6749 2835 6783
rect 2777 6743 2835 6749
rect 3878 6740 3884 6792
rect 3936 6780 3942 6792
rect 4157 6783 4215 6789
rect 4157 6780 4169 6783
rect 3936 6752 4169 6780
rect 3936 6740 3942 6752
rect 4157 6749 4169 6752
rect 4203 6749 4215 6783
rect 4157 6743 4215 6749
rect 4433 6783 4491 6789
rect 4433 6749 4445 6783
rect 4479 6780 4491 6783
rect 4522 6780 4528 6792
rect 4479 6752 4528 6780
rect 4479 6749 4491 6752
rect 4433 6743 4491 6749
rect 4522 6740 4528 6752
rect 4580 6740 4586 6792
rect 5261 6783 5319 6789
rect 5261 6749 5273 6783
rect 5307 6749 5319 6783
rect 5261 6743 5319 6749
rect 5997 6783 6055 6789
rect 5997 6749 6009 6783
rect 6043 6749 6055 6783
rect 5997 6743 6055 6749
rect 6181 6783 6239 6789
rect 6181 6749 6193 6783
rect 6227 6780 6239 6783
rect 6822 6780 6828 6792
rect 6227 6752 6828 6780
rect 6227 6749 6239 6752
rect 6181 6743 6239 6749
rect 2240 6712 2268 6740
rect 5276 6712 5304 6743
rect 5626 6712 5632 6724
rect 2240 6684 5632 6712
rect 5626 6672 5632 6684
rect 5684 6672 5690 6724
rect 6012 6712 6040 6743
rect 6822 6740 6828 6752
rect 6880 6740 6886 6792
rect 8202 6780 8208 6792
rect 8163 6752 8208 6780
rect 8202 6740 8208 6752
rect 8260 6740 8266 6792
rect 8294 6740 8300 6792
rect 8352 6780 8358 6792
rect 9122 6780 9128 6792
rect 8352 6752 8397 6780
rect 9083 6752 9128 6780
rect 8352 6740 8358 6752
rect 9122 6740 9128 6752
rect 9180 6740 9186 6792
rect 9217 6783 9275 6789
rect 9217 6749 9229 6783
rect 9263 6780 9275 6783
rect 9398 6780 9404 6792
rect 9263 6752 9404 6780
rect 9263 6749 9275 6752
rect 9217 6743 9275 6749
rect 9398 6740 9404 6752
rect 9456 6740 9462 6792
rect 5736 6684 6040 6712
rect 1305 6647 1363 6653
rect 1305 6613 1317 6647
rect 1351 6644 1363 6647
rect 1394 6644 1400 6656
rect 1351 6616 1400 6644
rect 1351 6613 1363 6616
rect 1305 6607 1363 6613
rect 1394 6604 1400 6616
rect 1452 6604 1458 6656
rect 1578 6644 1584 6656
rect 1539 6616 1584 6644
rect 1578 6604 1584 6616
rect 1636 6604 1642 6656
rect 1949 6647 2007 6653
rect 1949 6613 1961 6647
rect 1995 6644 2007 6647
rect 2038 6644 2044 6656
rect 1995 6616 2044 6644
rect 1995 6613 2007 6616
rect 1949 6607 2007 6613
rect 2038 6604 2044 6616
rect 2096 6604 2102 6656
rect 2222 6644 2228 6656
rect 2183 6616 2228 6644
rect 2222 6604 2228 6616
rect 2280 6604 2286 6656
rect 2501 6647 2559 6653
rect 2501 6613 2513 6647
rect 2547 6644 2559 6647
rect 2682 6644 2688 6656
rect 2547 6616 2688 6644
rect 2547 6613 2559 6616
rect 2501 6607 2559 6613
rect 2682 6604 2688 6616
rect 2740 6604 2746 6656
rect 2866 6604 2872 6656
rect 2924 6644 2930 6656
rect 3329 6647 3387 6653
rect 3329 6644 3341 6647
rect 2924 6616 3341 6644
rect 2924 6604 2930 6616
rect 3329 6613 3341 6616
rect 3375 6613 3387 6647
rect 3329 6607 3387 6613
rect 3510 6604 3516 6656
rect 3568 6644 3574 6656
rect 3605 6647 3663 6653
rect 3605 6644 3617 6647
rect 3568 6616 3617 6644
rect 3568 6604 3574 6616
rect 3605 6613 3617 6616
rect 3651 6613 3663 6647
rect 3605 6607 3663 6613
rect 3694 6604 3700 6656
rect 3752 6644 3758 6656
rect 3789 6647 3847 6653
rect 3789 6644 3801 6647
rect 3752 6616 3801 6644
rect 3752 6604 3758 6616
rect 3789 6613 3801 6616
rect 3835 6613 3847 6647
rect 3789 6607 3847 6613
rect 3973 6647 4031 6653
rect 3973 6613 3985 6647
rect 4019 6644 4031 6647
rect 5258 6644 5264 6656
rect 4019 6616 5264 6644
rect 4019 6613 4031 6616
rect 3973 6607 4031 6613
rect 5258 6604 5264 6616
rect 5316 6604 5322 6656
rect 5442 6604 5448 6656
rect 5500 6644 5506 6656
rect 5736 6644 5764 6684
rect 8110 6672 8116 6724
rect 8168 6712 8174 6724
rect 9582 6712 9588 6724
rect 8168 6684 9588 6712
rect 8168 6672 8174 6684
rect 9582 6672 9588 6684
rect 9640 6672 9646 6724
rect 5500 6616 5764 6644
rect 5813 6647 5871 6653
rect 5500 6604 5506 6616
rect 5813 6613 5825 6647
rect 5859 6644 5871 6647
rect 5902 6644 5908 6656
rect 5859 6616 5908 6644
rect 5859 6613 5871 6616
rect 5813 6607 5871 6613
rect 5902 6604 5908 6616
rect 5960 6604 5966 6656
rect 7650 6604 7656 6656
rect 7708 6644 7714 6656
rect 8021 6647 8079 6653
rect 8021 6644 8033 6647
rect 7708 6616 8033 6644
rect 7708 6604 7714 6616
rect 8021 6613 8033 6616
rect 8067 6613 8079 6647
rect 8021 6607 8079 6613
rect 8481 6647 8539 6653
rect 8481 6613 8493 6647
rect 8527 6644 8539 6647
rect 8527 6616 10456 6644
rect 8527 6613 8539 6616
rect 8481 6607 8539 6613
rect 920 6554 9844 6576
rect 920 6502 4116 6554
rect 4168 6502 4180 6554
rect 4232 6502 4244 6554
rect 4296 6502 4308 6554
rect 4360 6502 4372 6554
rect 4424 6502 7216 6554
rect 7268 6502 7280 6554
rect 7332 6502 7344 6554
rect 7396 6502 7408 6554
rect 7460 6502 7472 6554
rect 7524 6502 9844 6554
rect 920 6480 9844 6502
rect 1578 6440 1584 6452
rect 1539 6412 1584 6440
rect 1578 6400 1584 6412
rect 1636 6400 1642 6452
rect 2222 6440 2228 6452
rect 2183 6412 2228 6440
rect 2222 6400 2228 6412
rect 2280 6400 2286 6452
rect 3142 6400 3148 6452
rect 3200 6440 3206 6452
rect 3418 6440 3424 6452
rect 3200 6412 3424 6440
rect 3200 6400 3206 6412
rect 3418 6400 3424 6412
rect 3476 6400 3482 6452
rect 5166 6440 5172 6452
rect 3620 6412 5172 6440
rect 2130 6332 2136 6384
rect 2188 6372 2194 6384
rect 2866 6372 2872 6384
rect 2188 6344 2872 6372
rect 2188 6332 2194 6344
rect 2866 6332 2872 6344
rect 2924 6332 2930 6384
rect 3620 6381 3648 6412
rect 5166 6400 5172 6412
rect 5224 6400 5230 6452
rect 5258 6400 5264 6452
rect 5316 6440 5322 6452
rect 10321 6443 10379 6449
rect 10321 6440 10333 6443
rect 5316 6412 10333 6440
rect 5316 6400 5322 6412
rect 10321 6409 10333 6412
rect 10367 6409 10379 6443
rect 10321 6403 10379 6409
rect 3605 6375 3663 6381
rect 3605 6341 3617 6375
rect 3651 6341 3663 6375
rect 5074 6372 5080 6384
rect 4830 6344 5080 6372
rect 3605 6335 3663 6341
rect 5074 6332 5080 6344
rect 5132 6332 5138 6384
rect 5445 6375 5503 6381
rect 5445 6341 5457 6375
rect 5491 6372 5503 6375
rect 5534 6372 5540 6384
rect 5491 6344 5540 6372
rect 5491 6341 5503 6344
rect 5445 6335 5503 6341
rect 5534 6332 5540 6344
rect 5592 6332 5598 6384
rect 6454 6332 6460 6384
rect 6512 6332 6518 6384
rect 6914 6332 6920 6384
rect 6972 6372 6978 6384
rect 7377 6375 7435 6381
rect 7377 6372 7389 6375
rect 6972 6344 7389 6372
rect 6972 6332 6978 6344
rect 7377 6341 7389 6344
rect 7423 6341 7435 6375
rect 7742 6372 7748 6384
rect 7703 6344 7748 6372
rect 7377 6335 7435 6341
rect 7742 6332 7748 6344
rect 7800 6372 7806 6384
rect 10428 6372 10456 6616
rect 10505 6443 10563 6449
rect 10505 6409 10517 6443
rect 10551 6440 10563 6443
rect 13630 6440 13636 6452
rect 10551 6412 13636 6440
rect 10551 6409 10563 6412
rect 10505 6403 10563 6409
rect 13630 6400 13636 6412
rect 13688 6400 13694 6452
rect 13814 6372 13820 6384
rect 7800 6344 8340 6372
rect 10428 6344 13820 6372
rect 7800 6332 7806 6344
rect 3326 6304 3332 6316
rect 3287 6276 3332 6304
rect 3326 6264 3332 6276
rect 3384 6264 3390 6316
rect 1762 6196 1768 6248
rect 1820 6236 1826 6248
rect 3142 6236 3148 6248
rect 1820 6208 3148 6236
rect 1820 6196 1826 6208
rect 3142 6196 3148 6208
rect 3200 6236 3206 6248
rect 3694 6236 3700 6248
rect 3200 6208 3700 6236
rect 3200 6196 3206 6208
rect 3694 6196 3700 6208
rect 3752 6196 3758 6248
rect 5166 6236 5172 6248
rect 5127 6208 5172 6236
rect 5166 6196 5172 6208
rect 5224 6196 5230 6248
rect 6472 6236 6500 6332
rect 7006 6304 7012 6316
rect 6967 6276 7012 6304
rect 7006 6264 7012 6276
rect 7064 6264 7070 6316
rect 7193 6307 7251 6313
rect 7193 6273 7205 6307
rect 7239 6273 7251 6307
rect 7193 6267 7251 6273
rect 7208 6236 7236 6267
rect 7466 6264 7472 6316
rect 7524 6304 7530 6316
rect 8312 6313 8340 6344
rect 13814 6332 13820 6344
rect 13872 6332 13878 6384
rect 7653 6307 7711 6313
rect 7524 6302 7604 6304
rect 7653 6302 7665 6307
rect 7524 6276 7665 6302
rect 7524 6264 7530 6276
rect 7576 6274 7665 6276
rect 7653 6273 7665 6274
rect 7699 6273 7711 6307
rect 7653 6267 7711 6273
rect 7929 6307 7987 6313
rect 7929 6273 7941 6307
rect 7975 6273 7987 6307
rect 7929 6267 7987 6273
rect 8297 6307 8355 6313
rect 8297 6273 8309 6307
rect 8343 6273 8355 6307
rect 8849 6307 8907 6313
rect 8849 6304 8861 6307
rect 8297 6267 8355 6273
rect 8588 6276 8861 6304
rect 7944 6236 7972 6267
rect 8386 6236 8392 6248
rect 6472 6208 8392 6236
rect 8386 6196 8392 6208
rect 8444 6196 8450 6248
rect 7282 6128 7288 6180
rect 7340 6168 7346 6180
rect 7340 6140 7880 6168
rect 7340 6128 7346 6140
rect 3602 6060 3608 6112
rect 3660 6100 3666 6112
rect 5077 6103 5135 6109
rect 5077 6100 5089 6103
rect 3660 6072 5089 6100
rect 3660 6060 3666 6072
rect 5077 6069 5089 6072
rect 5123 6069 5135 6103
rect 5077 6063 5135 6069
rect 6086 6060 6092 6112
rect 6144 6100 6150 6112
rect 6917 6103 6975 6109
rect 6917 6100 6929 6103
rect 6144 6072 6929 6100
rect 6144 6060 6150 6072
rect 6917 6069 6929 6072
rect 6963 6069 6975 6103
rect 6917 6063 6975 6069
rect 7469 6103 7527 6109
rect 7469 6069 7481 6103
rect 7515 6100 7527 6103
rect 7558 6100 7564 6112
rect 7515 6072 7564 6100
rect 7515 6069 7527 6072
rect 7469 6063 7527 6069
rect 7558 6060 7564 6072
rect 7616 6060 7622 6112
rect 7852 6100 7880 6140
rect 7926 6128 7932 6180
rect 7984 6168 7990 6180
rect 8588 6168 8616 6276
rect 8849 6273 8861 6276
rect 8895 6273 8907 6307
rect 8849 6267 8907 6273
rect 7984 6140 8616 6168
rect 8757 6171 8815 6177
rect 7984 6128 7990 6140
rect 8757 6137 8769 6171
rect 8803 6168 8815 6171
rect 9490 6168 9496 6180
rect 8803 6140 9496 6168
rect 8803 6137 8815 6140
rect 8757 6131 8815 6137
rect 9490 6128 9496 6140
rect 9548 6128 9554 6180
rect 8113 6103 8171 6109
rect 8113 6100 8125 6103
rect 7852 6072 8125 6100
rect 8113 6069 8125 6072
rect 8159 6069 8171 6103
rect 8386 6100 8392 6112
rect 8347 6072 8392 6100
rect 8113 6063 8171 6069
rect 8386 6060 8392 6072
rect 8444 6060 8450 6112
rect 8478 6060 8484 6112
rect 8536 6100 8542 6112
rect 8941 6103 8999 6109
rect 8941 6100 8953 6103
rect 8536 6072 8953 6100
rect 8536 6060 8542 6072
rect 8941 6069 8953 6072
rect 8987 6100 8999 6103
rect 9122 6100 9128 6112
rect 8987 6072 9128 6100
rect 8987 6069 8999 6072
rect 8941 6063 8999 6069
rect 9122 6060 9128 6072
rect 9180 6060 9186 6112
rect 9309 6103 9367 6109
rect 9309 6069 9321 6103
rect 9355 6100 9367 6103
rect 9398 6100 9404 6112
rect 9355 6072 9404 6100
rect 9355 6069 9367 6072
rect 9309 6063 9367 6069
rect 9398 6060 9404 6072
rect 9456 6060 9462 6112
rect 3036 6010 9844 6032
rect 1486 5924 1492 5976
rect 1544 5964 1550 5976
rect 2498 5964 2504 5976
rect 1544 5936 2504 5964
rect 1544 5924 1550 5936
rect 2498 5924 2504 5936
rect 2556 5924 2562 5976
rect 3036 5958 5666 6010
rect 5718 5958 5730 6010
rect 5782 5958 5794 6010
rect 5846 5958 5858 6010
rect 5910 5958 5922 6010
rect 5974 5958 8766 6010
rect 8818 5958 8830 6010
rect 8882 5958 8894 6010
rect 8946 5958 8958 6010
rect 9010 5958 9022 6010
rect 9074 5958 9844 6010
rect 3036 5936 9844 5958
rect 1854 5856 1860 5908
rect 1912 5896 1918 5908
rect 2685 5899 2743 5905
rect 2685 5896 2697 5899
rect 1912 5868 2697 5896
rect 1912 5856 1918 5868
rect 2685 5865 2697 5868
rect 2731 5865 2743 5899
rect 2685 5859 2743 5865
rect 2961 5899 3019 5905
rect 2961 5865 2973 5899
rect 3007 5896 3019 5899
rect 6638 5896 6644 5908
rect 3007 5868 6644 5896
rect 3007 5865 3019 5868
rect 2961 5859 3019 5865
rect 6638 5856 6644 5868
rect 6696 5856 6702 5908
rect 7466 5856 7472 5908
rect 7524 5856 7530 5908
rect 7926 5856 7932 5908
rect 7984 5896 7990 5908
rect 8021 5899 8079 5905
rect 8021 5896 8033 5899
rect 7984 5868 8033 5896
rect 7984 5856 7990 5868
rect 8021 5865 8033 5868
rect 8067 5865 8079 5899
rect 8021 5859 8079 5865
rect 8113 5899 8171 5905
rect 8113 5865 8125 5899
rect 8159 5896 8171 5899
rect 13722 5896 13728 5908
rect 8159 5868 13728 5896
rect 8159 5865 8171 5868
rect 8113 5859 8171 5865
rect 13722 5856 13728 5868
rect 13780 5856 13786 5908
rect 1670 5788 1676 5840
rect 1728 5828 1734 5840
rect 2590 5828 2596 5840
rect 1728 5800 2596 5828
rect 1728 5788 1734 5800
rect 2590 5788 2596 5800
rect 2648 5788 2654 5840
rect 5074 5788 5080 5840
rect 5132 5788 5138 5840
rect 7484 5828 7512 5856
rect 8849 5831 8907 5837
rect 8849 5828 8861 5831
rect 7484 5800 8861 5828
rect 8849 5797 8861 5800
rect 8895 5797 8907 5831
rect 8849 5791 8907 5797
rect 9401 5831 9459 5837
rect 9401 5797 9413 5831
rect 9447 5828 9459 5831
rect 12802 5828 12808 5840
rect 9447 5800 12808 5828
rect 9447 5797 9459 5800
rect 9401 5791 9459 5797
rect 12802 5788 12808 5800
rect 12860 5788 12866 5840
rect 5092 5760 5120 5788
rect 6086 5760 6092 5772
rect 4724 5732 5120 5760
rect 6047 5732 6092 5760
rect 1581 5695 1639 5701
rect 1581 5661 1593 5695
rect 1627 5692 1639 5695
rect 2869 5695 2927 5701
rect 2869 5692 2881 5695
rect 1627 5664 2881 5692
rect 1627 5661 1639 5664
rect 1581 5655 1639 5661
rect 2869 5661 2881 5664
rect 2915 5661 2927 5695
rect 3326 5692 3332 5704
rect 3287 5664 3332 5692
rect 2869 5655 2927 5661
rect 3326 5652 3332 5664
rect 3384 5652 3390 5704
rect 4724 5678 4752 5732
rect 6086 5720 6092 5732
rect 6144 5720 6150 5772
rect 8389 5763 8447 5769
rect 8389 5729 8401 5763
rect 8435 5760 8447 5763
rect 8481 5763 8539 5769
rect 8481 5760 8493 5763
rect 8435 5732 8493 5760
rect 8435 5729 8447 5732
rect 8389 5723 8447 5729
rect 8481 5729 8493 5732
rect 8527 5760 8539 5763
rect 9674 5760 9680 5772
rect 8527 5732 9680 5760
rect 8527 5729 8539 5732
rect 8481 5723 8539 5729
rect 9674 5720 9680 5732
rect 9732 5720 9738 5772
rect 5074 5652 5080 5704
rect 5132 5692 5138 5704
rect 5442 5692 5448 5704
rect 5132 5664 5448 5692
rect 5132 5652 5138 5664
rect 5442 5652 5448 5664
rect 5500 5692 5506 5704
rect 5537 5695 5595 5701
rect 5537 5692 5549 5695
rect 5500 5664 5549 5692
rect 5500 5652 5506 5664
rect 5537 5661 5549 5664
rect 5583 5661 5595 5695
rect 5537 5655 5595 5661
rect 5626 5652 5632 5704
rect 5684 5692 5690 5704
rect 5721 5695 5779 5701
rect 5721 5692 5733 5695
rect 5684 5664 5733 5692
rect 5684 5652 5690 5664
rect 5721 5661 5733 5664
rect 5767 5661 5779 5695
rect 5721 5655 5779 5661
rect 7561 5695 7619 5701
rect 7561 5661 7573 5695
rect 7607 5692 7619 5695
rect 7926 5692 7932 5704
rect 7607 5664 7932 5692
rect 7607 5661 7619 5664
rect 7561 5655 7619 5661
rect 7926 5652 7932 5664
rect 7984 5652 7990 5704
rect 8662 5692 8668 5704
rect 8623 5664 8668 5692
rect 8662 5652 8668 5664
rect 8720 5652 8726 5704
rect 9122 5692 9128 5704
rect 9083 5664 9128 5692
rect 9122 5652 9128 5664
rect 9180 5652 9186 5704
rect 9217 5695 9275 5701
rect 9217 5661 9229 5695
rect 9263 5661 9275 5695
rect 9217 5655 9275 5661
rect 1394 5584 1400 5636
rect 1452 5624 1458 5636
rect 2682 5624 2688 5636
rect 1452 5596 2688 5624
rect 1452 5584 1458 5596
rect 2682 5584 2688 5596
rect 2740 5584 2746 5636
rect 3602 5624 3608 5636
rect 3563 5596 3608 5624
rect 3602 5584 3608 5596
rect 3660 5584 3666 5636
rect 4982 5584 4988 5636
rect 5040 5624 5046 5636
rect 7650 5624 7656 5636
rect 5040 5596 5488 5624
rect 7222 5596 7656 5624
rect 5040 5584 5046 5596
rect 2225 5559 2283 5565
rect 2225 5525 2237 5559
rect 2271 5556 2283 5559
rect 2961 5559 3019 5565
rect 2961 5556 2973 5559
rect 2271 5528 2973 5556
rect 2271 5525 2283 5528
rect 2225 5519 2283 5525
rect 2961 5525 2973 5528
rect 3007 5525 3019 5559
rect 2961 5519 3019 5525
rect 3786 5516 3792 5568
rect 3844 5556 3850 5568
rect 5077 5559 5135 5565
rect 5077 5556 5089 5559
rect 3844 5528 5089 5556
rect 3844 5516 3850 5528
rect 5077 5525 5089 5528
rect 5123 5525 5135 5559
rect 5350 5556 5356 5568
rect 5311 5528 5356 5556
rect 5077 5519 5135 5525
rect 5350 5516 5356 5528
rect 5408 5516 5414 5568
rect 5460 5556 5488 5596
rect 7650 5584 7656 5596
rect 7708 5584 7714 5636
rect 8386 5584 8392 5636
rect 8444 5624 8450 5636
rect 9232 5624 9260 5655
rect 8444 5596 9260 5624
rect 8444 5584 8450 5596
rect 8113 5559 8171 5565
rect 8113 5556 8125 5559
rect 5460 5528 8125 5556
rect 8113 5525 8125 5528
rect 8159 5525 8171 5559
rect 8113 5519 8171 5525
rect 8941 5559 8999 5565
rect 8941 5525 8953 5559
rect 8987 5556 8999 5559
rect 9214 5556 9220 5568
rect 8987 5528 9220 5556
rect 8987 5525 8999 5528
rect 8941 5519 8999 5525
rect 9214 5516 9220 5528
rect 9272 5516 9278 5568
rect 3036 5466 9844 5488
rect 3036 5414 4116 5466
rect 4168 5414 4180 5466
rect 4232 5414 4244 5466
rect 4296 5414 4308 5466
rect 4360 5414 4372 5466
rect 4424 5414 7216 5466
rect 7268 5414 7280 5466
rect 7332 5414 7344 5466
rect 7396 5414 7408 5466
rect 7460 5414 7472 5466
rect 7524 5414 9844 5466
rect 3036 5392 9844 5414
rect 2869 5355 2927 5361
rect 2869 5321 2881 5355
rect 2915 5352 2927 5355
rect 5074 5352 5080 5364
rect 2915 5324 5080 5352
rect 2915 5321 2927 5324
rect 2869 5315 2927 5321
rect 5074 5312 5080 5324
rect 5132 5312 5138 5364
rect 7653 5355 7711 5361
rect 6656 5324 7420 5352
rect 4706 5244 4712 5296
rect 4764 5244 4770 5296
rect 6086 5244 6092 5296
rect 6144 5284 6150 5296
rect 6181 5287 6239 5293
rect 6181 5284 6193 5287
rect 6144 5256 6193 5284
rect 6144 5244 6150 5256
rect 6181 5253 6193 5256
rect 6227 5253 6239 5287
rect 6181 5247 6239 5253
rect 6454 5244 6460 5296
rect 6512 5284 6518 5296
rect 6656 5284 6684 5324
rect 6512 5270 6684 5284
rect 7392 5284 7420 5324
rect 7653 5321 7665 5355
rect 7699 5352 7711 5355
rect 7742 5352 7748 5364
rect 7699 5324 7748 5352
rect 7699 5321 7711 5324
rect 7653 5315 7711 5321
rect 7742 5312 7748 5324
rect 7800 5352 7806 5364
rect 8662 5352 8668 5364
rect 7800 5324 8668 5352
rect 7800 5312 7806 5324
rect 8662 5312 8668 5324
rect 8720 5312 8726 5364
rect 8754 5312 8760 5364
rect 8812 5312 8818 5364
rect 9122 5352 9128 5364
rect 9083 5324 9128 5352
rect 9122 5312 9128 5324
rect 9180 5312 9186 5364
rect 9217 5355 9275 5361
rect 9217 5321 9229 5355
rect 9263 5352 9275 5355
rect 9582 5352 9588 5364
rect 9263 5324 9588 5352
rect 9263 5321 9275 5324
rect 9217 5315 9275 5321
rect 9582 5312 9588 5324
rect 9640 5312 9646 5364
rect 7929 5287 7987 5293
rect 7929 5284 7941 5287
rect 7392 5270 7941 5284
rect 6512 5256 6670 5270
rect 7406 5256 7941 5270
rect 6512 5244 6518 5256
rect 7929 5253 7941 5256
rect 7975 5253 7987 5287
rect 7929 5247 7987 5253
rect 3234 5176 3240 5228
rect 3292 5216 3298 5228
rect 3421 5219 3479 5225
rect 3421 5216 3433 5219
rect 3292 5188 3433 5216
rect 3292 5176 3298 5188
rect 3421 5185 3433 5188
rect 3467 5185 3479 5219
rect 3421 5179 3479 5185
rect 3602 5176 3608 5228
rect 3660 5216 3666 5228
rect 3789 5219 3847 5225
rect 3789 5216 3801 5219
rect 3660 5188 3801 5216
rect 3660 5176 3666 5188
rect 3789 5185 3801 5188
rect 3835 5185 3847 5219
rect 3789 5179 3847 5185
rect 4798 5176 4804 5228
rect 4856 5216 4862 5228
rect 5261 5219 5319 5225
rect 5261 5216 5273 5219
rect 4856 5188 5273 5216
rect 4856 5176 4862 5188
rect 5261 5185 5273 5188
rect 5307 5185 5319 5219
rect 5261 5179 5319 5185
rect 7745 5219 7803 5225
rect 7745 5185 7757 5219
rect 7791 5185 7803 5219
rect 7745 5179 7803 5185
rect 2774 5108 2780 5160
rect 2832 5108 2838 5160
rect 5442 5108 5448 5160
rect 5500 5148 5506 5160
rect 5905 5151 5963 5157
rect 5905 5148 5917 5151
rect 5500 5120 5917 5148
rect 5500 5108 5506 5120
rect 5905 5117 5917 5120
rect 5951 5117 5963 5151
rect 5905 5111 5963 5117
rect 6638 5108 6644 5160
rect 6696 5148 6702 5160
rect 7760 5148 7788 5179
rect 6696 5120 7788 5148
rect 6696 5108 6702 5120
rect 2792 5080 2820 5108
rect 3234 5080 3240 5092
rect 2792 5052 3240 5080
rect 3234 5040 3240 5052
rect 3292 5040 3298 5092
rect 7944 5080 7972 5247
rect 8662 5216 8668 5228
rect 8623 5188 8668 5216
rect 8662 5176 8668 5188
rect 8720 5176 8726 5228
rect 8772 5225 8800 5312
rect 8772 5219 8833 5225
rect 8772 5188 8787 5219
rect 8775 5185 8787 5188
rect 8821 5185 8833 5219
rect 8941 5219 8999 5225
rect 8941 5216 8953 5219
rect 8775 5179 8833 5185
rect 8864 5188 8953 5216
rect 8864 5080 8892 5188
rect 8941 5185 8953 5188
rect 8987 5185 8999 5219
rect 8941 5179 8999 5185
rect 9401 5219 9459 5225
rect 9401 5185 9413 5219
rect 9447 5216 9459 5219
rect 9490 5216 9496 5228
rect 9447 5188 9496 5216
rect 9447 5185 9459 5188
rect 9401 5179 9459 5185
rect 9490 5176 9496 5188
rect 9548 5176 9554 5228
rect 9490 5080 9496 5092
rect 7944 5052 9496 5080
rect 9490 5040 9496 5052
rect 9548 5040 9554 5092
rect 2774 4972 2780 5024
rect 2832 5012 2838 5024
rect 5258 5012 5264 5024
rect 2832 4984 5264 5012
rect 2832 4972 2838 4984
rect 5258 4972 5264 4984
rect 5316 4972 5322 5024
rect 5721 5015 5779 5021
rect 5721 4981 5733 5015
rect 5767 5012 5779 5015
rect 7834 5012 7840 5024
rect 5767 4984 7840 5012
rect 5767 4981 5779 4984
rect 5721 4975 5779 4981
rect 7834 4972 7840 4984
rect 7892 4972 7898 5024
rect 8110 5012 8116 5024
rect 8071 4984 8116 5012
rect 8110 4972 8116 4984
rect 8168 4972 8174 5024
rect 8478 5012 8484 5024
rect 8439 4984 8484 5012
rect 8478 4972 8484 4984
rect 8536 4972 8542 5024
rect 3036 4922 9844 4944
rect 2685 4879 2743 4885
rect 2685 4845 2697 4879
rect 2731 4876 2743 4879
rect 2774 4876 2780 4888
rect 2731 4848 2780 4876
rect 2731 4845 2743 4848
rect 2685 4839 2743 4845
rect 2774 4836 2780 4848
rect 2832 4836 2838 4888
rect 3036 4870 5666 4922
rect 5718 4870 5730 4922
rect 5782 4870 5794 4922
rect 5846 4870 5858 4922
rect 5910 4870 5922 4922
rect 5974 4870 8766 4922
rect 8818 4870 8830 4922
rect 8882 4870 8894 4922
rect 8946 4870 8958 4922
rect 9010 4870 9022 4922
rect 9074 4870 9844 4922
rect 3036 4848 9844 4870
rect 3050 4768 3056 4820
rect 3108 4808 3114 4820
rect 3329 4811 3387 4817
rect 3329 4808 3341 4811
rect 3108 4780 3341 4808
rect 3108 4768 3114 4780
rect 3329 4777 3341 4780
rect 3375 4777 3387 4811
rect 4338 4808 4344 4820
rect 3329 4771 3387 4777
rect 3528 4780 4344 4808
rect 3528 4613 3556 4780
rect 4338 4768 4344 4780
rect 4396 4768 4402 4820
rect 4430 4768 4436 4820
rect 4488 4808 4494 4820
rect 4488 4780 4533 4808
rect 4488 4768 4494 4780
rect 4614 4768 4620 4820
rect 4672 4808 4678 4820
rect 6089 4811 6147 4817
rect 4672 4780 4717 4808
rect 4672 4768 4678 4780
rect 6089 4777 6101 4811
rect 6135 4808 6147 4811
rect 6362 4808 6368 4820
rect 6135 4780 6368 4808
rect 6135 4777 6147 4780
rect 6089 4771 6147 4777
rect 6362 4768 6368 4780
rect 6420 4768 6426 4820
rect 6454 4768 6460 4820
rect 6512 4808 6518 4820
rect 6733 4811 6791 4817
rect 6733 4808 6745 4811
rect 6512 4780 6745 4808
rect 6512 4768 6518 4780
rect 6733 4777 6745 4780
rect 6779 4777 6791 4811
rect 6733 4771 6791 4777
rect 7101 4811 7159 4817
rect 7101 4777 7113 4811
rect 7147 4808 7159 4811
rect 8202 4808 8208 4820
rect 7147 4780 8208 4808
rect 7147 4777 7159 4780
rect 7101 4771 7159 4777
rect 8202 4768 8208 4780
rect 8260 4768 8266 4820
rect 9122 4768 9128 4820
rect 9180 4808 9186 4820
rect 9493 4811 9551 4817
rect 9493 4808 9505 4811
rect 9180 4780 9505 4808
rect 9180 4768 9186 4780
rect 9493 4777 9505 4780
rect 9539 4777 9551 4811
rect 9493 4771 9551 4777
rect 3605 4743 3663 4749
rect 3605 4709 3617 4743
rect 3651 4740 3663 4743
rect 5534 4740 5540 4752
rect 3651 4712 5540 4740
rect 3651 4709 3663 4712
rect 3605 4703 3663 4709
rect 5534 4700 5540 4712
rect 5592 4700 5598 4752
rect 5350 4672 5356 4684
rect 4080 4644 5356 4672
rect 4080 4613 4108 4644
rect 5350 4632 5356 4644
rect 5408 4632 5414 4684
rect 7193 4675 7251 4681
rect 7193 4641 7205 4675
rect 7239 4672 7251 4675
rect 7466 4672 7472 4684
rect 7239 4644 7472 4672
rect 7239 4641 7251 4644
rect 7193 4635 7251 4641
rect 7466 4632 7472 4644
rect 7524 4632 7530 4684
rect 7561 4675 7619 4681
rect 7561 4641 7573 4675
rect 7607 4672 7619 4675
rect 7742 4672 7748 4684
rect 7607 4644 7748 4672
rect 7607 4641 7619 4644
rect 7561 4635 7619 4641
rect 7742 4632 7748 4644
rect 7800 4632 7806 4684
rect 3513 4607 3571 4613
rect 3513 4573 3525 4607
rect 3559 4573 3571 4607
rect 3513 4567 3571 4573
rect 3789 4607 3847 4613
rect 3789 4573 3801 4607
rect 3835 4573 3847 4607
rect 3789 4567 3847 4573
rect 4065 4607 4123 4613
rect 4065 4573 4077 4607
rect 4111 4573 4123 4607
rect 4065 4567 4123 4573
rect 3804 4536 3832 4567
rect 4154 4564 4160 4616
rect 4212 4604 4218 4616
rect 4212 4576 4257 4604
rect 4212 4564 4218 4576
rect 4338 4564 4344 4616
rect 4396 4604 4402 4616
rect 4709 4607 4767 4613
rect 4709 4604 4721 4607
rect 4396 4576 4721 4604
rect 4396 4564 4402 4576
rect 4709 4573 4721 4576
rect 4755 4573 4767 4607
rect 4982 4604 4988 4616
rect 4943 4576 4988 4604
rect 4709 4567 4767 4573
rect 4982 4564 4988 4576
rect 5040 4564 5046 4616
rect 5166 4564 5172 4616
rect 5224 4604 5230 4616
rect 5442 4604 5448 4616
rect 5224 4576 5448 4604
rect 5224 4564 5230 4576
rect 5442 4564 5448 4576
rect 5500 4604 5506 4616
rect 6457 4607 6515 4613
rect 6457 4604 6469 4607
rect 5500 4576 6469 4604
rect 5500 4564 5506 4576
rect 6457 4573 6469 4576
rect 6503 4573 6515 4607
rect 6638 4604 6644 4616
rect 6599 4576 6644 4604
rect 6457 4567 6515 4573
rect 6638 4564 6644 4576
rect 6696 4564 6702 4616
rect 9033 4607 9091 4613
rect 9033 4573 9045 4607
rect 9079 4604 9091 4607
rect 9214 4604 9220 4616
rect 9079 4576 9220 4604
rect 9079 4573 9091 4576
rect 9033 4567 9091 4573
rect 9214 4564 9220 4576
rect 9272 4564 9278 4616
rect 5718 4536 5724 4548
rect 3804 4508 4844 4536
rect 5679 4508 5724 4536
rect 3881 4471 3939 4477
rect 3881 4437 3893 4471
rect 3927 4468 3939 4471
rect 4706 4468 4712 4480
rect 3927 4440 4712 4468
rect 3927 4437 3939 4440
rect 3881 4431 3939 4437
rect 4706 4428 4712 4440
rect 4764 4428 4770 4480
rect 4816 4468 4844 4508
rect 5718 4496 5724 4508
rect 5776 4496 5782 4548
rect 5902 4496 5908 4548
rect 5960 4536 5966 4548
rect 6273 4539 6331 4545
rect 5960 4508 6132 4536
rect 5960 4496 5966 4508
rect 5994 4468 6000 4480
rect 4816 4440 6000 4468
rect 5994 4428 6000 4440
rect 6052 4428 6058 4480
rect 6104 4468 6132 4508
rect 6273 4505 6285 4539
rect 6319 4536 6331 4539
rect 7098 4536 7104 4548
rect 6319 4508 7104 4536
rect 6319 4505 6331 4508
rect 6273 4499 6331 4505
rect 7098 4496 7104 4508
rect 7156 4496 7162 4548
rect 8478 4496 8484 4548
rect 8536 4496 8542 4548
rect 6454 4468 6460 4480
rect 6104 4440 6460 4468
rect 6454 4428 6460 4440
rect 6512 4428 6518 4480
rect 8110 4428 8116 4480
rect 8168 4468 8174 4480
rect 9214 4468 9220 4480
rect 8168 4440 9220 4468
rect 8168 4428 8174 4440
rect 9214 4428 9220 4440
rect 9272 4428 9278 4480
rect 3036 4378 9844 4400
rect 3036 4326 4116 4378
rect 4168 4326 4180 4378
rect 4232 4326 4244 4378
rect 4296 4326 4308 4378
rect 4360 4326 4372 4378
rect 4424 4326 7216 4378
rect 7268 4326 7280 4378
rect 7332 4326 7344 4378
rect 7396 4326 7408 4378
rect 7460 4326 7472 4378
rect 7524 4326 9844 4378
rect 3036 4304 9844 4326
rect 8018 4224 8024 4276
rect 8076 4264 8082 4276
rect 8297 4267 8355 4273
rect 8297 4264 8309 4267
rect 8076 4236 8309 4264
rect 8076 4224 8082 4236
rect 8297 4233 8309 4236
rect 8343 4233 8355 4267
rect 8297 4227 8355 4233
rect 8662 4224 8668 4276
rect 8720 4264 8726 4276
rect 9033 4267 9091 4273
rect 9033 4264 9045 4267
rect 8720 4236 9045 4264
rect 8720 4224 8726 4236
rect 9033 4233 9045 4236
rect 9079 4233 9091 4267
rect 9033 4227 9091 4233
rect 4154 4156 4160 4208
rect 4212 4156 4218 4208
rect 8202 4196 8208 4208
rect 7314 4168 8208 4196
rect 8202 4156 8208 4168
rect 8260 4156 8266 4208
rect 2958 4088 2964 4140
rect 3016 4128 3022 4140
rect 3421 4131 3479 4137
rect 3421 4128 3433 4131
rect 3016 4100 3433 4128
rect 3016 4088 3022 4100
rect 3421 4097 3433 4100
rect 3467 4097 3479 4131
rect 3786 4128 3792 4140
rect 3747 4100 3792 4128
rect 3421 4091 3479 4097
rect 3786 4088 3792 4100
rect 3844 4088 3850 4140
rect 5258 4128 5264 4140
rect 5219 4100 5264 4128
rect 5258 4088 5264 4100
rect 5316 4088 5322 4140
rect 6178 4128 6184 4140
rect 6139 4100 6184 4128
rect 6178 4088 6184 4100
rect 6236 4088 6242 4140
rect 7650 4128 7656 4140
rect 7611 4100 7656 4128
rect 7650 4088 7656 4100
rect 7708 4088 7714 4140
rect 8481 4131 8539 4137
rect 8481 4128 8493 4131
rect 7760 4100 8493 4128
rect 5813 4063 5871 4069
rect 5813 4029 5825 4063
rect 5859 4029 5871 4063
rect 5813 4023 5871 4029
rect 5828 3992 5856 4023
rect 4724 3964 5856 3992
rect 4724 3924 4752 3964
rect 7098 3952 7104 4004
rect 7156 3992 7162 4004
rect 7760 3992 7788 4100
rect 8481 4097 8493 4100
rect 8527 4097 8539 4131
rect 8481 4091 8539 4097
rect 8573 4131 8631 4137
rect 8573 4097 8585 4131
rect 8619 4128 8631 4131
rect 8754 4128 8760 4140
rect 8619 4100 8760 4128
rect 8619 4097 8631 4100
rect 8573 4091 8631 4097
rect 8754 4088 8760 4100
rect 8812 4088 8818 4140
rect 9214 4088 9220 4140
rect 9272 4128 9278 4140
rect 9309 4131 9367 4137
rect 9309 4128 9321 4131
rect 9272 4100 9321 4128
rect 9272 4088 9278 4100
rect 9309 4097 9321 4100
rect 9355 4097 9367 4131
rect 9309 4091 9367 4097
rect 7926 4020 7932 4072
rect 7984 4060 7990 4072
rect 7984 4032 9168 4060
rect 7984 4020 7990 4032
rect 9140 4001 9168 4032
rect 7156 3964 7788 3992
rect 9125 3995 9183 4001
rect 7156 3952 7162 3964
rect 9125 3961 9137 3995
rect 9171 3961 9183 3995
rect 9125 3955 9183 3961
rect 2608 3896 4752 3924
rect 5721 3927 5779 3933
rect 2608 3652 2636 3896
rect 5721 3893 5733 3927
rect 5767 3924 5779 3927
rect 6730 3924 6736 3936
rect 5767 3896 6736 3924
rect 5767 3893 5779 3896
rect 5721 3887 5779 3893
rect 6730 3884 6736 3896
rect 6788 3884 6794 3936
rect 8113 3927 8171 3933
rect 8113 3893 8125 3927
rect 8159 3924 8171 3927
rect 8570 3924 8576 3936
rect 8159 3896 8576 3924
rect 8159 3893 8171 3896
rect 8113 3887 8171 3893
rect 8570 3884 8576 3896
rect 8628 3884 8634 3936
rect 8662 3884 8668 3936
rect 8720 3924 8726 3936
rect 8849 3927 8907 3933
rect 8849 3924 8861 3927
rect 8720 3896 8861 3924
rect 8720 3884 8726 3896
rect 8849 3893 8861 3896
rect 8895 3924 8907 3927
rect 9490 3924 9496 3936
rect 8895 3896 9496 3924
rect 8895 3893 8907 3896
rect 8849 3887 8907 3893
rect 9490 3884 9496 3896
rect 9548 3884 9554 3936
rect 3036 3834 9844 3856
rect 3036 3782 5666 3834
rect 5718 3782 5730 3834
rect 5782 3782 5794 3834
rect 5846 3782 5858 3834
rect 5910 3782 5922 3834
rect 5974 3782 8766 3834
rect 8818 3782 8830 3834
rect 8882 3782 8894 3834
rect 8946 3782 8958 3834
rect 9010 3782 9022 3834
rect 9074 3782 9844 3834
rect 3036 3760 9844 3782
rect 2682 3680 2688 3732
rect 2740 3720 2746 3732
rect 5994 3720 6000 3732
rect 2740 3692 5764 3720
rect 5955 3692 6000 3720
rect 2740 3680 2746 3692
rect 5442 3652 5448 3664
rect 2608 3624 2728 3652
rect 2700 3596 2728 3624
rect 4724 3624 5448 3652
rect 2682 3544 2688 3596
rect 2740 3544 2746 3596
rect 3326 3584 3332 3596
rect 3287 3556 3332 3584
rect 3326 3544 3332 3556
rect 3384 3544 3390 3596
rect 3605 3587 3663 3593
rect 3605 3553 3617 3587
rect 3651 3584 3663 3587
rect 3694 3584 3700 3596
rect 3651 3556 3700 3584
rect 3651 3553 3663 3556
rect 3605 3547 3663 3553
rect 3694 3544 3700 3556
rect 3752 3544 3758 3596
rect 3970 3544 3976 3596
rect 4028 3584 4034 3596
rect 4724 3584 4752 3624
rect 5442 3612 5448 3624
rect 5500 3612 5506 3664
rect 5736 3652 5764 3692
rect 5994 3680 6000 3692
rect 6052 3680 6058 3732
rect 8018 3720 8024 3732
rect 6380 3692 8024 3720
rect 6380 3652 6408 3692
rect 8018 3680 8024 3692
rect 8076 3680 8082 3732
rect 8294 3680 8300 3732
rect 8352 3720 8358 3732
rect 8573 3723 8631 3729
rect 8573 3720 8585 3723
rect 8352 3692 8585 3720
rect 8352 3680 8358 3692
rect 8573 3689 8585 3692
rect 8619 3689 8631 3723
rect 8573 3683 8631 3689
rect 9217 3723 9275 3729
rect 9217 3689 9229 3723
rect 9263 3720 9275 3723
rect 9306 3720 9312 3732
rect 9263 3692 9312 3720
rect 9263 3689 9275 3692
rect 9217 3683 9275 3689
rect 9306 3680 9312 3692
rect 9364 3680 9370 3732
rect 5736 3624 6408 3652
rect 7650 3612 7656 3664
rect 7708 3652 7714 3664
rect 8941 3655 8999 3661
rect 8941 3652 8953 3655
rect 7708 3624 8953 3652
rect 7708 3612 7714 3624
rect 8941 3621 8953 3624
rect 8987 3621 8999 3655
rect 8941 3615 8999 3621
rect 4028 3556 4752 3584
rect 4028 3544 4034 3556
rect 4724 3502 4752 3556
rect 4982 3544 4988 3596
rect 5040 3584 5046 3596
rect 6273 3587 6331 3593
rect 6273 3584 6285 3587
rect 5040 3556 6285 3584
rect 5040 3544 5046 3556
rect 6273 3553 6285 3556
rect 6319 3584 6331 3587
rect 7098 3584 7104 3596
rect 6319 3556 7104 3584
rect 6319 3553 6331 3556
rect 6273 3547 6331 3553
rect 7098 3544 7104 3556
rect 7156 3544 7162 3596
rect 5721 3519 5779 3525
rect 5721 3516 5733 3519
rect 5184 3488 5733 3516
rect 5184 3457 5212 3488
rect 5721 3485 5733 3488
rect 5767 3485 5779 3519
rect 5721 3479 5779 3485
rect 6454 3476 6460 3528
rect 6512 3516 6518 3528
rect 6641 3519 6699 3525
rect 6641 3516 6653 3519
rect 6512 3488 6653 3516
rect 6512 3476 6518 3488
rect 6641 3485 6653 3488
rect 6687 3485 6699 3519
rect 8110 3516 8116 3528
rect 8071 3488 8116 3516
rect 6641 3479 6699 3485
rect 8110 3476 8116 3488
rect 8168 3476 8174 3528
rect 8754 3476 8760 3528
rect 8812 3516 8818 3528
rect 8849 3519 8907 3525
rect 8849 3516 8861 3519
rect 8812 3488 8861 3516
rect 8812 3476 8818 3488
rect 8849 3485 8861 3488
rect 8895 3485 8907 3519
rect 9122 3516 9128 3528
rect 9083 3488 9128 3516
rect 8849 3479 8907 3485
rect 9122 3476 9128 3488
rect 9180 3476 9186 3528
rect 9398 3516 9404 3528
rect 9359 3488 9404 3516
rect 9398 3476 9404 3488
rect 9456 3476 9462 3528
rect 5169 3451 5227 3457
rect 5169 3448 5181 3451
rect 4908 3420 5181 3448
rect 4908 3380 4936 3420
rect 5169 3417 5181 3420
rect 5215 3417 5227 3451
rect 5169 3411 5227 3417
rect 5353 3451 5411 3457
rect 5353 3417 5365 3451
rect 5399 3448 5411 3451
rect 5442 3448 5448 3460
rect 5399 3420 5448 3448
rect 5399 3417 5411 3420
rect 5353 3411 5411 3417
rect 5442 3408 5448 3420
rect 5500 3448 5506 3460
rect 5994 3448 6000 3460
rect 5500 3420 6000 3448
rect 5500 3408 5506 3420
rect 5994 3408 6000 3420
rect 6052 3408 6058 3460
rect 7926 3448 7932 3460
rect 7774 3420 7932 3448
rect 7926 3408 7932 3420
rect 7984 3408 7990 3460
rect 5074 3380 5080 3392
rect 2608 3352 4936 3380
rect 5035 3352 5080 3380
rect 2608 2972 2636 3352
rect 5074 3340 5080 3352
rect 5132 3340 5138 3392
rect 5534 3380 5540 3392
rect 5495 3352 5540 3380
rect 5534 3340 5540 3352
rect 5592 3340 5598 3392
rect 6181 3383 6239 3389
rect 6181 3349 6193 3383
rect 6227 3380 6239 3383
rect 6546 3380 6552 3392
rect 6227 3352 6552 3380
rect 6227 3349 6239 3352
rect 6181 3343 6239 3349
rect 6546 3340 6552 3352
rect 6604 3340 6610 3392
rect 8202 3340 8208 3392
rect 8260 3380 8266 3392
rect 8665 3383 8723 3389
rect 8665 3380 8677 3383
rect 8260 3352 8677 3380
rect 8260 3340 8266 3352
rect 8665 3349 8677 3352
rect 8711 3349 8723 3383
rect 8665 3343 8723 3349
rect 3036 3290 9844 3312
rect 3036 3238 4116 3290
rect 4168 3238 4180 3290
rect 4232 3238 4244 3290
rect 4296 3238 4308 3290
rect 4360 3238 4372 3290
rect 4424 3238 7216 3290
rect 7268 3238 7280 3290
rect 7332 3238 7344 3290
rect 7396 3238 7408 3290
rect 7460 3238 7472 3290
rect 7524 3238 9844 3290
rect 3036 3216 9844 3238
rect 3329 3179 3387 3185
rect 3329 3145 3341 3179
rect 3375 3176 3387 3179
rect 4617 3179 4675 3185
rect 4617 3176 4629 3179
rect 3375 3148 4629 3176
rect 3375 3145 3387 3148
rect 3329 3139 3387 3145
rect 4617 3145 4629 3148
rect 4663 3145 4675 3179
rect 4617 3139 4675 3145
rect 5534 3136 5540 3188
rect 5592 3176 5598 3188
rect 7193 3179 7251 3185
rect 5592 3148 7144 3176
rect 5592 3136 5598 3148
rect 2682 3068 2688 3120
rect 2740 3108 2746 3120
rect 3697 3111 3755 3117
rect 3697 3108 3709 3111
rect 2740 3080 3709 3108
rect 2740 3068 2746 3080
rect 3697 3077 3709 3080
rect 3743 3108 3755 3111
rect 3743 3080 4200 3108
rect 3743 3077 3755 3080
rect 3697 3071 3755 3077
rect 3329 3043 3387 3049
rect 3329 3009 3341 3043
rect 3375 3040 3387 3043
rect 3605 3043 3663 3049
rect 3605 3040 3617 3043
rect 3375 3012 3617 3040
rect 3375 3009 3387 3012
rect 3329 3003 3387 3009
rect 3605 3009 3617 3012
rect 3651 3009 3663 3043
rect 3878 3040 3884 3052
rect 3839 3012 3884 3040
rect 3605 3003 3663 3009
rect 3878 3000 3884 3012
rect 3936 3000 3942 3052
rect 4172 3049 4200 3080
rect 6178 3068 6184 3120
rect 6236 3068 6242 3120
rect 7116 3108 7144 3148
rect 7193 3145 7205 3179
rect 7239 3176 7251 3179
rect 8110 3176 8116 3188
rect 7239 3148 8116 3176
rect 7239 3145 7251 3148
rect 7193 3139 7251 3145
rect 8110 3136 8116 3148
rect 8168 3136 8174 3188
rect 8754 3176 8760 3188
rect 8715 3148 8760 3176
rect 8754 3136 8760 3148
rect 8812 3136 8818 3188
rect 9125 3179 9183 3185
rect 9125 3145 9137 3179
rect 9171 3176 9183 3179
rect 9217 3179 9275 3185
rect 9217 3176 9229 3179
rect 9171 3148 9229 3176
rect 9171 3145 9183 3148
rect 9125 3139 9183 3145
rect 9217 3145 9229 3148
rect 9263 3176 9275 3179
rect 9674 3176 9680 3188
rect 9263 3148 9680 3176
rect 9263 3145 9275 3148
rect 9217 3139 9275 3145
rect 9674 3136 9680 3148
rect 9732 3136 9738 3188
rect 9490 3108 9496 3120
rect 7116 3080 9496 3108
rect 9490 3068 9496 3080
rect 9548 3068 9554 3120
rect 4157 3043 4215 3049
rect 4157 3009 4169 3043
rect 4203 3009 4215 3043
rect 4157 3003 4215 3009
rect 4338 3000 4344 3052
rect 4396 3040 4402 3052
rect 5074 3040 5080 3052
rect 4396 3012 5080 3040
rect 4396 3000 4402 3012
rect 5074 3000 5080 3012
rect 5132 3000 5138 3052
rect 6549 3043 6607 3049
rect 6549 3009 6561 3043
rect 6595 3009 6607 3043
rect 7374 3040 7380 3052
rect 7335 3012 7380 3040
rect 6549 3003 6607 3009
rect 2682 2972 2688 2984
rect 2608 2944 2688 2972
rect 2682 2932 2688 2944
rect 2740 2932 2746 2984
rect 3896 2972 3924 3000
rect 4706 2972 4712 2984
rect 3896 2944 4292 2972
rect 4667 2944 4712 2972
rect 3421 2907 3479 2913
rect 3421 2873 3433 2907
rect 3467 2904 3479 2907
rect 3970 2904 3976 2916
rect 3467 2876 3976 2904
rect 3467 2873 3479 2876
rect 3421 2867 3479 2873
rect 3970 2864 3976 2876
rect 4028 2864 4034 2916
rect 3694 2796 3700 2848
rect 3752 2836 3758 2848
rect 4264 2845 4292 2944
rect 4706 2932 4712 2944
rect 4764 2932 4770 2984
rect 6564 2904 6592 3003
rect 7374 3000 7380 3012
rect 7432 3000 7438 3052
rect 7466 3000 7472 3052
rect 7524 3040 7530 3052
rect 7524 3012 7569 3040
rect 7524 3000 7530 3012
rect 8018 3000 8024 3052
rect 8076 3040 8082 3052
rect 8297 3043 8355 3049
rect 8297 3040 8309 3043
rect 8076 3012 8309 3040
rect 8076 3000 8082 3012
rect 8297 3009 8309 3012
rect 8343 3040 8355 3043
rect 8478 3040 8484 3052
rect 8343 3012 8484 3040
rect 8343 3009 8355 3012
rect 8297 3003 8355 3009
rect 8478 3000 8484 3012
rect 8536 3000 8542 3052
rect 7009 2975 7067 2981
rect 7009 2941 7021 2975
rect 7055 2972 7067 2975
rect 8386 2972 8392 2984
rect 7055 2944 8392 2972
rect 7055 2941 7067 2944
rect 7009 2935 7067 2941
rect 8386 2932 8392 2944
rect 8444 2932 8450 2984
rect 9306 2904 9312 2916
rect 6564 2876 9312 2904
rect 9306 2864 9312 2876
rect 9364 2864 9370 2916
rect 4065 2839 4123 2845
rect 4065 2836 4077 2839
rect 3752 2808 4077 2836
rect 3752 2796 3758 2808
rect 4065 2805 4077 2808
rect 4111 2805 4123 2839
rect 4065 2799 4123 2805
rect 4249 2839 4307 2845
rect 4249 2805 4261 2839
rect 4295 2836 4307 2839
rect 4522 2836 4528 2848
rect 4295 2808 4528 2836
rect 4295 2805 4307 2808
rect 4249 2799 4307 2805
rect 4522 2796 4528 2808
rect 4580 2796 4586 2848
rect 4982 2796 4988 2848
rect 5040 2836 5046 2848
rect 7466 2836 7472 2848
rect 5040 2808 7472 2836
rect 5040 2796 5046 2808
rect 7466 2796 7472 2808
rect 7524 2796 7530 2848
rect 7558 2796 7564 2848
rect 7616 2836 7622 2848
rect 7929 2839 7987 2845
rect 7616 2808 7661 2836
rect 7616 2796 7622 2808
rect 7929 2805 7941 2839
rect 7975 2836 7987 2839
rect 8110 2836 8116 2848
rect 7975 2808 8116 2836
rect 7975 2805 7987 2808
rect 7929 2799 7987 2805
rect 8110 2796 8116 2808
rect 8168 2796 8174 2848
rect 8389 2839 8447 2845
rect 8389 2805 8401 2839
rect 8435 2836 8447 2839
rect 8662 2836 8668 2848
rect 8435 2808 8668 2836
rect 8435 2805 8447 2808
rect 8389 2799 8447 2805
rect 8662 2796 8668 2808
rect 8720 2796 8726 2848
rect 9401 2839 9459 2845
rect 9401 2805 9413 2839
rect 9447 2836 9459 2839
rect 13814 2836 13820 2848
rect 9447 2808 13820 2836
rect 9447 2805 9459 2808
rect 9401 2799 9459 2805
rect 13814 2796 13820 2808
rect 13872 2796 13878 2848
rect 3036 2746 9844 2768
rect 3036 2694 5666 2746
rect 5718 2694 5730 2746
rect 5782 2694 5794 2746
rect 5846 2694 5858 2746
rect 5910 2694 5922 2746
rect 5974 2694 8766 2746
rect 8818 2694 8830 2746
rect 8882 2694 8894 2746
rect 8946 2694 8958 2746
rect 9010 2694 9022 2746
rect 9074 2694 9844 2746
rect 3036 2672 9844 2694
rect 3513 2635 3571 2641
rect 3513 2601 3525 2635
rect 3559 2632 3571 2635
rect 5258 2632 5264 2644
rect 3559 2604 5264 2632
rect 3559 2601 3571 2604
rect 3513 2595 3571 2601
rect 5258 2592 5264 2604
rect 5316 2592 5322 2644
rect 6178 2592 6184 2644
rect 6236 2632 6242 2644
rect 7561 2635 7619 2641
rect 7561 2632 7573 2635
rect 6236 2604 7573 2632
rect 6236 2592 6242 2604
rect 7561 2601 7573 2604
rect 7607 2601 7619 2635
rect 7926 2632 7932 2644
rect 7887 2604 7932 2632
rect 7561 2595 7619 2601
rect 7926 2592 7932 2604
rect 7984 2592 7990 2644
rect 9122 2592 9128 2644
rect 9180 2632 9186 2644
rect 9217 2635 9275 2641
rect 9217 2632 9229 2635
rect 9180 2604 9229 2632
rect 9180 2592 9186 2604
rect 9217 2601 9229 2604
rect 9263 2601 9275 2635
rect 9217 2595 9275 2601
rect 9306 2592 9312 2644
rect 9364 2632 9370 2644
rect 9364 2604 9409 2632
rect 9364 2592 9370 2604
rect 5166 2524 5172 2576
rect 5224 2524 5230 2576
rect 5537 2567 5595 2573
rect 5537 2533 5549 2567
rect 5583 2564 5595 2567
rect 5583 2536 5856 2564
rect 5583 2533 5595 2536
rect 5537 2527 5595 2533
rect 3326 2456 3332 2508
rect 3384 2496 3390 2508
rect 3789 2499 3847 2505
rect 3789 2496 3801 2499
rect 3384 2468 3801 2496
rect 3384 2456 3390 2468
rect 3789 2465 3801 2468
rect 3835 2496 3847 2499
rect 5184 2496 5212 2524
rect 5721 2499 5779 2505
rect 5721 2496 5733 2499
rect 3835 2468 5733 2496
rect 3835 2465 3847 2468
rect 3789 2459 3847 2465
rect 5721 2465 5733 2468
rect 5767 2465 5779 2499
rect 5828 2496 5856 2536
rect 7374 2524 7380 2576
rect 7432 2564 7438 2576
rect 8665 2567 8723 2573
rect 8665 2564 8677 2567
rect 7432 2536 8677 2564
rect 7432 2524 7438 2536
rect 8665 2533 8677 2536
rect 8711 2533 8723 2567
rect 8665 2527 8723 2533
rect 5997 2499 6055 2505
rect 5997 2496 6009 2499
rect 5828 2468 6009 2496
rect 5721 2459 5779 2465
rect 5997 2465 6009 2468
rect 6043 2496 6055 2499
rect 6454 2496 6460 2508
rect 6043 2468 6460 2496
rect 6043 2465 6055 2468
rect 5997 2459 6055 2465
rect 6454 2456 6460 2468
rect 6512 2456 6518 2508
rect 6546 2456 6552 2508
rect 6604 2496 6610 2508
rect 6604 2468 7788 2496
rect 6604 2456 6610 2468
rect 3694 2428 3700 2440
rect 3655 2400 3700 2428
rect 3694 2388 3700 2400
rect 3752 2388 3758 2440
rect 7760 2437 7788 2468
rect 7745 2431 7803 2437
rect 7745 2397 7757 2431
rect 7791 2397 7803 2431
rect 8110 2428 8116 2440
rect 8071 2400 8116 2428
rect 7745 2391 7803 2397
rect 8110 2388 8116 2400
rect 8168 2388 8174 2440
rect 8294 2428 8300 2440
rect 8255 2400 8300 2428
rect 8294 2388 8300 2400
rect 8352 2388 8358 2440
rect 8386 2388 8392 2440
rect 8444 2428 8450 2440
rect 8849 2431 8907 2437
rect 8849 2428 8861 2431
rect 8444 2400 8861 2428
rect 8444 2388 8450 2400
rect 8849 2397 8861 2400
rect 8895 2397 8907 2431
rect 9490 2428 9496 2440
rect 9451 2400 9496 2428
rect 8849 2391 8907 2397
rect 9490 2388 9496 2400
rect 9548 2388 9554 2440
rect 4065 2363 4123 2369
rect 4065 2329 4077 2363
rect 4111 2360 4123 2363
rect 4338 2360 4344 2372
rect 4111 2332 4344 2360
rect 4111 2329 4123 2332
rect 4065 2323 4123 2329
rect 4338 2320 4344 2332
rect 4396 2320 4402 2372
rect 4522 2320 4528 2372
rect 4580 2320 4586 2372
rect 7558 2360 7564 2372
rect 7222 2332 7564 2360
rect 7558 2320 7564 2332
rect 7616 2360 7622 2372
rect 8481 2363 8539 2369
rect 8481 2360 8493 2363
rect 7616 2332 8493 2360
rect 7616 2320 7622 2332
rect 8481 2329 8493 2332
rect 8527 2360 8539 2363
rect 8662 2360 8668 2372
rect 8527 2332 8668 2360
rect 8527 2329 8539 2332
rect 8481 2323 8539 2329
rect 8662 2320 8668 2332
rect 8720 2360 8726 2372
rect 9033 2363 9091 2369
rect 9033 2360 9045 2363
rect 8720 2332 9045 2360
rect 8720 2320 8726 2332
rect 9033 2329 9045 2332
rect 9079 2329 9091 2363
rect 9033 2323 9091 2329
rect 6086 2252 6092 2304
rect 6144 2292 6150 2304
rect 7469 2295 7527 2301
rect 7469 2292 7481 2295
rect 6144 2264 7481 2292
rect 6144 2252 6150 2264
rect 7469 2261 7481 2264
rect 7515 2261 7527 2295
rect 7469 2255 7527 2261
rect 3036 2202 9844 2224
rect 3036 2150 4116 2202
rect 4168 2150 4180 2202
rect 4232 2150 4244 2202
rect 4296 2150 4308 2202
rect 4360 2150 4372 2202
rect 4424 2150 7216 2202
rect 7268 2150 7280 2202
rect 7332 2150 7344 2202
rect 7396 2150 7408 2202
rect 7460 2150 7472 2202
rect 7524 2150 9844 2202
rect 3036 2128 9844 2150
<< via1 >>
rect 1216 11772 1268 11824
rect 4988 11772 5040 11824
rect 3424 11704 3476 11756
rect 7656 11704 7708 11756
rect 3240 11636 3292 11688
rect 5080 11636 5132 11688
rect 6276 11636 6328 11688
rect 1860 11568 1912 11620
rect 16580 11568 16632 11620
rect 1308 11500 1360 11552
rect 8576 11500 8628 11552
rect 2566 11398 2618 11450
rect 2630 11398 2682 11450
rect 2694 11398 2746 11450
rect 2758 11398 2810 11450
rect 2822 11398 2874 11450
rect 5666 11398 5718 11450
rect 5730 11398 5782 11450
rect 5794 11398 5846 11450
rect 5858 11398 5910 11450
rect 5922 11398 5974 11450
rect 8766 11398 8818 11450
rect 8830 11398 8882 11450
rect 8894 11398 8946 11450
rect 8958 11398 9010 11450
rect 9022 11398 9074 11450
rect 1308 11339 1360 11348
rect 1308 11305 1317 11339
rect 1317 11305 1351 11339
rect 1351 11305 1360 11339
rect 1308 11296 1360 11305
rect 1860 11339 1912 11348
rect 1860 11305 1869 11339
rect 1869 11305 1903 11339
rect 1903 11305 1912 11339
rect 1860 11296 1912 11305
rect 6460 11296 6512 11348
rect 9680 11296 9732 11348
rect 3056 11228 3108 11280
rect 6000 11228 6052 11280
rect 6276 11271 6328 11280
rect 6276 11237 6285 11271
rect 6285 11237 6319 11271
rect 6319 11237 6328 11271
rect 6276 11228 6328 11237
rect 9496 11228 9548 11280
rect 1860 11092 1912 11144
rect 2412 11092 2464 11144
rect 3148 11135 3200 11144
rect 3148 11101 3157 11135
rect 3157 11101 3191 11135
rect 3191 11101 3200 11135
rect 3148 11092 3200 11101
rect 3424 11135 3476 11144
rect 3424 11101 3433 11135
rect 3433 11101 3467 11135
rect 3467 11101 3476 11135
rect 3424 11092 3476 11101
rect 3608 11135 3660 11144
rect 3608 11101 3617 11135
rect 3617 11101 3651 11135
rect 3651 11101 3660 11135
rect 3608 11092 3660 11101
rect 5264 11092 5316 11144
rect 7104 11160 7156 11212
rect 7932 11203 7984 11212
rect 7932 11169 7941 11203
rect 7941 11169 7975 11203
rect 7975 11169 7984 11203
rect 7932 11160 7984 11169
rect 6184 11135 6236 11144
rect 6184 11101 6193 11135
rect 6193 11101 6227 11135
rect 6227 11101 6236 11135
rect 6184 11092 6236 11101
rect 6828 11135 6880 11144
rect 2412 10956 2464 11008
rect 3976 11024 4028 11076
rect 4344 11024 4396 11076
rect 6828 11101 6837 11135
rect 6837 11101 6871 11135
rect 6871 11101 6880 11135
rect 6828 11092 6880 11101
rect 8300 11092 8352 11144
rect 9220 11135 9272 11144
rect 9220 11101 9229 11135
rect 9229 11101 9263 11135
rect 9263 11101 9272 11135
rect 9220 11092 9272 11101
rect 6184 10956 6236 11008
rect 6368 10956 6420 11008
rect 13820 11024 13872 11076
rect 9404 10999 9456 11008
rect 9404 10965 9413 10999
rect 9413 10965 9447 10999
rect 9447 10965 9456 10999
rect 9404 10956 9456 10965
rect 4116 10854 4168 10906
rect 4180 10854 4232 10906
rect 4244 10854 4296 10906
rect 4308 10854 4360 10906
rect 4372 10854 4424 10906
rect 7216 10854 7268 10906
rect 7280 10854 7332 10906
rect 7344 10854 7396 10906
rect 7408 10854 7460 10906
rect 7472 10854 7524 10906
rect 2320 10659 2372 10668
rect 2320 10625 2329 10659
rect 2329 10625 2363 10659
rect 2363 10625 2372 10659
rect 2320 10616 2372 10625
rect 3424 10684 3476 10736
rect 4804 10659 4856 10668
rect 4804 10625 4813 10659
rect 4813 10625 4847 10659
rect 4847 10625 4856 10659
rect 4804 10616 4856 10625
rect 5080 10659 5132 10668
rect 5080 10625 5089 10659
rect 5089 10625 5123 10659
rect 5123 10625 5132 10659
rect 5080 10616 5132 10625
rect 5540 10616 5592 10668
rect 1492 10523 1544 10532
rect 1492 10489 1501 10523
rect 1501 10489 1535 10523
rect 1535 10489 1544 10523
rect 1492 10480 1544 10489
rect 2412 10523 2464 10532
rect 2412 10489 2421 10523
rect 2421 10489 2455 10523
rect 2455 10489 2464 10523
rect 2412 10480 2464 10489
rect 2136 10455 2188 10464
rect 2136 10421 2145 10455
rect 2145 10421 2179 10455
rect 2179 10421 2188 10455
rect 2136 10412 2188 10421
rect 3516 10548 3568 10600
rect 3976 10548 4028 10600
rect 4344 10548 4396 10600
rect 6000 10548 6052 10600
rect 6276 10548 6328 10600
rect 5264 10480 5316 10532
rect 6092 10480 6144 10532
rect 6920 10684 6972 10736
rect 6552 10659 6604 10668
rect 6552 10625 6561 10659
rect 6561 10625 6595 10659
rect 6595 10625 6604 10659
rect 6552 10616 6604 10625
rect 7932 10616 7984 10668
rect 8208 10616 8260 10668
rect 8484 10659 8536 10668
rect 8484 10625 8493 10659
rect 8493 10625 8527 10659
rect 8527 10625 8536 10659
rect 8484 10616 8536 10625
rect 6460 10548 6512 10600
rect 6920 10548 6972 10600
rect 9128 10616 9180 10668
rect 16764 10548 16816 10600
rect 3056 10412 3108 10464
rect 3608 10412 3660 10464
rect 3700 10412 3752 10464
rect 5080 10412 5132 10464
rect 5356 10412 5408 10464
rect 6460 10412 6512 10464
rect 6552 10412 6604 10464
rect 8300 10455 8352 10464
rect 8300 10421 8309 10455
rect 8309 10421 8343 10455
rect 8343 10421 8352 10455
rect 8300 10412 8352 10421
rect 13544 10412 13596 10464
rect 2566 10310 2618 10362
rect 2630 10310 2682 10362
rect 2694 10310 2746 10362
rect 2758 10310 2810 10362
rect 2822 10310 2874 10362
rect 5666 10310 5718 10362
rect 5730 10310 5782 10362
rect 5794 10310 5846 10362
rect 5858 10310 5910 10362
rect 5922 10310 5974 10362
rect 8766 10310 8818 10362
rect 8830 10310 8882 10362
rect 8894 10310 8946 10362
rect 8958 10310 9010 10362
rect 9022 10310 9074 10362
rect 3792 10208 3844 10260
rect 4068 10208 4120 10260
rect 9220 10208 9272 10260
rect 2412 10140 2464 10192
rect 3608 10183 3660 10192
rect 3608 10149 3617 10183
rect 3617 10149 3651 10183
rect 3651 10149 3660 10183
rect 3608 10140 3660 10149
rect 2136 10072 2188 10124
rect 5264 10140 5316 10192
rect 6092 10140 6144 10192
rect 6368 10140 6420 10192
rect 7840 10140 7892 10192
rect 8392 10140 8444 10192
rect 4344 10115 4396 10124
rect 4344 10081 4353 10115
rect 4353 10081 4387 10115
rect 4387 10081 4396 10115
rect 4344 10072 4396 10081
rect 6736 10072 6788 10124
rect 9312 10115 9364 10124
rect 9312 10081 9321 10115
rect 9321 10081 9355 10115
rect 9355 10081 9364 10115
rect 9312 10072 9364 10081
rect 2964 10004 3016 10056
rect 3240 10004 3292 10056
rect 3884 10047 3936 10056
rect 3884 10013 3893 10047
rect 3893 10013 3927 10047
rect 3927 10013 3936 10047
rect 3884 10004 3936 10013
rect 5356 10004 5408 10056
rect 6368 10047 6420 10056
rect 6368 10013 6377 10047
rect 6377 10013 6411 10047
rect 6411 10013 6420 10047
rect 6368 10004 6420 10013
rect 7932 10004 7984 10056
rect 8576 10004 8628 10056
rect 2136 9936 2188 9988
rect 2964 9868 3016 9920
rect 3424 9868 3476 9920
rect 3700 9868 3752 9920
rect 4620 9936 4672 9988
rect 6184 9936 6236 9988
rect 6736 9936 6788 9988
rect 8208 9979 8260 9988
rect 5632 9868 5684 9920
rect 6460 9868 6512 9920
rect 7012 9868 7064 9920
rect 8208 9945 8217 9979
rect 8217 9945 8251 9979
rect 8251 9945 8260 9979
rect 8208 9936 8260 9945
rect 9220 9911 9272 9920
rect 9220 9877 9229 9911
rect 9229 9877 9263 9911
rect 9263 9877 9272 9911
rect 9220 9868 9272 9877
rect 4116 9766 4168 9818
rect 4180 9766 4232 9818
rect 4244 9766 4296 9818
rect 4308 9766 4360 9818
rect 4372 9766 4424 9818
rect 7216 9766 7268 9818
rect 7280 9766 7332 9818
rect 7344 9766 7396 9818
rect 7408 9766 7460 9818
rect 7472 9766 7524 9818
rect 13820 9732 13872 9784
rect 2964 9664 3016 9716
rect 3240 9664 3292 9716
rect 1032 9528 1084 9580
rect 2412 9571 2464 9580
rect 1124 9460 1176 9512
rect 2412 9537 2421 9571
rect 2421 9537 2455 9571
rect 2455 9537 2464 9571
rect 2412 9528 2464 9537
rect 2780 9596 2832 9648
rect 4528 9664 4580 9716
rect 4804 9664 4856 9716
rect 3700 9596 3752 9648
rect 4436 9596 4488 9648
rect 5632 9664 5684 9716
rect 7932 9664 7984 9716
rect 9128 9664 9180 9716
rect 9312 9707 9364 9716
rect 9312 9673 9321 9707
rect 9321 9673 9355 9707
rect 9355 9673 9364 9707
rect 9312 9664 9364 9673
rect 4344 9528 4396 9580
rect 5080 9528 5132 9580
rect 3056 9460 3108 9512
rect 4068 9460 4120 9512
rect 5816 9571 5868 9580
rect 5816 9537 5825 9571
rect 5825 9537 5859 9571
rect 5859 9537 5868 9571
rect 5816 9528 5868 9537
rect 6000 9571 6052 9580
rect 6000 9537 6009 9571
rect 6009 9537 6043 9571
rect 6043 9537 6052 9571
rect 6000 9528 6052 9537
rect 6920 9528 6972 9580
rect 7380 9571 7432 9580
rect 7380 9537 7389 9571
rect 7389 9537 7423 9571
rect 7423 9537 7432 9571
rect 7380 9528 7432 9537
rect 1952 9392 2004 9444
rect 2688 9392 2740 9444
rect 4160 9392 4212 9444
rect 7104 9460 7156 9512
rect 5816 9392 5868 9444
rect 1400 9324 1452 9376
rect 1584 9367 1636 9376
rect 1584 9333 1593 9367
rect 1593 9333 1627 9367
rect 1627 9333 1636 9367
rect 1584 9324 1636 9333
rect 1768 9324 1820 9376
rect 3608 9324 3660 9376
rect 4344 9324 4396 9376
rect 4528 9367 4580 9376
rect 4528 9333 4537 9367
rect 4537 9333 4571 9367
rect 4571 9333 4580 9367
rect 4528 9324 4580 9333
rect 4712 9324 4764 9376
rect 6460 9367 6512 9376
rect 6460 9333 6469 9367
rect 6469 9333 6503 9367
rect 6503 9333 6512 9367
rect 6460 9324 6512 9333
rect 6736 9324 6788 9376
rect 2566 9222 2618 9274
rect 2630 9222 2682 9274
rect 2694 9222 2746 9274
rect 2758 9222 2810 9274
rect 2822 9222 2874 9274
rect 5666 9222 5718 9274
rect 5730 9222 5782 9274
rect 5794 9222 5846 9274
rect 5858 9222 5910 9274
rect 5922 9222 5974 9274
rect 8766 9222 8818 9274
rect 8830 9222 8882 9274
rect 8894 9222 8946 9274
rect 8958 9222 9010 9274
rect 9022 9222 9074 9274
rect 1860 9095 1912 9104
rect 1860 9061 1869 9095
rect 1869 9061 1903 9095
rect 1903 9061 1912 9095
rect 1860 9052 1912 9061
rect 2044 9095 2096 9104
rect 2044 9061 2053 9095
rect 2053 9061 2087 9095
rect 2087 9061 2096 9095
rect 2044 9052 2096 9061
rect 2320 9120 2372 9172
rect 3516 9120 3568 9172
rect 3792 9120 3844 9172
rect 4620 9120 4672 9172
rect 4804 9120 4856 9172
rect 6828 9120 6880 9172
rect 8208 9163 8260 9172
rect 8208 9129 8217 9163
rect 8217 9129 8251 9163
rect 8251 9129 8260 9163
rect 8208 9120 8260 9129
rect 8484 9120 8536 9172
rect 1676 8959 1728 8968
rect 1676 8925 1685 8959
rect 1685 8925 1719 8959
rect 1719 8925 1728 8959
rect 1676 8916 1728 8925
rect 2320 8984 2372 9036
rect 2228 8959 2280 8968
rect 2228 8925 2237 8959
rect 2237 8925 2271 8959
rect 2271 8925 2280 8959
rect 2228 8916 2280 8925
rect 3332 8984 3384 9036
rect 3148 8959 3200 8968
rect 3148 8925 3157 8959
rect 3157 8925 3191 8959
rect 3191 8925 3200 8959
rect 3148 8916 3200 8925
rect 3608 8916 3660 8968
rect 3056 8848 3108 8900
rect 3332 8848 3384 8900
rect 4068 8959 4120 8968
rect 4068 8925 4077 8959
rect 4077 8925 4111 8959
rect 4111 8925 4120 8959
rect 4068 8916 4120 8925
rect 4252 8848 4304 8900
rect 4896 8916 4948 8968
rect 5172 9027 5224 9036
rect 5172 8993 5187 9027
rect 5187 8993 5221 9027
rect 5221 8993 5224 9027
rect 5172 8984 5224 8993
rect 6184 8984 6236 9036
rect 10140 9052 10192 9104
rect 8668 8984 8720 9036
rect 9312 9027 9364 9036
rect 9312 8993 9321 9027
rect 9321 8993 9355 9027
rect 9355 8993 9364 9027
rect 9312 8984 9364 8993
rect 5632 8916 5684 8968
rect 7012 8959 7064 8968
rect 7012 8925 7021 8959
rect 7021 8925 7055 8959
rect 7055 8925 7064 8959
rect 7012 8916 7064 8925
rect 7748 8959 7800 8968
rect 7748 8925 7757 8959
rect 7757 8925 7791 8959
rect 7791 8925 7800 8959
rect 7748 8916 7800 8925
rect 7840 8916 7892 8968
rect 8208 8916 8260 8968
rect 5172 8848 5224 8900
rect 5908 8848 5960 8900
rect 6920 8848 6972 8900
rect 13452 8848 13504 8900
rect 22376 8848 22428 8900
rect 2964 8823 3016 8832
rect 2964 8789 2973 8823
rect 2973 8789 3007 8823
rect 3007 8789 3016 8823
rect 2964 8780 3016 8789
rect 3700 8780 3752 8832
rect 3884 8823 3936 8832
rect 3884 8789 3893 8823
rect 3893 8789 3927 8823
rect 3927 8789 3936 8823
rect 3884 8780 3936 8789
rect 3976 8780 4028 8832
rect 4712 8780 4764 8832
rect 5816 8780 5868 8832
rect 6276 8780 6328 8832
rect 6552 8780 6604 8832
rect 8392 8780 8444 8832
rect 4116 8678 4168 8730
rect 4180 8678 4232 8730
rect 4244 8678 4296 8730
rect 4308 8678 4360 8730
rect 4372 8678 4424 8730
rect 7216 8678 7268 8730
rect 7280 8678 7332 8730
rect 7344 8678 7396 8730
rect 7408 8678 7460 8730
rect 7472 8678 7524 8730
rect 1492 8619 1544 8628
rect 1492 8585 1501 8619
rect 1501 8585 1535 8619
rect 1535 8585 1544 8619
rect 1492 8576 1544 8585
rect 1860 8576 1912 8628
rect 2044 8576 2096 8628
rect 2872 8576 2924 8628
rect 4896 8576 4948 8628
rect 5080 8576 5132 8628
rect 5356 8576 5408 8628
rect 6368 8576 6420 8628
rect 9588 8576 9640 8628
rect 1216 8508 1268 8560
rect 2228 8508 2280 8560
rect 2320 8440 2372 8492
rect 3056 8508 3108 8560
rect 4804 8508 4856 8560
rect 6000 8508 6052 8560
rect 6184 8508 6236 8560
rect 2964 8483 3016 8492
rect 2964 8449 2973 8483
rect 2973 8449 3007 8483
rect 3007 8449 3016 8483
rect 2964 8440 3016 8449
rect 2688 8372 2740 8424
rect 5080 8467 5132 8476
rect 5080 8433 5089 8467
rect 5089 8433 5123 8467
rect 5123 8433 5132 8467
rect 5080 8424 5132 8433
rect 3884 8372 3936 8424
rect 4528 8372 4580 8424
rect 1768 8347 1820 8356
rect 1768 8313 1777 8347
rect 1777 8313 1811 8347
rect 1811 8313 1820 8347
rect 1768 8304 1820 8313
rect 4436 8304 4488 8356
rect 1216 8279 1268 8288
rect 1216 8245 1225 8279
rect 1225 8245 1259 8279
rect 1259 8245 1268 8279
rect 1216 8236 1268 8245
rect 4528 8236 4580 8288
rect 5172 8236 5224 8288
rect 7104 8508 7156 8560
rect 8208 8508 8260 8560
rect 6460 8483 6512 8492
rect 6460 8449 6469 8483
rect 6469 8449 6503 8483
rect 6503 8449 6512 8483
rect 6736 8483 6788 8492
rect 6460 8440 6512 8449
rect 6736 8449 6745 8483
rect 6745 8449 6779 8483
rect 6779 8449 6788 8483
rect 6736 8440 6788 8449
rect 6828 8440 6880 8492
rect 8300 8440 8352 8492
rect 8392 8483 8444 8492
rect 8392 8449 8401 8483
rect 8401 8449 8435 8483
rect 8435 8449 8444 8483
rect 8576 8483 8628 8492
rect 8392 8440 8444 8449
rect 8576 8449 8585 8483
rect 8585 8449 8619 8483
rect 8619 8449 8628 8483
rect 8576 8440 8628 8449
rect 8668 8483 8720 8492
rect 8668 8449 8677 8483
rect 8677 8449 8711 8483
rect 8711 8449 8720 8483
rect 8668 8440 8720 8449
rect 6276 8372 6328 8424
rect 7012 8372 7064 8424
rect 7840 8372 7892 8424
rect 10876 8372 10928 8424
rect 5724 8304 5776 8356
rect 6368 8304 6420 8356
rect 6552 8304 6604 8356
rect 13820 8508 13872 8560
rect 5448 8236 5500 8288
rect 8484 8236 8536 8288
rect 2566 8134 2618 8186
rect 2630 8134 2682 8186
rect 2694 8134 2746 8186
rect 2758 8134 2810 8186
rect 2822 8134 2874 8186
rect 5666 8134 5718 8186
rect 5730 8134 5782 8186
rect 5794 8134 5846 8186
rect 5858 8134 5910 8186
rect 5922 8134 5974 8186
rect 8766 8134 8818 8186
rect 8830 8134 8882 8186
rect 8894 8134 8946 8186
rect 8958 8134 9010 8186
rect 9022 8134 9074 8186
rect 3056 8032 3108 8084
rect 3148 8032 3200 8084
rect 6184 8032 6236 8084
rect 7748 8032 7800 8084
rect 8024 8075 8076 8084
rect 8024 8041 8033 8075
rect 8033 8041 8067 8075
rect 8067 8041 8076 8075
rect 8024 8032 8076 8041
rect 2136 7964 2188 8016
rect 2412 7964 2464 8016
rect 3700 7964 3752 8016
rect 2964 7896 3016 7948
rect 4436 7964 4488 8016
rect 4896 7964 4948 8016
rect 9220 8032 9272 8084
rect 1768 7871 1820 7880
rect 1768 7837 1777 7871
rect 1777 7837 1811 7871
rect 1811 7837 1820 7871
rect 1768 7828 1820 7837
rect 2044 7871 2096 7880
rect 2044 7837 2053 7871
rect 2053 7837 2087 7871
rect 2087 7837 2096 7871
rect 2044 7828 2096 7837
rect 2688 7871 2740 7880
rect 1032 7760 1084 7812
rect 2688 7837 2697 7871
rect 2697 7837 2731 7871
rect 2731 7837 2740 7871
rect 2688 7828 2740 7837
rect 3792 7828 3844 7880
rect 4528 7896 4580 7948
rect 5448 7896 5500 7948
rect 5172 7871 5224 7880
rect 5172 7837 5181 7871
rect 5181 7837 5215 7871
rect 5215 7837 5224 7871
rect 5172 7828 5224 7837
rect 6644 7871 6696 7880
rect 6644 7837 6653 7871
rect 6653 7837 6687 7871
rect 6687 7837 6696 7871
rect 6644 7828 6696 7837
rect 7932 7896 7984 7948
rect 7748 7871 7800 7880
rect 7748 7837 7757 7871
rect 7757 7837 7791 7871
rect 7791 7837 7800 7871
rect 7748 7828 7800 7837
rect 8392 7828 8444 7880
rect 13544 7964 13596 8016
rect 9312 7939 9364 7948
rect 9312 7905 9321 7939
rect 9321 7905 9355 7939
rect 9355 7905 9364 7939
rect 9312 7896 9364 7905
rect 13636 7828 13688 7880
rect 1124 7692 1176 7744
rect 2228 7692 2280 7744
rect 3148 7692 3200 7744
rect 3424 7735 3476 7744
rect 3424 7701 3433 7735
rect 3433 7701 3467 7735
rect 3467 7701 3476 7735
rect 3424 7692 3476 7701
rect 3516 7692 3568 7744
rect 4528 7735 4580 7744
rect 4528 7701 4537 7735
rect 4537 7701 4571 7735
rect 4571 7701 4580 7735
rect 4528 7692 4580 7701
rect 5540 7760 5592 7812
rect 6828 7760 6880 7812
rect 8484 7692 8536 7744
rect 9128 7735 9180 7744
rect 9128 7701 9137 7735
rect 9137 7701 9171 7735
rect 9171 7701 9180 7735
rect 9128 7692 9180 7701
rect 9220 7735 9272 7744
rect 9220 7701 9229 7735
rect 9229 7701 9263 7735
rect 9263 7701 9272 7735
rect 9220 7692 9272 7701
rect 13728 7692 13780 7744
rect 4116 7590 4168 7642
rect 4180 7590 4232 7642
rect 4244 7590 4296 7642
rect 4308 7590 4360 7642
rect 4372 7590 4424 7642
rect 7216 7590 7268 7642
rect 7280 7590 7332 7642
rect 7344 7590 7396 7642
rect 7408 7590 7460 7642
rect 7472 7590 7524 7642
rect 13452 7624 13504 7676
rect 22284 7624 22336 7676
rect 2136 7488 2188 7540
rect 3056 7488 3108 7540
rect 3240 7488 3292 7540
rect 4896 7488 4948 7540
rect 4988 7488 5040 7540
rect 5908 7488 5960 7540
rect 7748 7488 7800 7540
rect 7840 7488 7892 7540
rect 8024 7488 8076 7540
rect 8484 7488 8536 7540
rect 1768 7420 1820 7472
rect 4344 7420 4396 7472
rect 8116 7420 8168 7472
rect 8576 7420 8628 7472
rect 2780 7395 2832 7404
rect 2320 7284 2372 7336
rect 2412 7216 2464 7268
rect 2780 7361 2789 7395
rect 2789 7361 2823 7395
rect 2823 7361 2832 7395
rect 2780 7352 2832 7361
rect 3056 7395 3108 7404
rect 3056 7361 3065 7395
rect 3065 7361 3099 7395
rect 3099 7361 3108 7395
rect 3056 7352 3108 7361
rect 4068 7395 4120 7404
rect 3516 7284 3568 7336
rect 4068 7361 4077 7395
rect 4077 7361 4111 7395
rect 4111 7361 4120 7395
rect 4068 7352 4120 7361
rect 6000 7352 6052 7404
rect 6184 7395 6236 7404
rect 6184 7361 6193 7395
rect 6193 7361 6227 7395
rect 6227 7361 6236 7395
rect 6184 7352 6236 7361
rect 8668 7395 8720 7404
rect 8668 7361 8677 7395
rect 8677 7361 8711 7395
rect 8711 7361 8720 7395
rect 8668 7352 8720 7361
rect 4528 7284 4580 7336
rect 1400 7191 1452 7200
rect 1400 7157 1409 7191
rect 1409 7157 1443 7191
rect 1443 7157 1452 7191
rect 1400 7148 1452 7157
rect 3608 7216 3660 7268
rect 5080 7216 5132 7268
rect 5356 7216 5408 7268
rect 3240 7148 3292 7200
rect 5632 7216 5684 7268
rect 7564 7284 7616 7336
rect 13820 7284 13872 7336
rect 19432 7284 19484 7336
rect 9036 7216 9088 7268
rect 6460 7191 6512 7200
rect 6460 7157 6469 7191
rect 6469 7157 6503 7191
rect 6503 7157 6512 7191
rect 6460 7148 6512 7157
rect 6644 7191 6696 7200
rect 6644 7157 6653 7191
rect 6653 7157 6687 7191
rect 6687 7157 6696 7191
rect 6644 7148 6696 7157
rect 13728 7148 13780 7200
rect 2566 7046 2618 7098
rect 2630 7046 2682 7098
rect 2694 7046 2746 7098
rect 2758 7046 2810 7098
rect 2822 7046 2874 7098
rect 5666 7046 5718 7098
rect 5730 7046 5782 7098
rect 5794 7046 5846 7098
rect 5858 7046 5910 7098
rect 5922 7046 5974 7098
rect 8766 7046 8818 7098
rect 8830 7046 8882 7098
rect 8894 7046 8946 7098
rect 8958 7046 9010 7098
rect 9022 7046 9074 7098
rect 2044 6944 2096 6996
rect 4252 6944 4304 6996
rect 5080 6944 5132 6996
rect 6460 6944 6512 6996
rect 7104 6944 7156 6996
rect 9220 6944 9272 6996
rect 3516 6876 3568 6928
rect 3700 6876 3752 6928
rect 6644 6876 6696 6928
rect 8208 6876 8260 6928
rect 1676 6808 1728 6860
rect 1768 6783 1820 6792
rect 1768 6749 1777 6783
rect 1777 6749 1811 6783
rect 1811 6749 1820 6783
rect 1768 6740 1820 6749
rect 2136 6783 2188 6792
rect 2136 6749 2145 6783
rect 2145 6749 2179 6783
rect 2179 6749 2188 6783
rect 2136 6740 2188 6749
rect 2228 6740 2280 6792
rect 4252 6808 4304 6860
rect 4988 6808 5040 6860
rect 5356 6808 5408 6860
rect 5816 6808 5868 6860
rect 9312 6851 9364 6860
rect 9312 6817 9321 6851
rect 9321 6817 9355 6851
rect 9355 6817 9364 6851
rect 9312 6808 9364 6817
rect 3884 6740 3936 6792
rect 4528 6740 4580 6792
rect 5632 6672 5684 6724
rect 6828 6740 6880 6792
rect 8208 6783 8260 6792
rect 8208 6749 8217 6783
rect 8217 6749 8251 6783
rect 8251 6749 8260 6783
rect 8208 6740 8260 6749
rect 8300 6783 8352 6792
rect 8300 6749 8309 6783
rect 8309 6749 8343 6783
rect 8343 6749 8352 6783
rect 9128 6783 9180 6792
rect 8300 6740 8352 6749
rect 9128 6749 9137 6783
rect 9137 6749 9171 6783
rect 9171 6749 9180 6783
rect 9128 6740 9180 6749
rect 9404 6740 9456 6792
rect 1400 6604 1452 6656
rect 1584 6647 1636 6656
rect 1584 6613 1593 6647
rect 1593 6613 1627 6647
rect 1627 6613 1636 6647
rect 1584 6604 1636 6613
rect 2044 6604 2096 6656
rect 2228 6647 2280 6656
rect 2228 6613 2237 6647
rect 2237 6613 2271 6647
rect 2271 6613 2280 6647
rect 2228 6604 2280 6613
rect 2688 6604 2740 6656
rect 2872 6604 2924 6656
rect 3516 6604 3568 6656
rect 3700 6604 3752 6656
rect 5264 6604 5316 6656
rect 5448 6604 5500 6656
rect 8116 6672 8168 6724
rect 9588 6672 9640 6724
rect 5908 6604 5960 6656
rect 7656 6604 7708 6656
rect 4116 6502 4168 6554
rect 4180 6502 4232 6554
rect 4244 6502 4296 6554
rect 4308 6502 4360 6554
rect 4372 6502 4424 6554
rect 7216 6502 7268 6554
rect 7280 6502 7332 6554
rect 7344 6502 7396 6554
rect 7408 6502 7460 6554
rect 7472 6502 7524 6554
rect 1584 6443 1636 6452
rect 1584 6409 1593 6443
rect 1593 6409 1627 6443
rect 1627 6409 1636 6443
rect 1584 6400 1636 6409
rect 2228 6443 2280 6452
rect 2228 6409 2237 6443
rect 2237 6409 2271 6443
rect 2271 6409 2280 6443
rect 2228 6400 2280 6409
rect 3148 6400 3200 6452
rect 3424 6400 3476 6452
rect 2136 6332 2188 6384
rect 2872 6332 2924 6384
rect 5172 6400 5224 6452
rect 5264 6400 5316 6452
rect 5080 6332 5132 6384
rect 5540 6332 5592 6384
rect 6460 6332 6512 6384
rect 6920 6332 6972 6384
rect 7748 6375 7800 6384
rect 7748 6341 7757 6375
rect 7757 6341 7791 6375
rect 7791 6341 7800 6375
rect 13636 6400 13688 6452
rect 7748 6332 7800 6341
rect 3332 6307 3384 6316
rect 3332 6273 3341 6307
rect 3341 6273 3375 6307
rect 3375 6273 3384 6307
rect 3332 6264 3384 6273
rect 1768 6196 1820 6248
rect 3148 6196 3200 6248
rect 3700 6196 3752 6248
rect 5172 6239 5224 6248
rect 5172 6205 5181 6239
rect 5181 6205 5215 6239
rect 5215 6205 5224 6239
rect 5172 6196 5224 6205
rect 7012 6307 7064 6316
rect 7012 6273 7021 6307
rect 7021 6273 7055 6307
rect 7055 6273 7064 6307
rect 7012 6264 7064 6273
rect 7472 6264 7524 6316
rect 13820 6332 13872 6384
rect 8392 6196 8444 6248
rect 7288 6128 7340 6180
rect 3608 6060 3660 6112
rect 6092 6060 6144 6112
rect 7564 6060 7616 6112
rect 7932 6128 7984 6180
rect 9496 6128 9548 6180
rect 8392 6103 8444 6112
rect 8392 6069 8401 6103
rect 8401 6069 8435 6103
rect 8435 6069 8444 6103
rect 8392 6060 8444 6069
rect 8484 6060 8536 6112
rect 9128 6060 9180 6112
rect 9404 6060 9456 6112
rect 1492 5924 1544 5976
rect 2504 5924 2556 5976
rect 5666 5958 5718 6010
rect 5730 5958 5782 6010
rect 5794 5958 5846 6010
rect 5858 5958 5910 6010
rect 5922 5958 5974 6010
rect 8766 5958 8818 6010
rect 8830 5958 8882 6010
rect 8894 5958 8946 6010
rect 8958 5958 9010 6010
rect 9022 5958 9074 6010
rect 1860 5856 1912 5908
rect 6644 5856 6696 5908
rect 7472 5856 7524 5908
rect 7932 5856 7984 5908
rect 13728 5856 13780 5908
rect 1676 5788 1728 5840
rect 2596 5788 2648 5840
rect 5080 5788 5132 5840
rect 12808 5788 12860 5840
rect 6092 5763 6144 5772
rect 3332 5695 3384 5704
rect 3332 5661 3341 5695
rect 3341 5661 3375 5695
rect 3375 5661 3384 5695
rect 3332 5652 3384 5661
rect 6092 5729 6101 5763
rect 6101 5729 6135 5763
rect 6135 5729 6144 5763
rect 6092 5720 6144 5729
rect 9680 5720 9732 5772
rect 5080 5652 5132 5704
rect 5448 5652 5500 5704
rect 5632 5652 5684 5704
rect 7932 5652 7984 5704
rect 8668 5695 8720 5704
rect 8668 5661 8677 5695
rect 8677 5661 8711 5695
rect 8711 5661 8720 5695
rect 8668 5652 8720 5661
rect 9128 5695 9180 5704
rect 9128 5661 9137 5695
rect 9137 5661 9171 5695
rect 9171 5661 9180 5695
rect 9128 5652 9180 5661
rect 1400 5584 1452 5636
rect 2688 5584 2740 5636
rect 3608 5627 3660 5636
rect 3608 5593 3617 5627
rect 3617 5593 3651 5627
rect 3651 5593 3660 5627
rect 3608 5584 3660 5593
rect 4988 5584 5040 5636
rect 3792 5516 3844 5568
rect 5356 5559 5408 5568
rect 5356 5525 5365 5559
rect 5365 5525 5399 5559
rect 5399 5525 5408 5559
rect 5356 5516 5408 5525
rect 7656 5584 7708 5636
rect 8392 5584 8444 5636
rect 9220 5516 9272 5568
rect 4116 5414 4168 5466
rect 4180 5414 4232 5466
rect 4244 5414 4296 5466
rect 4308 5414 4360 5466
rect 4372 5414 4424 5466
rect 7216 5414 7268 5466
rect 7280 5414 7332 5466
rect 7344 5414 7396 5466
rect 7408 5414 7460 5466
rect 7472 5414 7524 5466
rect 5080 5312 5132 5364
rect 4712 5244 4764 5296
rect 6092 5244 6144 5296
rect 6460 5244 6512 5296
rect 7748 5312 7800 5364
rect 8668 5312 8720 5364
rect 8760 5312 8812 5364
rect 9128 5355 9180 5364
rect 9128 5321 9137 5355
rect 9137 5321 9171 5355
rect 9171 5321 9180 5355
rect 9128 5312 9180 5321
rect 9588 5312 9640 5364
rect 3240 5176 3292 5228
rect 3608 5176 3660 5228
rect 4804 5176 4856 5228
rect 2780 5108 2832 5160
rect 5448 5108 5500 5160
rect 6644 5108 6696 5160
rect 3240 5040 3292 5092
rect 8668 5219 8720 5228
rect 8668 5185 8677 5219
rect 8677 5185 8711 5219
rect 8711 5185 8720 5219
rect 8668 5176 8720 5185
rect 9496 5176 9548 5228
rect 9496 5040 9548 5092
rect 2780 4972 2832 5024
rect 5264 4972 5316 5024
rect 7840 4972 7892 5024
rect 8116 5015 8168 5024
rect 8116 4981 8125 5015
rect 8125 4981 8159 5015
rect 8159 4981 8168 5015
rect 8116 4972 8168 4981
rect 8484 5015 8536 5024
rect 8484 4981 8493 5015
rect 8493 4981 8527 5015
rect 8527 4981 8536 5015
rect 8484 4972 8536 4981
rect 2780 4836 2832 4888
rect 5666 4870 5718 4922
rect 5730 4870 5782 4922
rect 5794 4870 5846 4922
rect 5858 4870 5910 4922
rect 5922 4870 5974 4922
rect 8766 4870 8818 4922
rect 8830 4870 8882 4922
rect 8894 4870 8946 4922
rect 8958 4870 9010 4922
rect 9022 4870 9074 4922
rect 3056 4768 3108 4820
rect 4344 4768 4396 4820
rect 4436 4811 4488 4820
rect 4436 4777 4445 4811
rect 4445 4777 4479 4811
rect 4479 4777 4488 4811
rect 4436 4768 4488 4777
rect 4620 4811 4672 4820
rect 4620 4777 4629 4811
rect 4629 4777 4663 4811
rect 4663 4777 4672 4811
rect 4620 4768 4672 4777
rect 6368 4768 6420 4820
rect 6460 4768 6512 4820
rect 8208 4768 8260 4820
rect 9128 4768 9180 4820
rect 5540 4700 5592 4752
rect 5356 4632 5408 4684
rect 7472 4632 7524 4684
rect 7748 4632 7800 4684
rect 4160 4607 4212 4616
rect 4160 4573 4169 4607
rect 4169 4573 4203 4607
rect 4203 4573 4212 4607
rect 4160 4564 4212 4573
rect 4344 4564 4396 4616
rect 4988 4607 5040 4616
rect 4988 4573 4997 4607
rect 4997 4573 5031 4607
rect 5031 4573 5040 4607
rect 4988 4564 5040 4573
rect 5172 4564 5224 4616
rect 5448 4564 5500 4616
rect 6644 4607 6696 4616
rect 6644 4573 6653 4607
rect 6653 4573 6687 4607
rect 6687 4573 6696 4607
rect 6644 4564 6696 4573
rect 9220 4564 9272 4616
rect 5724 4539 5776 4548
rect 4712 4428 4764 4480
rect 5724 4505 5733 4539
rect 5733 4505 5767 4539
rect 5767 4505 5776 4539
rect 5724 4496 5776 4505
rect 5908 4539 5960 4548
rect 5908 4505 5917 4539
rect 5917 4505 5951 4539
rect 5951 4505 5960 4539
rect 5908 4496 5960 4505
rect 6000 4428 6052 4480
rect 7104 4496 7156 4548
rect 8484 4496 8536 4548
rect 6460 4428 6512 4480
rect 8116 4428 8168 4480
rect 9220 4428 9272 4480
rect 4116 4326 4168 4378
rect 4180 4326 4232 4378
rect 4244 4326 4296 4378
rect 4308 4326 4360 4378
rect 4372 4326 4424 4378
rect 7216 4326 7268 4378
rect 7280 4326 7332 4378
rect 7344 4326 7396 4378
rect 7408 4326 7460 4378
rect 7472 4326 7524 4378
rect 8024 4224 8076 4276
rect 8668 4224 8720 4276
rect 4160 4156 4212 4208
rect 8208 4156 8260 4208
rect 2964 4088 3016 4140
rect 3792 4131 3844 4140
rect 3792 4097 3801 4131
rect 3801 4097 3835 4131
rect 3835 4097 3844 4131
rect 3792 4088 3844 4097
rect 5264 4131 5316 4140
rect 5264 4097 5273 4131
rect 5273 4097 5307 4131
rect 5307 4097 5316 4131
rect 5264 4088 5316 4097
rect 6184 4131 6236 4140
rect 6184 4097 6193 4131
rect 6193 4097 6227 4131
rect 6227 4097 6236 4131
rect 6184 4088 6236 4097
rect 7656 4131 7708 4140
rect 7656 4097 7665 4131
rect 7665 4097 7699 4131
rect 7699 4097 7708 4131
rect 7656 4088 7708 4097
rect 7104 3952 7156 4004
rect 8760 4088 8812 4140
rect 9220 4088 9272 4140
rect 7932 4020 7984 4072
rect 6736 3884 6788 3936
rect 8576 3884 8628 3936
rect 8668 3884 8720 3936
rect 9496 3884 9548 3936
rect 5666 3782 5718 3834
rect 5730 3782 5782 3834
rect 5794 3782 5846 3834
rect 5858 3782 5910 3834
rect 5922 3782 5974 3834
rect 8766 3782 8818 3834
rect 8830 3782 8882 3834
rect 8894 3782 8946 3834
rect 8958 3782 9010 3834
rect 9022 3782 9074 3834
rect 2688 3680 2740 3732
rect 6000 3723 6052 3732
rect 2688 3544 2740 3596
rect 3332 3587 3384 3596
rect 3332 3553 3341 3587
rect 3341 3553 3375 3587
rect 3375 3553 3384 3587
rect 3332 3544 3384 3553
rect 3700 3544 3752 3596
rect 3976 3544 4028 3596
rect 5448 3612 5500 3664
rect 6000 3689 6009 3723
rect 6009 3689 6043 3723
rect 6043 3689 6052 3723
rect 6000 3680 6052 3689
rect 8024 3680 8076 3732
rect 8300 3680 8352 3732
rect 9312 3680 9364 3732
rect 7656 3612 7708 3664
rect 4988 3544 5040 3596
rect 7104 3544 7156 3596
rect 6460 3476 6512 3528
rect 8116 3519 8168 3528
rect 8116 3485 8125 3519
rect 8125 3485 8159 3519
rect 8159 3485 8168 3519
rect 8116 3476 8168 3485
rect 8760 3476 8812 3528
rect 9128 3519 9180 3528
rect 9128 3485 9137 3519
rect 9137 3485 9171 3519
rect 9171 3485 9180 3519
rect 9128 3476 9180 3485
rect 9404 3519 9456 3528
rect 9404 3485 9413 3519
rect 9413 3485 9447 3519
rect 9447 3485 9456 3519
rect 9404 3476 9456 3485
rect 5448 3408 5500 3460
rect 6000 3408 6052 3460
rect 7932 3408 7984 3460
rect 5080 3383 5132 3392
rect 5080 3349 5089 3383
rect 5089 3349 5123 3383
rect 5123 3349 5132 3383
rect 5080 3340 5132 3349
rect 5540 3383 5592 3392
rect 5540 3349 5549 3383
rect 5549 3349 5583 3383
rect 5583 3349 5592 3383
rect 5540 3340 5592 3349
rect 6552 3340 6604 3392
rect 8208 3340 8260 3392
rect 4116 3238 4168 3290
rect 4180 3238 4232 3290
rect 4244 3238 4296 3290
rect 4308 3238 4360 3290
rect 4372 3238 4424 3290
rect 7216 3238 7268 3290
rect 7280 3238 7332 3290
rect 7344 3238 7396 3290
rect 7408 3238 7460 3290
rect 7472 3238 7524 3290
rect 5540 3136 5592 3188
rect 2688 3068 2740 3120
rect 3884 3043 3936 3052
rect 3884 3009 3893 3043
rect 3893 3009 3927 3043
rect 3927 3009 3936 3043
rect 3884 3000 3936 3009
rect 6184 3068 6236 3120
rect 8116 3136 8168 3188
rect 8760 3179 8812 3188
rect 8760 3145 8769 3179
rect 8769 3145 8803 3179
rect 8803 3145 8812 3179
rect 8760 3136 8812 3145
rect 9680 3136 9732 3188
rect 9496 3068 9548 3120
rect 4344 3000 4396 3052
rect 5080 3043 5132 3052
rect 5080 3009 5089 3043
rect 5089 3009 5123 3043
rect 5123 3009 5132 3043
rect 5080 3000 5132 3009
rect 7380 3043 7432 3052
rect 2688 2932 2740 2984
rect 4712 2975 4764 2984
rect 3976 2864 4028 2916
rect 3700 2796 3752 2848
rect 4712 2941 4721 2975
rect 4721 2941 4755 2975
rect 4755 2941 4764 2975
rect 4712 2932 4764 2941
rect 7380 3009 7389 3043
rect 7389 3009 7423 3043
rect 7423 3009 7432 3043
rect 7380 3000 7432 3009
rect 7472 3043 7524 3052
rect 7472 3009 7481 3043
rect 7481 3009 7515 3043
rect 7515 3009 7524 3043
rect 7472 3000 7524 3009
rect 8024 3000 8076 3052
rect 8484 3000 8536 3052
rect 8392 2932 8444 2984
rect 9312 2864 9364 2916
rect 4528 2796 4580 2848
rect 4988 2796 5040 2848
rect 7472 2796 7524 2848
rect 7564 2839 7616 2848
rect 7564 2805 7573 2839
rect 7573 2805 7607 2839
rect 7607 2805 7616 2839
rect 7564 2796 7616 2805
rect 8116 2796 8168 2848
rect 8668 2796 8720 2848
rect 13820 2796 13872 2848
rect 5666 2694 5718 2746
rect 5730 2694 5782 2746
rect 5794 2694 5846 2746
rect 5858 2694 5910 2746
rect 5922 2694 5974 2746
rect 8766 2694 8818 2746
rect 8830 2694 8882 2746
rect 8894 2694 8946 2746
rect 8958 2694 9010 2746
rect 9022 2694 9074 2746
rect 5264 2592 5316 2644
rect 6184 2592 6236 2644
rect 7932 2635 7984 2644
rect 7932 2601 7941 2635
rect 7941 2601 7975 2635
rect 7975 2601 7984 2635
rect 7932 2592 7984 2601
rect 9128 2592 9180 2644
rect 9312 2635 9364 2644
rect 9312 2601 9321 2635
rect 9321 2601 9355 2635
rect 9355 2601 9364 2635
rect 9312 2592 9364 2601
rect 5172 2524 5224 2576
rect 3332 2456 3384 2508
rect 7380 2524 7432 2576
rect 6460 2456 6512 2508
rect 6552 2456 6604 2508
rect 3700 2431 3752 2440
rect 3700 2397 3709 2431
rect 3709 2397 3743 2431
rect 3743 2397 3752 2431
rect 3700 2388 3752 2397
rect 8116 2431 8168 2440
rect 8116 2397 8125 2431
rect 8125 2397 8159 2431
rect 8159 2397 8168 2431
rect 8116 2388 8168 2397
rect 8300 2431 8352 2440
rect 8300 2397 8309 2431
rect 8309 2397 8343 2431
rect 8343 2397 8352 2431
rect 8300 2388 8352 2397
rect 8392 2388 8444 2440
rect 9496 2431 9548 2440
rect 9496 2397 9505 2431
rect 9505 2397 9539 2431
rect 9539 2397 9548 2431
rect 9496 2388 9548 2397
rect 4344 2320 4396 2372
rect 4528 2320 4580 2372
rect 7564 2320 7616 2372
rect 8668 2320 8720 2372
rect 6092 2252 6144 2304
rect 4116 2150 4168 2202
rect 4180 2150 4232 2202
rect 4244 2150 4296 2202
rect 4308 2150 4360 2202
rect 4372 2150 4424 2202
rect 7216 2150 7268 2202
rect 7280 2150 7332 2202
rect 7344 2150 7396 2202
rect 7408 2150 7460 2202
rect 7472 2150 7524 2202
<< metal2 >>
rect 16578 13832 16634 13841
rect 16578 13767 16634 13776
rect 2410 13424 2466 13433
rect 2410 13359 2466 13368
rect 2318 12472 2374 12481
rect 2318 12407 2374 12416
rect 1216 11824 1268 11830
rect 1216 11766 1268 11772
rect 1032 9580 1084 9586
rect 1032 9522 1084 9528
rect 1044 7818 1072 9522
rect 1124 9512 1176 9518
rect 1124 9454 1176 9460
rect 1032 7812 1084 7818
rect 1032 7754 1084 7760
rect 1136 7750 1164 9454
rect 1228 8566 1256 11766
rect 1860 11620 1912 11626
rect 1860 11562 1912 11568
rect 1308 11552 1360 11558
rect 1308 11494 1360 11500
rect 1320 11354 1348 11494
rect 1872 11354 1900 11562
rect 1308 11348 1360 11354
rect 1308 11290 1360 11296
rect 1860 11348 1912 11354
rect 1860 11290 1912 11296
rect 1872 11150 1900 11290
rect 1860 11144 1912 11150
rect 1860 11086 1912 11092
rect 2226 10840 2282 10849
rect 2226 10775 2282 10784
rect 1490 10568 1546 10577
rect 1490 10503 1492 10512
rect 1544 10503 1546 10512
rect 1492 10474 1544 10480
rect 2136 10464 2188 10470
rect 2136 10406 2188 10412
rect 2148 10130 2176 10406
rect 2136 10124 2188 10130
rect 2136 10066 2188 10072
rect 2136 9988 2188 9994
rect 2136 9930 2188 9936
rect 1674 9616 1730 9625
rect 1674 9551 1730 9560
rect 1400 9376 1452 9382
rect 1400 9318 1452 9324
rect 1584 9376 1636 9382
rect 1584 9318 1636 9324
rect 1306 8800 1362 8809
rect 1306 8735 1362 8744
rect 1216 8560 1268 8566
rect 1216 8502 1268 8508
rect 1216 8288 1268 8294
rect 1216 8230 1268 8236
rect 1124 7744 1176 7750
rect 1124 7686 1176 7692
rect 1136 1465 1164 7686
rect 1228 6089 1256 8230
rect 1320 6633 1348 8735
rect 1412 7290 1440 9318
rect 1492 8628 1544 8634
rect 1492 8570 1544 8576
rect 1504 8537 1532 8570
rect 1490 8528 1546 8537
rect 1490 8463 1546 8472
rect 1412 7262 1532 7290
rect 1400 7200 1452 7206
rect 1400 7142 1452 7148
rect 1412 6905 1440 7142
rect 1398 6896 1454 6905
rect 1398 6831 1454 6840
rect 1400 6656 1452 6662
rect 1306 6624 1362 6633
rect 1400 6598 1452 6604
rect 1306 6559 1362 6568
rect 1214 6080 1270 6089
rect 1214 6015 1270 6024
rect 1412 5642 1440 6598
rect 1504 5982 1532 7262
rect 1596 6746 1624 9318
rect 1688 8974 1716 9551
rect 1858 9480 1914 9489
rect 1858 9415 1914 9424
rect 1952 9444 2004 9450
rect 1768 9376 1820 9382
rect 1768 9318 1820 9324
rect 1676 8968 1728 8974
rect 1676 8910 1728 8916
rect 1780 8480 1808 9318
rect 1872 9110 1900 9415
rect 1952 9386 2004 9392
rect 1860 9104 1912 9110
rect 1860 9046 1912 9052
rect 1860 8628 1912 8634
rect 1860 8570 1912 8576
rect 1688 8452 1808 8480
rect 1688 7585 1716 8452
rect 1766 8392 1822 8401
rect 1766 8327 1768 8336
rect 1820 8327 1822 8336
rect 1768 8298 1820 8304
rect 1768 7880 1820 7886
rect 1768 7822 1820 7828
rect 1674 7576 1730 7585
rect 1674 7511 1730 7520
rect 1688 6866 1716 7511
rect 1780 7478 1808 7822
rect 1768 7472 1820 7478
rect 1768 7414 1820 7420
rect 1676 6860 1728 6866
rect 1676 6802 1728 6808
rect 1768 6792 1820 6798
rect 1596 6718 1716 6746
rect 1768 6734 1820 6740
rect 1584 6656 1636 6662
rect 1584 6598 1636 6604
rect 1596 6458 1624 6598
rect 1584 6452 1636 6458
rect 1584 6394 1636 6400
rect 1492 5976 1544 5982
rect 1492 5918 1544 5924
rect 1688 5846 1716 6718
rect 1780 6254 1808 6734
rect 1768 6248 1820 6254
rect 1768 6190 1820 6196
rect 1872 5914 1900 8570
rect 1860 5908 1912 5914
rect 1860 5850 1912 5856
rect 1676 5840 1728 5846
rect 1676 5782 1728 5788
rect 1400 5636 1452 5642
rect 1400 5578 1452 5584
rect 1964 5522 1992 9386
rect 2044 9104 2096 9110
rect 2042 9072 2044 9081
rect 2096 9072 2098 9081
rect 2042 9007 2098 9016
rect 2148 8922 2176 9930
rect 2240 8974 2268 10775
rect 2332 10674 2360 12407
rect 2424 11150 2452 13359
rect 6090 13152 6146 13161
rect 6090 13087 6146 13096
rect 5998 12200 6054 12209
rect 5998 12135 6054 12144
rect 3146 11928 3202 11937
rect 3146 11863 3202 11872
rect 2566 11452 2874 11472
rect 2566 11450 2572 11452
rect 2628 11450 2652 11452
rect 2708 11450 2732 11452
rect 2788 11450 2812 11452
rect 2868 11450 2874 11452
rect 2628 11398 2630 11450
rect 2810 11398 2812 11450
rect 2566 11396 2572 11398
rect 2628 11396 2652 11398
rect 2708 11396 2732 11398
rect 2788 11396 2812 11398
rect 2868 11396 2874 11398
rect 2566 11376 2874 11396
rect 2962 11384 3018 11393
rect 2962 11319 3018 11328
rect 2412 11144 2464 11150
rect 2412 11086 2464 11092
rect 2412 11008 2464 11014
rect 2412 10950 2464 10956
rect 2320 10668 2372 10674
rect 2320 10610 2372 10616
rect 2424 10538 2452 10950
rect 2412 10532 2464 10538
rect 2412 10474 2464 10480
rect 2566 10364 2874 10384
rect 2566 10362 2572 10364
rect 2628 10362 2652 10364
rect 2708 10362 2732 10364
rect 2788 10362 2812 10364
rect 2868 10362 2874 10364
rect 2628 10310 2630 10362
rect 2810 10310 2812 10362
rect 2566 10308 2572 10310
rect 2628 10308 2652 10310
rect 2708 10308 2732 10310
rect 2788 10308 2812 10310
rect 2868 10308 2874 10310
rect 2566 10288 2874 10308
rect 2412 10192 2464 10198
rect 2318 10160 2374 10169
rect 2412 10134 2464 10140
rect 2318 10095 2374 10104
rect 2332 9178 2360 10095
rect 2424 9586 2452 10134
rect 2976 10062 3004 11319
rect 3056 11280 3108 11286
rect 3056 11222 3108 11228
rect 3068 11121 3096 11222
rect 3160 11150 3188 11863
rect 4988 11824 5040 11830
rect 4988 11766 5040 11772
rect 3424 11756 3476 11762
rect 3424 11698 3476 11704
rect 3240 11688 3292 11694
rect 3240 11630 3292 11636
rect 3148 11144 3200 11150
rect 3054 11112 3110 11121
rect 3148 11086 3200 11092
rect 3054 11047 3110 11056
rect 3056 10464 3108 10470
rect 3056 10406 3108 10412
rect 2964 10056 3016 10062
rect 2964 9998 3016 10004
rect 2964 9920 3016 9926
rect 2778 9888 2834 9897
rect 2964 9862 3016 9868
rect 2778 9823 2834 9832
rect 2792 9654 2820 9823
rect 2976 9722 3004 9862
rect 2964 9716 3016 9722
rect 2964 9658 3016 9664
rect 2780 9648 2832 9654
rect 2780 9590 2832 9596
rect 2412 9580 2464 9586
rect 2412 9522 2464 9528
rect 3068 9518 3096 10406
rect 3252 10062 3280 11630
rect 3436 11150 3464 11698
rect 3514 11248 3570 11257
rect 3514 11183 3570 11192
rect 4342 11248 4398 11257
rect 4342 11183 4398 11192
rect 4710 11248 4766 11257
rect 4710 11183 4766 11192
rect 3424 11144 3476 11150
rect 3424 11086 3476 11092
rect 3424 10736 3476 10742
rect 3330 10704 3386 10713
rect 3528 10724 3556 11183
rect 3608 11144 3660 11150
rect 3608 11086 3660 11092
rect 3476 10696 3556 10724
rect 3424 10678 3476 10684
rect 3330 10639 3386 10648
rect 3240 10056 3292 10062
rect 3240 9998 3292 10004
rect 3252 9874 3280 9998
rect 3160 9846 3280 9874
rect 3056 9512 3108 9518
rect 3056 9454 3108 9460
rect 2688 9444 2740 9450
rect 2740 9404 3004 9432
rect 2688 9386 2740 9392
rect 2566 9276 2874 9296
rect 2566 9274 2572 9276
rect 2628 9274 2652 9276
rect 2708 9274 2732 9276
rect 2788 9274 2812 9276
rect 2868 9274 2874 9276
rect 2628 9222 2630 9274
rect 2810 9222 2812 9274
rect 2566 9220 2572 9222
rect 2628 9220 2652 9222
rect 2708 9220 2732 9222
rect 2788 9220 2812 9222
rect 2868 9220 2874 9222
rect 2566 9200 2874 9220
rect 2976 9217 3004 9404
rect 2962 9208 3018 9217
rect 2320 9172 2372 9178
rect 2962 9143 3018 9152
rect 2320 9114 2372 9120
rect 2332 9042 2360 9114
rect 2320 9036 2372 9042
rect 2320 8978 2372 8984
rect 2056 8894 2176 8922
rect 2228 8968 2280 8974
rect 2228 8910 2280 8916
rect 2410 8936 2466 8945
rect 2056 8634 2084 8894
rect 3068 8906 3096 9454
rect 3160 8974 3188 9846
rect 3240 9716 3292 9722
rect 3240 9658 3292 9664
rect 3148 8968 3200 8974
rect 3148 8910 3200 8916
rect 2410 8871 2466 8880
rect 3056 8900 3108 8906
rect 2044 8628 2096 8634
rect 2044 8570 2096 8576
rect 2228 8560 2280 8566
rect 2148 8508 2228 8514
rect 2148 8502 2280 8508
rect 2148 8486 2268 8502
rect 2320 8492 2372 8498
rect 2148 8022 2176 8486
rect 2320 8434 2372 8440
rect 2136 8016 2188 8022
rect 2332 7993 2360 8434
rect 2424 8022 2452 8871
rect 3056 8842 3108 8848
rect 2964 8832 3016 8838
rect 2964 8774 3016 8780
rect 2872 8628 2924 8634
rect 2872 8570 2924 8576
rect 2688 8424 2740 8430
rect 2688 8366 2740 8372
rect 2700 8276 2728 8366
rect 2884 8344 2912 8570
rect 2976 8498 3004 8774
rect 3068 8566 3096 8842
rect 3160 8809 3188 8910
rect 3146 8800 3202 8809
rect 3146 8735 3202 8744
rect 3056 8560 3108 8566
rect 3056 8502 3108 8508
rect 2964 8492 3016 8498
rect 2964 8434 3016 8440
rect 2884 8316 3188 8344
rect 2700 8248 3004 8276
rect 2566 8188 2874 8208
rect 2566 8186 2572 8188
rect 2628 8186 2652 8188
rect 2708 8186 2732 8188
rect 2788 8186 2812 8188
rect 2868 8186 2874 8188
rect 2628 8134 2630 8186
rect 2810 8134 2812 8186
rect 2566 8132 2572 8134
rect 2628 8132 2652 8134
rect 2708 8132 2732 8134
rect 2788 8132 2812 8134
rect 2868 8132 2874 8134
rect 2566 8112 2874 8132
rect 2412 8016 2464 8022
rect 2136 7958 2188 7964
rect 2318 7984 2374 7993
rect 2044 7880 2096 7886
rect 2148 7857 2176 7958
rect 2412 7958 2464 7964
rect 2976 7954 3004 8248
rect 3054 8256 3110 8265
rect 3054 8191 3110 8200
rect 3068 8090 3096 8191
rect 3160 8090 3188 8316
rect 3056 8084 3108 8090
rect 3056 8026 3108 8032
rect 3148 8084 3200 8090
rect 3148 8026 3200 8032
rect 2318 7919 2374 7928
rect 2964 7948 3016 7954
rect 2964 7890 3016 7896
rect 2688 7880 2740 7886
rect 2044 7822 2096 7828
rect 2134 7848 2190 7857
rect 2056 7002 2084 7822
rect 2688 7822 2740 7828
rect 2134 7783 2190 7792
rect 2228 7744 2280 7750
rect 2228 7686 2280 7692
rect 2136 7540 2188 7546
rect 2136 7482 2188 7488
rect 2044 6996 2096 7002
rect 2044 6938 2096 6944
rect 2148 6882 2176 7482
rect 2056 6854 2176 6882
rect 2056 6769 2084 6854
rect 2240 6798 2268 7686
rect 2320 7336 2372 7342
rect 2320 7278 2372 7284
rect 2136 6792 2188 6798
rect 2042 6760 2098 6769
rect 2136 6734 2188 6740
rect 2228 6792 2280 6798
rect 2228 6734 2280 6740
rect 2042 6695 2098 6704
rect 2044 6656 2096 6662
rect 2044 6598 2096 6604
rect 2056 6225 2084 6598
rect 2148 6390 2176 6734
rect 2228 6656 2280 6662
rect 2228 6598 2280 6604
rect 2240 6458 2268 6598
rect 2228 6452 2280 6458
rect 2228 6394 2280 6400
rect 2136 6384 2188 6390
rect 2136 6326 2188 6332
rect 2042 6216 2098 6225
rect 2042 6151 2098 6160
rect 2332 5817 2360 7278
rect 2412 7268 2464 7274
rect 2412 7210 2464 7216
rect 2318 5808 2374 5817
rect 2318 5743 2374 5752
rect 1964 5494 2360 5522
rect 2332 3618 2360 5494
rect 2424 5273 2452 7210
rect 2700 7188 2728 7822
rect 3148 7744 3200 7750
rect 2778 7712 2834 7721
rect 3148 7686 3200 7692
rect 2778 7647 2834 7656
rect 2792 7410 2820 7647
rect 2870 7576 2926 7585
rect 2870 7511 2926 7520
rect 3054 7576 3110 7585
rect 3054 7511 3056 7520
rect 2780 7404 2832 7410
rect 2780 7346 2832 7352
rect 2884 7313 2912 7511
rect 3108 7511 3110 7520
rect 3056 7482 3108 7488
rect 3056 7404 3108 7410
rect 3056 7346 3108 7352
rect 2870 7304 2926 7313
rect 2870 7239 2926 7248
rect 2700 7160 3004 7188
rect 2566 7100 2874 7120
rect 2566 7098 2572 7100
rect 2628 7098 2652 7100
rect 2708 7098 2732 7100
rect 2788 7098 2812 7100
rect 2868 7098 2874 7100
rect 2628 7046 2630 7098
rect 2810 7046 2812 7098
rect 2566 7044 2572 7046
rect 2628 7044 2652 7046
rect 2708 7044 2732 7046
rect 2788 7044 2812 7046
rect 2868 7044 2874 7046
rect 2566 7024 2874 7044
rect 2976 6984 3004 7160
rect 2792 6956 3004 6984
rect 2688 6656 2740 6662
rect 2688 6598 2740 6604
rect 2504 5976 2556 5982
rect 2700 5953 2728 6598
rect 2504 5918 2556 5924
rect 2686 5944 2742 5953
rect 2410 5264 2466 5273
rect 2410 5199 2466 5208
rect 2410 3632 2466 3641
rect 2332 3590 2410 3618
rect 2410 3567 2466 3576
rect 2516 2938 2544 5918
rect 2686 5879 2742 5888
rect 2596 5840 2648 5846
rect 2596 5782 2648 5788
rect 2608 3482 2636 5782
rect 2688 5636 2740 5642
rect 2688 5578 2740 5584
rect 2700 3738 2728 5578
rect 2792 5166 2820 6956
rect 2962 6760 3018 6769
rect 2962 6695 3018 6704
rect 2872 6656 2924 6662
rect 2872 6598 2924 6604
rect 2884 6390 2912 6598
rect 2872 6384 2924 6390
rect 2872 6326 2924 6332
rect 2780 5160 2832 5166
rect 2780 5102 2832 5108
rect 2780 5024 2832 5030
rect 2778 4992 2780 5001
rect 2832 4992 2834 5001
rect 2778 4927 2834 4936
rect 2780 4888 2832 4894
rect 2780 4830 2832 4836
rect 2688 3732 2740 3738
rect 2688 3674 2740 3680
rect 2686 3632 2742 3641
rect 2686 3567 2688 3576
rect 2740 3567 2742 3576
rect 2688 3538 2740 3544
rect 2608 3454 2728 3482
rect 2700 3126 2728 3454
rect 2688 3120 2740 3126
rect 2688 3062 2740 3068
rect 2688 2984 2740 2990
rect 2516 2932 2688 2938
rect 2516 2926 2740 2932
rect 2516 2910 2728 2926
rect 1122 1456 1178 1465
rect 1122 1391 1178 1400
rect 2792 1057 2820 4830
rect 2884 4049 2912 6326
rect 2976 4146 3004 6695
rect 3068 4826 3096 7346
rect 3160 6458 3188 7686
rect 3252 7546 3280 9658
rect 3344 9042 3372 10639
rect 3436 9926 3464 10678
rect 3516 10600 3568 10606
rect 3516 10542 3568 10548
rect 3528 10441 3556 10542
rect 3620 10470 3648 11086
rect 4356 11082 4384 11183
rect 3976 11076 4028 11082
rect 3976 11018 4028 11024
rect 4344 11076 4396 11082
rect 4344 11018 4396 11024
rect 3882 10840 3938 10849
rect 3882 10775 3938 10784
rect 3608 10464 3660 10470
rect 3514 10432 3570 10441
rect 3608 10406 3660 10412
rect 3700 10464 3752 10470
rect 3752 10412 3832 10418
rect 3700 10406 3832 10412
rect 3712 10390 3832 10406
rect 3514 10367 3570 10376
rect 3804 10266 3832 10390
rect 3792 10260 3844 10266
rect 3896 10248 3924 10775
rect 3988 10606 4016 11018
rect 4116 10908 4424 10928
rect 4116 10906 4122 10908
rect 4178 10906 4202 10908
rect 4258 10906 4282 10908
rect 4338 10906 4362 10908
rect 4418 10906 4424 10908
rect 4178 10854 4180 10906
rect 4360 10854 4362 10906
rect 4116 10852 4122 10854
rect 4178 10852 4202 10854
rect 4258 10852 4282 10854
rect 4338 10852 4362 10854
rect 4418 10852 4424 10854
rect 4116 10832 4424 10852
rect 3976 10600 4028 10606
rect 3976 10542 4028 10548
rect 4344 10600 4396 10606
rect 4344 10542 4396 10548
rect 4068 10260 4120 10266
rect 3896 10220 4068 10248
rect 3792 10202 3844 10208
rect 4068 10202 4120 10208
rect 3608 10192 3660 10198
rect 3606 10160 3608 10169
rect 3660 10160 3662 10169
rect 4356 10130 4384 10542
rect 3606 10095 3662 10104
rect 4344 10124 4396 10130
rect 4344 10066 4396 10072
rect 3884 10056 3936 10062
rect 3514 10024 3570 10033
rect 3884 9998 3936 10004
rect 3514 9959 3570 9968
rect 3424 9920 3476 9926
rect 3424 9862 3476 9868
rect 3528 9178 3556 9959
rect 3700 9920 3752 9926
rect 3700 9862 3752 9868
rect 3790 9888 3846 9897
rect 3712 9654 3740 9862
rect 3790 9823 3846 9832
rect 3700 9648 3752 9654
rect 3700 9590 3752 9596
rect 3804 9489 3832 9823
rect 3790 9480 3846 9489
rect 3790 9415 3846 9424
rect 3608 9376 3660 9382
rect 3608 9318 3660 9324
rect 3516 9172 3568 9178
rect 3516 9114 3568 9120
rect 3332 9036 3384 9042
rect 3332 8978 3384 8984
rect 3620 8974 3648 9318
rect 3792 9172 3844 9178
rect 3896 9160 3924 9998
rect 4620 9988 4672 9994
rect 4620 9930 4672 9936
rect 4116 9820 4424 9840
rect 4116 9818 4122 9820
rect 4178 9818 4202 9820
rect 4258 9818 4282 9820
rect 4338 9818 4362 9820
rect 4418 9818 4424 9820
rect 4178 9766 4180 9818
rect 4360 9766 4362 9818
rect 4116 9764 4122 9766
rect 4178 9764 4202 9766
rect 4258 9764 4282 9766
rect 4338 9764 4362 9766
rect 4418 9764 4424 9766
rect 4116 9744 4424 9764
rect 4526 9752 4582 9761
rect 4526 9687 4528 9696
rect 4580 9687 4582 9696
rect 4528 9658 4580 9664
rect 4436 9648 4488 9654
rect 4436 9590 4488 9596
rect 4344 9580 4396 9586
rect 4264 9540 4344 9568
rect 4068 9512 4120 9518
rect 4068 9454 4120 9460
rect 3844 9132 3924 9160
rect 3792 9114 3844 9120
rect 4080 9058 4108 9454
rect 4160 9444 4212 9450
rect 4160 9386 4212 9392
rect 3896 9030 4108 9058
rect 3608 8968 3660 8974
rect 3608 8910 3660 8916
rect 3698 8936 3754 8945
rect 3332 8900 3384 8906
rect 3896 8922 3924 9030
rect 3754 8894 3924 8922
rect 4068 8968 4120 8974
rect 4172 8956 4200 9386
rect 4120 8928 4200 8956
rect 4068 8910 4120 8916
rect 4264 8906 4292 9540
rect 4344 9522 4396 9528
rect 4344 9376 4396 9382
rect 4448 9364 4476 9590
rect 4396 9336 4476 9364
rect 4528 9376 4580 9382
rect 4344 9318 4396 9324
rect 4528 9318 4580 9324
rect 4252 8900 4304 8906
rect 3698 8871 3754 8880
rect 3332 8842 3384 8848
rect 4252 8842 4304 8848
rect 3344 8616 3372 8842
rect 3700 8832 3752 8838
rect 3884 8832 3936 8838
rect 3700 8774 3752 8780
rect 3882 8800 3884 8809
rect 3976 8832 4028 8838
rect 3936 8800 3938 8809
rect 3344 8588 3464 8616
rect 3436 8464 3464 8588
rect 3344 8436 3464 8464
rect 3240 7540 3292 7546
rect 3240 7482 3292 7488
rect 3240 7200 3292 7206
rect 3240 7142 3292 7148
rect 3148 6452 3200 6458
rect 3148 6394 3200 6400
rect 3148 6248 3200 6254
rect 3148 6190 3200 6196
rect 3056 4820 3108 4826
rect 3056 4762 3108 4768
rect 2964 4140 3016 4146
rect 2964 4082 3016 4088
rect 2870 4040 2926 4049
rect 2870 3975 2926 3984
rect 3160 2009 3188 6190
rect 3252 5234 3280 7142
rect 3344 6769 3372 8436
rect 3712 8242 3740 8774
rect 3976 8774 4028 8780
rect 3882 8735 3938 8744
rect 3884 8424 3936 8430
rect 3884 8366 3936 8372
rect 3712 8214 3832 8242
rect 3698 8120 3754 8129
rect 3698 8055 3754 8064
rect 3712 8022 3740 8055
rect 3700 8016 3752 8022
rect 3606 7984 3662 7993
rect 3700 7958 3752 7964
rect 3606 7919 3662 7928
rect 3424 7744 3476 7750
rect 3424 7686 3476 7692
rect 3516 7744 3568 7750
rect 3516 7686 3568 7692
rect 3436 7177 3464 7686
rect 3528 7342 3556 7686
rect 3620 7562 3648 7919
rect 3804 7886 3832 8214
rect 3792 7880 3844 7886
rect 3792 7822 3844 7828
rect 3804 7721 3832 7822
rect 3790 7712 3846 7721
rect 3790 7647 3846 7656
rect 3620 7534 3740 7562
rect 3516 7336 3568 7342
rect 3516 7278 3568 7284
rect 3608 7268 3660 7274
rect 3608 7210 3660 7216
rect 3422 7168 3478 7177
rect 3422 7103 3478 7112
rect 3516 6928 3568 6934
rect 3516 6870 3568 6876
rect 3330 6760 3386 6769
rect 3330 6695 3386 6704
rect 3344 6322 3372 6695
rect 3528 6662 3556 6870
rect 3516 6656 3568 6662
rect 3516 6598 3568 6604
rect 3424 6452 3476 6458
rect 3424 6394 3476 6400
rect 3332 6316 3384 6322
rect 3332 6258 3384 6264
rect 3332 5704 3384 5710
rect 3332 5646 3384 5652
rect 3240 5228 3292 5234
rect 3240 5170 3292 5176
rect 3240 5092 3292 5098
rect 3240 5034 3292 5040
rect 3252 2961 3280 5034
rect 3344 3602 3372 5646
rect 3332 3596 3384 3602
rect 3332 3538 3384 3544
rect 3238 2952 3294 2961
rect 3238 2887 3294 2896
rect 3344 2514 3372 3538
rect 3332 2508 3384 2514
rect 3332 2450 3384 2456
rect 3146 2000 3202 2009
rect 3146 1935 3202 1944
rect 3436 1737 3464 6394
rect 3422 1728 3478 1737
rect 3422 1663 3478 1672
rect 2778 1048 2834 1057
rect 2778 983 2834 992
rect 3528 513 3556 6598
rect 3620 6361 3648 7210
rect 3712 6934 3740 7534
rect 3804 7392 3832 7647
rect 3896 7528 3924 8366
rect 3988 7993 4016 8774
rect 4116 8732 4424 8752
rect 4116 8730 4122 8732
rect 4178 8730 4202 8732
rect 4258 8730 4282 8732
rect 4338 8730 4362 8732
rect 4418 8730 4424 8732
rect 4178 8678 4180 8730
rect 4360 8678 4362 8730
rect 4116 8676 4122 8678
rect 4178 8676 4202 8678
rect 4258 8676 4282 8678
rect 4338 8676 4362 8678
rect 4418 8676 4424 8678
rect 4116 8656 4424 8676
rect 4540 8430 4568 9318
rect 4632 9178 4660 9930
rect 4724 9382 4752 11183
rect 4804 10668 4856 10674
rect 4804 10610 4856 10616
rect 4816 9722 4844 10610
rect 4894 10296 4950 10305
rect 4894 10231 4950 10240
rect 4804 9716 4856 9722
rect 4804 9658 4856 9664
rect 4908 9602 4936 10231
rect 4816 9574 4936 9602
rect 4712 9376 4764 9382
rect 4712 9318 4764 9324
rect 4620 9172 4672 9178
rect 4620 9114 4672 9120
rect 4724 8922 4752 9318
rect 4816 9178 4844 9574
rect 4804 9172 4856 9178
rect 4804 9114 4856 9120
rect 4896 8968 4948 8974
rect 4724 8894 4844 8922
rect 4896 8910 4948 8916
rect 4712 8832 4764 8838
rect 4618 8800 4674 8809
rect 4712 8774 4764 8780
rect 4618 8735 4674 8744
rect 4528 8424 4580 8430
rect 4528 8366 4580 8372
rect 4436 8356 4488 8362
rect 4436 8298 4488 8304
rect 4448 8022 4476 8298
rect 4528 8288 4580 8294
rect 4528 8230 4580 8236
rect 4436 8016 4488 8022
rect 3974 7984 4030 7993
rect 4436 7958 4488 7964
rect 4540 7954 4568 8230
rect 3974 7919 4030 7928
rect 4528 7948 4580 7954
rect 4528 7890 4580 7896
rect 4528 7744 4580 7750
rect 4528 7686 4580 7692
rect 4116 7644 4424 7664
rect 4116 7642 4122 7644
rect 4178 7642 4202 7644
rect 4258 7642 4282 7644
rect 4338 7642 4362 7644
rect 4418 7642 4424 7644
rect 4178 7590 4180 7642
rect 4360 7590 4362 7642
rect 4116 7588 4122 7590
rect 4178 7588 4202 7590
rect 4258 7588 4282 7590
rect 4338 7588 4362 7590
rect 4418 7588 4424 7590
rect 4116 7568 4424 7588
rect 3896 7500 4108 7528
rect 4080 7410 4108 7500
rect 4344 7472 4396 7478
rect 4344 7414 4396 7420
rect 4068 7404 4120 7410
rect 3804 7364 3924 7392
rect 3896 7041 3924 7364
rect 4068 7346 4120 7352
rect 4356 7154 4384 7414
rect 4540 7342 4568 7686
rect 4528 7336 4580 7342
rect 4528 7278 4580 7284
rect 3988 7126 4384 7154
rect 3882 7032 3938 7041
rect 3882 6967 3938 6976
rect 3700 6928 3752 6934
rect 3988 6916 4016 7126
rect 4526 7032 4582 7041
rect 4252 6996 4304 7002
rect 4526 6967 4582 6976
rect 4252 6938 4304 6944
rect 3700 6870 3752 6876
rect 3804 6888 4016 6916
rect 3700 6656 3752 6662
rect 3700 6598 3752 6604
rect 3606 6352 3662 6361
rect 3606 6287 3662 6296
rect 3712 6254 3740 6598
rect 3700 6248 3752 6254
rect 3700 6190 3752 6196
rect 3608 6112 3660 6118
rect 3608 6054 3660 6060
rect 3620 5642 3648 6054
rect 3804 5658 3832 6888
rect 4264 6866 4292 6938
rect 4252 6860 4304 6866
rect 4252 6802 4304 6808
rect 4540 6798 4568 6967
rect 3884 6792 3936 6798
rect 3884 6734 3936 6740
rect 4528 6792 4580 6798
rect 4528 6734 4580 6740
rect 3896 6633 3924 6734
rect 3882 6624 3938 6633
rect 3882 6559 3938 6568
rect 3896 6100 3924 6559
rect 4116 6556 4424 6576
rect 4116 6554 4122 6556
rect 4178 6554 4202 6556
rect 4258 6554 4282 6556
rect 4338 6554 4362 6556
rect 4418 6554 4424 6556
rect 4178 6502 4180 6554
rect 4360 6502 4362 6554
rect 4116 6500 4122 6502
rect 4178 6500 4202 6502
rect 4258 6500 4282 6502
rect 4338 6500 4362 6502
rect 4418 6500 4424 6502
rect 4116 6480 4424 6500
rect 3896 6072 4016 6100
rect 3608 5636 3660 5642
rect 3804 5630 3924 5658
rect 3608 5578 3660 5584
rect 3620 5234 3648 5578
rect 3792 5568 3844 5574
rect 3792 5510 3844 5516
rect 3608 5228 3660 5234
rect 3608 5170 3660 5176
rect 3804 4146 3832 5510
rect 3896 5284 3924 5630
rect 3988 5352 4016 6072
rect 4116 5468 4424 5488
rect 4116 5466 4122 5468
rect 4178 5466 4202 5468
rect 4258 5466 4282 5468
rect 4338 5466 4362 5468
rect 4418 5466 4424 5468
rect 4178 5414 4180 5466
rect 4360 5414 4362 5466
rect 4116 5412 4122 5414
rect 4178 5412 4202 5414
rect 4258 5412 4282 5414
rect 4338 5412 4362 5414
rect 4418 5412 4424 5414
rect 4116 5392 4424 5412
rect 4540 5352 4568 6734
rect 3988 5324 4292 5352
rect 3896 5256 4200 5284
rect 4172 4622 4200 5256
rect 4160 4616 4212 4622
rect 4158 4584 4160 4593
rect 4264 4604 4292 5324
rect 4356 5324 4568 5352
rect 4356 4826 4384 5324
rect 4632 4826 4660 8735
rect 4724 5302 4752 8774
rect 4816 8566 4844 8894
rect 4908 8809 4936 8910
rect 4894 8800 4950 8809
rect 4894 8735 4950 8744
rect 4896 8628 4948 8634
rect 4896 8570 4948 8576
rect 4804 8560 4856 8566
rect 4804 8502 4856 8508
rect 4908 8129 4936 8570
rect 4894 8120 4950 8129
rect 4894 8055 4950 8064
rect 4896 8016 4948 8022
rect 4802 7984 4858 7993
rect 4896 7958 4948 7964
rect 4802 7919 4858 7928
rect 4712 5296 4764 5302
rect 4712 5238 4764 5244
rect 4816 5234 4844 7919
rect 4908 7546 4936 7958
rect 5000 7721 5028 11766
rect 5080 11688 5132 11694
rect 5080 11630 5132 11636
rect 5092 10674 5120 11630
rect 5666 11452 5974 11472
rect 5666 11450 5672 11452
rect 5728 11450 5752 11452
rect 5808 11450 5832 11452
rect 5888 11450 5912 11452
rect 5968 11450 5974 11452
rect 5728 11398 5730 11450
rect 5910 11398 5912 11450
rect 5666 11396 5672 11398
rect 5728 11396 5752 11398
rect 5808 11396 5832 11398
rect 5888 11396 5912 11398
rect 5968 11396 5974 11398
rect 5666 11376 5974 11396
rect 6012 11286 6040 12135
rect 6000 11280 6052 11286
rect 6000 11222 6052 11228
rect 5264 11144 5316 11150
rect 5264 11086 5316 11092
rect 5080 10668 5132 10674
rect 5080 10610 5132 10616
rect 5276 10538 5304 11086
rect 5540 10668 5592 10674
rect 5540 10610 5592 10616
rect 5264 10532 5316 10538
rect 5264 10474 5316 10480
rect 5080 10464 5132 10470
rect 5356 10464 5408 10470
rect 5080 10406 5132 10412
rect 5262 10432 5318 10441
rect 5092 9738 5120 10406
rect 5356 10406 5408 10412
rect 5262 10367 5318 10376
rect 5276 10198 5304 10367
rect 5264 10192 5316 10198
rect 5264 10134 5316 10140
rect 5368 10062 5396 10406
rect 5356 10056 5408 10062
rect 5356 9998 5408 10004
rect 5552 10010 5580 10610
rect 6000 10600 6052 10606
rect 6000 10542 6052 10548
rect 5666 10364 5974 10384
rect 5666 10362 5672 10364
rect 5728 10362 5752 10364
rect 5808 10362 5832 10364
rect 5888 10362 5912 10364
rect 5968 10362 5974 10364
rect 5728 10310 5730 10362
rect 5910 10310 5912 10362
rect 5666 10308 5672 10310
rect 5728 10308 5752 10310
rect 5808 10308 5832 10310
rect 5888 10308 5912 10310
rect 5968 10308 5974 10310
rect 5666 10288 5974 10308
rect 5552 9982 5948 10010
rect 5632 9920 5684 9926
rect 5632 9862 5684 9868
rect 5092 9710 5212 9738
rect 5644 9722 5672 9862
rect 5080 9580 5132 9586
rect 5080 9522 5132 9528
rect 5092 8634 5120 9522
rect 5184 9042 5212 9710
rect 5632 9716 5684 9722
rect 5632 9658 5684 9664
rect 5816 9580 5868 9586
rect 5816 9522 5868 9528
rect 5828 9450 5856 9522
rect 5816 9444 5868 9450
rect 5816 9386 5868 9392
rect 5920 9364 5948 9982
rect 6012 9586 6040 10542
rect 6104 10538 6132 13087
rect 7656 11756 7708 11762
rect 7656 11698 7708 11704
rect 6276 11688 6328 11694
rect 6276 11630 6328 11636
rect 6288 11286 6316 11630
rect 6460 11348 6512 11354
rect 6460 11290 6512 11296
rect 6276 11280 6328 11286
rect 6182 11248 6238 11257
rect 6276 11222 6328 11228
rect 6182 11183 6238 11192
rect 6196 11150 6224 11183
rect 6184 11144 6236 11150
rect 6184 11086 6236 11092
rect 6184 11008 6236 11014
rect 6184 10950 6236 10956
rect 6368 11008 6420 11014
rect 6368 10950 6420 10956
rect 6092 10532 6144 10538
rect 6092 10474 6144 10480
rect 6092 10192 6144 10198
rect 6092 10134 6144 10140
rect 6000 9580 6052 9586
rect 6000 9522 6052 9528
rect 5446 9344 5502 9353
rect 5920 9336 6040 9364
rect 5446 9279 5502 9288
rect 5262 9208 5318 9217
rect 5262 9143 5318 9152
rect 5172 9036 5224 9042
rect 5172 8978 5224 8984
rect 5172 8900 5224 8906
rect 5172 8842 5224 8848
rect 5080 8628 5132 8634
rect 5080 8570 5132 8576
rect 5184 8548 5212 8842
rect 5276 8673 5304 9143
rect 5460 8882 5488 9279
rect 5666 9276 5974 9296
rect 5666 9274 5672 9276
rect 5728 9274 5752 9276
rect 5808 9274 5832 9276
rect 5888 9274 5912 9276
rect 5968 9274 5974 9276
rect 5728 9222 5730 9274
rect 5910 9222 5912 9274
rect 5666 9220 5672 9222
rect 5728 9220 5752 9222
rect 5808 9220 5832 9222
rect 5888 9220 5912 9222
rect 5968 9220 5974 9222
rect 5666 9200 5974 9220
rect 5632 8968 5684 8974
rect 5684 8928 5764 8956
rect 5632 8910 5684 8916
rect 5460 8854 5672 8882
rect 5644 8809 5672 8854
rect 5630 8800 5686 8809
rect 5630 8735 5686 8744
rect 5262 8664 5318 8673
rect 5262 8599 5318 8608
rect 5356 8628 5408 8634
rect 5356 8570 5408 8576
rect 5184 8520 5304 8548
rect 5080 8476 5132 8482
rect 5080 8418 5132 8424
rect 4986 7712 5042 7721
rect 4986 7647 5042 7656
rect 4896 7540 4948 7546
rect 4896 7482 4948 7488
rect 4988 7540 5040 7546
rect 4988 7482 5040 7488
rect 5000 7041 5028 7482
rect 5092 7274 5120 8418
rect 5172 8288 5224 8294
rect 5172 8230 5224 8236
rect 5184 7886 5212 8230
rect 5172 7880 5224 7886
rect 5172 7822 5224 7828
rect 5080 7268 5132 7274
rect 5080 7210 5132 7216
rect 4986 7032 5042 7041
rect 4986 6967 5042 6976
rect 5080 6996 5132 7002
rect 5080 6938 5132 6944
rect 4988 6860 5040 6866
rect 4988 6802 5040 6808
rect 5000 5642 5028 6802
rect 5092 6390 5120 6938
rect 5184 6458 5212 7822
rect 5276 7585 5304 8520
rect 5262 7576 5318 7585
rect 5262 7511 5318 7520
rect 5368 7392 5396 8570
rect 5538 8392 5594 8401
rect 5736 8362 5764 8928
rect 5906 8936 5962 8945
rect 5906 8871 5908 8880
rect 5960 8871 5962 8880
rect 5908 8842 5960 8848
rect 5816 8832 5868 8838
rect 5816 8774 5868 8780
rect 5538 8327 5594 8336
rect 5724 8356 5776 8362
rect 5448 8288 5500 8294
rect 5446 8256 5448 8265
rect 5500 8256 5502 8265
rect 5446 8191 5502 8200
rect 5448 7948 5500 7954
rect 5448 7890 5500 7896
rect 5276 7364 5396 7392
rect 5276 6769 5304 7364
rect 5356 7268 5408 7274
rect 5356 7210 5408 7216
rect 5368 6866 5396 7210
rect 5356 6860 5408 6866
rect 5356 6802 5408 6808
rect 5262 6760 5318 6769
rect 5262 6695 5318 6704
rect 5460 6662 5488 7890
rect 5552 7818 5580 8327
rect 5724 8298 5776 8304
rect 5828 8276 5856 8774
rect 6012 8566 6040 9336
rect 6000 8560 6052 8566
rect 6000 8502 6052 8508
rect 5828 8248 6040 8276
rect 5666 8188 5974 8208
rect 5666 8186 5672 8188
rect 5728 8186 5752 8188
rect 5808 8186 5832 8188
rect 5888 8186 5912 8188
rect 5968 8186 5974 8188
rect 5728 8134 5730 8186
rect 5910 8134 5912 8186
rect 5666 8132 5672 8134
rect 5728 8132 5752 8134
rect 5808 8132 5832 8134
rect 5888 8132 5912 8134
rect 5968 8132 5974 8134
rect 5666 8112 5974 8132
rect 5906 7984 5962 7993
rect 5906 7919 5962 7928
rect 5540 7812 5592 7818
rect 5540 7754 5592 7760
rect 5920 7546 5948 7919
rect 5908 7540 5960 7546
rect 5908 7482 5960 7488
rect 6012 7410 6040 8248
rect 6000 7404 6052 7410
rect 6000 7346 6052 7352
rect 5632 7268 5684 7274
rect 5552 7228 5632 7256
rect 5264 6656 5316 6662
rect 5448 6656 5500 6662
rect 5264 6598 5316 6604
rect 5354 6624 5410 6633
rect 5276 6458 5304 6598
rect 5448 6598 5500 6604
rect 5354 6559 5410 6568
rect 5172 6452 5224 6458
rect 5172 6394 5224 6400
rect 5264 6452 5316 6458
rect 5264 6394 5316 6400
rect 5080 6384 5132 6390
rect 5080 6326 5132 6332
rect 5092 5846 5120 6326
rect 5172 6248 5224 6254
rect 5172 6190 5224 6196
rect 5080 5840 5132 5846
rect 5080 5782 5132 5788
rect 5080 5704 5132 5710
rect 5080 5646 5132 5652
rect 4988 5636 5040 5642
rect 4988 5578 5040 5584
rect 5092 5522 5120 5646
rect 5000 5494 5120 5522
rect 4804 5228 4856 5234
rect 4804 5170 4856 5176
rect 4344 4820 4396 4826
rect 4344 4762 4396 4768
rect 4436 4820 4488 4826
rect 4436 4762 4488 4768
rect 4620 4820 4672 4826
rect 4620 4762 4672 4768
rect 4448 4729 4476 4762
rect 4434 4720 4490 4729
rect 4434 4655 4490 4664
rect 5000 4622 5028 5494
rect 5080 5364 5132 5370
rect 5080 5306 5132 5312
rect 4344 4616 4396 4622
rect 4212 4584 4214 4593
rect 4264 4576 4344 4604
rect 4344 4558 4396 4564
rect 4988 4616 5040 4622
rect 4988 4558 5040 4564
rect 4158 4519 4214 4528
rect 4712 4480 4764 4486
rect 4712 4422 4764 4428
rect 4116 4380 4424 4400
rect 4116 4378 4122 4380
rect 4178 4378 4202 4380
rect 4258 4378 4282 4380
rect 4338 4378 4362 4380
rect 4418 4378 4424 4380
rect 4178 4326 4180 4378
rect 4360 4326 4362 4378
rect 4116 4324 4122 4326
rect 4178 4324 4202 4326
rect 4258 4324 4282 4326
rect 4338 4324 4362 4326
rect 4418 4324 4424 4326
rect 4116 4304 4424 4324
rect 4160 4208 4212 4214
rect 4160 4150 4212 4156
rect 3792 4140 3844 4146
rect 3792 4082 3844 4088
rect 3700 3596 3752 3602
rect 3804 3584 3832 4082
rect 3976 3596 4028 3602
rect 3752 3556 3832 3584
rect 3896 3556 3976 3584
rect 3700 3538 3752 3544
rect 3896 3058 3924 3556
rect 3976 3538 4028 3544
rect 4172 3482 4200 4150
rect 3988 3454 4200 3482
rect 3884 3052 3936 3058
rect 3884 2994 3936 3000
rect 3988 2922 4016 3454
rect 4116 3292 4424 3312
rect 4116 3290 4122 3292
rect 4178 3290 4202 3292
rect 4258 3290 4282 3292
rect 4338 3290 4362 3292
rect 4418 3290 4424 3292
rect 4178 3238 4180 3290
rect 4360 3238 4362 3290
rect 4116 3236 4122 3238
rect 4178 3236 4202 3238
rect 4258 3236 4282 3238
rect 4338 3236 4362 3238
rect 4418 3236 4424 3238
rect 4116 3216 4424 3236
rect 4344 3052 4396 3058
rect 4344 2994 4396 3000
rect 3976 2916 4028 2922
rect 3976 2858 4028 2864
rect 3700 2848 3752 2854
rect 3700 2790 3752 2796
rect 3712 2446 3740 2790
rect 3700 2440 3752 2446
rect 3700 2382 3752 2388
rect 4356 2378 4384 2994
rect 4724 2990 4752 4422
rect 5000 3602 5028 4558
rect 4988 3596 5040 3602
rect 4988 3538 5040 3544
rect 5092 3482 5120 5306
rect 5184 4622 5212 6190
rect 5368 5658 5396 6559
rect 5460 5710 5488 6598
rect 5552 6390 5580 7228
rect 5632 7210 5684 7216
rect 5666 7100 5974 7120
rect 5666 7098 5672 7100
rect 5728 7098 5752 7100
rect 5808 7098 5832 7100
rect 5888 7098 5912 7100
rect 5968 7098 5974 7100
rect 5728 7046 5730 7098
rect 5910 7046 5912 7098
rect 5666 7044 5672 7046
rect 5728 7044 5752 7046
rect 5808 7044 5832 7046
rect 5888 7044 5912 7046
rect 5968 7044 5974 7046
rect 5666 7024 5974 7044
rect 5816 6860 5868 6866
rect 5816 6802 5868 6808
rect 5632 6724 5684 6730
rect 5632 6666 5684 6672
rect 5644 6497 5672 6666
rect 5630 6488 5686 6497
rect 5630 6423 5686 6432
rect 5540 6384 5592 6390
rect 5540 6326 5592 6332
rect 5828 6236 5856 6802
rect 5908 6656 5960 6662
rect 5908 6598 5960 6604
rect 5552 6208 5856 6236
rect 5552 6089 5580 6208
rect 5920 6100 5948 6598
rect 6104 6202 6132 10134
rect 6196 9994 6224 10950
rect 6276 10600 6328 10606
rect 6276 10542 6328 10548
rect 6184 9988 6236 9994
rect 6184 9930 6236 9936
rect 6196 9042 6224 9930
rect 6184 9036 6236 9042
rect 6184 8978 6236 8984
rect 6288 8838 6316 10542
rect 6380 10198 6408 10950
rect 6472 10606 6500 11290
rect 7104 11212 7156 11218
rect 7104 11154 7156 11160
rect 6828 11144 6880 11150
rect 6828 11086 6880 11092
rect 6552 10668 6604 10674
rect 6552 10610 6604 10616
rect 6460 10600 6512 10606
rect 6460 10542 6512 10548
rect 6564 10470 6592 10610
rect 6460 10464 6512 10470
rect 6460 10406 6512 10412
rect 6552 10464 6604 10470
rect 6552 10406 6604 10412
rect 6368 10192 6420 10198
rect 6368 10134 6420 10140
rect 6368 10056 6420 10062
rect 6368 9998 6420 10004
rect 6380 9738 6408 9998
rect 6472 9926 6500 10406
rect 6460 9920 6512 9926
rect 6460 9862 6512 9868
rect 6564 9738 6592 10406
rect 6734 10160 6790 10169
rect 6734 10095 6736 10104
rect 6788 10095 6790 10104
rect 6736 10066 6788 10072
rect 6736 9988 6788 9994
rect 6380 9710 6592 9738
rect 6656 9948 6736 9976
rect 6276 8832 6328 8838
rect 6276 8774 6328 8780
rect 6380 8634 6408 9710
rect 6460 9376 6512 9382
rect 6656 9364 6684 9948
rect 6736 9930 6788 9936
rect 6512 9336 6684 9364
rect 6736 9376 6788 9382
rect 6460 9318 6512 9324
rect 6736 9318 6788 9324
rect 6368 8628 6420 8634
rect 6368 8570 6420 8576
rect 6184 8560 6236 8566
rect 6184 8502 6236 8508
rect 6196 8090 6224 8502
rect 6472 8498 6500 9318
rect 6748 9081 6776 9318
rect 6840 9178 6868 11086
rect 6920 10736 6972 10742
rect 6920 10678 6972 10684
rect 6932 10606 6960 10678
rect 6920 10600 6972 10606
rect 6920 10542 6972 10548
rect 7012 9920 7064 9926
rect 7012 9862 7064 9868
rect 6918 9752 6974 9761
rect 6918 9687 6974 9696
rect 6932 9586 6960 9687
rect 6920 9580 6972 9586
rect 6920 9522 6972 9528
rect 6828 9172 6880 9178
rect 6828 9114 6880 9120
rect 6734 9072 6790 9081
rect 6734 9007 6790 9016
rect 7024 8974 7052 9862
rect 7116 9518 7144 11154
rect 7216 10908 7524 10928
rect 7216 10906 7222 10908
rect 7278 10906 7302 10908
rect 7358 10906 7382 10908
rect 7438 10906 7462 10908
rect 7518 10906 7524 10908
rect 7278 10854 7280 10906
rect 7460 10854 7462 10906
rect 7216 10852 7222 10854
rect 7278 10852 7302 10854
rect 7358 10852 7382 10854
rect 7438 10852 7462 10854
rect 7518 10852 7524 10854
rect 7216 10832 7524 10852
rect 7562 10160 7618 10169
rect 7562 10095 7618 10104
rect 7216 9820 7524 9840
rect 7216 9818 7222 9820
rect 7278 9818 7302 9820
rect 7358 9818 7382 9820
rect 7438 9818 7462 9820
rect 7518 9818 7524 9820
rect 7278 9766 7280 9818
rect 7460 9766 7462 9818
rect 7216 9764 7222 9766
rect 7278 9764 7302 9766
rect 7358 9764 7382 9766
rect 7438 9764 7462 9766
rect 7518 9764 7524 9766
rect 7216 9744 7524 9764
rect 7380 9580 7432 9586
rect 7380 9522 7432 9528
rect 7104 9512 7156 9518
rect 7104 9454 7156 9460
rect 7392 9353 7420 9522
rect 7378 9344 7434 9353
rect 7378 9279 7434 9288
rect 7012 8968 7064 8974
rect 7012 8910 7064 8916
rect 6920 8900 6972 8906
rect 6920 8842 6972 8848
rect 6552 8832 6604 8838
rect 6552 8774 6604 8780
rect 6826 8800 6882 8809
rect 6460 8492 6512 8498
rect 6460 8434 6512 8440
rect 6276 8424 6328 8430
rect 6276 8366 6328 8372
rect 6184 8084 6236 8090
rect 6184 8026 6236 8032
rect 6196 7410 6224 8026
rect 6288 7721 6316 8366
rect 6368 8356 6420 8362
rect 6368 8298 6420 8304
rect 6274 7712 6330 7721
rect 6274 7647 6330 7656
rect 6184 7404 6236 7410
rect 6184 7346 6236 7352
rect 6274 6896 6330 6905
rect 6274 6831 6330 6840
rect 6104 6174 6224 6202
rect 6092 6112 6144 6118
rect 5538 6080 5594 6089
rect 5920 6072 6040 6100
rect 5538 6015 5594 6024
rect 5666 6012 5974 6032
rect 5666 6010 5672 6012
rect 5728 6010 5752 6012
rect 5808 6010 5832 6012
rect 5888 6010 5912 6012
rect 5968 6010 5974 6012
rect 5728 5958 5730 6010
rect 5910 5958 5912 6010
rect 5666 5956 5672 5958
rect 5728 5956 5752 5958
rect 5808 5956 5832 5958
rect 5888 5956 5912 5958
rect 5968 5956 5974 5958
rect 5666 5936 5974 5956
rect 5276 5630 5396 5658
rect 5448 5704 5500 5710
rect 5448 5646 5500 5652
rect 5632 5704 5684 5710
rect 5632 5646 5684 5652
rect 5276 5030 5304 5630
rect 5356 5568 5408 5574
rect 5356 5510 5408 5516
rect 5264 5024 5316 5030
rect 5264 4966 5316 4972
rect 5368 4690 5396 5510
rect 5448 5160 5500 5166
rect 5644 5114 5672 5646
rect 5448 5102 5500 5108
rect 5356 4684 5408 4690
rect 5356 4626 5408 4632
rect 5460 4622 5488 5102
rect 5552 5086 5672 5114
rect 5552 4758 5580 5086
rect 5666 4924 5974 4944
rect 5666 4922 5672 4924
rect 5728 4922 5752 4924
rect 5808 4922 5832 4924
rect 5888 4922 5912 4924
rect 5968 4922 5974 4924
rect 5728 4870 5730 4922
rect 5910 4870 5912 4922
rect 5666 4868 5672 4870
rect 5728 4868 5752 4870
rect 5808 4868 5832 4870
rect 5888 4868 5912 4870
rect 5968 4868 5974 4870
rect 5666 4848 5974 4868
rect 5540 4752 5592 4758
rect 5540 4694 5592 4700
rect 5906 4720 5962 4729
rect 5906 4655 5962 4664
rect 5172 4616 5224 4622
rect 5172 4558 5224 4564
rect 5448 4616 5500 4622
rect 5448 4558 5500 4564
rect 5722 4584 5778 4593
rect 5000 3454 5120 3482
rect 4712 2984 4764 2990
rect 4712 2926 4764 2932
rect 5000 2854 5028 3454
rect 5080 3392 5132 3398
rect 5080 3334 5132 3340
rect 5092 3058 5120 3334
rect 5080 3052 5132 3058
rect 5080 2994 5132 3000
rect 4528 2848 4580 2854
rect 4528 2790 4580 2796
rect 4988 2848 5040 2854
rect 4988 2790 5040 2796
rect 4540 2378 4568 2790
rect 5184 2582 5212 4558
rect 5920 4554 5948 4655
rect 5722 4519 5724 4528
rect 5776 4519 5778 4528
rect 5908 4548 5960 4554
rect 5724 4490 5776 4496
rect 5908 4490 5960 4496
rect 5920 4264 5948 4490
rect 6012 4486 6040 6072
rect 6092 6054 6144 6060
rect 6104 5778 6132 6054
rect 6092 5772 6144 5778
rect 6092 5714 6144 5720
rect 6104 5302 6132 5714
rect 6092 5296 6144 5302
rect 6092 5238 6144 5244
rect 6000 4480 6052 4486
rect 6000 4422 6052 4428
rect 5920 4236 6040 4264
rect 5264 4140 5316 4146
rect 5264 4082 5316 4088
rect 5276 2650 5304 4082
rect 5666 3836 5974 3856
rect 5666 3834 5672 3836
rect 5728 3834 5752 3836
rect 5808 3834 5832 3836
rect 5888 3834 5912 3836
rect 5968 3834 5974 3836
rect 5728 3782 5730 3834
rect 5910 3782 5912 3834
rect 5666 3780 5672 3782
rect 5728 3780 5752 3782
rect 5808 3780 5832 3782
rect 5888 3780 5912 3782
rect 5968 3780 5974 3782
rect 5666 3760 5974 3780
rect 6012 3738 6040 4236
rect 6196 4146 6224 6174
rect 6184 4140 6236 4146
rect 6104 4100 6184 4128
rect 6000 3732 6052 3738
rect 6000 3674 6052 3680
rect 5448 3664 5500 3670
rect 5448 3606 5500 3612
rect 5460 3466 5488 3606
rect 6012 3466 6040 3674
rect 5448 3460 5500 3466
rect 5448 3402 5500 3408
rect 6000 3460 6052 3466
rect 6000 3402 6052 3408
rect 5540 3392 5592 3398
rect 5540 3334 5592 3340
rect 5552 3194 5580 3334
rect 5540 3188 5592 3194
rect 5540 3130 5592 3136
rect 5666 2748 5974 2768
rect 5666 2746 5672 2748
rect 5728 2746 5752 2748
rect 5808 2746 5832 2748
rect 5888 2746 5912 2748
rect 5968 2746 5974 2748
rect 5728 2694 5730 2746
rect 5910 2694 5912 2746
rect 5666 2692 5672 2694
rect 5728 2692 5752 2694
rect 5808 2692 5832 2694
rect 5888 2692 5912 2694
rect 5968 2692 5974 2694
rect 5666 2672 5974 2692
rect 5264 2644 5316 2650
rect 5264 2586 5316 2592
rect 5172 2576 5224 2582
rect 5172 2518 5224 2524
rect 4344 2372 4396 2378
rect 4344 2314 4396 2320
rect 4528 2372 4580 2378
rect 4528 2314 4580 2320
rect 6104 2310 6132 4100
rect 6184 4082 6236 4088
rect 6184 3120 6236 3126
rect 6288 3097 6316 6831
rect 6380 4826 6408 8298
rect 6472 7206 6500 8434
rect 6564 8362 6592 8774
rect 6826 8735 6882 8744
rect 6642 8528 6698 8537
rect 6840 8498 6868 8735
rect 6932 8673 6960 8842
rect 7216 8732 7524 8752
rect 7216 8730 7222 8732
rect 7278 8730 7302 8732
rect 7358 8730 7382 8732
rect 7438 8730 7462 8732
rect 7518 8730 7524 8732
rect 7278 8678 7280 8730
rect 7460 8678 7462 8730
rect 7216 8676 7222 8678
rect 7278 8676 7302 8678
rect 7358 8676 7382 8678
rect 7438 8676 7462 8678
rect 7518 8676 7524 8678
rect 6918 8664 6974 8673
rect 7216 8656 7524 8676
rect 6918 8599 6974 8608
rect 7104 8560 7156 8566
rect 7104 8502 7156 8508
rect 6642 8463 6698 8472
rect 6736 8492 6788 8498
rect 6552 8356 6604 8362
rect 6552 8298 6604 8304
rect 6656 7886 6684 8463
rect 6736 8434 6788 8440
rect 6828 8492 6880 8498
rect 6828 8434 6880 8440
rect 6644 7880 6696 7886
rect 6644 7822 6696 7828
rect 6460 7200 6512 7206
rect 6460 7142 6512 7148
rect 6644 7200 6696 7206
rect 6644 7142 6696 7148
rect 6472 7002 6500 7142
rect 6460 6996 6512 7002
rect 6460 6938 6512 6944
rect 6472 6390 6500 6938
rect 6656 6934 6684 7142
rect 6644 6928 6696 6934
rect 6644 6870 6696 6876
rect 6460 6384 6512 6390
rect 6460 6326 6512 6332
rect 6472 5302 6500 6326
rect 6644 5908 6696 5914
rect 6644 5850 6696 5856
rect 6460 5296 6512 5302
rect 6460 5238 6512 5244
rect 6472 4826 6500 5238
rect 6656 5166 6684 5850
rect 6644 5160 6696 5166
rect 6644 5102 6696 5108
rect 6368 4820 6420 4826
rect 6368 4762 6420 4768
rect 6460 4820 6512 4826
rect 6460 4762 6512 4768
rect 6472 4486 6500 4762
rect 6656 4622 6684 5102
rect 6644 4616 6696 4622
rect 6644 4558 6696 4564
rect 6460 4480 6512 4486
rect 6460 4422 6512 4428
rect 6748 3942 6776 8434
rect 7012 8424 7064 8430
rect 7012 8366 7064 8372
rect 6828 7812 6880 7818
rect 6828 7754 6880 7760
rect 6840 6798 6868 7754
rect 6918 7576 6974 7585
rect 6918 7511 6974 7520
rect 6828 6792 6880 6798
rect 6828 6734 6880 6740
rect 6932 6390 6960 7511
rect 7024 6769 7052 8366
rect 7116 7002 7144 8502
rect 7216 7644 7524 7664
rect 7216 7642 7222 7644
rect 7278 7642 7302 7644
rect 7358 7642 7382 7644
rect 7438 7642 7462 7644
rect 7518 7642 7524 7644
rect 7278 7590 7280 7642
rect 7460 7590 7462 7642
rect 7216 7588 7222 7590
rect 7278 7588 7302 7590
rect 7358 7588 7382 7590
rect 7438 7588 7462 7590
rect 7518 7588 7524 7590
rect 7216 7568 7524 7588
rect 7576 7342 7604 10095
rect 7564 7336 7616 7342
rect 7564 7278 7616 7284
rect 7104 6996 7156 7002
rect 7104 6938 7156 6944
rect 7010 6760 7066 6769
rect 7010 6695 7066 6704
rect 7010 6488 7066 6497
rect 7010 6423 7066 6432
rect 6920 6384 6972 6390
rect 6920 6326 6972 6332
rect 7024 6322 7052 6423
rect 7012 6316 7064 6322
rect 7012 6258 7064 6264
rect 7116 4554 7144 6938
rect 7668 6746 7696 11698
rect 16592 11626 16620 13767
rect 16762 12880 16818 12889
rect 16762 12815 16818 12824
rect 16580 11620 16632 11626
rect 16580 11562 16632 11568
rect 8576 11552 8628 11558
rect 8576 11494 8628 11500
rect 13450 11520 13506 11529
rect 7932 11212 7984 11218
rect 7932 11154 7984 11160
rect 7944 10674 7972 11154
rect 8300 11144 8352 11150
rect 8114 11112 8170 11121
rect 8300 11086 8352 11092
rect 8114 11047 8170 11056
rect 8022 10704 8078 10713
rect 7932 10668 7984 10674
rect 8022 10639 8078 10648
rect 7932 10610 7984 10616
rect 7840 10192 7892 10198
rect 7838 10160 7840 10169
rect 7892 10160 7894 10169
rect 7838 10095 7894 10104
rect 7932 10056 7984 10062
rect 7838 10024 7894 10033
rect 7894 10004 7932 10010
rect 8036 10033 8064 10639
rect 7894 9998 7984 10004
rect 8022 10024 8078 10033
rect 7894 9982 7972 9998
rect 7838 9959 7894 9968
rect 8022 9959 8078 9968
rect 7852 8974 7880 9959
rect 7932 9716 7984 9722
rect 7932 9658 7984 9664
rect 7944 9330 7972 9658
rect 7944 9302 8064 9330
rect 7748 8968 7800 8974
rect 7748 8910 7800 8916
rect 7840 8968 7892 8974
rect 7840 8910 7892 8916
rect 7760 8090 7788 8910
rect 7840 8424 7892 8430
rect 7840 8366 7892 8372
rect 7748 8084 7800 8090
rect 7748 8026 7800 8032
rect 7748 7880 7800 7886
rect 7852 7868 7880 8366
rect 8036 8090 8064 9302
rect 8128 8956 8156 11047
rect 8312 10713 8340 11086
rect 8298 10704 8354 10713
rect 8208 10668 8260 10674
rect 8298 10639 8354 10648
rect 8484 10668 8536 10674
rect 8208 10610 8260 10616
rect 8484 10610 8536 10616
rect 8220 9994 8248 10610
rect 8300 10464 8352 10470
rect 8300 10406 8352 10412
rect 8208 9988 8260 9994
rect 8208 9930 8260 9936
rect 8220 9178 8248 9930
rect 8312 9353 8340 10406
rect 8392 10192 8444 10198
rect 8392 10134 8444 10140
rect 8298 9344 8354 9353
rect 8298 9279 8354 9288
rect 8208 9172 8260 9178
rect 8208 9114 8260 9120
rect 8208 8968 8260 8974
rect 8128 8928 8208 8956
rect 8208 8910 8260 8916
rect 8404 8838 8432 10134
rect 8496 9178 8524 10610
rect 8588 10062 8616 11494
rect 8766 11452 9074 11472
rect 13450 11455 13506 11464
rect 8766 11450 8772 11452
rect 8828 11450 8852 11452
rect 8908 11450 8932 11452
rect 8988 11450 9012 11452
rect 9068 11450 9074 11452
rect 8828 11398 8830 11450
rect 9010 11398 9012 11450
rect 8766 11396 8772 11398
rect 8828 11396 8852 11398
rect 8908 11396 8932 11398
rect 8988 11396 9012 11398
rect 9068 11396 9074 11398
rect 8766 11376 9074 11396
rect 9680 11348 9732 11354
rect 9680 11290 9732 11296
rect 9496 11280 9548 11286
rect 9496 11222 9548 11228
rect 9220 11144 9272 11150
rect 9220 11086 9272 11092
rect 9128 10668 9180 10674
rect 9128 10610 9180 10616
rect 8766 10364 9074 10384
rect 8766 10362 8772 10364
rect 8828 10362 8852 10364
rect 8908 10362 8932 10364
rect 8988 10362 9012 10364
rect 9068 10362 9074 10364
rect 8828 10310 8830 10362
rect 9010 10310 9012 10362
rect 8766 10308 8772 10310
rect 8828 10308 8852 10310
rect 8908 10308 8932 10310
rect 8988 10308 9012 10310
rect 9068 10308 9074 10310
rect 8766 10288 9074 10308
rect 8576 10056 8628 10062
rect 8576 9998 8628 10004
rect 9140 9722 9168 10610
rect 9232 10266 9260 11086
rect 9404 11008 9456 11014
rect 9508 10985 9536 11222
rect 9404 10950 9456 10956
rect 9494 10976 9550 10985
rect 9220 10260 9272 10266
rect 9220 10202 9272 10208
rect 9312 10124 9364 10130
rect 9312 10066 9364 10072
rect 9220 9920 9272 9926
rect 9220 9862 9272 9868
rect 9128 9716 9180 9722
rect 9128 9658 9180 9664
rect 8574 9480 8630 9489
rect 8574 9415 8630 9424
rect 8484 9172 8536 9178
rect 8484 9114 8536 9120
rect 8392 8832 8444 8838
rect 8392 8774 8444 8780
rect 8208 8560 8260 8566
rect 8208 8502 8260 8508
rect 8024 8084 8076 8090
rect 8024 8026 8076 8032
rect 7932 7948 7984 7954
rect 7932 7890 7984 7896
rect 7800 7840 7880 7868
rect 7748 7822 7800 7828
rect 7760 7546 7788 7822
rect 7748 7540 7800 7546
rect 7748 7482 7800 7488
rect 7840 7540 7892 7546
rect 7840 7482 7892 7488
rect 7576 6718 7696 6746
rect 7216 6556 7524 6576
rect 7216 6554 7222 6556
rect 7278 6554 7302 6556
rect 7358 6554 7382 6556
rect 7438 6554 7462 6556
rect 7518 6554 7524 6556
rect 7278 6502 7280 6554
rect 7460 6502 7462 6554
rect 7216 6500 7222 6502
rect 7278 6500 7302 6502
rect 7358 6500 7382 6502
rect 7438 6500 7462 6502
rect 7518 6500 7524 6502
rect 7216 6480 7524 6500
rect 7286 6352 7342 6361
rect 7286 6287 7342 6296
rect 7470 6352 7526 6361
rect 7470 6287 7472 6296
rect 7300 6186 7328 6287
rect 7524 6287 7526 6296
rect 7472 6258 7524 6264
rect 7576 6202 7604 6718
rect 7656 6656 7708 6662
rect 7656 6598 7708 6604
rect 7288 6180 7340 6186
rect 7288 6122 7340 6128
rect 7484 6174 7604 6202
rect 7484 5914 7512 6174
rect 7564 6112 7616 6118
rect 7564 6054 7616 6060
rect 7472 5908 7524 5914
rect 7472 5850 7524 5856
rect 7216 5468 7524 5488
rect 7216 5466 7222 5468
rect 7278 5466 7302 5468
rect 7358 5466 7382 5468
rect 7438 5466 7462 5468
rect 7518 5466 7524 5468
rect 7278 5414 7280 5466
rect 7460 5414 7462 5466
rect 7216 5412 7222 5414
rect 7278 5412 7302 5414
rect 7358 5412 7382 5414
rect 7438 5412 7462 5414
rect 7518 5412 7524 5414
rect 7216 5392 7524 5412
rect 7576 4706 7604 6054
rect 7668 5642 7696 6598
rect 7748 6384 7800 6390
rect 7748 6326 7800 6332
rect 7760 5817 7788 6326
rect 7746 5808 7802 5817
rect 7746 5743 7802 5752
rect 7656 5636 7708 5642
rect 7656 5578 7708 5584
rect 7748 5364 7800 5370
rect 7748 5306 7800 5312
rect 7484 4690 7604 4706
rect 7760 4690 7788 5306
rect 7852 5030 7880 7482
rect 7944 6186 7972 7890
rect 8036 7546 8064 8026
rect 8024 7540 8076 7546
rect 8024 7482 8076 7488
rect 8116 7472 8168 7478
rect 8116 7414 8168 7420
rect 8128 6730 8156 7414
rect 8220 6934 8248 8502
rect 8588 8498 8616 9415
rect 8766 9276 9074 9296
rect 8766 9274 8772 9276
rect 8828 9274 8852 9276
rect 8908 9274 8932 9276
rect 8988 9274 9012 9276
rect 9068 9274 9074 9276
rect 8828 9222 8830 9274
rect 9010 9222 9012 9274
rect 8766 9220 8772 9222
rect 8828 9220 8852 9222
rect 8908 9220 8932 9222
rect 8988 9220 9012 9222
rect 9068 9220 9074 9222
rect 8766 9200 9074 9220
rect 8668 9036 8720 9042
rect 8668 8978 8720 8984
rect 8680 8498 8708 8978
rect 8300 8492 8352 8498
rect 8300 8434 8352 8440
rect 8392 8492 8444 8498
rect 8392 8434 8444 8440
rect 8576 8492 8628 8498
rect 8576 8434 8628 8440
rect 8668 8492 8720 8498
rect 8668 8434 8720 8440
rect 8208 6928 8260 6934
rect 8208 6870 8260 6876
rect 8312 6882 8340 8434
rect 8404 7993 8432 8434
rect 8484 8288 8536 8294
rect 8484 8230 8536 8236
rect 8390 7984 8446 7993
rect 8390 7919 8446 7928
rect 8392 7880 8444 7886
rect 8392 7822 8444 7828
rect 8404 7562 8432 7822
rect 8496 7750 8524 8230
rect 8766 8188 9074 8208
rect 8766 8186 8772 8188
rect 8828 8186 8852 8188
rect 8908 8186 8932 8188
rect 8988 8186 9012 8188
rect 9068 8186 9074 8188
rect 8828 8134 8830 8186
rect 9010 8134 9012 8186
rect 8766 8132 8772 8134
rect 8828 8132 8852 8134
rect 8908 8132 8932 8134
rect 8988 8132 9012 8134
rect 9068 8132 9074 8134
rect 8766 8112 9074 8132
rect 9232 8090 9260 9862
rect 9324 9722 9352 10066
rect 9312 9716 9364 9722
rect 9312 9658 9364 9664
rect 9324 9042 9352 9658
rect 9416 9353 9444 10950
rect 9494 10911 9550 10920
rect 9692 10305 9720 11290
rect 13464 10577 13492 11455
rect 13726 11248 13782 11257
rect 13726 11183 13782 11192
rect 13450 10568 13506 10577
rect 13450 10503 13506 10512
rect 13544 10464 13596 10470
rect 13544 10406 13596 10412
rect 9678 10296 9734 10305
rect 9678 10231 9734 10240
rect 9402 9344 9458 9353
rect 9402 9279 9458 9288
rect 10140 9104 10192 9110
rect 13556 9081 13584 10406
rect 13634 10024 13690 10033
rect 13634 9959 13690 9968
rect 10140 9046 10192 9052
rect 13542 9072 13598 9081
rect 9312 9036 9364 9042
rect 9312 8978 9364 8984
rect 9588 8628 9640 8634
rect 9588 8570 9640 8576
rect 9600 8265 9628 8570
rect 9586 8256 9642 8265
rect 9586 8191 9642 8200
rect 9220 8084 9272 8090
rect 9220 8026 9272 8032
rect 10152 7993 10180 9046
rect 13542 9007 13598 9016
rect 13450 8936 13506 8945
rect 13450 8871 13452 8880
rect 13504 8871 13506 8880
rect 13452 8842 13504 8848
rect 13648 8673 13676 9959
rect 13634 8664 13690 8673
rect 13634 8599 13690 8608
rect 10876 8424 10928 8430
rect 10876 8366 10928 8372
rect 9310 7984 9366 7993
rect 9310 7919 9312 7928
rect 9364 7919 9366 7928
rect 10138 7984 10194 7993
rect 10138 7919 10194 7928
rect 9312 7890 9364 7896
rect 9140 7806 9444 7834
rect 9140 7750 9168 7806
rect 8484 7744 8536 7750
rect 8484 7686 8536 7692
rect 9128 7744 9180 7750
rect 9128 7686 9180 7692
rect 9220 7744 9272 7750
rect 9220 7686 9272 7692
rect 8404 7546 8524 7562
rect 8404 7540 8536 7546
rect 8404 7534 8484 7540
rect 8484 7482 8536 7488
rect 8576 7472 8628 7478
rect 8576 7414 8628 7420
rect 8312 6854 8524 6882
rect 8208 6792 8260 6798
rect 8208 6734 8260 6740
rect 8300 6792 8352 6798
rect 8300 6734 8352 6740
rect 8116 6724 8168 6730
rect 8116 6666 8168 6672
rect 8022 6352 8078 6361
rect 8022 6287 8078 6296
rect 7932 6180 7984 6186
rect 7932 6122 7984 6128
rect 7944 5914 7972 6122
rect 7932 5908 7984 5914
rect 7932 5850 7984 5856
rect 7932 5704 7984 5710
rect 7932 5646 7984 5652
rect 7840 5024 7892 5030
rect 7840 4966 7892 4972
rect 7472 4684 7604 4690
rect 7524 4678 7604 4684
rect 7748 4684 7800 4690
rect 7472 4626 7524 4632
rect 7748 4626 7800 4632
rect 7104 4548 7156 4554
rect 7104 4490 7156 4496
rect 7216 4380 7524 4400
rect 7216 4378 7222 4380
rect 7278 4378 7302 4380
rect 7358 4378 7382 4380
rect 7438 4378 7462 4380
rect 7518 4378 7524 4380
rect 7278 4326 7280 4378
rect 7460 4326 7462 4378
rect 7216 4324 7222 4326
rect 7278 4324 7302 4326
rect 7358 4324 7382 4326
rect 7438 4324 7462 4326
rect 7518 4324 7524 4326
rect 7216 4304 7524 4324
rect 7656 4140 7708 4146
rect 7656 4082 7708 4088
rect 7104 4004 7156 4010
rect 7104 3946 7156 3952
rect 6736 3936 6788 3942
rect 6736 3878 6788 3884
rect 7116 3602 7144 3946
rect 7668 3670 7696 4082
rect 7944 4078 7972 5646
rect 8036 4282 8064 6287
rect 8116 5024 8168 5030
rect 8116 4966 8168 4972
rect 8128 4486 8156 4966
rect 8220 4826 8248 6734
rect 8208 4820 8260 4826
rect 8208 4762 8260 4768
rect 8116 4480 8168 4486
rect 8116 4422 8168 4428
rect 8024 4276 8076 4282
rect 8024 4218 8076 4224
rect 8208 4208 8260 4214
rect 8208 4150 8260 4156
rect 7932 4072 7984 4078
rect 7932 4014 7984 4020
rect 8024 3732 8076 3738
rect 8024 3674 8076 3680
rect 7656 3664 7708 3670
rect 7656 3606 7708 3612
rect 7104 3596 7156 3602
rect 7104 3538 7156 3544
rect 6460 3528 6512 3534
rect 6460 3470 6512 3476
rect 6184 3062 6236 3068
rect 6274 3088 6330 3097
rect 6196 2650 6224 3062
rect 6274 3023 6330 3032
rect 6184 2644 6236 2650
rect 6184 2586 6236 2592
rect 6472 2514 6500 3470
rect 7932 3460 7984 3466
rect 7932 3402 7984 3408
rect 6552 3392 6604 3398
rect 6552 3334 6604 3340
rect 6564 2514 6592 3334
rect 7216 3292 7524 3312
rect 7216 3290 7222 3292
rect 7278 3290 7302 3292
rect 7358 3290 7382 3292
rect 7438 3290 7462 3292
rect 7518 3290 7524 3292
rect 7278 3238 7280 3290
rect 7460 3238 7462 3290
rect 7216 3236 7222 3238
rect 7278 3236 7302 3238
rect 7358 3236 7382 3238
rect 7438 3236 7462 3238
rect 7518 3236 7524 3238
rect 7216 3216 7524 3236
rect 7380 3052 7432 3058
rect 7380 2994 7432 3000
rect 7472 3052 7524 3058
rect 7472 2994 7524 3000
rect 7392 2582 7420 2994
rect 7484 2854 7512 2994
rect 7472 2848 7524 2854
rect 7470 2816 7472 2825
rect 7564 2848 7616 2854
rect 7524 2816 7526 2825
rect 7564 2790 7616 2796
rect 7470 2751 7526 2760
rect 7380 2576 7432 2582
rect 7380 2518 7432 2524
rect 6460 2508 6512 2514
rect 6460 2450 6512 2456
rect 6552 2508 6604 2514
rect 6552 2450 6604 2456
rect 7576 2378 7604 2790
rect 7944 2650 7972 3402
rect 8036 3058 8064 3674
rect 8116 3528 8168 3534
rect 8116 3470 8168 3476
rect 8128 3194 8156 3470
rect 8220 3398 8248 4150
rect 8312 3738 8340 6734
rect 8392 6248 8444 6254
rect 8392 6190 8444 6196
rect 8404 6118 8432 6190
rect 8496 6118 8524 6854
rect 8392 6112 8444 6118
rect 8392 6054 8444 6060
rect 8484 6112 8536 6118
rect 8484 6054 8536 6060
rect 8392 5636 8444 5642
rect 8392 5578 8444 5584
rect 8300 3732 8352 3738
rect 8300 3674 8352 3680
rect 8208 3392 8260 3398
rect 8208 3334 8260 3340
rect 8116 3188 8168 3194
rect 8116 3130 8168 3136
rect 8024 3052 8076 3058
rect 8024 2994 8076 3000
rect 8404 2990 8432 5578
rect 8484 5024 8536 5030
rect 8484 4966 8536 4972
rect 8496 4554 8524 4966
rect 8484 4548 8536 4554
rect 8484 4490 8536 4496
rect 8588 3942 8616 7414
rect 8668 7404 8720 7410
rect 8668 7346 8720 7352
rect 8680 7313 8708 7346
rect 8666 7304 8722 7313
rect 8666 7239 8722 7248
rect 9036 7268 9088 7274
rect 9088 7228 9168 7256
rect 9036 7210 9088 7216
rect 8766 7100 9074 7120
rect 8766 7098 8772 7100
rect 8828 7098 8852 7100
rect 8908 7098 8932 7100
rect 8988 7098 9012 7100
rect 9068 7098 9074 7100
rect 8828 7046 8830 7098
rect 9010 7046 9012 7098
rect 8766 7044 8772 7046
rect 8828 7044 8852 7046
rect 8908 7044 8932 7046
rect 8988 7044 9012 7046
rect 9068 7044 9074 7046
rect 8766 7024 9074 7044
rect 9140 6798 9168 7228
rect 9232 7002 9260 7686
rect 9220 6996 9272 7002
rect 9220 6938 9272 6944
rect 9312 6860 9364 6866
rect 9312 6802 9364 6808
rect 9128 6792 9180 6798
rect 9128 6734 9180 6740
rect 8666 6216 8722 6225
rect 8666 6151 8722 6160
rect 8680 5794 8708 6151
rect 9128 6112 9180 6118
rect 9128 6054 9180 6060
rect 8766 6012 9074 6032
rect 8766 6010 8772 6012
rect 8828 6010 8852 6012
rect 8908 6010 8932 6012
rect 8988 6010 9012 6012
rect 9068 6010 9074 6012
rect 8828 5958 8830 6010
rect 9010 5958 9012 6010
rect 8766 5956 8772 5958
rect 8828 5956 8852 5958
rect 8908 5956 8932 5958
rect 8988 5956 9012 5958
rect 9068 5956 9074 5958
rect 8766 5936 9074 5956
rect 9140 5794 9168 6054
rect 8680 5766 8800 5794
rect 8668 5704 8720 5710
rect 8668 5646 8720 5652
rect 8680 5370 8708 5646
rect 8772 5370 8800 5766
rect 9048 5766 9168 5794
rect 8668 5364 8720 5370
rect 8668 5306 8720 5312
rect 8760 5364 8812 5370
rect 8812 5324 8892 5352
rect 8760 5306 8812 5312
rect 8668 5228 8720 5234
rect 8668 5170 8720 5176
rect 8680 4282 8708 5170
rect 8864 5137 8892 5324
rect 8850 5128 8906 5137
rect 9048 5114 9076 5766
rect 9128 5704 9180 5710
rect 9128 5646 9180 5652
rect 9140 5370 9168 5646
rect 9220 5568 9272 5574
rect 9220 5510 9272 5516
rect 9128 5364 9180 5370
rect 9128 5306 9180 5312
rect 9048 5086 9168 5114
rect 8850 5063 8906 5072
rect 8766 4924 9074 4944
rect 8766 4922 8772 4924
rect 8828 4922 8852 4924
rect 8908 4922 8932 4924
rect 8988 4922 9012 4924
rect 9068 4922 9074 4924
rect 8828 4870 8830 4922
rect 9010 4870 9012 4922
rect 8766 4868 8772 4870
rect 8828 4868 8852 4870
rect 8908 4868 8932 4870
rect 8988 4868 9012 4870
rect 9068 4868 9074 4870
rect 8766 4848 9074 4868
rect 9140 4826 9168 5086
rect 9128 4820 9180 4826
rect 9128 4762 9180 4768
rect 8758 4720 8814 4729
rect 8758 4655 8814 4664
rect 8668 4276 8720 4282
rect 8668 4218 8720 4224
rect 8772 4146 8800 4655
rect 9232 4622 9260 5510
rect 9220 4616 9272 4622
rect 9220 4558 9272 4564
rect 9220 4480 9272 4486
rect 9220 4422 9272 4428
rect 9232 4146 9260 4422
rect 8760 4140 8812 4146
rect 8760 4082 8812 4088
rect 9220 4140 9272 4146
rect 9220 4082 9272 4088
rect 8576 3936 8628 3942
rect 8576 3878 8628 3884
rect 8668 3936 8720 3942
rect 8668 3878 8720 3884
rect 8484 3052 8536 3058
rect 8484 2994 8536 3000
rect 8392 2984 8444 2990
rect 8392 2926 8444 2932
rect 8116 2848 8168 2854
rect 8116 2790 8168 2796
rect 8298 2816 8354 2825
rect 7932 2644 7984 2650
rect 7932 2586 7984 2592
rect 8128 2446 8156 2790
rect 8496 2774 8524 2994
rect 8680 2854 8708 3878
rect 8766 3836 9074 3856
rect 8766 3834 8772 3836
rect 8828 3834 8852 3836
rect 8908 3834 8932 3836
rect 8988 3834 9012 3836
rect 9068 3834 9074 3836
rect 8828 3782 8830 3834
rect 9010 3782 9012 3834
rect 8766 3780 8772 3782
rect 8828 3780 8852 3782
rect 8908 3780 8932 3782
rect 8988 3780 9012 3782
rect 9068 3780 9074 3782
rect 8766 3760 9074 3780
rect 9324 3738 9352 6802
rect 9416 6798 9444 7806
rect 9404 6792 9456 6798
rect 9404 6734 9456 6740
rect 9588 6724 9640 6730
rect 9588 6666 9640 6672
rect 9496 6180 9548 6186
rect 9496 6122 9548 6128
rect 9404 6112 9456 6118
rect 9404 6054 9456 6060
rect 9312 3732 9364 3738
rect 9312 3674 9364 3680
rect 9416 3534 9444 6054
rect 9508 5234 9536 6122
rect 9600 5370 9628 6666
rect 9680 5772 9732 5778
rect 9680 5714 9732 5720
rect 9588 5364 9640 5370
rect 9588 5306 9640 5312
rect 9496 5228 9548 5234
rect 9496 5170 9548 5176
rect 9496 5092 9548 5098
rect 9496 5034 9548 5040
rect 9508 3942 9536 5034
rect 9692 4729 9720 5714
rect 10888 5001 10916 8366
rect 13544 8016 13596 8022
rect 13544 7958 13596 7964
rect 13450 7712 13506 7721
rect 13450 7647 13452 7656
rect 13504 7647 13506 7656
rect 13452 7618 13504 7624
rect 13556 7313 13584 7958
rect 13636 7880 13688 7886
rect 13636 7822 13688 7828
rect 13542 7304 13598 7313
rect 13542 7239 13598 7248
rect 13648 7041 13676 7822
rect 13740 7750 13768 11183
rect 13820 11076 13872 11082
rect 13820 11018 13872 11024
rect 13832 9897 13860 11018
rect 16776 10606 16804 12815
rect 16764 10600 16816 10606
rect 16764 10542 16816 10548
rect 13818 9888 13874 9897
rect 13818 9823 13874 9832
rect 13820 9784 13872 9790
rect 13820 9726 13872 9732
rect 13832 9625 13860 9726
rect 13818 9616 13874 9625
rect 13818 9551 13874 9560
rect 22376 8900 22428 8906
rect 22376 8842 22428 8848
rect 13820 8560 13872 8566
rect 13820 8502 13872 8508
rect 13832 7857 13860 8502
rect 13818 7848 13874 7857
rect 13818 7783 13874 7792
rect 13728 7744 13780 7750
rect 13728 7686 13780 7692
rect 22284 7676 22336 7682
rect 22284 7618 22336 7624
rect 13818 7440 13874 7449
rect 13818 7375 13874 7384
rect 13832 7342 13860 7375
rect 13820 7336 13872 7342
rect 13820 7278 13872 7284
rect 19432 7336 19484 7342
rect 19432 7278 19484 7284
rect 13728 7200 13780 7206
rect 13728 7142 13780 7148
rect 13634 7032 13690 7041
rect 13634 6967 13690 6976
rect 13636 6452 13688 6458
rect 13636 6394 13688 6400
rect 12806 6080 12862 6089
rect 12806 6015 12862 6024
rect 12820 5846 12848 6015
rect 12808 5840 12860 5846
rect 12808 5782 12860 5788
rect 10874 4992 10930 5001
rect 10874 4927 10930 4936
rect 9678 4720 9734 4729
rect 9678 4655 9734 4664
rect 9496 3936 9548 3942
rect 9496 3878 9548 3884
rect 8760 3528 8812 3534
rect 8760 3470 8812 3476
rect 9128 3528 9180 3534
rect 9128 3470 9180 3476
rect 9404 3528 9456 3534
rect 9404 3470 9456 3476
rect 8772 3194 8800 3470
rect 8760 3188 8812 3194
rect 8760 3130 8812 3136
rect 8668 2848 8720 2854
rect 8668 2790 8720 2796
rect 8298 2751 8354 2760
rect 8312 2446 8340 2751
rect 8404 2746 8524 2774
rect 8404 2446 8432 2746
rect 8116 2440 8168 2446
rect 8116 2382 8168 2388
rect 8300 2440 8352 2446
rect 8300 2382 8352 2388
rect 8392 2440 8444 2446
rect 8392 2382 8444 2388
rect 8680 2378 8708 2790
rect 8766 2748 9074 2768
rect 8766 2746 8772 2748
rect 8828 2746 8852 2748
rect 8908 2746 8932 2748
rect 8988 2746 9012 2748
rect 9068 2746 9074 2748
rect 8828 2694 8830 2746
rect 9010 2694 9012 2746
rect 8766 2692 8772 2694
rect 8828 2692 8852 2694
rect 8908 2692 8932 2694
rect 8988 2692 9012 2694
rect 9068 2692 9074 2694
rect 8766 2672 9074 2692
rect 9140 2650 9168 3470
rect 9692 3194 9720 4655
rect 13648 3777 13676 6394
rect 13740 6361 13768 7142
rect 13818 6624 13874 6633
rect 13818 6559 13874 6568
rect 13832 6390 13860 6559
rect 13820 6384 13872 6390
rect 13726 6352 13782 6361
rect 13820 6326 13872 6332
rect 13726 6287 13782 6296
rect 13728 5908 13780 5914
rect 13728 5850 13780 5856
rect 13634 3768 13690 3777
rect 13634 3703 13690 3712
rect 13740 3369 13768 5850
rect 13818 4448 13874 4457
rect 13818 4383 13874 4392
rect 13726 3360 13782 3369
rect 13726 3295 13782 3304
rect 9680 3188 9732 3194
rect 9680 3130 9732 3136
rect 9496 3120 9548 3126
rect 9496 3062 9548 3068
rect 9312 2916 9364 2922
rect 9312 2858 9364 2864
rect 9324 2650 9352 2858
rect 9128 2644 9180 2650
rect 9128 2586 9180 2592
rect 9312 2644 9364 2650
rect 9312 2586 9364 2592
rect 9508 2446 9536 3062
rect 13832 2854 13860 4383
rect 13820 2848 13872 2854
rect 13820 2790 13872 2796
rect 9496 2440 9548 2446
rect 19444 2417 19472 7278
rect 9496 2382 9548 2388
rect 19430 2408 19486 2417
rect 7564 2372 7616 2378
rect 7564 2314 7616 2320
rect 8668 2372 8720 2378
rect 19430 2343 19486 2352
rect 8668 2314 8720 2320
rect 6092 2304 6144 2310
rect 6092 2246 6144 2252
rect 4116 2204 4424 2224
rect 4116 2202 4122 2204
rect 4178 2202 4202 2204
rect 4258 2202 4282 2204
rect 4338 2202 4362 2204
rect 4418 2202 4424 2204
rect 4178 2150 4180 2202
rect 4360 2150 4362 2202
rect 4116 2148 4122 2150
rect 4178 2148 4202 2150
rect 4258 2148 4282 2150
rect 4338 2148 4362 2150
rect 4418 2148 4424 2150
rect 4116 2128 4424 2148
rect 7216 2204 7524 2224
rect 7216 2202 7222 2204
rect 7278 2202 7302 2204
rect 7358 2202 7382 2204
rect 7438 2202 7462 2204
rect 7518 2202 7524 2204
rect 7278 2150 7280 2202
rect 7460 2150 7462 2202
rect 7216 2148 7222 2150
rect 7278 2148 7302 2150
rect 7358 2148 7382 2150
rect 7438 2148 7462 2150
rect 7518 2148 7524 2150
rect 7216 2128 7524 2148
rect 22296 785 22324 7618
rect 22282 776 22338 785
rect 22282 711 22338 720
rect 3514 504 3570 513
rect 3514 439 3570 448
rect 22388 241 22416 8842
rect 22374 232 22430 241
rect 22374 167 22430 176
<< via2 >>
rect 16578 13776 16634 13832
rect 2410 13368 2466 13424
rect 2318 12416 2374 12472
rect 2226 10784 2282 10840
rect 1490 10532 1546 10568
rect 1490 10512 1492 10532
rect 1492 10512 1544 10532
rect 1544 10512 1546 10532
rect 1674 9560 1730 9616
rect 1306 8744 1362 8800
rect 1490 8472 1546 8528
rect 1398 6840 1454 6896
rect 1306 6568 1362 6624
rect 1214 6024 1270 6080
rect 1858 9424 1914 9480
rect 1766 8356 1822 8392
rect 1766 8336 1768 8356
rect 1768 8336 1820 8356
rect 1820 8336 1822 8356
rect 1674 7520 1730 7576
rect 2042 9052 2044 9072
rect 2044 9052 2096 9072
rect 2096 9052 2098 9072
rect 2042 9016 2098 9052
rect 6090 13096 6146 13152
rect 5998 12144 6054 12200
rect 3146 11872 3202 11928
rect 2572 11450 2628 11452
rect 2652 11450 2708 11452
rect 2732 11450 2788 11452
rect 2812 11450 2868 11452
rect 2572 11398 2618 11450
rect 2618 11398 2628 11450
rect 2652 11398 2682 11450
rect 2682 11398 2694 11450
rect 2694 11398 2708 11450
rect 2732 11398 2746 11450
rect 2746 11398 2758 11450
rect 2758 11398 2788 11450
rect 2812 11398 2822 11450
rect 2822 11398 2868 11450
rect 2572 11396 2628 11398
rect 2652 11396 2708 11398
rect 2732 11396 2788 11398
rect 2812 11396 2868 11398
rect 2962 11328 3018 11384
rect 2572 10362 2628 10364
rect 2652 10362 2708 10364
rect 2732 10362 2788 10364
rect 2812 10362 2868 10364
rect 2572 10310 2618 10362
rect 2618 10310 2628 10362
rect 2652 10310 2682 10362
rect 2682 10310 2694 10362
rect 2694 10310 2708 10362
rect 2732 10310 2746 10362
rect 2746 10310 2758 10362
rect 2758 10310 2788 10362
rect 2812 10310 2822 10362
rect 2822 10310 2868 10362
rect 2572 10308 2628 10310
rect 2652 10308 2708 10310
rect 2732 10308 2788 10310
rect 2812 10308 2868 10310
rect 2318 10104 2374 10160
rect 3054 11056 3110 11112
rect 2778 9832 2834 9888
rect 3514 11192 3570 11248
rect 4342 11192 4398 11248
rect 4710 11192 4766 11248
rect 3330 10648 3386 10704
rect 2572 9274 2628 9276
rect 2652 9274 2708 9276
rect 2732 9274 2788 9276
rect 2812 9274 2868 9276
rect 2572 9222 2618 9274
rect 2618 9222 2628 9274
rect 2652 9222 2682 9274
rect 2682 9222 2694 9274
rect 2694 9222 2708 9274
rect 2732 9222 2746 9274
rect 2746 9222 2758 9274
rect 2758 9222 2788 9274
rect 2812 9222 2822 9274
rect 2822 9222 2868 9274
rect 2572 9220 2628 9222
rect 2652 9220 2708 9222
rect 2732 9220 2788 9222
rect 2812 9220 2868 9222
rect 2962 9152 3018 9208
rect 2410 8880 2466 8936
rect 3146 8744 3202 8800
rect 2572 8186 2628 8188
rect 2652 8186 2708 8188
rect 2732 8186 2788 8188
rect 2812 8186 2868 8188
rect 2572 8134 2618 8186
rect 2618 8134 2628 8186
rect 2652 8134 2682 8186
rect 2682 8134 2694 8186
rect 2694 8134 2708 8186
rect 2732 8134 2746 8186
rect 2746 8134 2758 8186
rect 2758 8134 2788 8186
rect 2812 8134 2822 8186
rect 2822 8134 2868 8186
rect 2572 8132 2628 8134
rect 2652 8132 2708 8134
rect 2732 8132 2788 8134
rect 2812 8132 2868 8134
rect 2318 7928 2374 7984
rect 3054 8200 3110 8256
rect 2134 7792 2190 7848
rect 2042 6704 2098 6760
rect 2042 6160 2098 6216
rect 2318 5752 2374 5808
rect 2778 7656 2834 7712
rect 2870 7520 2926 7576
rect 3054 7540 3110 7576
rect 3054 7520 3056 7540
rect 3056 7520 3108 7540
rect 3108 7520 3110 7540
rect 2870 7248 2926 7304
rect 2572 7098 2628 7100
rect 2652 7098 2708 7100
rect 2732 7098 2788 7100
rect 2812 7098 2868 7100
rect 2572 7046 2618 7098
rect 2618 7046 2628 7098
rect 2652 7046 2682 7098
rect 2682 7046 2694 7098
rect 2694 7046 2708 7098
rect 2732 7046 2746 7098
rect 2746 7046 2758 7098
rect 2758 7046 2788 7098
rect 2812 7046 2822 7098
rect 2822 7046 2868 7098
rect 2572 7044 2628 7046
rect 2652 7044 2708 7046
rect 2732 7044 2788 7046
rect 2812 7044 2868 7046
rect 2410 5208 2466 5264
rect 2410 3576 2466 3632
rect 2686 5888 2742 5944
rect 2962 6704 3018 6760
rect 2778 4972 2780 4992
rect 2780 4972 2832 4992
rect 2832 4972 2834 4992
rect 2778 4936 2834 4972
rect 2686 3596 2742 3632
rect 2686 3576 2688 3596
rect 2688 3576 2740 3596
rect 2740 3576 2742 3596
rect 1122 1400 1178 1456
rect 3882 10784 3938 10840
rect 3514 10376 3570 10432
rect 4122 10906 4178 10908
rect 4202 10906 4258 10908
rect 4282 10906 4338 10908
rect 4362 10906 4418 10908
rect 4122 10854 4168 10906
rect 4168 10854 4178 10906
rect 4202 10854 4232 10906
rect 4232 10854 4244 10906
rect 4244 10854 4258 10906
rect 4282 10854 4296 10906
rect 4296 10854 4308 10906
rect 4308 10854 4338 10906
rect 4362 10854 4372 10906
rect 4372 10854 4418 10906
rect 4122 10852 4178 10854
rect 4202 10852 4258 10854
rect 4282 10852 4338 10854
rect 4362 10852 4418 10854
rect 3606 10140 3608 10160
rect 3608 10140 3660 10160
rect 3660 10140 3662 10160
rect 3606 10104 3662 10140
rect 3514 9968 3570 10024
rect 3790 9832 3846 9888
rect 3790 9424 3846 9480
rect 4122 9818 4178 9820
rect 4202 9818 4258 9820
rect 4282 9818 4338 9820
rect 4362 9818 4418 9820
rect 4122 9766 4168 9818
rect 4168 9766 4178 9818
rect 4202 9766 4232 9818
rect 4232 9766 4244 9818
rect 4244 9766 4258 9818
rect 4282 9766 4296 9818
rect 4296 9766 4308 9818
rect 4308 9766 4338 9818
rect 4362 9766 4372 9818
rect 4372 9766 4418 9818
rect 4122 9764 4178 9766
rect 4202 9764 4258 9766
rect 4282 9764 4338 9766
rect 4362 9764 4418 9766
rect 4526 9716 4582 9752
rect 4526 9696 4528 9716
rect 4528 9696 4580 9716
rect 4580 9696 4582 9716
rect 3698 8880 3754 8936
rect 3882 8780 3884 8800
rect 3884 8780 3936 8800
rect 3936 8780 3938 8800
rect 2870 3984 2926 4040
rect 3882 8744 3938 8780
rect 3698 8064 3754 8120
rect 3606 7928 3662 7984
rect 3790 7656 3846 7712
rect 3422 7112 3478 7168
rect 3330 6704 3386 6760
rect 3238 2896 3294 2952
rect 3146 1944 3202 2000
rect 3422 1672 3478 1728
rect 2778 992 2834 1048
rect 4122 8730 4178 8732
rect 4202 8730 4258 8732
rect 4282 8730 4338 8732
rect 4362 8730 4418 8732
rect 4122 8678 4168 8730
rect 4168 8678 4178 8730
rect 4202 8678 4232 8730
rect 4232 8678 4244 8730
rect 4244 8678 4258 8730
rect 4282 8678 4296 8730
rect 4296 8678 4308 8730
rect 4308 8678 4338 8730
rect 4362 8678 4372 8730
rect 4372 8678 4418 8730
rect 4122 8676 4178 8678
rect 4202 8676 4258 8678
rect 4282 8676 4338 8678
rect 4362 8676 4418 8678
rect 4894 10240 4950 10296
rect 4618 8744 4674 8800
rect 3974 7928 4030 7984
rect 4122 7642 4178 7644
rect 4202 7642 4258 7644
rect 4282 7642 4338 7644
rect 4362 7642 4418 7644
rect 4122 7590 4168 7642
rect 4168 7590 4178 7642
rect 4202 7590 4232 7642
rect 4232 7590 4244 7642
rect 4244 7590 4258 7642
rect 4282 7590 4296 7642
rect 4296 7590 4308 7642
rect 4308 7590 4338 7642
rect 4362 7590 4372 7642
rect 4372 7590 4418 7642
rect 4122 7588 4178 7590
rect 4202 7588 4258 7590
rect 4282 7588 4338 7590
rect 4362 7588 4418 7590
rect 3882 6976 3938 7032
rect 4526 6976 4582 7032
rect 3606 6296 3662 6352
rect 3882 6568 3938 6624
rect 4122 6554 4178 6556
rect 4202 6554 4258 6556
rect 4282 6554 4338 6556
rect 4362 6554 4418 6556
rect 4122 6502 4168 6554
rect 4168 6502 4178 6554
rect 4202 6502 4232 6554
rect 4232 6502 4244 6554
rect 4244 6502 4258 6554
rect 4282 6502 4296 6554
rect 4296 6502 4308 6554
rect 4308 6502 4338 6554
rect 4362 6502 4372 6554
rect 4372 6502 4418 6554
rect 4122 6500 4178 6502
rect 4202 6500 4258 6502
rect 4282 6500 4338 6502
rect 4362 6500 4418 6502
rect 4122 5466 4178 5468
rect 4202 5466 4258 5468
rect 4282 5466 4338 5468
rect 4362 5466 4418 5468
rect 4122 5414 4168 5466
rect 4168 5414 4178 5466
rect 4202 5414 4232 5466
rect 4232 5414 4244 5466
rect 4244 5414 4258 5466
rect 4282 5414 4296 5466
rect 4296 5414 4308 5466
rect 4308 5414 4338 5466
rect 4362 5414 4372 5466
rect 4372 5414 4418 5466
rect 4122 5412 4178 5414
rect 4202 5412 4258 5414
rect 4282 5412 4338 5414
rect 4362 5412 4418 5414
rect 4894 8744 4950 8800
rect 4894 8064 4950 8120
rect 4802 7928 4858 7984
rect 5672 11450 5728 11452
rect 5752 11450 5808 11452
rect 5832 11450 5888 11452
rect 5912 11450 5968 11452
rect 5672 11398 5718 11450
rect 5718 11398 5728 11450
rect 5752 11398 5782 11450
rect 5782 11398 5794 11450
rect 5794 11398 5808 11450
rect 5832 11398 5846 11450
rect 5846 11398 5858 11450
rect 5858 11398 5888 11450
rect 5912 11398 5922 11450
rect 5922 11398 5968 11450
rect 5672 11396 5728 11398
rect 5752 11396 5808 11398
rect 5832 11396 5888 11398
rect 5912 11396 5968 11398
rect 5262 10376 5318 10432
rect 5672 10362 5728 10364
rect 5752 10362 5808 10364
rect 5832 10362 5888 10364
rect 5912 10362 5968 10364
rect 5672 10310 5718 10362
rect 5718 10310 5728 10362
rect 5752 10310 5782 10362
rect 5782 10310 5794 10362
rect 5794 10310 5808 10362
rect 5832 10310 5846 10362
rect 5846 10310 5858 10362
rect 5858 10310 5888 10362
rect 5912 10310 5922 10362
rect 5922 10310 5968 10362
rect 5672 10308 5728 10310
rect 5752 10308 5808 10310
rect 5832 10308 5888 10310
rect 5912 10308 5968 10310
rect 6182 11192 6238 11248
rect 5446 9288 5502 9344
rect 5262 9152 5318 9208
rect 5672 9274 5728 9276
rect 5752 9274 5808 9276
rect 5832 9274 5888 9276
rect 5912 9274 5968 9276
rect 5672 9222 5718 9274
rect 5718 9222 5728 9274
rect 5752 9222 5782 9274
rect 5782 9222 5794 9274
rect 5794 9222 5808 9274
rect 5832 9222 5846 9274
rect 5846 9222 5858 9274
rect 5858 9222 5888 9274
rect 5912 9222 5922 9274
rect 5922 9222 5968 9274
rect 5672 9220 5728 9222
rect 5752 9220 5808 9222
rect 5832 9220 5888 9222
rect 5912 9220 5968 9222
rect 5630 8744 5686 8800
rect 5262 8608 5318 8664
rect 4986 7656 5042 7712
rect 4986 6976 5042 7032
rect 5262 7520 5318 7576
rect 5538 8336 5594 8392
rect 5906 8900 5962 8936
rect 5906 8880 5908 8900
rect 5908 8880 5960 8900
rect 5960 8880 5962 8900
rect 5446 8236 5448 8256
rect 5448 8236 5500 8256
rect 5500 8236 5502 8256
rect 5446 8200 5502 8236
rect 5262 6704 5318 6760
rect 5672 8186 5728 8188
rect 5752 8186 5808 8188
rect 5832 8186 5888 8188
rect 5912 8186 5968 8188
rect 5672 8134 5718 8186
rect 5718 8134 5728 8186
rect 5752 8134 5782 8186
rect 5782 8134 5794 8186
rect 5794 8134 5808 8186
rect 5832 8134 5846 8186
rect 5846 8134 5858 8186
rect 5858 8134 5888 8186
rect 5912 8134 5922 8186
rect 5922 8134 5968 8186
rect 5672 8132 5728 8134
rect 5752 8132 5808 8134
rect 5832 8132 5888 8134
rect 5912 8132 5968 8134
rect 5906 7928 5962 7984
rect 5354 6568 5410 6624
rect 4434 4664 4490 4720
rect 4158 4564 4160 4584
rect 4160 4564 4212 4584
rect 4212 4564 4214 4584
rect 4158 4528 4214 4564
rect 4122 4378 4178 4380
rect 4202 4378 4258 4380
rect 4282 4378 4338 4380
rect 4362 4378 4418 4380
rect 4122 4326 4168 4378
rect 4168 4326 4178 4378
rect 4202 4326 4232 4378
rect 4232 4326 4244 4378
rect 4244 4326 4258 4378
rect 4282 4326 4296 4378
rect 4296 4326 4308 4378
rect 4308 4326 4338 4378
rect 4362 4326 4372 4378
rect 4372 4326 4418 4378
rect 4122 4324 4178 4326
rect 4202 4324 4258 4326
rect 4282 4324 4338 4326
rect 4362 4324 4418 4326
rect 4122 3290 4178 3292
rect 4202 3290 4258 3292
rect 4282 3290 4338 3292
rect 4362 3290 4418 3292
rect 4122 3238 4168 3290
rect 4168 3238 4178 3290
rect 4202 3238 4232 3290
rect 4232 3238 4244 3290
rect 4244 3238 4258 3290
rect 4282 3238 4296 3290
rect 4296 3238 4308 3290
rect 4308 3238 4338 3290
rect 4362 3238 4372 3290
rect 4372 3238 4418 3290
rect 4122 3236 4178 3238
rect 4202 3236 4258 3238
rect 4282 3236 4338 3238
rect 4362 3236 4418 3238
rect 5672 7098 5728 7100
rect 5752 7098 5808 7100
rect 5832 7098 5888 7100
rect 5912 7098 5968 7100
rect 5672 7046 5718 7098
rect 5718 7046 5728 7098
rect 5752 7046 5782 7098
rect 5782 7046 5794 7098
rect 5794 7046 5808 7098
rect 5832 7046 5846 7098
rect 5846 7046 5858 7098
rect 5858 7046 5888 7098
rect 5912 7046 5922 7098
rect 5922 7046 5968 7098
rect 5672 7044 5728 7046
rect 5752 7044 5808 7046
rect 5832 7044 5888 7046
rect 5912 7044 5968 7046
rect 5630 6432 5686 6488
rect 6734 10124 6790 10160
rect 6734 10104 6736 10124
rect 6736 10104 6788 10124
rect 6788 10104 6790 10124
rect 6918 9696 6974 9752
rect 6734 9016 6790 9072
rect 7222 10906 7278 10908
rect 7302 10906 7358 10908
rect 7382 10906 7438 10908
rect 7462 10906 7518 10908
rect 7222 10854 7268 10906
rect 7268 10854 7278 10906
rect 7302 10854 7332 10906
rect 7332 10854 7344 10906
rect 7344 10854 7358 10906
rect 7382 10854 7396 10906
rect 7396 10854 7408 10906
rect 7408 10854 7438 10906
rect 7462 10854 7472 10906
rect 7472 10854 7518 10906
rect 7222 10852 7278 10854
rect 7302 10852 7358 10854
rect 7382 10852 7438 10854
rect 7462 10852 7518 10854
rect 7562 10104 7618 10160
rect 7222 9818 7278 9820
rect 7302 9818 7358 9820
rect 7382 9818 7438 9820
rect 7462 9818 7518 9820
rect 7222 9766 7268 9818
rect 7268 9766 7278 9818
rect 7302 9766 7332 9818
rect 7332 9766 7344 9818
rect 7344 9766 7358 9818
rect 7382 9766 7396 9818
rect 7396 9766 7408 9818
rect 7408 9766 7438 9818
rect 7462 9766 7472 9818
rect 7472 9766 7518 9818
rect 7222 9764 7278 9766
rect 7302 9764 7358 9766
rect 7382 9764 7438 9766
rect 7462 9764 7518 9766
rect 7378 9288 7434 9344
rect 6274 7656 6330 7712
rect 6274 6840 6330 6896
rect 5538 6024 5594 6080
rect 5672 6010 5728 6012
rect 5752 6010 5808 6012
rect 5832 6010 5888 6012
rect 5912 6010 5968 6012
rect 5672 5958 5718 6010
rect 5718 5958 5728 6010
rect 5752 5958 5782 6010
rect 5782 5958 5794 6010
rect 5794 5958 5808 6010
rect 5832 5958 5846 6010
rect 5846 5958 5858 6010
rect 5858 5958 5888 6010
rect 5912 5958 5922 6010
rect 5922 5958 5968 6010
rect 5672 5956 5728 5958
rect 5752 5956 5808 5958
rect 5832 5956 5888 5958
rect 5912 5956 5968 5958
rect 5672 4922 5728 4924
rect 5752 4922 5808 4924
rect 5832 4922 5888 4924
rect 5912 4922 5968 4924
rect 5672 4870 5718 4922
rect 5718 4870 5728 4922
rect 5752 4870 5782 4922
rect 5782 4870 5794 4922
rect 5794 4870 5808 4922
rect 5832 4870 5846 4922
rect 5846 4870 5858 4922
rect 5858 4870 5888 4922
rect 5912 4870 5922 4922
rect 5922 4870 5968 4922
rect 5672 4868 5728 4870
rect 5752 4868 5808 4870
rect 5832 4868 5888 4870
rect 5912 4868 5968 4870
rect 5906 4664 5962 4720
rect 5722 4548 5778 4584
rect 5722 4528 5724 4548
rect 5724 4528 5776 4548
rect 5776 4528 5778 4548
rect 5672 3834 5728 3836
rect 5752 3834 5808 3836
rect 5832 3834 5888 3836
rect 5912 3834 5968 3836
rect 5672 3782 5718 3834
rect 5718 3782 5728 3834
rect 5752 3782 5782 3834
rect 5782 3782 5794 3834
rect 5794 3782 5808 3834
rect 5832 3782 5846 3834
rect 5846 3782 5858 3834
rect 5858 3782 5888 3834
rect 5912 3782 5922 3834
rect 5922 3782 5968 3834
rect 5672 3780 5728 3782
rect 5752 3780 5808 3782
rect 5832 3780 5888 3782
rect 5912 3780 5968 3782
rect 5672 2746 5728 2748
rect 5752 2746 5808 2748
rect 5832 2746 5888 2748
rect 5912 2746 5968 2748
rect 5672 2694 5718 2746
rect 5718 2694 5728 2746
rect 5752 2694 5782 2746
rect 5782 2694 5794 2746
rect 5794 2694 5808 2746
rect 5832 2694 5846 2746
rect 5846 2694 5858 2746
rect 5858 2694 5888 2746
rect 5912 2694 5922 2746
rect 5922 2694 5968 2746
rect 5672 2692 5728 2694
rect 5752 2692 5808 2694
rect 5832 2692 5888 2694
rect 5912 2692 5968 2694
rect 6826 8744 6882 8800
rect 6642 8472 6698 8528
rect 7222 8730 7278 8732
rect 7302 8730 7358 8732
rect 7382 8730 7438 8732
rect 7462 8730 7518 8732
rect 7222 8678 7268 8730
rect 7268 8678 7278 8730
rect 7302 8678 7332 8730
rect 7332 8678 7344 8730
rect 7344 8678 7358 8730
rect 7382 8678 7396 8730
rect 7396 8678 7408 8730
rect 7408 8678 7438 8730
rect 7462 8678 7472 8730
rect 7472 8678 7518 8730
rect 7222 8676 7278 8678
rect 7302 8676 7358 8678
rect 7382 8676 7438 8678
rect 7462 8676 7518 8678
rect 6918 8608 6974 8664
rect 6918 7520 6974 7576
rect 7222 7642 7278 7644
rect 7302 7642 7358 7644
rect 7382 7642 7438 7644
rect 7462 7642 7518 7644
rect 7222 7590 7268 7642
rect 7268 7590 7278 7642
rect 7302 7590 7332 7642
rect 7332 7590 7344 7642
rect 7344 7590 7358 7642
rect 7382 7590 7396 7642
rect 7396 7590 7408 7642
rect 7408 7590 7438 7642
rect 7462 7590 7472 7642
rect 7472 7590 7518 7642
rect 7222 7588 7278 7590
rect 7302 7588 7358 7590
rect 7382 7588 7438 7590
rect 7462 7588 7518 7590
rect 7010 6704 7066 6760
rect 7010 6432 7066 6488
rect 16762 12824 16818 12880
rect 8114 11056 8170 11112
rect 8022 10648 8078 10704
rect 7838 10140 7840 10160
rect 7840 10140 7892 10160
rect 7892 10140 7894 10160
rect 7838 10104 7894 10140
rect 7838 9968 7894 10024
rect 8022 9968 8078 10024
rect 8298 10648 8354 10704
rect 8298 9288 8354 9344
rect 13450 11464 13506 11520
rect 8772 11450 8828 11452
rect 8852 11450 8908 11452
rect 8932 11450 8988 11452
rect 9012 11450 9068 11452
rect 8772 11398 8818 11450
rect 8818 11398 8828 11450
rect 8852 11398 8882 11450
rect 8882 11398 8894 11450
rect 8894 11398 8908 11450
rect 8932 11398 8946 11450
rect 8946 11398 8958 11450
rect 8958 11398 8988 11450
rect 9012 11398 9022 11450
rect 9022 11398 9068 11450
rect 8772 11396 8828 11398
rect 8852 11396 8908 11398
rect 8932 11396 8988 11398
rect 9012 11396 9068 11398
rect 8772 10362 8828 10364
rect 8852 10362 8908 10364
rect 8932 10362 8988 10364
rect 9012 10362 9068 10364
rect 8772 10310 8818 10362
rect 8818 10310 8828 10362
rect 8852 10310 8882 10362
rect 8882 10310 8894 10362
rect 8894 10310 8908 10362
rect 8932 10310 8946 10362
rect 8946 10310 8958 10362
rect 8958 10310 8988 10362
rect 9012 10310 9022 10362
rect 9022 10310 9068 10362
rect 8772 10308 8828 10310
rect 8852 10308 8908 10310
rect 8932 10308 8988 10310
rect 9012 10308 9068 10310
rect 8574 9424 8630 9480
rect 7222 6554 7278 6556
rect 7302 6554 7358 6556
rect 7382 6554 7438 6556
rect 7462 6554 7518 6556
rect 7222 6502 7268 6554
rect 7268 6502 7278 6554
rect 7302 6502 7332 6554
rect 7332 6502 7344 6554
rect 7344 6502 7358 6554
rect 7382 6502 7396 6554
rect 7396 6502 7408 6554
rect 7408 6502 7438 6554
rect 7462 6502 7472 6554
rect 7472 6502 7518 6554
rect 7222 6500 7278 6502
rect 7302 6500 7358 6502
rect 7382 6500 7438 6502
rect 7462 6500 7518 6502
rect 7286 6296 7342 6352
rect 7470 6316 7526 6352
rect 7470 6296 7472 6316
rect 7472 6296 7524 6316
rect 7524 6296 7526 6316
rect 7222 5466 7278 5468
rect 7302 5466 7358 5468
rect 7382 5466 7438 5468
rect 7462 5466 7518 5468
rect 7222 5414 7268 5466
rect 7268 5414 7278 5466
rect 7302 5414 7332 5466
rect 7332 5414 7344 5466
rect 7344 5414 7358 5466
rect 7382 5414 7396 5466
rect 7396 5414 7408 5466
rect 7408 5414 7438 5466
rect 7462 5414 7472 5466
rect 7472 5414 7518 5466
rect 7222 5412 7278 5414
rect 7302 5412 7358 5414
rect 7382 5412 7438 5414
rect 7462 5412 7518 5414
rect 7746 5752 7802 5808
rect 8772 9274 8828 9276
rect 8852 9274 8908 9276
rect 8932 9274 8988 9276
rect 9012 9274 9068 9276
rect 8772 9222 8818 9274
rect 8818 9222 8828 9274
rect 8852 9222 8882 9274
rect 8882 9222 8894 9274
rect 8894 9222 8908 9274
rect 8932 9222 8946 9274
rect 8946 9222 8958 9274
rect 8958 9222 8988 9274
rect 9012 9222 9022 9274
rect 9022 9222 9068 9274
rect 8772 9220 8828 9222
rect 8852 9220 8908 9222
rect 8932 9220 8988 9222
rect 9012 9220 9068 9222
rect 8390 7928 8446 7984
rect 8772 8186 8828 8188
rect 8852 8186 8908 8188
rect 8932 8186 8988 8188
rect 9012 8186 9068 8188
rect 8772 8134 8818 8186
rect 8818 8134 8828 8186
rect 8852 8134 8882 8186
rect 8882 8134 8894 8186
rect 8894 8134 8908 8186
rect 8932 8134 8946 8186
rect 8946 8134 8958 8186
rect 8958 8134 8988 8186
rect 9012 8134 9022 8186
rect 9022 8134 9068 8186
rect 8772 8132 8828 8134
rect 8852 8132 8908 8134
rect 8932 8132 8988 8134
rect 9012 8132 9068 8134
rect 9494 10920 9550 10976
rect 13726 11192 13782 11248
rect 13450 10512 13506 10568
rect 9678 10240 9734 10296
rect 9402 9288 9458 9344
rect 13634 9968 13690 10024
rect 9586 8200 9642 8256
rect 13542 9016 13598 9072
rect 13450 8900 13506 8936
rect 13450 8880 13452 8900
rect 13452 8880 13504 8900
rect 13504 8880 13506 8900
rect 13634 8608 13690 8664
rect 9310 7948 9366 7984
rect 9310 7928 9312 7948
rect 9312 7928 9364 7948
rect 9364 7928 9366 7948
rect 10138 7928 10194 7984
rect 8022 6296 8078 6352
rect 7222 4378 7278 4380
rect 7302 4378 7358 4380
rect 7382 4378 7438 4380
rect 7462 4378 7518 4380
rect 7222 4326 7268 4378
rect 7268 4326 7278 4378
rect 7302 4326 7332 4378
rect 7332 4326 7344 4378
rect 7344 4326 7358 4378
rect 7382 4326 7396 4378
rect 7396 4326 7408 4378
rect 7408 4326 7438 4378
rect 7462 4326 7472 4378
rect 7472 4326 7518 4378
rect 7222 4324 7278 4326
rect 7302 4324 7358 4326
rect 7382 4324 7438 4326
rect 7462 4324 7518 4326
rect 6274 3032 6330 3088
rect 7222 3290 7278 3292
rect 7302 3290 7358 3292
rect 7382 3290 7438 3292
rect 7462 3290 7518 3292
rect 7222 3238 7268 3290
rect 7268 3238 7278 3290
rect 7302 3238 7332 3290
rect 7332 3238 7344 3290
rect 7344 3238 7358 3290
rect 7382 3238 7396 3290
rect 7396 3238 7408 3290
rect 7408 3238 7438 3290
rect 7462 3238 7472 3290
rect 7472 3238 7518 3290
rect 7222 3236 7278 3238
rect 7302 3236 7358 3238
rect 7382 3236 7438 3238
rect 7462 3236 7518 3238
rect 7470 2796 7472 2816
rect 7472 2796 7524 2816
rect 7524 2796 7526 2816
rect 7470 2760 7526 2796
rect 8666 7248 8722 7304
rect 8772 7098 8828 7100
rect 8852 7098 8908 7100
rect 8932 7098 8988 7100
rect 9012 7098 9068 7100
rect 8772 7046 8818 7098
rect 8818 7046 8828 7098
rect 8852 7046 8882 7098
rect 8882 7046 8894 7098
rect 8894 7046 8908 7098
rect 8932 7046 8946 7098
rect 8946 7046 8958 7098
rect 8958 7046 8988 7098
rect 9012 7046 9022 7098
rect 9022 7046 9068 7098
rect 8772 7044 8828 7046
rect 8852 7044 8908 7046
rect 8932 7044 8988 7046
rect 9012 7044 9068 7046
rect 8666 6160 8722 6216
rect 8772 6010 8828 6012
rect 8852 6010 8908 6012
rect 8932 6010 8988 6012
rect 9012 6010 9068 6012
rect 8772 5958 8818 6010
rect 8818 5958 8828 6010
rect 8852 5958 8882 6010
rect 8882 5958 8894 6010
rect 8894 5958 8908 6010
rect 8932 5958 8946 6010
rect 8946 5958 8958 6010
rect 8958 5958 8988 6010
rect 9012 5958 9022 6010
rect 9022 5958 9068 6010
rect 8772 5956 8828 5958
rect 8852 5956 8908 5958
rect 8932 5956 8988 5958
rect 9012 5956 9068 5958
rect 8850 5072 8906 5128
rect 8772 4922 8828 4924
rect 8852 4922 8908 4924
rect 8932 4922 8988 4924
rect 9012 4922 9068 4924
rect 8772 4870 8818 4922
rect 8818 4870 8828 4922
rect 8852 4870 8882 4922
rect 8882 4870 8894 4922
rect 8894 4870 8908 4922
rect 8932 4870 8946 4922
rect 8946 4870 8958 4922
rect 8958 4870 8988 4922
rect 9012 4870 9022 4922
rect 9022 4870 9068 4922
rect 8772 4868 8828 4870
rect 8852 4868 8908 4870
rect 8932 4868 8988 4870
rect 9012 4868 9068 4870
rect 8758 4664 8814 4720
rect 8298 2760 8354 2816
rect 8772 3834 8828 3836
rect 8852 3834 8908 3836
rect 8932 3834 8988 3836
rect 9012 3834 9068 3836
rect 8772 3782 8818 3834
rect 8818 3782 8828 3834
rect 8852 3782 8882 3834
rect 8882 3782 8894 3834
rect 8894 3782 8908 3834
rect 8932 3782 8946 3834
rect 8946 3782 8958 3834
rect 8958 3782 8988 3834
rect 9012 3782 9022 3834
rect 9022 3782 9068 3834
rect 8772 3780 8828 3782
rect 8852 3780 8908 3782
rect 8932 3780 8988 3782
rect 9012 3780 9068 3782
rect 13450 7676 13506 7712
rect 13450 7656 13452 7676
rect 13452 7656 13504 7676
rect 13504 7656 13506 7676
rect 13542 7248 13598 7304
rect 13818 9832 13874 9888
rect 13818 9560 13874 9616
rect 13818 7792 13874 7848
rect 13818 7384 13874 7440
rect 13634 6976 13690 7032
rect 12806 6024 12862 6080
rect 10874 4936 10930 4992
rect 9678 4664 9734 4720
rect 8772 2746 8828 2748
rect 8852 2746 8908 2748
rect 8932 2746 8988 2748
rect 9012 2746 9068 2748
rect 8772 2694 8818 2746
rect 8818 2694 8828 2746
rect 8852 2694 8882 2746
rect 8882 2694 8894 2746
rect 8894 2694 8908 2746
rect 8932 2694 8946 2746
rect 8946 2694 8958 2746
rect 8958 2694 8988 2746
rect 9012 2694 9022 2746
rect 9022 2694 9068 2746
rect 8772 2692 8828 2694
rect 8852 2692 8908 2694
rect 8932 2692 8988 2694
rect 9012 2692 9068 2694
rect 13818 6568 13874 6624
rect 13726 6296 13782 6352
rect 13634 3712 13690 3768
rect 13818 4392 13874 4448
rect 13726 3304 13782 3360
rect 19430 2352 19486 2408
rect 4122 2202 4178 2204
rect 4202 2202 4258 2204
rect 4282 2202 4338 2204
rect 4362 2202 4418 2204
rect 4122 2150 4168 2202
rect 4168 2150 4178 2202
rect 4202 2150 4232 2202
rect 4232 2150 4244 2202
rect 4244 2150 4258 2202
rect 4282 2150 4296 2202
rect 4296 2150 4308 2202
rect 4308 2150 4338 2202
rect 4362 2150 4372 2202
rect 4372 2150 4418 2202
rect 4122 2148 4178 2150
rect 4202 2148 4258 2150
rect 4282 2148 4338 2150
rect 4362 2148 4418 2150
rect 7222 2202 7278 2204
rect 7302 2202 7358 2204
rect 7382 2202 7438 2204
rect 7462 2202 7518 2204
rect 7222 2150 7268 2202
rect 7268 2150 7278 2202
rect 7302 2150 7332 2202
rect 7332 2150 7344 2202
rect 7344 2150 7358 2202
rect 7382 2150 7396 2202
rect 7396 2150 7408 2202
rect 7408 2150 7438 2202
rect 7462 2150 7472 2202
rect 7472 2150 7518 2202
rect 7222 2148 7278 2150
rect 7302 2148 7358 2150
rect 7382 2148 7438 2150
rect 7462 2148 7518 2150
rect 22282 720 22338 776
rect 3514 448 3570 504
rect 22374 176 22430 232
<< metal3 >>
rect 14000 13832 34000 13864
rect 14000 13776 16578 13832
rect 16634 13776 34000 13832
rect 14000 13744 34000 13776
rect 14000 13562 34000 13592
rect 6870 13502 34000 13562
rect 2405 13426 2471 13429
rect 6870 13426 6930 13502
rect 14000 13472 34000 13502
rect 2405 13424 6930 13426
rect 2405 13368 2410 13424
rect 2466 13368 6930 13424
rect 2405 13366 6930 13368
rect 2405 13363 2471 13366
rect 6085 13154 6151 13157
rect 14000 13154 34000 13184
rect 6085 13152 34000 13154
rect 6085 13096 6090 13152
rect 6146 13096 34000 13152
rect 6085 13094 34000 13096
rect 6085 13091 6151 13094
rect 14000 13064 34000 13094
rect 14000 12880 34000 12912
rect 14000 12824 16762 12880
rect 16818 12824 34000 12880
rect 14000 12792 34000 12824
rect 14000 12610 34000 12640
rect 6870 12550 34000 12610
rect 2313 12474 2379 12477
rect 6870 12474 6930 12550
rect 14000 12520 34000 12550
rect 2313 12472 6930 12474
rect 2313 12416 2318 12472
rect 2374 12416 6930 12472
rect 2313 12414 6930 12416
rect 2313 12411 2379 12414
rect 5993 12202 6059 12205
rect 14000 12202 34000 12232
rect 5993 12200 34000 12202
rect 5993 12144 5998 12200
rect 6054 12144 34000 12200
rect 5993 12142 34000 12144
rect 5993 12139 6059 12142
rect 14000 12112 34000 12142
rect 3141 11930 3207 11933
rect 14000 11930 34000 11960
rect 3141 11928 34000 11930
rect 3141 11872 3146 11928
rect 3202 11872 34000 11928
rect 3141 11870 34000 11872
rect 3141 11867 3207 11870
rect 14000 11840 34000 11870
rect 13445 11522 13511 11525
rect 14000 11522 34000 11552
rect 13445 11520 34000 11522
rect 13445 11464 13450 11520
rect 13506 11464 34000 11520
rect 13445 11462 34000 11464
rect 13445 11459 13511 11462
rect 2560 11456 2880 11457
rect 2560 11392 2568 11456
rect 2632 11392 2648 11456
rect 2712 11392 2728 11456
rect 2792 11392 2808 11456
rect 2872 11392 2880 11456
rect 2560 11391 2880 11392
rect 5660 11456 5980 11457
rect 5660 11392 5668 11456
rect 5732 11392 5748 11456
rect 5812 11392 5828 11456
rect 5892 11392 5908 11456
rect 5972 11392 5980 11456
rect 5660 11391 5980 11392
rect 8760 11456 9080 11457
rect 8760 11392 8768 11456
rect 8832 11392 8848 11456
rect 8912 11392 8928 11456
rect 8992 11392 9008 11456
rect 9072 11392 9080 11456
rect 14000 11432 34000 11462
rect 8760 11391 9080 11392
rect 2957 11386 3023 11389
rect 2957 11384 4906 11386
rect 2957 11328 2962 11384
rect 3018 11328 4906 11384
rect 2957 11326 4906 11328
rect 2957 11323 3023 11326
rect 3509 11250 3575 11253
rect 4337 11250 4403 11253
rect 4705 11250 4771 11253
rect 3509 11248 4771 11250
rect 3509 11192 3514 11248
rect 3570 11192 4342 11248
rect 4398 11192 4710 11248
rect 4766 11192 4771 11248
rect 3509 11190 4771 11192
rect 4846 11250 4906 11326
rect 6177 11250 6243 11253
rect 4846 11248 6243 11250
rect 4846 11192 6182 11248
rect 6238 11192 6243 11248
rect 4846 11190 6243 11192
rect 3509 11187 3575 11190
rect 4337 11187 4403 11190
rect 4705 11187 4771 11190
rect 6177 11187 6243 11190
rect 13721 11250 13787 11253
rect 14000 11250 34000 11280
rect 13721 11248 34000 11250
rect 13721 11192 13726 11248
rect 13782 11192 34000 11248
rect 13721 11190 34000 11192
rect 13721 11187 13787 11190
rect 14000 11160 34000 11190
rect 3049 11114 3115 11117
rect 8109 11114 8175 11117
rect 3049 11112 8175 11114
rect 3049 11056 3054 11112
rect 3110 11056 8114 11112
rect 8170 11056 8175 11112
rect 3049 11054 8175 11056
rect 3049 11051 3115 11054
rect 8109 11051 8175 11054
rect 9489 10978 9555 10981
rect 14000 10978 34000 11008
rect 9489 10976 34000 10978
rect 9489 10920 9494 10976
rect 9550 10920 34000 10976
rect 9489 10918 34000 10920
rect 9489 10915 9555 10918
rect 4110 10912 4430 10913
rect 4110 10848 4118 10912
rect 4182 10848 4198 10912
rect 4262 10848 4278 10912
rect 4342 10848 4358 10912
rect 4422 10848 4430 10912
rect 4110 10847 4430 10848
rect 7210 10912 7530 10913
rect 7210 10848 7218 10912
rect 7282 10848 7298 10912
rect 7362 10848 7378 10912
rect 7442 10848 7458 10912
rect 7522 10848 7530 10912
rect 14000 10888 34000 10918
rect 7210 10847 7530 10848
rect 2221 10842 2287 10845
rect 3877 10842 3943 10845
rect 2221 10840 3943 10842
rect 2221 10784 2226 10840
rect 2282 10784 3882 10840
rect 3938 10784 3943 10840
rect 2221 10782 3943 10784
rect 2221 10779 2287 10782
rect 3877 10779 3943 10782
rect 3325 10706 3391 10709
rect 8017 10706 8083 10709
rect 3325 10704 8083 10706
rect 3325 10648 3330 10704
rect 3386 10648 8022 10704
rect 8078 10648 8083 10704
rect 3325 10646 8083 10648
rect 3325 10643 3391 10646
rect 8017 10643 8083 10646
rect 8293 10706 8359 10709
rect 8293 10704 13922 10706
rect 8293 10648 8298 10704
rect 8354 10648 13922 10704
rect 8293 10646 13922 10648
rect 8293 10643 8359 10646
rect 1485 10570 1551 10573
rect 13445 10570 13511 10573
rect 1485 10568 13511 10570
rect 1485 10512 1490 10568
rect 1546 10512 13450 10568
rect 13506 10512 13511 10568
rect 1485 10510 13511 10512
rect 13862 10570 13922 10646
rect 14000 10570 34000 10600
rect 13862 10510 34000 10570
rect 1485 10507 1551 10510
rect 13445 10507 13511 10510
rect 14000 10480 34000 10510
rect 3509 10434 3575 10437
rect 5257 10434 5323 10437
rect 3509 10432 5323 10434
rect 3509 10376 3514 10432
rect 3570 10376 5262 10432
rect 5318 10376 5323 10432
rect 3509 10374 5323 10376
rect 3509 10371 3575 10374
rect 5257 10371 5323 10374
rect 2560 10368 2880 10369
rect 2560 10304 2568 10368
rect 2632 10304 2648 10368
rect 2712 10304 2728 10368
rect 2792 10304 2808 10368
rect 2872 10304 2880 10368
rect 2560 10303 2880 10304
rect 5660 10368 5980 10369
rect 5660 10304 5668 10368
rect 5732 10304 5748 10368
rect 5812 10304 5828 10368
rect 5892 10304 5908 10368
rect 5972 10304 5980 10368
rect 5660 10303 5980 10304
rect 8760 10368 9080 10369
rect 8760 10304 8768 10368
rect 8832 10304 8848 10368
rect 8912 10304 8928 10368
rect 8992 10304 9008 10368
rect 9072 10304 9080 10368
rect 8760 10303 9080 10304
rect 4889 10298 4955 10301
rect 2960 10296 4955 10298
rect 2960 10240 4894 10296
rect 4950 10240 4955 10296
rect 2960 10238 4955 10240
rect 2313 10162 2379 10165
rect 2960 10162 3020 10238
rect 4889 10235 4955 10238
rect 9673 10298 9739 10301
rect 14000 10298 34000 10328
rect 9673 10296 34000 10298
rect 9673 10240 9678 10296
rect 9734 10240 34000 10296
rect 9673 10238 34000 10240
rect 9673 10235 9739 10238
rect 14000 10208 34000 10238
rect 2313 10160 3020 10162
rect 2313 10104 2318 10160
rect 2374 10104 3020 10160
rect 2313 10102 3020 10104
rect 3601 10162 3667 10165
rect 6729 10162 6795 10165
rect 3601 10160 6795 10162
rect 3601 10104 3606 10160
rect 3662 10104 6734 10160
rect 6790 10104 6795 10160
rect 3601 10102 6795 10104
rect 2313 10099 2379 10102
rect 3601 10099 3667 10102
rect 6729 10099 6795 10102
rect 7557 10162 7623 10165
rect 7833 10162 7899 10165
rect 7557 10160 7899 10162
rect 7557 10104 7562 10160
rect 7618 10104 7838 10160
rect 7894 10104 7899 10160
rect 7557 10102 7899 10104
rect 7557 10099 7623 10102
rect 7833 10099 7899 10102
rect 3509 10026 3575 10029
rect 7833 10026 7899 10029
rect 3509 10024 7899 10026
rect 3509 9968 3514 10024
rect 3570 9968 7838 10024
rect 7894 9968 7899 10024
rect 3509 9966 7899 9968
rect 3509 9963 3575 9966
rect 7833 9963 7899 9966
rect 8017 10026 8083 10029
rect 13629 10026 13695 10029
rect 8017 10024 13695 10026
rect 8017 9968 8022 10024
rect 8078 9968 13634 10024
rect 13690 9968 13695 10024
rect 8017 9966 13695 9968
rect 8017 9963 8083 9966
rect 13629 9963 13695 9966
rect 2773 9890 2839 9893
rect 3785 9890 3851 9893
rect 2773 9888 3851 9890
rect 2773 9832 2778 9888
rect 2834 9832 3790 9888
rect 3846 9832 3851 9888
rect 2773 9830 3851 9832
rect 2773 9827 2839 9830
rect 3785 9827 3851 9830
rect 13813 9890 13879 9893
rect 14000 9890 34000 9920
rect 13813 9888 34000 9890
rect 13813 9832 13818 9888
rect 13874 9832 34000 9888
rect 13813 9830 34000 9832
rect 13813 9827 13879 9830
rect 4110 9824 4430 9825
rect 4110 9760 4118 9824
rect 4182 9760 4198 9824
rect 4262 9760 4278 9824
rect 4342 9760 4358 9824
rect 4422 9760 4430 9824
rect 4110 9759 4430 9760
rect 7210 9824 7530 9825
rect 7210 9760 7218 9824
rect 7282 9760 7298 9824
rect 7362 9760 7378 9824
rect 7442 9760 7458 9824
rect 7522 9760 7530 9824
rect 14000 9800 34000 9830
rect 7210 9759 7530 9760
rect 4521 9754 4587 9757
rect 6913 9754 6979 9757
rect 4521 9752 6979 9754
rect 4521 9696 4526 9752
rect 4582 9696 6918 9752
rect 6974 9696 6979 9752
rect 4521 9694 6979 9696
rect 4521 9691 4587 9694
rect 6913 9691 6979 9694
rect 1669 9618 1735 9621
rect 13813 9618 13879 9621
rect 14000 9618 34000 9648
rect 1669 9616 9322 9618
rect 1669 9560 1674 9616
rect 1730 9560 9322 9616
rect 1669 9558 9322 9560
rect 1669 9555 1735 9558
rect 1853 9482 1919 9485
rect 3785 9482 3851 9485
rect 8569 9482 8635 9485
rect 1853 9480 3618 9482
rect 1853 9424 1858 9480
rect 1914 9424 3618 9480
rect 1853 9422 3618 9424
rect 1853 9419 1919 9422
rect 3558 9346 3618 9422
rect 3785 9480 8635 9482
rect 3785 9424 3790 9480
rect 3846 9424 8574 9480
rect 8630 9424 8635 9480
rect 3785 9422 8635 9424
rect 3785 9419 3851 9422
rect 8569 9419 8635 9422
rect 5441 9346 5507 9349
rect 3558 9344 5507 9346
rect 3558 9288 5446 9344
rect 5502 9288 5507 9344
rect 3558 9286 5507 9288
rect 5441 9283 5507 9286
rect 7373 9346 7439 9349
rect 8293 9346 8359 9349
rect 7373 9344 8359 9346
rect 7373 9288 7378 9344
rect 7434 9288 8298 9344
rect 8354 9288 8359 9344
rect 7373 9286 8359 9288
rect 7373 9283 7439 9286
rect 8293 9283 8359 9286
rect 2560 9280 2880 9281
rect 2560 9216 2568 9280
rect 2632 9216 2648 9280
rect 2712 9216 2728 9280
rect 2792 9216 2808 9280
rect 2872 9216 2880 9280
rect 2560 9215 2880 9216
rect 5660 9280 5980 9281
rect 5660 9216 5668 9280
rect 5732 9216 5748 9280
rect 5812 9216 5828 9280
rect 5892 9216 5908 9280
rect 5972 9216 5980 9280
rect 5660 9215 5980 9216
rect 8760 9280 9080 9281
rect 8760 9216 8768 9280
rect 8832 9216 8848 9280
rect 8912 9216 8928 9280
rect 8992 9216 9008 9280
rect 9072 9216 9080 9280
rect 8760 9215 9080 9216
rect 2957 9210 3023 9213
rect 5257 9210 5323 9213
rect 2957 9208 5323 9210
rect 2957 9152 2962 9208
rect 3018 9152 5262 9208
rect 5318 9152 5323 9208
rect 2957 9150 5323 9152
rect 9262 9210 9322 9558
rect 13813 9616 34000 9618
rect 13813 9560 13818 9616
rect 13874 9560 34000 9616
rect 13813 9558 34000 9560
rect 13813 9555 13879 9558
rect 14000 9528 34000 9558
rect 9397 9346 9463 9349
rect 14000 9346 34000 9376
rect 9397 9344 34000 9346
rect 9397 9288 9402 9344
rect 9458 9288 34000 9344
rect 9397 9286 34000 9288
rect 9397 9283 9463 9286
rect 14000 9256 34000 9286
rect 9262 9150 12450 9210
rect 2957 9147 3023 9150
rect 5257 9147 5323 9150
rect 2037 9074 2103 9077
rect 6729 9074 6795 9077
rect 2037 9072 6795 9074
rect 2037 9016 2042 9072
rect 2098 9016 6734 9072
rect 6790 9016 6795 9072
rect 2037 9014 6795 9016
rect 2037 9011 2103 9014
rect 6729 9011 6795 9014
rect 2405 8938 2471 8941
rect 3693 8938 3759 8941
rect 5901 8938 5967 8941
rect 2405 8936 3759 8938
rect 2405 8880 2410 8936
rect 2466 8880 3698 8936
rect 3754 8880 3759 8936
rect 2405 8878 3759 8880
rect 2405 8875 2471 8878
rect 3693 8875 3759 8878
rect 3880 8936 5967 8938
rect 3880 8880 5906 8936
rect 5962 8880 5967 8936
rect 3880 8878 5967 8880
rect 12390 8938 12450 9150
rect 13537 9074 13603 9077
rect 13537 9072 13922 9074
rect 13537 9016 13542 9072
rect 13598 9016 13922 9072
rect 13537 9014 13922 9016
rect 13537 9011 13603 9014
rect 13445 8938 13511 8941
rect 12390 8936 13511 8938
rect 12390 8880 13450 8936
rect 13506 8880 13511 8936
rect 12390 8878 13511 8880
rect 13862 8938 13922 9014
rect 14000 8938 34000 8968
rect 13862 8878 34000 8938
rect 3880 8805 3940 8878
rect 5901 8875 5967 8878
rect 13445 8875 13511 8878
rect 14000 8848 34000 8878
rect 1301 8802 1367 8805
rect 3141 8802 3207 8805
rect 1301 8800 3207 8802
rect 1301 8744 1306 8800
rect 1362 8744 3146 8800
rect 3202 8744 3207 8800
rect 1301 8742 3207 8744
rect 1301 8739 1367 8742
rect 3141 8739 3207 8742
rect 3877 8800 3943 8805
rect 3877 8744 3882 8800
rect 3938 8744 3943 8800
rect 3877 8739 3943 8744
rect 4613 8802 4679 8805
rect 4889 8802 4955 8805
rect 4613 8800 4955 8802
rect 4613 8744 4618 8800
rect 4674 8744 4894 8800
rect 4950 8744 4955 8800
rect 4613 8742 4955 8744
rect 4613 8739 4679 8742
rect 4889 8739 4955 8742
rect 5625 8802 5691 8805
rect 6821 8802 6887 8805
rect 5625 8800 6887 8802
rect 5625 8744 5630 8800
rect 5686 8744 6826 8800
rect 6882 8744 6887 8800
rect 5625 8742 6887 8744
rect 5625 8739 5691 8742
rect 6821 8739 6887 8742
rect 4110 8736 4430 8737
rect 4110 8672 4118 8736
rect 4182 8672 4198 8736
rect 4262 8672 4278 8736
rect 4342 8672 4358 8736
rect 4422 8672 4430 8736
rect 4110 8671 4430 8672
rect 7210 8736 7530 8737
rect 7210 8672 7218 8736
rect 7282 8672 7298 8736
rect 7362 8672 7378 8736
rect 7442 8672 7458 8736
rect 7522 8672 7530 8736
rect 7210 8671 7530 8672
rect 5257 8666 5323 8669
rect 6913 8666 6979 8669
rect 5257 8664 6979 8666
rect 5257 8608 5262 8664
rect 5318 8608 6918 8664
rect 6974 8608 6979 8664
rect 5257 8606 6979 8608
rect 5257 8603 5323 8606
rect 6913 8603 6979 8606
rect 13629 8666 13695 8669
rect 14000 8666 34000 8696
rect 13629 8664 34000 8666
rect 13629 8608 13634 8664
rect 13690 8608 34000 8664
rect 13629 8606 34000 8608
rect 13629 8603 13695 8606
rect 14000 8576 34000 8606
rect 1485 8530 1551 8533
rect 6637 8530 6703 8533
rect 1485 8528 6703 8530
rect 1485 8472 1490 8528
rect 1546 8472 6642 8528
rect 6698 8472 6703 8528
rect 1485 8470 6703 8472
rect 1485 8467 1551 8470
rect 6637 8467 6703 8470
rect 1761 8394 1827 8397
rect 5533 8394 5599 8397
rect 1761 8392 5599 8394
rect 1761 8336 1766 8392
rect 1822 8336 5538 8392
rect 5594 8336 5599 8392
rect 1761 8334 5599 8336
rect 1761 8331 1827 8334
rect 5533 8331 5599 8334
rect 3049 8258 3115 8261
rect 5441 8258 5507 8261
rect 3049 8256 5507 8258
rect 3049 8200 3054 8256
rect 3110 8200 5446 8256
rect 5502 8200 5507 8256
rect 3049 8198 5507 8200
rect 3049 8195 3115 8198
rect 5441 8195 5507 8198
rect 9581 8258 9647 8261
rect 14000 8258 34000 8288
rect 9581 8256 34000 8258
rect 9581 8200 9586 8256
rect 9642 8200 34000 8256
rect 9581 8198 34000 8200
rect 9581 8195 9647 8198
rect 2560 8192 2880 8193
rect 2560 8128 2568 8192
rect 2632 8128 2648 8192
rect 2712 8128 2728 8192
rect 2792 8128 2808 8192
rect 2872 8128 2880 8192
rect 2560 8127 2880 8128
rect 5660 8192 5980 8193
rect 5660 8128 5668 8192
rect 5732 8128 5748 8192
rect 5812 8128 5828 8192
rect 5892 8128 5908 8192
rect 5972 8128 5980 8192
rect 5660 8127 5980 8128
rect 8760 8192 9080 8193
rect 8760 8128 8768 8192
rect 8832 8128 8848 8192
rect 8912 8128 8928 8192
rect 8992 8128 9008 8192
rect 9072 8128 9080 8192
rect 14000 8168 34000 8198
rect 8760 8127 9080 8128
rect 3693 8122 3759 8125
rect 4889 8122 4955 8125
rect 3693 8120 4955 8122
rect 3693 8064 3698 8120
rect 3754 8064 4894 8120
rect 4950 8064 4955 8120
rect 3693 8062 4955 8064
rect 3693 8059 3759 8062
rect 4889 8059 4955 8062
rect 2313 7986 2379 7989
rect 3601 7986 3667 7989
rect 2313 7984 3667 7986
rect 2313 7928 2318 7984
rect 2374 7928 3606 7984
rect 3662 7928 3667 7984
rect 2313 7926 3667 7928
rect 2313 7923 2379 7926
rect 3601 7923 3667 7926
rect 3969 7986 4035 7989
rect 4797 7986 4863 7989
rect 3969 7984 4863 7986
rect 3969 7928 3974 7984
rect 4030 7928 4802 7984
rect 4858 7928 4863 7984
rect 3969 7926 4863 7928
rect 3969 7923 4035 7926
rect 4797 7923 4863 7926
rect 5901 7986 5967 7989
rect 8385 7986 8451 7989
rect 9305 7986 9371 7989
rect 5901 7984 9371 7986
rect 5901 7928 5906 7984
rect 5962 7928 8390 7984
rect 8446 7928 9310 7984
rect 9366 7928 9371 7984
rect 5901 7926 9371 7928
rect 5901 7923 5967 7926
rect 8385 7923 8451 7926
rect 9305 7923 9371 7926
rect 10133 7986 10199 7989
rect 14000 7986 34000 8016
rect 10133 7984 34000 7986
rect 10133 7928 10138 7984
rect 10194 7928 34000 7984
rect 10133 7926 34000 7928
rect 10133 7923 10199 7926
rect 14000 7896 34000 7926
rect 2129 7850 2195 7853
rect 13813 7850 13879 7853
rect 2129 7848 12450 7850
rect 2129 7792 2134 7848
rect 2190 7792 12450 7848
rect 2129 7790 12450 7792
rect 2129 7787 2195 7790
rect 2773 7714 2839 7717
rect 3785 7714 3851 7717
rect 2773 7712 3851 7714
rect 2773 7656 2778 7712
rect 2834 7656 3790 7712
rect 3846 7656 3851 7712
rect 2773 7654 3851 7656
rect 2773 7651 2839 7654
rect 3785 7651 3851 7654
rect 4981 7714 5047 7717
rect 6269 7714 6335 7717
rect 4981 7712 6335 7714
rect 4981 7656 4986 7712
rect 5042 7656 6274 7712
rect 6330 7656 6335 7712
rect 4981 7654 6335 7656
rect 12390 7714 12450 7790
rect 13813 7848 13922 7850
rect 13813 7792 13818 7848
rect 13874 7792 13922 7848
rect 13813 7787 13922 7792
rect 13445 7714 13511 7717
rect 12390 7712 13511 7714
rect 12390 7656 13450 7712
rect 13506 7656 13511 7712
rect 12390 7654 13511 7656
rect 13862 7714 13922 7787
rect 14000 7714 34000 7744
rect 13862 7654 34000 7714
rect 4981 7651 5047 7654
rect 6269 7651 6335 7654
rect 13445 7651 13511 7654
rect 4110 7648 4430 7649
rect 4110 7584 4118 7648
rect 4182 7584 4198 7648
rect 4262 7584 4278 7648
rect 4342 7584 4358 7648
rect 4422 7584 4430 7648
rect 4110 7583 4430 7584
rect 7210 7648 7530 7649
rect 7210 7584 7218 7648
rect 7282 7584 7298 7648
rect 7362 7584 7378 7648
rect 7442 7584 7458 7648
rect 7522 7584 7530 7648
rect 14000 7624 34000 7654
rect 7210 7583 7530 7584
rect 1669 7578 1735 7581
rect 2865 7578 2931 7581
rect 3049 7578 3115 7581
rect 1669 7576 2790 7578
rect 1669 7520 1674 7576
rect 1730 7520 2790 7576
rect 1669 7518 2790 7520
rect 1669 7515 1735 7518
rect 2730 7442 2790 7518
rect 2865 7576 3115 7578
rect 2865 7520 2870 7576
rect 2926 7520 3054 7576
rect 3110 7520 3115 7576
rect 2865 7518 3115 7520
rect 2865 7515 2931 7518
rect 3049 7515 3115 7518
rect 5257 7578 5323 7581
rect 6913 7578 6979 7581
rect 5257 7576 6979 7578
rect 5257 7520 5262 7576
rect 5318 7520 6918 7576
rect 6974 7520 6979 7576
rect 5257 7518 6979 7520
rect 5257 7515 5323 7518
rect 6913 7515 6979 7518
rect 13813 7442 13879 7445
rect 2730 7440 13879 7442
rect 2730 7384 13818 7440
rect 13874 7384 13879 7440
rect 2730 7382 13879 7384
rect 13813 7379 13879 7382
rect 2865 7306 2931 7309
rect 8661 7306 8727 7309
rect 2865 7304 8727 7306
rect 2865 7248 2870 7304
rect 2926 7248 8666 7304
rect 8722 7248 8727 7304
rect 2865 7246 8727 7248
rect 2865 7243 2931 7246
rect 8661 7243 8727 7246
rect 13537 7306 13603 7309
rect 14000 7306 34000 7336
rect 13537 7304 34000 7306
rect 13537 7248 13542 7304
rect 13598 7248 34000 7304
rect 13537 7246 34000 7248
rect 13537 7243 13603 7246
rect 14000 7216 34000 7246
rect 3417 7170 3483 7173
rect 3417 7168 5274 7170
rect 3417 7112 3422 7168
rect 3478 7112 5274 7168
rect 3417 7110 5274 7112
rect 3417 7107 3483 7110
rect 2560 7104 2880 7105
rect 2560 7040 2568 7104
rect 2632 7040 2648 7104
rect 2712 7040 2728 7104
rect 2792 7040 2808 7104
rect 2872 7040 2880 7104
rect 2560 7039 2880 7040
rect 3877 7034 3943 7037
rect 4521 7034 4587 7037
rect 3877 7032 4587 7034
rect 3877 6976 3882 7032
rect 3938 6976 4526 7032
rect 4582 6976 4587 7032
rect 3877 6974 4587 6976
rect 3877 6971 3943 6974
rect 4521 6971 4587 6974
rect 4981 7032 5047 7037
rect 4981 6976 4986 7032
rect 5042 6976 5047 7032
rect 4981 6971 5047 6976
rect 1393 6898 1459 6901
rect 4984 6898 5044 6971
rect 1393 6896 5044 6898
rect 1393 6840 1398 6896
rect 1454 6840 5044 6896
rect 1393 6838 5044 6840
rect 5214 6898 5274 7110
rect 5660 7104 5980 7105
rect 5660 7040 5668 7104
rect 5732 7040 5748 7104
rect 5812 7040 5828 7104
rect 5892 7040 5908 7104
rect 5972 7040 5980 7104
rect 5660 7039 5980 7040
rect 8760 7104 9080 7105
rect 8760 7040 8768 7104
rect 8832 7040 8848 7104
rect 8912 7040 8928 7104
rect 8992 7040 9008 7104
rect 9072 7040 9080 7104
rect 8760 7039 9080 7040
rect 13629 7034 13695 7037
rect 14000 7034 34000 7064
rect 13629 7032 34000 7034
rect 13629 6976 13634 7032
rect 13690 6976 34000 7032
rect 13629 6974 34000 6976
rect 13629 6971 13695 6974
rect 14000 6944 34000 6974
rect 6269 6898 6335 6901
rect 5214 6896 6335 6898
rect 5214 6840 6274 6896
rect 6330 6840 6335 6896
rect 5214 6838 6335 6840
rect 1393 6835 1459 6838
rect 6269 6835 6335 6838
rect 2037 6762 2103 6765
rect 2957 6762 3023 6765
rect 2037 6760 3023 6762
rect 2037 6704 2042 6760
rect 2098 6704 2962 6760
rect 3018 6704 3023 6760
rect 2037 6702 3023 6704
rect 2037 6699 2103 6702
rect 2957 6699 3023 6702
rect 3325 6762 3391 6765
rect 5257 6762 5323 6765
rect 7005 6762 7071 6765
rect 3325 6760 5323 6762
rect 3325 6704 3330 6760
rect 3386 6704 5262 6760
rect 5318 6704 5323 6760
rect 3325 6702 5323 6704
rect 3325 6699 3391 6702
rect 5257 6699 5323 6702
rect 5766 6760 7071 6762
rect 5766 6704 7010 6760
rect 7066 6704 7071 6760
rect 5766 6702 7071 6704
rect 1301 6626 1367 6629
rect 3877 6626 3943 6629
rect 1301 6624 3943 6626
rect 1301 6568 1306 6624
rect 1362 6568 3882 6624
rect 3938 6568 3943 6624
rect 1301 6566 3943 6568
rect 1301 6563 1367 6566
rect 3877 6563 3943 6566
rect 5349 6626 5415 6629
rect 5766 6626 5826 6702
rect 7005 6699 7071 6702
rect 5349 6624 5826 6626
rect 5349 6568 5354 6624
rect 5410 6568 5826 6624
rect 5349 6566 5826 6568
rect 13813 6626 13879 6629
rect 14000 6626 34000 6656
rect 13813 6624 34000 6626
rect 13813 6568 13818 6624
rect 13874 6568 34000 6624
rect 13813 6566 34000 6568
rect 5349 6563 5415 6566
rect 13813 6563 13879 6566
rect 4110 6560 4430 6561
rect 4110 6496 4118 6560
rect 4182 6496 4198 6560
rect 4262 6496 4278 6560
rect 4342 6496 4358 6560
rect 4422 6496 4430 6560
rect 4110 6495 4430 6496
rect 7210 6560 7530 6561
rect 7210 6496 7218 6560
rect 7282 6496 7298 6560
rect 7362 6496 7378 6560
rect 7442 6496 7458 6560
rect 7522 6496 7530 6560
rect 14000 6536 34000 6566
rect 7210 6495 7530 6496
rect 5625 6490 5691 6493
rect 7005 6490 7071 6493
rect 5625 6488 7071 6490
rect 5625 6432 5630 6488
rect 5686 6432 7010 6488
rect 7066 6432 7071 6488
rect 5625 6430 7071 6432
rect 5625 6427 5691 6430
rect 7005 6427 7071 6430
rect 3601 6354 3667 6357
rect 7281 6354 7347 6357
rect 3601 6352 7347 6354
rect 3601 6296 3606 6352
rect 3662 6296 7286 6352
rect 7342 6296 7347 6352
rect 3601 6294 7347 6296
rect 3601 6291 3667 6294
rect 7281 6291 7347 6294
rect 7465 6354 7531 6357
rect 8017 6354 8083 6357
rect 7465 6352 8083 6354
rect 7465 6296 7470 6352
rect 7526 6296 8022 6352
rect 8078 6296 8083 6352
rect 7465 6294 8083 6296
rect 7465 6291 7531 6294
rect 8017 6291 8083 6294
rect 13721 6354 13787 6357
rect 14000 6354 34000 6384
rect 13721 6352 34000 6354
rect 13721 6296 13726 6352
rect 13782 6296 34000 6352
rect 13721 6294 34000 6296
rect 13721 6291 13787 6294
rect 14000 6264 34000 6294
rect 2037 6218 2103 6221
rect 8661 6218 8727 6221
rect 2037 6216 8727 6218
rect 2037 6160 2042 6216
rect 2098 6160 8666 6216
rect 8722 6160 8727 6216
rect 2037 6158 8727 6160
rect 2037 6155 2103 6158
rect 8661 6155 8727 6158
rect 1209 6082 1275 6085
rect 5533 6082 5599 6085
rect 1209 6080 5599 6082
rect 1209 6024 1214 6080
rect 1270 6024 5538 6080
rect 5594 6024 5599 6080
rect 1209 6022 5599 6024
rect 1209 6019 1275 6022
rect 5533 6019 5599 6022
rect 12801 6082 12867 6085
rect 14000 6082 34000 6112
rect 12801 6080 34000 6082
rect 12801 6024 12806 6080
rect 12862 6024 34000 6080
rect 12801 6022 34000 6024
rect 12801 6019 12867 6022
rect 5660 6016 5980 6017
rect 5660 5952 5668 6016
rect 5732 5952 5748 6016
rect 5812 5952 5828 6016
rect 5892 5952 5908 6016
rect 5972 5952 5980 6016
rect 5660 5951 5980 5952
rect 8760 6016 9080 6017
rect 8760 5952 8768 6016
rect 8832 5952 8848 6016
rect 8912 5952 8928 6016
rect 8992 5952 9008 6016
rect 9072 5952 9080 6016
rect 14000 5992 34000 6022
rect 8760 5951 9080 5952
rect 2681 5946 2747 5949
rect 2681 5944 5596 5946
rect 2681 5888 2686 5944
rect 2742 5888 5596 5944
rect 2681 5886 5596 5888
rect 2681 5883 2747 5886
rect 2313 5810 2379 5813
rect 5536 5810 5596 5886
rect 7741 5810 7807 5813
rect 2313 5808 2790 5810
rect 2313 5752 2318 5808
rect 2374 5752 2790 5808
rect 2313 5750 2790 5752
rect 5536 5808 7807 5810
rect 5536 5752 7746 5808
rect 7802 5752 7807 5808
rect 5536 5750 7807 5752
rect 2313 5747 2379 5750
rect 2730 5674 2790 5750
rect 7741 5747 7807 5750
rect 14000 5674 34000 5704
rect 2730 5614 34000 5674
rect 14000 5584 34000 5614
rect 4110 5472 4430 5473
rect 4110 5408 4118 5472
rect 4182 5408 4198 5472
rect 4262 5408 4278 5472
rect 4342 5408 4358 5472
rect 4422 5408 4430 5472
rect 4110 5407 4430 5408
rect 7210 5472 7530 5473
rect 7210 5408 7218 5472
rect 7282 5408 7298 5472
rect 7362 5408 7378 5472
rect 7442 5408 7458 5472
rect 7522 5408 7530 5472
rect 7210 5407 7530 5408
rect 14000 5402 34000 5432
rect 12390 5342 34000 5402
rect 2405 5266 2471 5269
rect 12390 5266 12450 5342
rect 14000 5312 34000 5342
rect 2405 5264 12450 5266
rect 2405 5208 2410 5264
rect 2466 5208 12450 5264
rect 2405 5206 12450 5208
rect 2405 5203 2471 5206
rect 8845 5130 8911 5133
rect 8572 5128 8911 5130
rect 8572 5072 8850 5128
rect 8906 5072 8911 5128
rect 8572 5070 8911 5072
rect 2773 4994 2839 4997
rect 2454 4992 2839 4994
rect 2454 4936 2778 4992
rect 2834 4936 2839 4992
rect 2454 4934 2839 4936
rect 2454 4420 2514 4934
rect 2773 4931 2839 4934
rect 5660 4928 5980 4929
rect 5660 4864 5668 4928
rect 5732 4864 5748 4928
rect 5812 4864 5828 4928
rect 5892 4864 5908 4928
rect 5972 4864 5980 4928
rect 5660 4863 5980 4864
rect 4429 4722 4495 4725
rect 5901 4722 5967 4725
rect 4429 4720 5967 4722
rect 4429 4664 4434 4720
rect 4490 4664 5906 4720
rect 5962 4664 5967 4720
rect 4429 4662 5967 4664
rect 8572 4722 8632 5070
rect 8845 5067 8911 5070
rect 10869 4994 10935 4997
rect 14000 4994 34000 5024
rect 10869 4992 34000 4994
rect 10869 4936 10874 4992
rect 10930 4936 34000 4992
rect 10869 4934 34000 4936
rect 10869 4931 10935 4934
rect 8760 4928 9080 4929
rect 8760 4864 8768 4928
rect 8832 4864 8848 4928
rect 8912 4864 8928 4928
rect 8992 4864 9008 4928
rect 9072 4864 9080 4928
rect 14000 4904 34000 4934
rect 8760 4863 9080 4864
rect 8753 4722 8819 4725
rect 8572 4720 8819 4722
rect 8572 4664 8758 4720
rect 8814 4664 8819 4720
rect 8572 4662 8819 4664
rect 4429 4659 4495 4662
rect 5901 4659 5967 4662
rect 8753 4659 8819 4662
rect 9673 4722 9739 4725
rect 14000 4722 34000 4752
rect 9673 4720 34000 4722
rect 9673 4664 9678 4720
rect 9734 4664 34000 4720
rect 9673 4662 34000 4664
rect 9673 4659 9739 4662
rect 14000 4632 34000 4662
rect 4153 4586 4219 4589
rect 5717 4586 5783 4589
rect 4153 4584 5783 4586
rect 4153 4528 4158 4584
rect 4214 4528 5722 4584
rect 5778 4528 5783 4584
rect 4153 4526 5783 4528
rect 4153 4523 4219 4526
rect 5717 4523 5783 4526
rect 13813 4450 13879 4453
rect 14000 4450 34000 4480
rect 13813 4448 34000 4450
rect 13813 4392 13818 4448
rect 13874 4392 34000 4448
rect 13813 4390 34000 4392
rect 13813 4387 13879 4390
rect 4110 4384 4430 4385
rect 4110 4320 4118 4384
rect 4182 4320 4198 4384
rect 4262 4320 4278 4384
rect 4342 4320 4358 4384
rect 4422 4320 4430 4384
rect 4110 4319 4430 4320
rect 7210 4384 7530 4385
rect 7210 4320 7218 4384
rect 7282 4320 7298 4384
rect 7362 4320 7378 4384
rect 7442 4320 7458 4384
rect 7522 4320 7530 4384
rect 14000 4360 34000 4390
rect 7210 4319 7530 4320
rect 2865 4042 2931 4045
rect 14000 4042 34000 4072
rect 2865 4040 34000 4042
rect 2865 3984 2870 4040
rect 2926 3984 34000 4040
rect 2865 3982 34000 3984
rect 2865 3979 2931 3982
rect 14000 3952 34000 3982
rect 5660 3840 5980 3841
rect 5660 3776 5668 3840
rect 5732 3776 5748 3840
rect 5812 3776 5828 3840
rect 5892 3776 5908 3840
rect 5972 3776 5980 3840
rect 5660 3775 5980 3776
rect 8760 3840 9080 3841
rect 8760 3776 8768 3840
rect 8832 3776 8848 3840
rect 8912 3776 8928 3840
rect 8992 3776 9008 3840
rect 9072 3776 9080 3840
rect 8760 3775 9080 3776
rect 13629 3770 13695 3773
rect 14000 3770 34000 3800
rect 13629 3768 34000 3770
rect 13629 3712 13634 3768
rect 13690 3712 34000 3768
rect 13629 3710 34000 3712
rect 13629 3707 13695 3710
rect 14000 3680 34000 3710
rect 2405 3634 2471 3637
rect 2681 3634 2747 3637
rect 2405 3632 2747 3634
rect 2405 3576 2410 3632
rect 2466 3576 2686 3632
rect 2742 3576 2747 3632
rect 2405 3574 2747 3576
rect 2405 3571 2471 3574
rect 2681 3571 2747 3574
rect 13721 3362 13787 3365
rect 14000 3362 34000 3392
rect 13721 3360 34000 3362
rect 13721 3304 13726 3360
rect 13782 3304 34000 3360
rect 13721 3302 34000 3304
rect 13721 3299 13787 3302
rect 4110 3296 4430 3297
rect 4110 3232 4118 3296
rect 4182 3232 4198 3296
rect 4262 3232 4278 3296
rect 4342 3232 4358 3296
rect 4422 3232 4430 3296
rect 4110 3231 4430 3232
rect 7210 3296 7530 3297
rect 7210 3232 7218 3296
rect 7282 3232 7298 3296
rect 7362 3232 7378 3296
rect 7442 3232 7458 3296
rect 7522 3232 7530 3296
rect 14000 3272 34000 3302
rect 7210 3231 7530 3232
rect 6269 3090 6335 3093
rect 14000 3090 34000 3120
rect 6269 3088 34000 3090
rect 6269 3032 6274 3088
rect 6330 3032 34000 3088
rect 6269 3030 34000 3032
rect 6269 3027 6335 3030
rect 14000 3000 34000 3030
rect 3233 2954 3299 2957
rect 3233 2952 12450 2954
rect 3233 2896 3238 2952
rect 3294 2896 12450 2952
rect 3233 2894 12450 2896
rect 3233 2891 3299 2894
rect 7465 2818 7531 2821
rect 8293 2818 8359 2821
rect 7465 2816 8359 2818
rect 7465 2760 7470 2816
rect 7526 2760 8298 2816
rect 8354 2760 8359 2816
rect 7465 2758 8359 2760
rect 12390 2818 12450 2894
rect 14000 2818 34000 2848
rect 12390 2758 34000 2818
rect 7465 2755 7531 2758
rect 8293 2755 8359 2758
rect 5660 2752 5980 2753
rect 5660 2688 5668 2752
rect 5732 2688 5748 2752
rect 5812 2688 5828 2752
rect 5892 2688 5908 2752
rect 5972 2688 5980 2752
rect 5660 2687 5980 2688
rect 8760 2752 9080 2753
rect 8760 2688 8768 2752
rect 8832 2688 8848 2752
rect 8912 2688 8928 2752
rect 8992 2688 9008 2752
rect 9072 2688 9080 2752
rect 14000 2728 34000 2758
rect 8760 2687 9080 2688
rect 14000 2408 34000 2440
rect 14000 2352 19430 2408
rect 19486 2352 34000 2408
rect 14000 2320 34000 2352
rect 4110 2208 4430 2209
rect 4110 2144 4118 2208
rect 4182 2144 4198 2208
rect 4262 2144 4278 2208
rect 4342 2144 4358 2208
rect 4422 2144 4430 2208
rect 4110 2143 4430 2144
rect 7210 2208 7530 2209
rect 7210 2144 7218 2208
rect 7282 2144 7298 2208
rect 7362 2144 7378 2208
rect 7442 2144 7458 2208
rect 7522 2144 7530 2208
rect 7210 2143 7530 2144
rect 14000 2138 34000 2168
rect 10366 2078 34000 2138
rect 3141 2002 3207 2005
rect 10366 2002 10426 2078
rect 14000 2048 34000 2078
rect 3141 2000 10426 2002
rect 3141 1944 3146 2000
rect 3202 1944 10426 2000
rect 3141 1942 10426 1944
rect 3141 1939 3207 1942
rect 3417 1730 3483 1733
rect 14000 1730 34000 1760
rect 3417 1728 34000 1730
rect 3417 1672 3422 1728
rect 3478 1672 34000 1728
rect 3417 1670 34000 1672
rect 3417 1667 3483 1670
rect 14000 1640 34000 1670
rect 1117 1458 1183 1461
rect 14000 1458 34000 1488
rect 1117 1456 34000 1458
rect 1117 1400 1122 1456
rect 1178 1400 34000 1456
rect 1117 1398 34000 1400
rect 1117 1395 1183 1398
rect 14000 1368 34000 1398
rect 14000 1186 34000 1216
rect 6870 1126 34000 1186
rect 2773 1050 2839 1053
rect 6870 1050 6930 1126
rect 14000 1096 34000 1126
rect 2773 1048 6930 1050
rect 2773 992 2778 1048
rect 2834 992 6930 1048
rect 2773 990 6930 992
rect 2773 987 2839 990
rect 14000 776 34000 808
rect 14000 720 22282 776
rect 22338 720 34000 776
rect 14000 688 34000 720
rect 3509 506 3575 509
rect 14000 506 34000 536
rect 3509 504 34000 506
rect 3509 448 3514 504
rect 3570 448 34000 504
rect 3509 446 34000 448
rect 3509 443 3575 446
rect 14000 416 34000 446
rect 14000 232 34000 264
rect 14000 176 22374 232
rect 22430 176 34000 232
rect 14000 144 34000 176
<< via3 >>
rect 2568 11452 2632 11456
rect 2568 11396 2572 11452
rect 2572 11396 2628 11452
rect 2628 11396 2632 11452
rect 2568 11392 2632 11396
rect 2648 11452 2712 11456
rect 2648 11396 2652 11452
rect 2652 11396 2708 11452
rect 2708 11396 2712 11452
rect 2648 11392 2712 11396
rect 2728 11452 2792 11456
rect 2728 11396 2732 11452
rect 2732 11396 2788 11452
rect 2788 11396 2792 11452
rect 2728 11392 2792 11396
rect 2808 11452 2872 11456
rect 2808 11396 2812 11452
rect 2812 11396 2868 11452
rect 2868 11396 2872 11452
rect 2808 11392 2872 11396
rect 5668 11452 5732 11456
rect 5668 11396 5672 11452
rect 5672 11396 5728 11452
rect 5728 11396 5732 11452
rect 5668 11392 5732 11396
rect 5748 11452 5812 11456
rect 5748 11396 5752 11452
rect 5752 11396 5808 11452
rect 5808 11396 5812 11452
rect 5748 11392 5812 11396
rect 5828 11452 5892 11456
rect 5828 11396 5832 11452
rect 5832 11396 5888 11452
rect 5888 11396 5892 11452
rect 5828 11392 5892 11396
rect 5908 11452 5972 11456
rect 5908 11396 5912 11452
rect 5912 11396 5968 11452
rect 5968 11396 5972 11452
rect 5908 11392 5972 11396
rect 8768 11452 8832 11456
rect 8768 11396 8772 11452
rect 8772 11396 8828 11452
rect 8828 11396 8832 11452
rect 8768 11392 8832 11396
rect 8848 11452 8912 11456
rect 8848 11396 8852 11452
rect 8852 11396 8908 11452
rect 8908 11396 8912 11452
rect 8848 11392 8912 11396
rect 8928 11452 8992 11456
rect 8928 11396 8932 11452
rect 8932 11396 8988 11452
rect 8988 11396 8992 11452
rect 8928 11392 8992 11396
rect 9008 11452 9072 11456
rect 9008 11396 9012 11452
rect 9012 11396 9068 11452
rect 9068 11396 9072 11452
rect 9008 11392 9072 11396
rect 4118 10908 4182 10912
rect 4118 10852 4122 10908
rect 4122 10852 4178 10908
rect 4178 10852 4182 10908
rect 4118 10848 4182 10852
rect 4198 10908 4262 10912
rect 4198 10852 4202 10908
rect 4202 10852 4258 10908
rect 4258 10852 4262 10908
rect 4198 10848 4262 10852
rect 4278 10908 4342 10912
rect 4278 10852 4282 10908
rect 4282 10852 4338 10908
rect 4338 10852 4342 10908
rect 4278 10848 4342 10852
rect 4358 10908 4422 10912
rect 4358 10852 4362 10908
rect 4362 10852 4418 10908
rect 4418 10852 4422 10908
rect 4358 10848 4422 10852
rect 7218 10908 7282 10912
rect 7218 10852 7222 10908
rect 7222 10852 7278 10908
rect 7278 10852 7282 10908
rect 7218 10848 7282 10852
rect 7298 10908 7362 10912
rect 7298 10852 7302 10908
rect 7302 10852 7358 10908
rect 7358 10852 7362 10908
rect 7298 10848 7362 10852
rect 7378 10908 7442 10912
rect 7378 10852 7382 10908
rect 7382 10852 7438 10908
rect 7438 10852 7442 10908
rect 7378 10848 7442 10852
rect 7458 10908 7522 10912
rect 7458 10852 7462 10908
rect 7462 10852 7518 10908
rect 7518 10852 7522 10908
rect 7458 10848 7522 10852
rect 2568 10364 2632 10368
rect 2568 10308 2572 10364
rect 2572 10308 2628 10364
rect 2628 10308 2632 10364
rect 2568 10304 2632 10308
rect 2648 10364 2712 10368
rect 2648 10308 2652 10364
rect 2652 10308 2708 10364
rect 2708 10308 2712 10364
rect 2648 10304 2712 10308
rect 2728 10364 2792 10368
rect 2728 10308 2732 10364
rect 2732 10308 2788 10364
rect 2788 10308 2792 10364
rect 2728 10304 2792 10308
rect 2808 10364 2872 10368
rect 2808 10308 2812 10364
rect 2812 10308 2868 10364
rect 2868 10308 2872 10364
rect 2808 10304 2872 10308
rect 5668 10364 5732 10368
rect 5668 10308 5672 10364
rect 5672 10308 5728 10364
rect 5728 10308 5732 10364
rect 5668 10304 5732 10308
rect 5748 10364 5812 10368
rect 5748 10308 5752 10364
rect 5752 10308 5808 10364
rect 5808 10308 5812 10364
rect 5748 10304 5812 10308
rect 5828 10364 5892 10368
rect 5828 10308 5832 10364
rect 5832 10308 5888 10364
rect 5888 10308 5892 10364
rect 5828 10304 5892 10308
rect 5908 10364 5972 10368
rect 5908 10308 5912 10364
rect 5912 10308 5968 10364
rect 5968 10308 5972 10364
rect 5908 10304 5972 10308
rect 8768 10364 8832 10368
rect 8768 10308 8772 10364
rect 8772 10308 8828 10364
rect 8828 10308 8832 10364
rect 8768 10304 8832 10308
rect 8848 10364 8912 10368
rect 8848 10308 8852 10364
rect 8852 10308 8908 10364
rect 8908 10308 8912 10364
rect 8848 10304 8912 10308
rect 8928 10364 8992 10368
rect 8928 10308 8932 10364
rect 8932 10308 8988 10364
rect 8988 10308 8992 10364
rect 8928 10304 8992 10308
rect 9008 10364 9072 10368
rect 9008 10308 9012 10364
rect 9012 10308 9068 10364
rect 9068 10308 9072 10364
rect 9008 10304 9072 10308
rect 4118 9820 4182 9824
rect 4118 9764 4122 9820
rect 4122 9764 4178 9820
rect 4178 9764 4182 9820
rect 4118 9760 4182 9764
rect 4198 9820 4262 9824
rect 4198 9764 4202 9820
rect 4202 9764 4258 9820
rect 4258 9764 4262 9820
rect 4198 9760 4262 9764
rect 4278 9820 4342 9824
rect 4278 9764 4282 9820
rect 4282 9764 4338 9820
rect 4338 9764 4342 9820
rect 4278 9760 4342 9764
rect 4358 9820 4422 9824
rect 4358 9764 4362 9820
rect 4362 9764 4418 9820
rect 4418 9764 4422 9820
rect 4358 9760 4422 9764
rect 7218 9820 7282 9824
rect 7218 9764 7222 9820
rect 7222 9764 7278 9820
rect 7278 9764 7282 9820
rect 7218 9760 7282 9764
rect 7298 9820 7362 9824
rect 7298 9764 7302 9820
rect 7302 9764 7358 9820
rect 7358 9764 7362 9820
rect 7298 9760 7362 9764
rect 7378 9820 7442 9824
rect 7378 9764 7382 9820
rect 7382 9764 7438 9820
rect 7438 9764 7442 9820
rect 7378 9760 7442 9764
rect 7458 9820 7522 9824
rect 7458 9764 7462 9820
rect 7462 9764 7518 9820
rect 7518 9764 7522 9820
rect 7458 9760 7522 9764
rect 2568 9276 2632 9280
rect 2568 9220 2572 9276
rect 2572 9220 2628 9276
rect 2628 9220 2632 9276
rect 2568 9216 2632 9220
rect 2648 9276 2712 9280
rect 2648 9220 2652 9276
rect 2652 9220 2708 9276
rect 2708 9220 2712 9276
rect 2648 9216 2712 9220
rect 2728 9276 2792 9280
rect 2728 9220 2732 9276
rect 2732 9220 2788 9276
rect 2788 9220 2792 9276
rect 2728 9216 2792 9220
rect 2808 9276 2872 9280
rect 2808 9220 2812 9276
rect 2812 9220 2868 9276
rect 2868 9220 2872 9276
rect 2808 9216 2872 9220
rect 5668 9276 5732 9280
rect 5668 9220 5672 9276
rect 5672 9220 5728 9276
rect 5728 9220 5732 9276
rect 5668 9216 5732 9220
rect 5748 9276 5812 9280
rect 5748 9220 5752 9276
rect 5752 9220 5808 9276
rect 5808 9220 5812 9276
rect 5748 9216 5812 9220
rect 5828 9276 5892 9280
rect 5828 9220 5832 9276
rect 5832 9220 5888 9276
rect 5888 9220 5892 9276
rect 5828 9216 5892 9220
rect 5908 9276 5972 9280
rect 5908 9220 5912 9276
rect 5912 9220 5968 9276
rect 5968 9220 5972 9276
rect 5908 9216 5972 9220
rect 8768 9276 8832 9280
rect 8768 9220 8772 9276
rect 8772 9220 8828 9276
rect 8828 9220 8832 9276
rect 8768 9216 8832 9220
rect 8848 9276 8912 9280
rect 8848 9220 8852 9276
rect 8852 9220 8908 9276
rect 8908 9220 8912 9276
rect 8848 9216 8912 9220
rect 8928 9276 8992 9280
rect 8928 9220 8932 9276
rect 8932 9220 8988 9276
rect 8988 9220 8992 9276
rect 8928 9216 8992 9220
rect 9008 9276 9072 9280
rect 9008 9220 9012 9276
rect 9012 9220 9068 9276
rect 9068 9220 9072 9276
rect 9008 9216 9072 9220
rect 4118 8732 4182 8736
rect 4118 8676 4122 8732
rect 4122 8676 4178 8732
rect 4178 8676 4182 8732
rect 4118 8672 4182 8676
rect 4198 8732 4262 8736
rect 4198 8676 4202 8732
rect 4202 8676 4258 8732
rect 4258 8676 4262 8732
rect 4198 8672 4262 8676
rect 4278 8732 4342 8736
rect 4278 8676 4282 8732
rect 4282 8676 4338 8732
rect 4338 8676 4342 8732
rect 4278 8672 4342 8676
rect 4358 8732 4422 8736
rect 4358 8676 4362 8732
rect 4362 8676 4418 8732
rect 4418 8676 4422 8732
rect 4358 8672 4422 8676
rect 7218 8732 7282 8736
rect 7218 8676 7222 8732
rect 7222 8676 7278 8732
rect 7278 8676 7282 8732
rect 7218 8672 7282 8676
rect 7298 8732 7362 8736
rect 7298 8676 7302 8732
rect 7302 8676 7358 8732
rect 7358 8676 7362 8732
rect 7298 8672 7362 8676
rect 7378 8732 7442 8736
rect 7378 8676 7382 8732
rect 7382 8676 7438 8732
rect 7438 8676 7442 8732
rect 7378 8672 7442 8676
rect 7458 8732 7522 8736
rect 7458 8676 7462 8732
rect 7462 8676 7518 8732
rect 7518 8676 7522 8732
rect 7458 8672 7522 8676
rect 2568 8188 2632 8192
rect 2568 8132 2572 8188
rect 2572 8132 2628 8188
rect 2628 8132 2632 8188
rect 2568 8128 2632 8132
rect 2648 8188 2712 8192
rect 2648 8132 2652 8188
rect 2652 8132 2708 8188
rect 2708 8132 2712 8188
rect 2648 8128 2712 8132
rect 2728 8188 2792 8192
rect 2728 8132 2732 8188
rect 2732 8132 2788 8188
rect 2788 8132 2792 8188
rect 2728 8128 2792 8132
rect 2808 8188 2872 8192
rect 2808 8132 2812 8188
rect 2812 8132 2868 8188
rect 2868 8132 2872 8188
rect 2808 8128 2872 8132
rect 5668 8188 5732 8192
rect 5668 8132 5672 8188
rect 5672 8132 5728 8188
rect 5728 8132 5732 8188
rect 5668 8128 5732 8132
rect 5748 8188 5812 8192
rect 5748 8132 5752 8188
rect 5752 8132 5808 8188
rect 5808 8132 5812 8188
rect 5748 8128 5812 8132
rect 5828 8188 5892 8192
rect 5828 8132 5832 8188
rect 5832 8132 5888 8188
rect 5888 8132 5892 8188
rect 5828 8128 5892 8132
rect 5908 8188 5972 8192
rect 5908 8132 5912 8188
rect 5912 8132 5968 8188
rect 5968 8132 5972 8188
rect 5908 8128 5972 8132
rect 8768 8188 8832 8192
rect 8768 8132 8772 8188
rect 8772 8132 8828 8188
rect 8828 8132 8832 8188
rect 8768 8128 8832 8132
rect 8848 8188 8912 8192
rect 8848 8132 8852 8188
rect 8852 8132 8908 8188
rect 8908 8132 8912 8188
rect 8848 8128 8912 8132
rect 8928 8188 8992 8192
rect 8928 8132 8932 8188
rect 8932 8132 8988 8188
rect 8988 8132 8992 8188
rect 8928 8128 8992 8132
rect 9008 8188 9072 8192
rect 9008 8132 9012 8188
rect 9012 8132 9068 8188
rect 9068 8132 9072 8188
rect 9008 8128 9072 8132
rect 4118 7644 4182 7648
rect 4118 7588 4122 7644
rect 4122 7588 4178 7644
rect 4178 7588 4182 7644
rect 4118 7584 4182 7588
rect 4198 7644 4262 7648
rect 4198 7588 4202 7644
rect 4202 7588 4258 7644
rect 4258 7588 4262 7644
rect 4198 7584 4262 7588
rect 4278 7644 4342 7648
rect 4278 7588 4282 7644
rect 4282 7588 4338 7644
rect 4338 7588 4342 7644
rect 4278 7584 4342 7588
rect 4358 7644 4422 7648
rect 4358 7588 4362 7644
rect 4362 7588 4418 7644
rect 4418 7588 4422 7644
rect 4358 7584 4422 7588
rect 7218 7644 7282 7648
rect 7218 7588 7222 7644
rect 7222 7588 7278 7644
rect 7278 7588 7282 7644
rect 7218 7584 7282 7588
rect 7298 7644 7362 7648
rect 7298 7588 7302 7644
rect 7302 7588 7358 7644
rect 7358 7588 7362 7644
rect 7298 7584 7362 7588
rect 7378 7644 7442 7648
rect 7378 7588 7382 7644
rect 7382 7588 7438 7644
rect 7438 7588 7442 7644
rect 7378 7584 7442 7588
rect 7458 7644 7522 7648
rect 7458 7588 7462 7644
rect 7462 7588 7518 7644
rect 7518 7588 7522 7644
rect 7458 7584 7522 7588
rect 2568 7100 2632 7104
rect 2568 7044 2572 7100
rect 2572 7044 2628 7100
rect 2628 7044 2632 7100
rect 2568 7040 2632 7044
rect 2648 7100 2712 7104
rect 2648 7044 2652 7100
rect 2652 7044 2708 7100
rect 2708 7044 2712 7100
rect 2648 7040 2712 7044
rect 2728 7100 2792 7104
rect 2728 7044 2732 7100
rect 2732 7044 2788 7100
rect 2788 7044 2792 7100
rect 2728 7040 2792 7044
rect 2808 7100 2872 7104
rect 2808 7044 2812 7100
rect 2812 7044 2868 7100
rect 2868 7044 2872 7100
rect 2808 7040 2872 7044
rect 5668 7100 5732 7104
rect 5668 7044 5672 7100
rect 5672 7044 5728 7100
rect 5728 7044 5732 7100
rect 5668 7040 5732 7044
rect 5748 7100 5812 7104
rect 5748 7044 5752 7100
rect 5752 7044 5808 7100
rect 5808 7044 5812 7100
rect 5748 7040 5812 7044
rect 5828 7100 5892 7104
rect 5828 7044 5832 7100
rect 5832 7044 5888 7100
rect 5888 7044 5892 7100
rect 5828 7040 5892 7044
rect 5908 7100 5972 7104
rect 5908 7044 5912 7100
rect 5912 7044 5968 7100
rect 5968 7044 5972 7100
rect 5908 7040 5972 7044
rect 8768 7100 8832 7104
rect 8768 7044 8772 7100
rect 8772 7044 8828 7100
rect 8828 7044 8832 7100
rect 8768 7040 8832 7044
rect 8848 7100 8912 7104
rect 8848 7044 8852 7100
rect 8852 7044 8908 7100
rect 8908 7044 8912 7100
rect 8848 7040 8912 7044
rect 8928 7100 8992 7104
rect 8928 7044 8932 7100
rect 8932 7044 8988 7100
rect 8988 7044 8992 7100
rect 8928 7040 8992 7044
rect 9008 7100 9072 7104
rect 9008 7044 9012 7100
rect 9012 7044 9068 7100
rect 9068 7044 9072 7100
rect 9008 7040 9072 7044
rect 4118 6556 4182 6560
rect 4118 6500 4122 6556
rect 4122 6500 4178 6556
rect 4178 6500 4182 6556
rect 4118 6496 4182 6500
rect 4198 6556 4262 6560
rect 4198 6500 4202 6556
rect 4202 6500 4258 6556
rect 4258 6500 4262 6556
rect 4198 6496 4262 6500
rect 4278 6556 4342 6560
rect 4278 6500 4282 6556
rect 4282 6500 4338 6556
rect 4338 6500 4342 6556
rect 4278 6496 4342 6500
rect 4358 6556 4422 6560
rect 4358 6500 4362 6556
rect 4362 6500 4418 6556
rect 4418 6500 4422 6556
rect 4358 6496 4422 6500
rect 7218 6556 7282 6560
rect 7218 6500 7222 6556
rect 7222 6500 7278 6556
rect 7278 6500 7282 6556
rect 7218 6496 7282 6500
rect 7298 6556 7362 6560
rect 7298 6500 7302 6556
rect 7302 6500 7358 6556
rect 7358 6500 7362 6556
rect 7298 6496 7362 6500
rect 7378 6556 7442 6560
rect 7378 6500 7382 6556
rect 7382 6500 7438 6556
rect 7438 6500 7442 6556
rect 7378 6496 7442 6500
rect 7458 6556 7522 6560
rect 7458 6500 7462 6556
rect 7462 6500 7518 6556
rect 7518 6500 7522 6556
rect 7458 6496 7522 6500
rect 5668 6012 5732 6016
rect 5668 5956 5672 6012
rect 5672 5956 5728 6012
rect 5728 5956 5732 6012
rect 5668 5952 5732 5956
rect 5748 6012 5812 6016
rect 5748 5956 5752 6012
rect 5752 5956 5808 6012
rect 5808 5956 5812 6012
rect 5748 5952 5812 5956
rect 5828 6012 5892 6016
rect 5828 5956 5832 6012
rect 5832 5956 5888 6012
rect 5888 5956 5892 6012
rect 5828 5952 5892 5956
rect 5908 6012 5972 6016
rect 5908 5956 5912 6012
rect 5912 5956 5968 6012
rect 5968 5956 5972 6012
rect 5908 5952 5972 5956
rect 8768 6012 8832 6016
rect 8768 5956 8772 6012
rect 8772 5956 8828 6012
rect 8828 5956 8832 6012
rect 8768 5952 8832 5956
rect 8848 6012 8912 6016
rect 8848 5956 8852 6012
rect 8852 5956 8908 6012
rect 8908 5956 8912 6012
rect 8848 5952 8912 5956
rect 8928 6012 8992 6016
rect 8928 5956 8932 6012
rect 8932 5956 8988 6012
rect 8988 5956 8992 6012
rect 8928 5952 8992 5956
rect 9008 6012 9072 6016
rect 9008 5956 9012 6012
rect 9012 5956 9068 6012
rect 9068 5956 9072 6012
rect 9008 5952 9072 5956
rect 4118 5468 4182 5472
rect 4118 5412 4122 5468
rect 4122 5412 4178 5468
rect 4178 5412 4182 5468
rect 4118 5408 4182 5412
rect 4198 5468 4262 5472
rect 4198 5412 4202 5468
rect 4202 5412 4258 5468
rect 4258 5412 4262 5468
rect 4198 5408 4262 5412
rect 4278 5468 4342 5472
rect 4278 5412 4282 5468
rect 4282 5412 4338 5468
rect 4338 5412 4342 5468
rect 4278 5408 4342 5412
rect 4358 5468 4422 5472
rect 4358 5412 4362 5468
rect 4362 5412 4418 5468
rect 4418 5412 4422 5468
rect 4358 5408 4422 5412
rect 7218 5468 7282 5472
rect 7218 5412 7222 5468
rect 7222 5412 7278 5468
rect 7278 5412 7282 5468
rect 7218 5408 7282 5412
rect 7298 5468 7362 5472
rect 7298 5412 7302 5468
rect 7302 5412 7358 5468
rect 7358 5412 7362 5468
rect 7298 5408 7362 5412
rect 7378 5468 7442 5472
rect 7378 5412 7382 5468
rect 7382 5412 7438 5468
rect 7438 5412 7442 5468
rect 7378 5408 7442 5412
rect 7458 5468 7522 5472
rect 7458 5412 7462 5468
rect 7462 5412 7518 5468
rect 7518 5412 7522 5468
rect 7458 5408 7522 5412
rect 5668 4924 5732 4928
rect 5668 4868 5672 4924
rect 5672 4868 5728 4924
rect 5728 4868 5732 4924
rect 5668 4864 5732 4868
rect 5748 4924 5812 4928
rect 5748 4868 5752 4924
rect 5752 4868 5808 4924
rect 5808 4868 5812 4924
rect 5748 4864 5812 4868
rect 5828 4924 5892 4928
rect 5828 4868 5832 4924
rect 5832 4868 5888 4924
rect 5888 4868 5892 4924
rect 5828 4864 5892 4868
rect 5908 4924 5972 4928
rect 5908 4868 5912 4924
rect 5912 4868 5968 4924
rect 5968 4868 5972 4924
rect 5908 4864 5972 4868
rect 8768 4924 8832 4928
rect 8768 4868 8772 4924
rect 8772 4868 8828 4924
rect 8828 4868 8832 4924
rect 8768 4864 8832 4868
rect 8848 4924 8912 4928
rect 8848 4868 8852 4924
rect 8852 4868 8908 4924
rect 8908 4868 8912 4924
rect 8848 4864 8912 4868
rect 8928 4924 8992 4928
rect 8928 4868 8932 4924
rect 8932 4868 8988 4924
rect 8988 4868 8992 4924
rect 8928 4864 8992 4868
rect 9008 4924 9072 4928
rect 9008 4868 9012 4924
rect 9012 4868 9068 4924
rect 9068 4868 9072 4924
rect 9008 4864 9072 4868
rect 4118 4380 4182 4384
rect 4118 4324 4122 4380
rect 4122 4324 4178 4380
rect 4178 4324 4182 4380
rect 4118 4320 4182 4324
rect 4198 4380 4262 4384
rect 4198 4324 4202 4380
rect 4202 4324 4258 4380
rect 4258 4324 4262 4380
rect 4198 4320 4262 4324
rect 4278 4380 4342 4384
rect 4278 4324 4282 4380
rect 4282 4324 4338 4380
rect 4338 4324 4342 4380
rect 4278 4320 4342 4324
rect 4358 4380 4422 4384
rect 4358 4324 4362 4380
rect 4362 4324 4418 4380
rect 4418 4324 4422 4380
rect 4358 4320 4422 4324
rect 7218 4380 7282 4384
rect 7218 4324 7222 4380
rect 7222 4324 7278 4380
rect 7278 4324 7282 4380
rect 7218 4320 7282 4324
rect 7298 4380 7362 4384
rect 7298 4324 7302 4380
rect 7302 4324 7358 4380
rect 7358 4324 7362 4380
rect 7298 4320 7362 4324
rect 7378 4380 7442 4384
rect 7378 4324 7382 4380
rect 7382 4324 7438 4380
rect 7438 4324 7442 4380
rect 7378 4320 7442 4324
rect 7458 4380 7522 4384
rect 7458 4324 7462 4380
rect 7462 4324 7518 4380
rect 7518 4324 7522 4380
rect 7458 4320 7522 4324
rect 5668 3836 5732 3840
rect 5668 3780 5672 3836
rect 5672 3780 5728 3836
rect 5728 3780 5732 3836
rect 5668 3776 5732 3780
rect 5748 3836 5812 3840
rect 5748 3780 5752 3836
rect 5752 3780 5808 3836
rect 5808 3780 5812 3836
rect 5748 3776 5812 3780
rect 5828 3836 5892 3840
rect 5828 3780 5832 3836
rect 5832 3780 5888 3836
rect 5888 3780 5892 3836
rect 5828 3776 5892 3780
rect 5908 3836 5972 3840
rect 5908 3780 5912 3836
rect 5912 3780 5968 3836
rect 5968 3780 5972 3836
rect 5908 3776 5972 3780
rect 8768 3836 8832 3840
rect 8768 3780 8772 3836
rect 8772 3780 8828 3836
rect 8828 3780 8832 3836
rect 8768 3776 8832 3780
rect 8848 3836 8912 3840
rect 8848 3780 8852 3836
rect 8852 3780 8908 3836
rect 8908 3780 8912 3836
rect 8848 3776 8912 3780
rect 8928 3836 8992 3840
rect 8928 3780 8932 3836
rect 8932 3780 8988 3836
rect 8988 3780 8992 3836
rect 8928 3776 8992 3780
rect 9008 3836 9072 3840
rect 9008 3780 9012 3836
rect 9012 3780 9068 3836
rect 9068 3780 9072 3836
rect 9008 3776 9072 3780
rect 4118 3292 4182 3296
rect 4118 3236 4122 3292
rect 4122 3236 4178 3292
rect 4178 3236 4182 3292
rect 4118 3232 4182 3236
rect 4198 3292 4262 3296
rect 4198 3236 4202 3292
rect 4202 3236 4258 3292
rect 4258 3236 4262 3292
rect 4198 3232 4262 3236
rect 4278 3292 4342 3296
rect 4278 3236 4282 3292
rect 4282 3236 4338 3292
rect 4338 3236 4342 3292
rect 4278 3232 4342 3236
rect 4358 3292 4422 3296
rect 4358 3236 4362 3292
rect 4362 3236 4418 3292
rect 4418 3236 4422 3292
rect 4358 3232 4422 3236
rect 7218 3292 7282 3296
rect 7218 3236 7222 3292
rect 7222 3236 7278 3292
rect 7278 3236 7282 3292
rect 7218 3232 7282 3236
rect 7298 3292 7362 3296
rect 7298 3236 7302 3292
rect 7302 3236 7358 3292
rect 7358 3236 7362 3292
rect 7298 3232 7362 3236
rect 7378 3292 7442 3296
rect 7378 3236 7382 3292
rect 7382 3236 7438 3292
rect 7438 3236 7442 3292
rect 7378 3232 7442 3236
rect 7458 3292 7522 3296
rect 7458 3236 7462 3292
rect 7462 3236 7518 3292
rect 7518 3236 7522 3292
rect 7458 3232 7522 3236
rect 5668 2748 5732 2752
rect 5668 2692 5672 2748
rect 5672 2692 5728 2748
rect 5728 2692 5732 2748
rect 5668 2688 5732 2692
rect 5748 2748 5812 2752
rect 5748 2692 5752 2748
rect 5752 2692 5808 2748
rect 5808 2692 5812 2748
rect 5748 2688 5812 2692
rect 5828 2748 5892 2752
rect 5828 2692 5832 2748
rect 5832 2692 5888 2748
rect 5888 2692 5892 2748
rect 5828 2688 5892 2692
rect 5908 2748 5972 2752
rect 5908 2692 5912 2748
rect 5912 2692 5968 2748
rect 5968 2692 5972 2748
rect 5908 2688 5972 2692
rect 8768 2748 8832 2752
rect 8768 2692 8772 2748
rect 8772 2692 8828 2748
rect 8828 2692 8832 2748
rect 8768 2688 8832 2692
rect 8848 2748 8912 2752
rect 8848 2692 8852 2748
rect 8852 2692 8908 2748
rect 8908 2692 8912 2748
rect 8848 2688 8912 2692
rect 8928 2748 8992 2752
rect 8928 2692 8932 2748
rect 8932 2692 8988 2748
rect 8988 2692 8992 2748
rect 8928 2688 8992 2692
rect 9008 2748 9072 2752
rect 9008 2692 9012 2748
rect 9012 2692 9068 2748
rect 9068 2692 9072 2748
rect 9008 2688 9072 2692
rect 4118 2204 4182 2208
rect 4118 2148 4122 2204
rect 4122 2148 4178 2204
rect 4178 2148 4182 2204
rect 4118 2144 4182 2148
rect 4198 2204 4262 2208
rect 4198 2148 4202 2204
rect 4202 2148 4258 2204
rect 4258 2148 4262 2204
rect 4198 2144 4262 2148
rect 4278 2204 4342 2208
rect 4278 2148 4282 2204
rect 4282 2148 4338 2204
rect 4338 2148 4342 2204
rect 4278 2144 4342 2148
rect 4358 2204 4422 2208
rect 4358 2148 4362 2204
rect 4362 2148 4418 2204
rect 4418 2148 4422 2204
rect 4358 2144 4422 2148
rect 7218 2204 7282 2208
rect 7218 2148 7222 2204
rect 7222 2148 7278 2204
rect 7278 2148 7282 2204
rect 7218 2144 7282 2148
rect 7298 2204 7362 2208
rect 7298 2148 7302 2204
rect 7302 2148 7358 2204
rect 7358 2148 7362 2204
rect 7298 2144 7362 2148
rect 7378 2204 7442 2208
rect 7378 2148 7382 2204
rect 7382 2148 7438 2204
rect 7438 2148 7442 2204
rect 7378 2144 7442 2148
rect 7458 2204 7522 2208
rect 7458 2148 7462 2204
rect 7462 2148 7518 2204
rect 7518 2148 7522 2204
rect 7458 2144 7522 2148
<< metal4 >>
rect -1620 13922 -1300 13964
rect -1620 13686 -1578 13922
rect -1342 13686 -1300 13922
rect -1620 8244 -1300 13686
rect 12064 13922 12384 13964
rect 12064 13686 12106 13922
rect 12342 13686 12384 13922
rect -1620 8008 -1578 8244
rect -1342 8008 -1300 8244
rect -1620 5144 -1300 8008
rect -1620 4908 -1578 5144
rect -1342 4908 -1300 5144
rect -1620 -86 -1300 4908
rect -960 13262 -640 13304
rect -960 13026 -918 13262
rect -682 13026 -640 13262
rect -960 9794 -640 13026
rect 11404 13262 11724 13304
rect 11404 13026 11446 13262
rect 11682 13026 11724 13262
rect -960 9558 -918 9794
rect -682 9558 -640 9794
rect -960 6694 -640 9558
rect -960 6458 -918 6694
rect -682 6458 -640 6694
rect -960 3594 -640 6458
rect -960 3358 -918 3594
rect -682 3358 -640 3594
rect -960 574 -640 3358
rect -300 12602 20 12644
rect -300 12366 -258 12602
rect -22 12366 20 12602
rect -300 10444 20 12366
rect -300 10208 -258 10444
rect -22 10208 20 10444
rect -300 7344 20 10208
rect -300 7108 -258 7344
rect -22 7108 20 7344
rect -300 4244 20 7108
rect -300 4008 -258 4244
rect -22 4008 20 4244
rect -300 1234 20 4008
rect 360 11942 680 11984
rect 360 11706 402 11942
rect 638 11706 680 11942
rect 360 8894 680 11706
rect 360 8658 402 8894
rect 638 8658 680 8894
rect 360 5794 680 8658
rect 360 5558 402 5794
rect 638 5558 680 5794
rect 360 2694 680 5558
rect 2560 11942 2880 12644
rect 2560 11706 2602 11942
rect 2838 11706 2880 11942
rect 2560 11456 2880 11706
rect 2560 11392 2568 11456
rect 2632 11392 2648 11456
rect 2712 11392 2728 11456
rect 2792 11392 2808 11456
rect 2872 11392 2880 11456
rect 2560 10368 2880 11392
rect 2560 10304 2568 10368
rect 2632 10304 2648 10368
rect 2712 10304 2728 10368
rect 2792 10304 2808 10368
rect 2872 10304 2880 10368
rect 2560 9280 2880 10304
rect 2560 9216 2568 9280
rect 2632 9216 2648 9280
rect 2712 9216 2728 9280
rect 2792 9216 2808 9280
rect 2872 9216 2880 9280
rect 2560 8894 2880 9216
rect 2560 8658 2602 8894
rect 2838 8658 2880 8894
rect 2560 8192 2880 8658
rect 2560 8128 2568 8192
rect 2632 8128 2648 8192
rect 2712 8128 2728 8192
rect 2792 8128 2808 8192
rect 2872 8128 2880 8192
rect 2560 7104 2880 8128
rect 2560 7040 2568 7104
rect 2632 7040 2648 7104
rect 2712 7040 2728 7104
rect 2792 7040 2808 7104
rect 2872 7040 2880 7104
rect 2560 5794 2880 7040
rect 2560 5558 2602 5794
rect 2838 5558 2880 5794
rect 1996 5144 2276 5186
rect 1996 4908 2018 5144
rect 2254 4908 2276 5144
rect 1996 4866 2276 4908
rect 1256 3594 1536 3636
rect 1256 3358 1278 3594
rect 1514 3358 1536 3594
rect 1256 3316 1536 3358
rect 360 2458 402 2694
rect 638 2458 680 2694
rect 360 1894 680 2458
rect 360 1658 402 1894
rect 638 1658 680 1894
rect 360 1616 680 1658
rect 2560 2694 2880 5558
rect 2560 2458 2602 2694
rect 2838 2458 2880 2694
rect 2560 1894 2880 2458
rect 2560 1658 2602 1894
rect 2838 1658 2880 1894
rect -300 998 -258 1234
rect -22 998 20 1234
rect -300 956 20 998
rect 2560 956 2880 1658
rect 4110 12602 4430 12644
rect 4110 12366 4152 12602
rect 4388 12366 4430 12602
rect 4110 10912 4430 12366
rect 4110 10848 4118 10912
rect 4182 10848 4198 10912
rect 4262 10848 4278 10912
rect 4342 10848 4358 10912
rect 4422 10848 4430 10912
rect 4110 10444 4430 10848
rect 4110 10208 4152 10444
rect 4388 10208 4430 10444
rect 4110 9824 4430 10208
rect 4110 9760 4118 9824
rect 4182 9760 4198 9824
rect 4262 9760 4278 9824
rect 4342 9760 4358 9824
rect 4422 9760 4430 9824
rect 4110 8736 4430 9760
rect 4110 8672 4118 8736
rect 4182 8672 4198 8736
rect 4262 8672 4278 8736
rect 4342 8672 4358 8736
rect 4422 8672 4430 8736
rect 4110 7648 4430 8672
rect 4110 7584 4118 7648
rect 4182 7584 4198 7648
rect 4262 7584 4278 7648
rect 4342 7584 4358 7648
rect 4422 7584 4430 7648
rect 4110 7344 4430 7584
rect 4110 7108 4152 7344
rect 4388 7108 4430 7344
rect 4110 6560 4430 7108
rect 4110 6496 4118 6560
rect 4182 6496 4198 6560
rect 4262 6496 4278 6560
rect 4342 6496 4358 6560
rect 4422 6496 4430 6560
rect 4110 5472 4430 6496
rect 4110 5408 4118 5472
rect 4182 5408 4198 5472
rect 4262 5408 4278 5472
rect 4342 5408 4358 5472
rect 4422 5408 4430 5472
rect 4110 4384 4430 5408
rect 4110 4320 4118 4384
rect 4182 4320 4198 4384
rect 4262 4320 4278 4384
rect 4342 4320 4358 4384
rect 4422 4320 4430 4384
rect 4110 4244 4430 4320
rect 4110 4008 4152 4244
rect 4388 4008 4430 4244
rect 4110 3296 4430 4008
rect 4110 3232 4118 3296
rect 4182 3232 4198 3296
rect 4262 3232 4278 3296
rect 4342 3232 4358 3296
rect 4422 3232 4430 3296
rect 4110 2208 4430 3232
rect 4110 2144 4118 2208
rect 4182 2144 4198 2208
rect 4262 2144 4278 2208
rect 4342 2144 4358 2208
rect 4422 2144 4430 2208
rect 4110 1234 4430 2144
rect 4110 998 4152 1234
rect 4388 998 4430 1234
rect 4110 956 4430 998
rect 5660 11942 5980 12644
rect 5660 11706 5702 11942
rect 5938 11706 5980 11942
rect 5660 11456 5980 11706
rect 5660 11392 5668 11456
rect 5732 11392 5748 11456
rect 5812 11392 5828 11456
rect 5892 11392 5908 11456
rect 5972 11392 5980 11456
rect 5660 10368 5980 11392
rect 5660 10304 5668 10368
rect 5732 10304 5748 10368
rect 5812 10304 5828 10368
rect 5892 10304 5908 10368
rect 5972 10304 5980 10368
rect 5660 9280 5980 10304
rect 5660 9216 5668 9280
rect 5732 9216 5748 9280
rect 5812 9216 5828 9280
rect 5892 9216 5908 9280
rect 5972 9216 5980 9280
rect 5660 8894 5980 9216
rect 5660 8658 5702 8894
rect 5938 8658 5980 8894
rect 5660 8192 5980 8658
rect 5660 8128 5668 8192
rect 5732 8128 5748 8192
rect 5812 8128 5828 8192
rect 5892 8128 5908 8192
rect 5972 8128 5980 8192
rect 5660 7104 5980 8128
rect 5660 7040 5668 7104
rect 5732 7040 5748 7104
rect 5812 7040 5828 7104
rect 5892 7040 5908 7104
rect 5972 7040 5980 7104
rect 5660 6016 5980 7040
rect 5660 5952 5668 6016
rect 5732 5952 5748 6016
rect 5812 5952 5828 6016
rect 5892 5952 5908 6016
rect 5972 5952 5980 6016
rect 5660 5794 5980 5952
rect 5660 5558 5702 5794
rect 5938 5558 5980 5794
rect 5660 4928 5980 5558
rect 5660 4864 5668 4928
rect 5732 4864 5748 4928
rect 5812 4864 5828 4928
rect 5892 4864 5908 4928
rect 5972 4864 5980 4928
rect 5660 3840 5980 4864
rect 5660 3776 5668 3840
rect 5732 3776 5748 3840
rect 5812 3776 5828 3840
rect 5892 3776 5908 3840
rect 5972 3776 5980 3840
rect 5660 2752 5980 3776
rect 5660 2688 5668 2752
rect 5732 2694 5748 2752
rect 5812 2694 5828 2752
rect 5892 2694 5908 2752
rect 5972 2688 5980 2752
rect 5660 2458 5702 2688
rect 5938 2458 5980 2688
rect 5660 1894 5980 2458
rect 5660 1658 5702 1894
rect 5938 1658 5980 1894
rect 5660 956 5980 1658
rect 7210 12602 7530 12644
rect 7210 12366 7252 12602
rect 7488 12366 7530 12602
rect 7210 10912 7530 12366
rect 7210 10848 7218 10912
rect 7282 10848 7298 10912
rect 7362 10848 7378 10912
rect 7442 10848 7458 10912
rect 7522 10848 7530 10912
rect 7210 10444 7530 10848
rect 7210 10208 7252 10444
rect 7488 10208 7530 10444
rect 7210 9824 7530 10208
rect 7210 9760 7218 9824
rect 7282 9760 7298 9824
rect 7362 9760 7378 9824
rect 7442 9760 7458 9824
rect 7522 9760 7530 9824
rect 7210 8736 7530 9760
rect 7210 8672 7218 8736
rect 7282 8672 7298 8736
rect 7362 8672 7378 8736
rect 7442 8672 7458 8736
rect 7522 8672 7530 8736
rect 7210 7648 7530 8672
rect 7210 7584 7218 7648
rect 7282 7584 7298 7648
rect 7362 7584 7378 7648
rect 7442 7584 7458 7648
rect 7522 7584 7530 7648
rect 7210 7344 7530 7584
rect 7210 7108 7252 7344
rect 7488 7108 7530 7344
rect 7210 6560 7530 7108
rect 7210 6496 7218 6560
rect 7282 6496 7298 6560
rect 7362 6496 7378 6560
rect 7442 6496 7458 6560
rect 7522 6496 7530 6560
rect 7210 5472 7530 6496
rect 7210 5408 7218 5472
rect 7282 5408 7298 5472
rect 7362 5408 7378 5472
rect 7442 5408 7458 5472
rect 7522 5408 7530 5472
rect 7210 4384 7530 5408
rect 7210 4320 7218 4384
rect 7282 4320 7298 4384
rect 7362 4320 7378 4384
rect 7442 4320 7458 4384
rect 7522 4320 7530 4384
rect 7210 4244 7530 4320
rect 7210 4008 7252 4244
rect 7488 4008 7530 4244
rect 7210 3296 7530 4008
rect 7210 3232 7218 3296
rect 7282 3232 7298 3296
rect 7362 3232 7378 3296
rect 7442 3232 7458 3296
rect 7522 3232 7530 3296
rect 7210 2208 7530 3232
rect 7210 2144 7218 2208
rect 7282 2144 7298 2208
rect 7362 2144 7378 2208
rect 7442 2144 7458 2208
rect 7522 2144 7530 2208
rect 7210 1234 7530 2144
rect 7210 998 7252 1234
rect 7488 998 7530 1234
rect 7210 956 7530 998
rect 8760 11942 9080 12644
rect 10744 12602 11064 12644
rect 10744 12366 10786 12602
rect 11022 12366 11064 12602
rect 8760 11706 8802 11942
rect 9038 11706 9080 11942
rect 8760 11456 9080 11706
rect 8760 11392 8768 11456
rect 8832 11392 8848 11456
rect 8912 11392 8928 11456
rect 8992 11392 9008 11456
rect 9072 11392 9080 11456
rect 8760 10368 9080 11392
rect 8760 10304 8768 10368
rect 8832 10304 8848 10368
rect 8912 10304 8928 10368
rect 8992 10304 9008 10368
rect 9072 10304 9080 10368
rect 8760 9280 9080 10304
rect 8760 9216 8768 9280
rect 8832 9216 8848 9280
rect 8912 9216 8928 9280
rect 8992 9216 9008 9280
rect 9072 9216 9080 9280
rect 8760 8894 9080 9216
rect 8760 8658 8802 8894
rect 9038 8658 9080 8894
rect 8760 8192 9080 8658
rect 8760 8128 8768 8192
rect 8832 8128 8848 8192
rect 8912 8128 8928 8192
rect 8992 8128 9008 8192
rect 9072 8128 9080 8192
rect 8760 7104 9080 8128
rect 8760 7040 8768 7104
rect 8832 7040 8848 7104
rect 8912 7040 8928 7104
rect 8992 7040 9008 7104
rect 9072 7040 9080 7104
rect 8760 6016 9080 7040
rect 8760 5952 8768 6016
rect 8832 5952 8848 6016
rect 8912 5952 8928 6016
rect 8992 5952 9008 6016
rect 9072 5952 9080 6016
rect 8760 5794 9080 5952
rect 8760 5558 8802 5794
rect 9038 5558 9080 5794
rect 8760 4928 9080 5558
rect 8760 4864 8768 4928
rect 8832 4864 8848 4928
rect 8912 4864 8928 4928
rect 8992 4864 9008 4928
rect 9072 4864 9080 4928
rect 8760 3840 9080 4864
rect 8760 3776 8768 3840
rect 8832 3776 8848 3840
rect 8912 3776 8928 3840
rect 8992 3776 9008 3840
rect 9072 3776 9080 3840
rect 8760 2752 9080 3776
rect 8760 2688 8768 2752
rect 8832 2694 8848 2752
rect 8912 2694 8928 2752
rect 8992 2694 9008 2752
rect 9072 2688 9080 2752
rect 8760 2458 8802 2688
rect 9038 2458 9080 2688
rect 8760 1894 9080 2458
rect 8760 1658 8802 1894
rect 9038 1658 9080 1894
rect 8760 956 9080 1658
rect 10084 11942 10404 11984
rect 10084 11706 10126 11942
rect 10362 11706 10404 11942
rect 10084 8894 10404 11706
rect 10084 8658 10126 8894
rect 10362 8658 10404 8894
rect 10084 5794 10404 8658
rect 10084 5558 10126 5794
rect 10362 5558 10404 5794
rect 10084 2694 10404 5558
rect 10084 2458 10126 2694
rect 10362 2458 10404 2694
rect 10084 1894 10404 2458
rect 10084 1658 10126 1894
rect 10362 1658 10404 1894
rect 10084 1616 10404 1658
rect 10744 10444 11064 12366
rect 10744 10208 10786 10444
rect 11022 10208 11064 10444
rect 10744 7344 11064 10208
rect 10744 7108 10786 7344
rect 11022 7108 11064 7344
rect 10744 4244 11064 7108
rect 10744 4008 10786 4244
rect 11022 4008 11064 4244
rect 10744 1234 11064 4008
rect 10744 998 10786 1234
rect 11022 998 11064 1234
rect 10744 956 11064 998
rect 11404 9794 11724 13026
rect 11404 9558 11446 9794
rect 11682 9558 11724 9794
rect 11404 6694 11724 9558
rect 11404 6458 11446 6694
rect 11682 6458 11724 6694
rect 11404 3594 11724 6458
rect 11404 3358 11446 3594
rect 11682 3358 11724 3594
rect -960 338 -918 574
rect -682 338 -640 574
rect -960 296 -640 338
rect 11404 574 11724 3358
rect 11404 338 11446 574
rect 11682 338 11724 574
rect 11404 296 11724 338
rect 12064 8244 12384 13686
rect 12064 8008 12106 8244
rect 12342 8008 12384 8244
rect 12064 5144 12384 8008
rect 12064 4908 12106 5144
rect 12342 4908 12384 5144
rect -1620 -322 -1578 -86
rect -1342 -322 -1300 -86
rect -1620 -364 -1300 -322
rect 12064 -86 12384 4908
rect 12064 -322 12106 -86
rect 12342 -322 12384 -86
rect 12064 -364 12384 -322
<< via4 >>
rect -1578 13686 -1342 13922
rect 12106 13686 12342 13922
rect -1578 8008 -1342 8244
rect -1578 4908 -1342 5144
rect -918 13026 -682 13262
rect 11446 13026 11682 13262
rect -918 9558 -682 9794
rect -918 6458 -682 6694
rect -918 3358 -682 3594
rect -258 12366 -22 12602
rect -258 10208 -22 10444
rect -258 7108 -22 7344
rect -258 4008 -22 4244
rect 402 11706 638 11942
rect 402 8658 638 8894
rect 402 5558 638 5794
rect 2602 11706 2838 11942
rect 2602 8658 2838 8894
rect 2602 5558 2838 5794
rect 2018 4908 2254 5144
rect 1278 3358 1514 3594
rect 402 2458 638 2694
rect 402 1658 638 1894
rect 2602 2458 2838 2694
rect 2602 1658 2838 1894
rect -258 998 -22 1234
rect 4152 12366 4388 12602
rect 4152 10208 4388 10444
rect 4152 7108 4388 7344
rect 4152 4008 4388 4244
rect 4152 998 4388 1234
rect 5702 11706 5938 11942
rect 5702 8658 5938 8894
rect 5702 5558 5938 5794
rect 5702 2688 5732 2694
rect 5732 2688 5748 2694
rect 5748 2688 5812 2694
rect 5812 2688 5828 2694
rect 5828 2688 5892 2694
rect 5892 2688 5908 2694
rect 5908 2688 5938 2694
rect 5702 2458 5938 2688
rect 5702 1658 5938 1894
rect 7252 12366 7488 12602
rect 7252 10208 7488 10444
rect 7252 7108 7488 7344
rect 7252 4008 7488 4244
rect 7252 998 7488 1234
rect 10786 12366 11022 12602
rect 8802 11706 9038 11942
rect 8802 8658 9038 8894
rect 8802 5558 9038 5794
rect 8802 2688 8832 2694
rect 8832 2688 8848 2694
rect 8848 2688 8912 2694
rect 8912 2688 8928 2694
rect 8928 2688 8992 2694
rect 8992 2688 9008 2694
rect 9008 2688 9038 2694
rect 8802 2458 9038 2688
rect 8802 1658 9038 1894
rect 10126 11706 10362 11942
rect 10126 8658 10362 8894
rect 10126 5558 10362 5794
rect 10126 2458 10362 2694
rect 10126 1658 10362 1894
rect 10786 10208 11022 10444
rect 10786 7108 11022 7344
rect 10786 4008 11022 4244
rect 10786 998 11022 1234
rect 11446 9558 11682 9794
rect 11446 6458 11682 6694
rect 11446 3358 11682 3594
rect -918 338 -682 574
rect 11446 338 11682 574
rect 12106 8008 12342 8244
rect 12106 4908 12342 5144
rect -1578 -322 -1342 -86
rect 12106 -322 12342 -86
<< metal5 >>
rect -1620 13922 12384 13964
rect -1620 13686 -1578 13922
rect -1342 13686 12106 13922
rect 12342 13686 12384 13922
rect -1620 13644 12384 13686
rect -960 13262 11724 13304
rect -960 13026 -918 13262
rect -682 13026 11446 13262
rect 11682 13026 11724 13262
rect -960 12984 11724 13026
rect -300 12602 11064 12644
rect -300 12366 -258 12602
rect -22 12366 4152 12602
rect 4388 12366 7252 12602
rect 7488 12366 10786 12602
rect 11022 12366 11064 12602
rect -300 12324 11064 12366
rect 360 11942 10404 11984
rect 360 11706 402 11942
rect 638 11706 2602 11942
rect 2838 11706 5702 11942
rect 5938 11706 8802 11942
rect 9038 11706 10126 11942
rect 10362 11706 10404 11942
rect 360 11664 10404 11706
rect -300 10444 11064 10486
rect -300 10208 -258 10444
rect -22 10208 4152 10444
rect 4388 10208 7252 10444
rect 7488 10208 10786 10444
rect 11022 10208 11064 10444
rect -300 10166 11064 10208
rect -1620 9794 12384 9836
rect -1620 9558 -918 9794
rect -682 9558 11446 9794
rect 11682 9558 12384 9794
rect -1620 9516 12384 9558
rect -300 8894 11064 8936
rect -300 8658 402 8894
rect 638 8658 2602 8894
rect 2838 8658 5702 8894
rect 5938 8658 8802 8894
rect 9038 8658 10126 8894
rect 10362 8658 11064 8894
rect -300 8616 11064 8658
rect -1620 8244 12384 8286
rect -1620 8008 -1578 8244
rect -1342 8008 12106 8244
rect 12342 8008 12384 8244
rect -1620 7966 12384 8008
rect -300 7344 11064 7386
rect -300 7108 -258 7344
rect -22 7108 4152 7344
rect 4388 7108 7252 7344
rect 7488 7108 10786 7344
rect 11022 7108 11064 7344
rect -300 7066 11064 7108
rect -1620 6694 12384 6736
rect -1620 6458 -918 6694
rect -682 6458 11446 6694
rect 11682 6458 12384 6694
rect -1620 6416 12384 6458
rect -300 5794 11064 5836
rect -300 5558 402 5794
rect 638 5558 2602 5794
rect 2838 5558 5702 5794
rect 5938 5558 8802 5794
rect 9038 5558 10126 5794
rect 10362 5558 11064 5794
rect -300 5516 11064 5558
rect -1620 5144 12384 5186
rect -1620 4908 -1578 5144
rect -1342 4908 2018 5144
rect 2254 4908 12106 5144
rect 12342 4908 12384 5144
rect -1620 4866 12384 4908
rect -300 4244 11064 4286
rect -300 4008 -258 4244
rect -22 4008 4152 4244
rect 4388 4008 7252 4244
rect 7488 4008 10786 4244
rect 11022 4008 11064 4244
rect -300 3966 11064 4008
rect -1620 3594 12384 3636
rect -1620 3358 -918 3594
rect -682 3358 1278 3594
rect 1514 3358 11446 3594
rect 11682 3358 12384 3594
rect -1620 3316 12384 3358
rect -300 2694 11064 2736
rect -300 2458 402 2694
rect 638 2458 2602 2694
rect 2838 2458 5702 2694
rect 5938 2458 8802 2694
rect 9038 2458 10126 2694
rect 10362 2458 11064 2694
rect -300 2416 11064 2458
rect 360 1894 10404 1936
rect 360 1658 402 1894
rect 638 1658 2602 1894
rect 2838 1658 5702 1894
rect 5938 1658 8802 1894
rect 9038 1658 10126 1894
rect 10362 1658 10404 1894
rect 360 1616 10404 1658
rect -300 1234 11064 1276
rect -300 998 -258 1234
rect -22 998 4152 1234
rect 4388 998 7252 1234
rect 7488 998 10786 1234
rect 11022 998 11064 1234
rect -300 956 11064 998
rect -960 574 11724 616
rect -960 338 -918 574
rect -682 338 11446 574
rect 11682 338 11724 574
rect -960 296 11724 338
rect -1620 -86 12384 -44
rect -1620 -322 -1578 -86
rect -1342 -322 12106 -86
rect 12342 -322 12384 -86
rect -1620 -364 12384 -322
use sky130_fd_sc_hd__dfrtp_1  _216_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 3312 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 3036 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1635271187
transform 1 0 3036 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1635271187
transform 1 0 3036 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_26 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 3312 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 3312 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _143_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 3312 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1635271187
transform 1 0 3036 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1635271187
transform 1 0 3036 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1635271187
transform 1 0 3036 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_26
timestamp 1635271187
transform 1 0 3312 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_26
timestamp 1635271187
transform 1 0 3312 0 -1 4352
box -38 -48 130 592
use gpio_logic_high  gpio_logic_high
timestamp 1636038210
transform 1 0 1196 0 1 2680
box -38 -48 1418 2768
use sky130_fd_sc_hd__dfrtp_1  _218_
timestamp 1635271187
transform 1 0 5704 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _217_
timestamp 1635271187
transform 1 0 3772 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfbbn_1  _208_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 4692 0 -1 3264
box -38 -48 2430 592
use sky130_fd_sc_hd__clkbuf_1  _148_
timestamp 1635271187
transform 1 0 3496 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _147_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 3680 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _146_
timestamp 1635271187
transform 1 0 3404 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _145_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 4140 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 5612 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _116_
timestamp 1635271187
transform 1 0 5152 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _114_
timestamp 1635271187
transform 1 0 5704 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1635271187
transform 1 0 5612 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__dfbbn_1  _210_
timestamp 1635271187
transform 1 0 5796 0 -1 4352
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbn_1  _203_
timestamp 1635271187
transform 1 0 3404 0 -1 4352
box -38 -48 2430 592
use sky130_fd_sc_hd__or2_1  _153_
timestamp 1635271187
transform 1 0 5704 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _151_
timestamp 1635271187
transform 1 0 4140 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _125_
timestamp 1635271187
transform 1 0 3588 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _113_
timestamp 1635271187
transform 1 0 3864 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _107_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 4692 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1635271187
transform 1 0 5612 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__dfbbn_1  _202_
timestamp 1635271187
transform 1 0 3404 0 -1 5440
box -38 -48 2430 592
use sky130_fd_sc_hd__fill_1  FILLER_5_53
timestamp 1635271187
transform 1 0 5796 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_67
timestamp 1635271187
transform 1 0 7084 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__or2b_1  _108_
timestamp 1635271187
transform 1 0 7452 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _111_
timestamp 1635271187
transform 1 0 7176 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _115_
timestamp 1635271187
transform 1 0 7544 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75
timestamp 1635271187
transform 1 0 7820 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_77
timestamp 1635271187
transform 1 0 8004 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1635271187
transform 1 0 8188 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1635271187
transform 1 0 8188 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__or2b_1  _102_
timestamp 1635271187
transform 1 0 8280 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _109_
timestamp 1635271187
transform 1 0 7912 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _110_
timestamp 1635271187
transform 1 0 8280 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__dfbbn_1  _209_
timestamp 1635271187
transform 1 0 6256 0 1 3264
box -38 -48 2430 592
use sky130_fd_sc_hd__clkbuf_1  _118_
timestamp 1635271187
transform 1 0 8280 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1635271187
transform 1 0 8188 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_serial_clock $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 6164 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dfbbn_1  _207_
timestamp 1635271187
transform 1 0 7176 0 1 4352
box -38 -48 2430 592
use sky130_fd_sc_hd__or2b_1  _126_
timestamp 1635271187
transform 1 0 6624 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_61
timestamp 1635271187
transform 1 0 6532 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _223_
timestamp 1635271187
transform 1 0 5888 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__or2_1  _128_
timestamp 1635271187
transform 1 0 7728 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1635271187
transform 1 0 8188 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_80
timestamp 1635271187
transform 1 0 8280 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__or2_1  _104_
timestamp 1635271187
transform 1 0 8832 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__fill_2  FILLER_1_86
timestamp 1635271187
transform 1 0 8832 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85
timestamp 1635271187
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  const_source $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 9200 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _117_
timestamp 1635271187
transform 1 0 9292 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1635271187
transform -1 0 9844 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1635271187
transform -1 0 9844 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_93
timestamp 1635271187
transform 1 0 9476 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 9016 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _105_
timestamp 1635271187
transform 1 0 8924 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _103_
timestamp 1635271187
transform 1 0 8648 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _184_
timestamp 1635271187
transform 1 0 9200 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1635271187
transform -1 0 9844 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_93
timestamp 1635271187
transform 1 0 9476 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__or2b_1  _120_
timestamp 1635271187
transform 1 0 8556 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _129_
timestamp 1635271187
transform 1 0 9108 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1635271187
transform -1 0 9844 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_92
timestamp 1635271187
transform 1 0 9384 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1635271187
transform -1 0 9844 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _122_
timestamp 1635271187
transform 1 0 8740 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _121_
timestamp 1635271187
transform 1 0 8464 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _133_
timestamp 1635271187
transform 1 0 9200 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1635271187
transform -1 0 9844 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_93
timestamp 1635271187
transform 1 0 9476 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _215_
timestamp 1635271187
transform 1 0 3312 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1635271187
transform 1 0 3036 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _214_
timestamp 1635271187
transform 1 0 3312 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1635271187
transform 1 0 3036 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3
timestamp 1635271187
transform 1 0 1196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1635271187
transform 1 0 920 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1635271187
transform 1 0 1564 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1635271187
transform 1 0 1288 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_10
timestamp 1635271187
transform 1 0 1840 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1635271187
transform 1 0 1932 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1635271187
transform 1 0 2208 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1635271187
transform 1 0 2484 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0
timestamp 1635271187
transform -1 0 3128 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_20
timestamp 1635271187
transform 1 0 2760 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1635271187
transform -1 0 3312 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1635271187
transform -1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1635271187
transform 1 0 1196 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1635271187
transform 1 0 920 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1635271187
transform 1 0 1380 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1635271187
transform -1 0 2024 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_8
timestamp 1635271187
transform 1 0 1656 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1635271187
transform -1 0 2208 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_14
timestamp 1635271187
transform 1 0 2208 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _150_
timestamp 1635271187
transform 1 0 2300 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _149_
timestamp 1635271187
transform 1 0 2576 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _144_
timestamp 1635271187
transform 1 0 2852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _135_
timestamp 1635271187
transform 1 0 3128 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1635271187
transform -1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1635271187
transform 1 0 920 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1635271187
transform -1 0 1564 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1635271187
transform 1 0 1564 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1635271187
transform 1 0 1840 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_13
timestamp 1635271187
transform 1 0 2116 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1635271187
transform 1 0 2208 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1635271187
transform 1 0 2484 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1635271187
transform -1 0 3128 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_20
timestamp 1635271187
transform 1 0 2760 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1635271187
transform -1 0 3312 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1635271187
transform -1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__dfbbn_1  _206_
timestamp 1635271187
transform 1 0 5704 0 1 5440
box -38 -48 2430 592
use sky130_fd_sc_hd__clkbuf_1  _112_
timestamp 1635271187
transform 1 0 5336 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1635271187
transform 1 0 5612 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_46
timestamp 1635271187
transform 1 0 5152 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_1  _222_
timestamp 1635271187
transform 1 0 5152 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__or2b_1  _139_
timestamp 1635271187
transform 1 0 5244 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _136_
timestamp 1635271187
transform 1 0 4140 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _124_
timestamp 1635271187
transform 1 0 5796 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1635271187
transform 1 0 3496 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_45
timestamp 1635271187
transform 1 0 5060 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_33
timestamp 1635271187
transform 1 0 3956 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1635271187
transform -1 0 3956 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1635271187
transform -1 0 3772 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__dfbbn_1  _204_
timestamp 1635271187
transform 1 0 3680 0 -1 7616
box -38 -48 2430 592
use sky130_fd_sc_hd__clkbuf_1  _131_
timestamp 1635271187
transform 1 0 3404 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dfbbn_1  _199_
timestamp 1635271187
transform 1 0 4784 0 1 7616
box -38 -48 2430 592
use sky130_fd_sc_hd__clkbuf_1  _138_
timestamp 1635271187
transform 1 0 4048 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _137_
timestamp 1635271187
transform 1 0 3772 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _130_
timestamp 1635271187
transform 1 0 4508 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1635271187
transform 1 0 3496 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_37
timestamp 1635271187
transform 1 0 4324 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1635271187
transform 1 0 3588 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_78
timestamp 1635271187
transform 1 0 8096 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1635271187
transform -1 0 8464 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__or2_1  _141_
timestamp 1635271187
transform 1 0 6992 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _134_
timestamp 1635271187
transform 1 0 7728 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _132_
timestamp 1635271187
transform 1 0 8280 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _119_
timestamp 1635271187
transform 1 0 7452 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1635271187
transform 1 0 8188 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output25 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 8280 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_serial_clock $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 6164 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  _127_
timestamp 1635271187
transform 1 0 8004 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1635271187
transform 1 0 6072 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__dfbbn_1  _205_
timestamp 1635271187
transform 1 0 6808 0 -1 7616
box -38 -48 2430 592
use sky130_fd_sc_hd__or2b_1  _169_
timestamp 1635271187
transform 1 0 6164 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1635271187
transform 1 0 6072 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_63
timestamp 1635271187
transform 1 0 6716 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 1635271187
transform 1 0 7360 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp 1635271187
transform 1 0 8280 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _179_
timestamp 1635271187
transform 1 0 7728 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_68
timestamp 1635271187
transform 1 0 7176 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 1635271187
transform 1 0 9200 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _186_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 8464 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _123_
timestamp 1635271187
transform 1 0 8924 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1635271187
transform -1 0 9844 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _183_
timestamp 1635271187
transform 1 0 8832 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1635271187
transform -1 0 9844 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_92
timestamp 1635271187
transform 1 0 9384 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _194_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 8740 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1635271187
transform 1 0 8648 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1635271187
transform -1 0 9844 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output24
timestamp 1635271187
transform 1 0 9200 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1635271187
transform -1 0 9844 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _195_
timestamp 1635271187
transform 1 0 8740 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1635271187
transform 1 0 8648 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1635271187
transform -1 0 9844 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_12
timestamp 1635271187
transform 1 0 2024 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1635271187
transform 1 0 920 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _170_
timestamp 1635271187
transform 1 0 1748 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _172_
timestamp 1635271187
transform 1 0 1472 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _180_
timestamp 1635271187
transform 1 0 1196 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1635271187
transform -1 0 2392 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_19
timestamp 1635271187
transform 1 0 2668 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _168_
timestamp 1635271187
transform 1 0 2760 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1635271187
transform 1 0 2392 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _213_
timestamp 1635271187
transform 1 0 3036 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_12_3
timestamp 1635271187
transform 1 0 1196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1635271187
transform 1 0 920 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1635271187
transform 1 0 1288 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1635271187
transform 1 0 1472 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _185_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 1748 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_15
timestamp 1635271187
transform 1 0 2300 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _178_
timestamp 1635271187
transform 1 0 2024 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1635271187
transform 1 0 2484 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1635271187
transform 1 0 2668 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _167_
timestamp 1635271187
transform 1 0 2944 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _164_
timestamp 1635271187
transform 1 0 3220 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1635271187
transform 1 0 1288 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1635271187
transform 1 0 1564 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _212_
timestamp 1635271187
transform 1 0 2760 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  _189_
timestamp 1635271187
transform 1 0 2208 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _182_
timestamp 1635271187
transform 1 0 2484 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1635271187
transform 1 0 920 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3
timestamp 1635271187
transform 1 0 1196 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_10
timestamp 1635271187
transform 1 0 1840 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1635271187
transform 1 0 2024 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1635271187
transform 1 0 1932 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 1196 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_3
timestamp 1635271187
transform 1 0 1196 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_9
timestamp 1635271187
transform 1 0 1748 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1635271187
transform 1 0 920 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1635271187
transform 1 0 920 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1635271187
transform 1 0 2116 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output37
timestamp 1635271187
transform 1 0 1472 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_15
timestamp 1635271187
transform 1 0 2300 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _176_
timestamp 1635271187
transform 1 0 3220 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _188_
timestamp 1635271187
transform 1 0 2944 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _190_
timestamp 1635271187
transform 1 0 2392 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _192_
timestamp 1635271187
transform 1 0 2668 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1635271187
transform 1 0 2392 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _219_
timestamp 1635271187
transform 1 0 2668 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_serial_clock
timestamp 1635271187
transform 1 0 5704 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _165_
timestamp 1635271187
transform 1 0 5244 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _140_
timestamp 1635271187
transform 1 0 4876 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_46
timestamp 1635271187
transform 1 0 5152 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__dfbbn_1  _201_
timestamp 1635271187
transform 1 0 5152 0 1 8704
box -38 -48 2430 592
use sky130_fd_sc_hd__clkbuf_1  _161_
timestamp 1635271187
transform 1 0 3588 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _158_
timestamp 1635271187
transform 1 0 3864 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _154_
timestamp 1635271187
transform 1 0 4140 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _152_
timestamp 1635271187
transform 1 0 4416 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _142_
timestamp 1635271187
transform 1 0 4876 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1635271187
transform 1 0 3496 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_41
timestamp 1635271187
transform 1 0 4692 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__or2b_1  _163_
timestamp 1635271187
transform 1 0 4876 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _159_
timestamp 1635271187
transform 1 0 5612 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _155_
timestamp 1635271187
transform 1 0 4600 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_49
timestamp 1635271187
transform 1 0 5428 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_29
timestamp 1635271187
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_39
timestamp 1635271187
transform 1 0 4508 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1635271187
transform 1 0 3496 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _156_
timestamp 1635271187
transform 1 0 4600 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _162_
timestamp 1635271187
transform 1 0 3680 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _160_
timestamp 1635271187
transform 1 0 5428 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _166_
timestamp 1635271187
transform 1 0 5152 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _173_
timestamp 1635271187
transform 1 0 4876 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output40
timestamp 1635271187
transform 1 0 5704 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dfbbn_1  _200_
timestamp 1635271187
transform 1 0 3956 0 1 9792
box -38 -48 2430 592
use sky130_fd_sc_hd__buf_2  output30
timestamp 1635271187
transform 1 0 6716 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output28
timestamp 1635271187
transform 1 0 7728 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_2  gpio_in_buf $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 7084 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _181_
timestamp 1635271187
transform 1 0 8188 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _171_
timestamp 1635271187
transform 1 0 6256 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1635271187
transform 1 0 6072 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_78
timestamp 1635271187
transform 1 0 8096 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_57
timestamp 1635271187
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output29
timestamp 1635271187
transform 1 0 7728 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _175_
timestamp 1635271187
transform 1 0 8096 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_72
timestamp 1635271187
transform 1 0 7544 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__dfbbn_1  _198_
timestamp 1635271187
transform 1 0 6992 0 -1 9792
box -38 -48 2430 592
use sky130_fd_sc_hd__or2b_1  _157_
timestamp 1635271187
transform 1 0 6348 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1635271187
transform 1 0 6072 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_65
timestamp 1635271187
transform 1 0 6900 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_57
timestamp 1635271187
transform 1 0 6164 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  output39
timestamp 1635271187
transform 1 0 6164 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _221_
timestamp 1635271187
transform 1 0 6348 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _211_
timestamp 1635271187
transform 1 0 6532 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__or2_1  _177_
timestamp 1635271187
transform 1 0 8188 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1635271187
transform 1 0 6072 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__ebufn_1  _197_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 8648 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1635271187
transform -1 0 9844 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_92
timestamp 1635271187
transform 1 0 9384 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _193_
timestamp 1635271187
transform 1 0 8740 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1635271187
transform 1 0 8648 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1635271187
transform -1 0 9844 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1635271187
transform -1 0 9844 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_92
timestamp 1635271187
transform 1 0 9384 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  output33
timestamp 1635271187
transform 1 0 8464 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp 1635271187
transform 1 0 9200 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _196_
timestamp 1635271187
transform 1 0 8740 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _191_
timestamp 1635271187
transform 1 0 8832 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1635271187
transform 1 0 8648 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_81
timestamp 1635271187
transform 1 0 8372 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1635271187
transform -1 0 9844 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1635271187
transform -1 0 9844 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1635271187
transform 1 0 1288 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1635271187
transform 1 0 920 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_7
timestamp 1635271187
transform 1 0 1564 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_3
timestamp 1635271187
transform 1 0 1196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1635271187
transform 1 0 2300 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_13
timestamp 1635271187
transform 1 0 2116 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1635271187
transform -1 0 1932 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1635271187
transform -1 0 2116 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1635271187
transform 1 0 2944 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_18
timestamp 1635271187
transform 1 0 2576 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1635271187
transform -1 0 2944 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _187_
timestamp 1635271187
transform 1 0 3220 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1635271187
transform 1 0 3496 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _174_
timestamp 1635271187
transform 1 0 5428 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _220_
timestamp 1635271187
transform 1 0 3588 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_2  output38
timestamp 1635271187
transform 1 0 5704 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1635271187
transform 1 0 6072 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _106_
timestamp 1635271187
transform 1 0 6164 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  input17 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 7176 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  output35
timestamp 1635271187
transform 1 0 6808 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output36
timestamp 1635271187
transform 1 0 6440 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_85
timestamp 1635271187
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1635271187
transform -1 0 9844 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1635271187
transform 1 0 8648 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output32
timestamp 1635271187
transform 1 0 9200 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp 1635271187
transform 1 0 8832 0 1 10880
box -38 -48 406 592
<< labels >>
rlabel metal3 s 14000 144 34000 264 6 gpio_defaults[0]
port 0 nsew signal input
rlabel metal3 s 14000 3272 34000 3392 6 gpio_defaults[10]
port 1 nsew signal input
rlabel metal3 s 14000 3680 34000 3800 6 gpio_defaults[11]
port 2 nsew signal input
rlabel metal3 s 14000 3952 34000 4072 6 gpio_defaults[12]
port 3 nsew signal input
rlabel metal3 s 14000 416 34000 536 6 gpio_defaults[1]
port 4 nsew signal input
rlabel metal3 s 14000 688 34000 808 6 gpio_defaults[2]
port 5 nsew signal input
rlabel metal3 s 14000 1096 34000 1216 6 gpio_defaults[3]
port 6 nsew signal input
rlabel metal3 s 14000 1368 34000 1488 6 gpio_defaults[4]
port 7 nsew signal input
rlabel metal3 s 14000 1640 34000 1760 6 gpio_defaults[5]
port 8 nsew signal input
rlabel metal3 s 14000 2048 34000 2168 6 gpio_defaults[6]
port 9 nsew signal input
rlabel metal3 s 14000 2320 34000 2440 6 gpio_defaults[7]
port 10 nsew signal input
rlabel metal3 s 14000 2728 34000 2848 6 gpio_defaults[8]
port 11 nsew signal input
rlabel metal3 s 14000 3000 34000 3120 6 gpio_defaults[9]
port 12 nsew signal input
rlabel metal3 s 14000 4904 34000 5024 6 mgmt_gpio_in
port 13 nsew signal tristate
rlabel metal3 s 14000 5312 34000 5432 6 mgmt_gpio_oeb
port 14 nsew signal input
rlabel metal3 s 14000 5584 34000 5704 6 mgmt_gpio_out
port 15 nsew signal input
rlabel metal3 s 14000 4632 34000 4752 6 one
port 16 nsew signal tristate
rlabel metal3 s 14000 5992 34000 6112 6 pad_gpio_ana_en
port 17 nsew signal tristate
rlabel metal3 s 14000 6264 34000 6384 6 pad_gpio_ana_pol
port 18 nsew signal tristate
rlabel metal3 s 14000 6536 34000 6656 6 pad_gpio_ana_sel
port 19 nsew signal tristate
rlabel metal3 s 14000 6944 34000 7064 6 pad_gpio_dm[0]
port 20 nsew signal tristate
rlabel metal3 s 14000 7216 34000 7336 6 pad_gpio_dm[1]
port 21 nsew signal tristate
rlabel metal3 s 14000 7624 34000 7744 6 pad_gpio_dm[2]
port 22 nsew signal tristate
rlabel metal3 s 14000 7896 34000 8016 6 pad_gpio_holdover
port 23 nsew signal tristate
rlabel metal3 s 14000 8168 34000 8288 6 pad_gpio_ib_mode_sel
port 24 nsew signal tristate
rlabel metal3 s 14000 8576 34000 8696 6 pad_gpio_in
port 25 nsew signal input
rlabel metal3 s 14000 8848 34000 8968 6 pad_gpio_inenb
port 26 nsew signal tristate
rlabel metal3 s 14000 9256 34000 9376 6 pad_gpio_out
port 27 nsew signal tristate
rlabel metal3 s 14000 9528 34000 9648 6 pad_gpio_outenb
port 28 nsew signal tristate
rlabel metal3 s 14000 9800 34000 9920 6 pad_gpio_slow_sel
port 29 nsew signal tristate
rlabel metal3 s 14000 10208 34000 10328 6 pad_gpio_vtrip_sel
port 30 nsew signal tristate
rlabel metal3 s 14000 10480 34000 10600 6 resetn
port 31 nsew signal input
rlabel metal3 s 14000 10888 34000 11008 6 resetn_out
port 32 nsew signal tristate
rlabel metal3 s 14000 11160 34000 11280 6 serial_clock
port 33 nsew signal input
rlabel metal3 s 14000 11432 34000 11552 6 serial_clock_out
port 34 nsew signal tristate
rlabel metal3 s 14000 11840 34000 11960 6 serial_data_in
port 35 nsew signal input
rlabel metal3 s 14000 12112 34000 12232 6 serial_data_out
port 36 nsew signal tristate
rlabel metal3 s 14000 12520 34000 12640 6 serial_load
port 37 nsew signal input
rlabel metal3 s 14000 12792 34000 12912 6 serial_load_out
port 38 nsew signal tristate
rlabel metal3 s 14000 13064 34000 13184 6 user_gpio_in
port 39 nsew signal tristate
rlabel metal3 s 14000 13472 34000 13592 6 user_gpio_oeb
port 40 nsew signal input
rlabel metal3 s 14000 13744 34000 13864 6 user_gpio_out
port 41 nsew signal input
rlabel metal5 s 360 1616 10404 1936 6 vccd
port 42 nsew power input
rlabel metal5 s -300 2416 11064 2736 6 vccd
port 42 nsew power input
rlabel metal5 s -300 5516 11064 5836 6 vccd
port 42 nsew power input
rlabel metal5 s -300 8616 11064 8936 6 vccd
port 42 nsew power input
rlabel metal5 s 360 11664 10404 11984 6 vccd
port 42 nsew power input
rlabel metal4 s 360 1616 680 11984 6 vccd
port 42 nsew power input
rlabel metal4 s 10084 1616 10404 11984 6 vccd
port 42 nsew power input
rlabel metal4 s 2560 956 2880 12644 6 vccd
port 42 nsew power input
rlabel metal4 s 5660 956 5980 12644 6 vccd
port 42 nsew power input
rlabel metal4 s 8760 956 9080 12644 6 vccd
port 42 nsew power input
rlabel metal5 s -960 296 11724 616 6 vccd1
port 43 nsew power input
rlabel metal5 s -1620 3316 12384 3636 6 vccd1
port 43 nsew power input
rlabel metal5 s -1620 6416 12384 6736 6 vccd1
port 43 nsew power input
rlabel metal5 s -1620 9516 12384 9836 6 vccd1
port 43 nsew power input
rlabel metal5 s -960 12984 11724 13304 6 vccd1
port 43 nsew power input
rlabel metal4 s -960 296 -640 13304 4 vccd1
port 43 nsew power input
rlabel metal4 s 11404 296 11724 13304 6 vccd1
port 43 nsew power input
rlabel metal5 s -300 956 11064 1276 6 vssd
port 44 nsew ground input
rlabel metal5 s -300 3966 11064 4286 6 vssd
port 44 nsew ground input
rlabel metal5 s -300 7066 11064 7386 6 vssd
port 44 nsew ground input
rlabel metal5 s -300 10166 11064 10486 6 vssd
port 44 nsew ground input
rlabel metal5 s -300 12324 11064 12644 6 vssd
port 44 nsew ground input
rlabel metal4 s -300 956 20 12644 4 vssd
port 44 nsew ground input
rlabel metal4 s 4110 956 4430 12644 6 vssd
port 44 nsew ground input
rlabel metal4 s 7210 956 7530 12644 6 vssd
port 44 nsew ground input
rlabel metal4 s 10744 956 11064 12644 6 vssd
port 44 nsew ground input
rlabel metal5 s -1620 -364 12384 -44 8 vssd1
port 45 nsew ground input
rlabel metal5 s -1620 4866 12384 5186 6 vssd1
port 45 nsew ground input
rlabel metal5 s -1620 7966 12384 8286 6 vssd1
port 45 nsew ground input
rlabel metal5 s -1620 13644 12384 13964 6 vssd1
port 45 nsew ground input
rlabel metal4 s -1620 -364 -1300 13964 4 vssd1
port 45 nsew ground input
rlabel metal4 s 12064 -364 12384 13964 6 vssd1
port 45 nsew ground input
rlabel metal3 s 14000 4360 34000 4480 6 zero
port 46 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 34000 14000
<< end >>
