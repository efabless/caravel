magic
tech sky130A
magscale 1 2
timestamp 1675162640
<< viali >>
rect 2145 7361 2179 7395
rect 7113 7361 7147 7395
rect 6469 6953 6503 6987
rect 1593 6817 1627 6851
rect 3341 6817 3375 6851
rect 5917 6817 5951 6851
rect 2145 6749 2179 6783
rect 2973 6749 3007 6783
rect 3157 6749 3191 6783
rect 6561 6749 6595 6783
rect 7021 6749 7055 6783
rect 1685 6273 1719 6307
rect 1961 6273 1995 6307
rect 3249 6273 3283 6307
rect 7113 6273 7147 6307
rect 1593 6205 1627 6239
rect 2421 6205 2455 6239
rect 7205 6069 7239 6103
rect 7205 5865 7239 5899
rect 6837 5729 6871 5763
rect 1593 5661 1627 5695
rect 6653 5593 6687 5627
rect 6745 5525 6779 5559
rect 6561 4981 6595 5015
rect 1961 4777 1995 4811
rect 7113 4777 7147 4811
rect 2421 4709 2455 4743
rect 6653 4709 6687 4743
rect 1777 4165 1811 4199
rect 1961 4165 1995 4199
rect 1685 4097 1719 4131
rect 7021 4097 7055 4131
rect 7297 4097 7331 4131
rect 6929 4029 6963 4063
rect 2237 3961 2271 3995
rect 2789 3893 2823 3927
rect 6469 3689 6503 3723
rect 7297 3689 7331 3723
rect 1593 3485 1627 3519
rect 3985 3145 4019 3179
rect 2329 3009 2363 3043
rect 3801 3009 3835 3043
rect 7297 3009 7331 3043
rect 1961 2941 1995 2975
rect 4261 2805 4295 2839
rect 7205 2805 7239 2839
rect 5181 2601 5215 2635
rect 5825 2601 5859 2635
rect 1961 2465 1995 2499
rect 2605 2397 2639 2431
rect 7297 2397 7331 2431
rect 4261 2057 4295 2091
rect 4077 1921 4111 1955
rect 5641 1921 5675 1955
rect 5825 1921 5859 1955
rect 6561 1921 6595 1955
rect 2237 1853 2271 1887
rect 2605 1853 2639 1887
rect 5917 1853 5951 1887
rect 1593 1717 1627 1751
rect 4537 1717 4571 1751
rect 5273 1513 5307 1547
rect 1593 1377 1627 1411
rect 3249 1377 3283 1411
rect 3985 1377 4019 1411
rect 7113 1309 7147 1343
rect 7205 1173 7239 1207
<< metal1 >>
rect 2866 7896 2872 7948
rect 2924 7936 2930 7948
rect 5718 7936 5724 7948
rect 2924 7908 5724 7936
rect 2924 7896 2930 7908
rect 5718 7896 5724 7908
rect 5776 7896 5782 7948
rect 1104 7642 7820 7664
rect 1104 7590 3150 7642
rect 3202 7590 3214 7642
rect 3266 7590 3278 7642
rect 3330 7590 3342 7642
rect 3394 7590 3406 7642
rect 3458 7590 7150 7642
rect 7202 7590 7214 7642
rect 7266 7590 7278 7642
rect 7330 7590 7342 7642
rect 7394 7590 7406 7642
rect 7458 7590 7820 7642
rect 1104 7568 7820 7590
rect 2130 7392 2136 7404
rect 2091 7364 2136 7392
rect 2130 7352 2136 7364
rect 2188 7352 2194 7404
rect 6822 7352 6828 7404
rect 6880 7392 6886 7404
rect 7101 7395 7159 7401
rect 7101 7392 7113 7395
rect 6880 7364 7113 7392
rect 6880 7352 6886 7364
rect 7101 7361 7113 7364
rect 7147 7392 7159 7395
rect 7558 7392 7564 7404
rect 7147 7364 7564 7392
rect 7147 7361 7159 7364
rect 7101 7355 7159 7361
rect 7558 7352 7564 7364
rect 7616 7352 7622 7404
rect 1104 7098 7820 7120
rect 1104 7046 1150 7098
rect 1202 7046 1214 7098
rect 1266 7046 1278 7098
rect 1330 7046 1342 7098
rect 1394 7046 1406 7098
rect 1458 7046 5150 7098
rect 5202 7046 5214 7098
rect 5266 7046 5278 7098
rect 5330 7046 5342 7098
rect 5394 7046 5406 7098
rect 5458 7046 7820 7098
rect 1104 7024 7820 7046
rect 14 6944 20 6996
rect 72 6984 78 6996
rect 6457 6987 6515 6993
rect 6457 6984 6469 6987
rect 72 6956 6469 6984
rect 72 6944 78 6956
rect 6457 6953 6469 6956
rect 6503 6953 6515 6987
rect 6457 6947 6515 6953
rect 1578 6848 1584 6860
rect 1539 6820 1584 6848
rect 1578 6808 1584 6820
rect 1636 6808 1642 6860
rect 3329 6851 3387 6857
rect 3329 6817 3341 6851
rect 3375 6848 3387 6851
rect 4246 6848 4252 6860
rect 3375 6820 4252 6848
rect 3375 6817 3387 6820
rect 3329 6811 3387 6817
rect 4246 6808 4252 6820
rect 4304 6808 4310 6860
rect 5905 6851 5963 6857
rect 5905 6817 5917 6851
rect 5951 6848 5963 6851
rect 6730 6848 6736 6860
rect 5951 6820 6736 6848
rect 5951 6817 5963 6820
rect 5905 6811 5963 6817
rect 6730 6808 6736 6820
rect 6788 6808 6794 6860
rect 2130 6780 2136 6792
rect 2091 6752 2136 6780
rect 2130 6740 2136 6752
rect 2188 6740 2194 6792
rect 2774 6740 2780 6792
rect 2832 6780 2838 6792
rect 2961 6783 3019 6789
rect 2961 6780 2973 6783
rect 2832 6752 2973 6780
rect 2832 6740 2838 6752
rect 2961 6749 2973 6752
rect 3007 6749 3019 6783
rect 2961 6743 3019 6749
rect 3050 6740 3056 6792
rect 3108 6780 3114 6792
rect 3145 6783 3203 6789
rect 3145 6780 3157 6783
rect 3108 6752 3157 6780
rect 3108 6740 3114 6752
rect 3145 6749 3157 6752
rect 3191 6749 3203 6783
rect 3145 6743 3203 6749
rect 6549 6783 6607 6789
rect 6549 6749 6561 6783
rect 6595 6780 6607 6783
rect 7009 6783 7067 6789
rect 7009 6780 7021 6783
rect 6595 6752 7021 6780
rect 6595 6749 6607 6752
rect 6549 6743 6607 6749
rect 7009 6749 7021 6752
rect 7055 6780 7067 6783
rect 8386 6780 8392 6792
rect 7055 6752 8392 6780
rect 7055 6749 7067 6752
rect 7009 6743 7067 6749
rect 8386 6740 8392 6752
rect 8444 6740 8450 6792
rect 1104 6554 7820 6576
rect 1104 6502 3150 6554
rect 3202 6502 3214 6554
rect 3266 6502 3278 6554
rect 3330 6502 3342 6554
rect 3394 6502 3406 6554
rect 3458 6502 7150 6554
rect 7202 6502 7214 6554
rect 7266 6502 7278 6554
rect 7330 6502 7342 6554
rect 7394 6502 7406 6554
rect 7458 6502 7820 6554
rect 1104 6480 7820 6502
rect 1673 6307 1731 6313
rect 1673 6273 1685 6307
rect 1719 6273 1731 6307
rect 1673 6267 1731 6273
rect 1949 6307 2007 6313
rect 1949 6273 1961 6307
rect 1995 6273 2007 6307
rect 1949 6267 2007 6273
rect 1578 6236 1584 6248
rect 1539 6208 1584 6236
rect 1578 6196 1584 6208
rect 1636 6196 1642 6248
rect 1688 6168 1716 6267
rect 1964 6236 1992 6267
rect 3050 6264 3056 6316
rect 3108 6304 3114 6316
rect 3237 6307 3295 6313
rect 3237 6304 3249 6307
rect 3108 6276 3249 6304
rect 3108 6264 3114 6276
rect 3237 6273 3249 6276
rect 3283 6273 3295 6307
rect 3237 6267 3295 6273
rect 6730 6264 6736 6316
rect 6788 6304 6794 6316
rect 7101 6307 7159 6313
rect 7101 6304 7113 6307
rect 6788 6276 7113 6304
rect 6788 6264 6794 6276
rect 7101 6273 7113 6276
rect 7147 6273 7159 6307
rect 7101 6267 7159 6273
rect 2409 6239 2467 6245
rect 2409 6236 2421 6239
rect 1964 6208 2421 6236
rect 2409 6205 2421 6208
rect 2455 6236 2467 6239
rect 4798 6236 4804 6248
rect 2455 6208 4804 6236
rect 2455 6205 2467 6208
rect 2409 6199 2467 6205
rect 4798 6196 4804 6208
rect 4856 6196 4862 6248
rect 1596 6140 1716 6168
rect 1596 6112 1624 6140
rect 1578 6060 1584 6112
rect 1636 6060 1642 6112
rect 7193 6103 7251 6109
rect 7193 6069 7205 6103
rect 7239 6100 7251 6103
rect 7558 6100 7564 6112
rect 7239 6072 7564 6100
rect 7239 6069 7251 6072
rect 7193 6063 7251 6069
rect 7558 6060 7564 6072
rect 7616 6060 7622 6112
rect 1104 6010 7820 6032
rect 1104 5958 1150 6010
rect 1202 5958 1214 6010
rect 1266 5958 1278 6010
rect 1330 5958 1342 6010
rect 1394 5958 1406 6010
rect 1458 5958 5150 6010
rect 5202 5958 5214 6010
rect 5266 5958 5278 6010
rect 5330 5958 5342 6010
rect 5394 5958 5406 6010
rect 5458 5958 7820 6010
rect 1104 5936 7820 5958
rect 7006 5856 7012 5908
rect 7064 5896 7070 5908
rect 7193 5899 7251 5905
rect 7193 5896 7205 5899
rect 7064 5868 7205 5896
rect 7064 5856 7070 5868
rect 7193 5865 7205 5868
rect 7239 5865 7251 5899
rect 7193 5859 7251 5865
rect 6822 5760 6828 5772
rect 6783 5732 6828 5760
rect 6822 5720 6828 5732
rect 6880 5720 6886 5772
rect 1578 5692 1584 5704
rect 1539 5664 1584 5692
rect 1578 5652 1584 5664
rect 1636 5652 1642 5704
rect 6641 5627 6699 5633
rect 6641 5593 6653 5627
rect 6687 5624 6699 5627
rect 6822 5624 6828 5636
rect 6687 5596 6828 5624
rect 6687 5593 6699 5596
rect 6641 5587 6699 5593
rect 6822 5584 6828 5596
rect 6880 5584 6886 5636
rect 6546 5516 6552 5568
rect 6604 5556 6610 5568
rect 6733 5559 6791 5565
rect 6733 5556 6745 5559
rect 6604 5528 6745 5556
rect 6604 5516 6610 5528
rect 6733 5525 6745 5528
rect 6779 5525 6791 5559
rect 6733 5519 6791 5525
rect 1104 5466 7820 5488
rect 1104 5414 3150 5466
rect 3202 5414 3214 5466
rect 3266 5414 3278 5466
rect 3330 5414 3342 5466
rect 3394 5414 3406 5466
rect 3458 5414 7150 5466
rect 7202 5414 7214 5466
rect 7266 5414 7278 5466
rect 7330 5414 7342 5466
rect 7394 5414 7406 5466
rect 7458 5414 7820 5466
rect 1104 5392 7820 5414
rect 6546 5012 6552 5024
rect 6507 4984 6552 5012
rect 6546 4972 6552 4984
rect 6604 4972 6610 5024
rect 1104 4922 7820 4944
rect 1104 4870 1150 4922
rect 1202 4870 1214 4922
rect 1266 4870 1278 4922
rect 1330 4870 1342 4922
rect 1394 4870 1406 4922
rect 1458 4870 5150 4922
rect 5202 4870 5214 4922
rect 5266 4870 5278 4922
rect 5330 4870 5342 4922
rect 5394 4870 5406 4922
rect 5458 4870 7820 4922
rect 1104 4848 7820 4870
rect 1946 4808 1952 4820
rect 1907 4780 1952 4808
rect 1946 4768 1952 4780
rect 2004 4768 2010 4820
rect 6822 4768 6828 4820
rect 6880 4808 6886 4820
rect 7101 4811 7159 4817
rect 7101 4808 7113 4811
rect 6880 4780 7113 4808
rect 6880 4768 6886 4780
rect 7101 4777 7113 4780
rect 7147 4777 7159 4811
rect 7101 4771 7159 4777
rect 1486 4700 1492 4752
rect 1544 4740 1550 4752
rect 2409 4743 2467 4749
rect 2409 4740 2421 4743
rect 1544 4712 2421 4740
rect 1544 4700 1550 4712
rect 2409 4709 2421 4712
rect 2455 4709 2467 4743
rect 2409 4703 2467 4709
rect 6641 4743 6699 4749
rect 6641 4709 6653 4743
rect 6687 4740 6699 4743
rect 7006 4740 7012 4752
rect 6687 4712 7012 4740
rect 6687 4709 6699 4712
rect 6641 4703 6699 4709
rect 7006 4700 7012 4712
rect 7064 4740 7070 4752
rect 7742 4740 7748 4752
rect 7064 4712 7748 4740
rect 7064 4700 7070 4712
rect 7742 4700 7748 4712
rect 7800 4700 7806 4752
rect 1104 4378 7820 4400
rect 1104 4326 3150 4378
rect 3202 4326 3214 4378
rect 3266 4326 3278 4378
rect 3330 4326 3342 4378
rect 3394 4326 3406 4378
rect 3458 4326 7150 4378
rect 7202 4326 7214 4378
rect 7266 4326 7278 4378
rect 7330 4326 7342 4378
rect 7394 4326 7406 4378
rect 7458 4326 7820 4378
rect 1104 4304 7820 4326
rect 1578 4156 1584 4208
rect 1636 4196 1642 4208
rect 1765 4199 1823 4205
rect 1765 4196 1777 4199
rect 1636 4168 1777 4196
rect 1636 4156 1642 4168
rect 1765 4165 1777 4168
rect 1811 4165 1823 4199
rect 1946 4196 1952 4208
rect 1907 4168 1952 4196
rect 1765 4159 1823 4165
rect 1946 4156 1952 4168
rect 2004 4156 2010 4208
rect 4062 4156 4068 4208
rect 4120 4196 4126 4208
rect 6454 4196 6460 4208
rect 4120 4168 6460 4196
rect 4120 4156 4126 4168
rect 6454 4156 6460 4168
rect 6512 4156 6518 4208
rect 1486 4088 1492 4140
rect 1544 4128 1550 4140
rect 1673 4131 1731 4137
rect 1673 4128 1685 4131
rect 1544 4100 1685 4128
rect 1544 4088 1550 4100
rect 1673 4097 1685 4100
rect 1719 4097 1731 4131
rect 7006 4128 7012 4140
rect 6967 4100 7012 4128
rect 1673 4091 1731 4097
rect 7006 4088 7012 4100
rect 7064 4088 7070 4140
rect 7282 4128 7288 4140
rect 7243 4100 7288 4128
rect 7282 4088 7288 4100
rect 7340 4088 7346 4140
rect 1026 4020 1032 4072
rect 1084 4060 1090 4072
rect 6917 4063 6975 4069
rect 6917 4060 6929 4063
rect 1084 4032 6929 4060
rect 1084 4020 1090 4032
rect 6917 4029 6929 4032
rect 6963 4029 6975 4063
rect 6917 4023 6975 4029
rect 2225 3995 2283 4001
rect 2225 3961 2237 3995
rect 2271 3992 2283 3995
rect 4982 3992 4988 4004
rect 2271 3964 4988 3992
rect 2271 3961 2283 3964
rect 2225 3955 2283 3961
rect 4982 3952 4988 3964
rect 5040 3952 5046 4004
rect 2774 3924 2780 3936
rect 2735 3896 2780 3924
rect 2774 3884 2780 3896
rect 2832 3884 2838 3936
rect 1104 3834 7820 3856
rect 1104 3782 1150 3834
rect 1202 3782 1214 3834
rect 1266 3782 1278 3834
rect 1330 3782 1342 3834
rect 1394 3782 1406 3834
rect 1458 3782 5150 3834
rect 5202 3782 5214 3834
rect 5266 3782 5278 3834
rect 5330 3782 5342 3834
rect 5394 3782 5406 3834
rect 5458 3782 7820 3834
rect 1104 3760 7820 3782
rect 6454 3720 6460 3732
rect 6415 3692 6460 3720
rect 6454 3680 6460 3692
rect 6512 3720 6518 3732
rect 7006 3720 7012 3732
rect 6512 3692 7012 3720
rect 6512 3680 6518 3692
rect 7006 3680 7012 3692
rect 7064 3680 7070 3732
rect 7282 3720 7288 3732
rect 7243 3692 7288 3720
rect 7282 3680 7288 3692
rect 7340 3680 7346 3732
rect 14 3612 20 3664
rect 72 3652 78 3664
rect 6546 3652 6552 3664
rect 72 3624 6552 3652
rect 72 3612 78 3624
rect 6546 3612 6552 3624
rect 6604 3612 6610 3664
rect 1578 3516 1584 3528
rect 1539 3488 1584 3516
rect 1578 3476 1584 3488
rect 1636 3476 1642 3528
rect 1104 3290 7820 3312
rect 1104 3238 3150 3290
rect 3202 3238 3214 3290
rect 3266 3238 3278 3290
rect 3330 3238 3342 3290
rect 3394 3238 3406 3290
rect 3458 3238 7150 3290
rect 7202 3238 7214 3290
rect 7266 3238 7278 3290
rect 7330 3238 7342 3290
rect 7394 3238 7406 3290
rect 7458 3238 7820 3290
rect 1104 3216 7820 3238
rect 3973 3179 4031 3185
rect 3973 3145 3985 3179
rect 4019 3176 4031 3179
rect 4522 3176 4528 3188
rect 4019 3148 4528 3176
rect 4019 3145 4031 3148
rect 3973 3139 4031 3145
rect 4522 3136 4528 3148
rect 4580 3136 4586 3188
rect 2590 3068 2596 3120
rect 2648 3108 2654 3120
rect 2648 3080 2714 3108
rect 2648 3068 2654 3080
rect 1486 3000 1492 3052
rect 1544 3040 1550 3052
rect 2317 3043 2375 3049
rect 2317 3040 2329 3043
rect 1544 3012 2329 3040
rect 1544 3000 1550 3012
rect 2317 3009 2329 3012
rect 2363 3009 2375 3043
rect 2317 3003 2375 3009
rect 3789 3043 3847 3049
rect 3789 3009 3801 3043
rect 3835 3040 3847 3043
rect 5074 3040 5080 3052
rect 3835 3012 5080 3040
rect 3835 3009 3847 3012
rect 3789 3003 3847 3009
rect 5074 3000 5080 3012
rect 5132 3000 5138 3052
rect 7282 3040 7288 3052
rect 7243 3012 7288 3040
rect 7282 3000 7288 3012
rect 7340 3000 7346 3052
rect 1946 2972 1952 2984
rect 1907 2944 1952 2972
rect 1946 2932 1952 2944
rect 2004 2932 2010 2984
rect 4154 2796 4160 2848
rect 4212 2836 4218 2848
rect 4249 2839 4307 2845
rect 4249 2836 4261 2839
rect 4212 2808 4261 2836
rect 4212 2796 4218 2808
rect 4249 2805 4261 2808
rect 4295 2805 4307 2839
rect 4249 2799 4307 2805
rect 7193 2839 7251 2845
rect 7193 2805 7205 2839
rect 7239 2836 7251 2839
rect 7834 2836 7840 2848
rect 7239 2808 7840 2836
rect 7239 2805 7251 2808
rect 7193 2799 7251 2805
rect 7834 2796 7840 2808
rect 7892 2796 7898 2848
rect 1104 2746 7820 2768
rect 1104 2694 1150 2746
rect 1202 2694 1214 2746
rect 1266 2694 1278 2746
rect 1330 2694 1342 2746
rect 1394 2694 1406 2746
rect 1458 2694 5150 2746
rect 5202 2694 5214 2746
rect 5266 2694 5278 2746
rect 5330 2694 5342 2746
rect 5394 2694 5406 2746
rect 5458 2694 7820 2746
rect 1104 2672 7820 2694
rect 5074 2592 5080 2644
rect 5132 2632 5138 2644
rect 5169 2635 5227 2641
rect 5169 2632 5181 2635
rect 5132 2604 5181 2632
rect 5132 2592 5138 2604
rect 5169 2601 5181 2604
rect 5215 2601 5227 2635
rect 5169 2595 5227 2601
rect 5718 2592 5724 2644
rect 5776 2632 5782 2644
rect 5813 2635 5871 2641
rect 5813 2632 5825 2635
rect 5776 2604 5825 2632
rect 5776 2592 5782 2604
rect 5813 2601 5825 2604
rect 5859 2601 5871 2635
rect 5813 2595 5871 2601
rect 1946 2496 1952 2508
rect 1859 2468 1952 2496
rect 1946 2456 1952 2468
rect 2004 2496 2010 2508
rect 4246 2496 4252 2508
rect 2004 2468 4252 2496
rect 2004 2456 2010 2468
rect 4246 2456 4252 2468
rect 4304 2456 4310 2508
rect 2590 2428 2596 2440
rect 2551 2400 2596 2428
rect 2590 2388 2596 2400
rect 2648 2388 2654 2440
rect 7282 2428 7288 2440
rect 7195 2400 7288 2428
rect 7282 2388 7288 2400
rect 7340 2428 7346 2440
rect 7742 2428 7748 2440
rect 7340 2400 7748 2428
rect 7340 2388 7346 2400
rect 7742 2388 7748 2400
rect 7800 2388 7806 2440
rect 1104 2202 7820 2224
rect 1104 2150 3150 2202
rect 3202 2150 3214 2202
rect 3266 2150 3278 2202
rect 3330 2150 3342 2202
rect 3394 2150 3406 2202
rect 3458 2150 7150 2202
rect 7202 2150 7214 2202
rect 7266 2150 7278 2202
rect 7330 2150 7342 2202
rect 7394 2150 7406 2202
rect 7458 2150 7820 2202
rect 1104 2128 7820 2150
rect 4249 2091 4307 2097
rect 4249 2057 4261 2091
rect 4295 2088 4307 2091
rect 4338 2088 4344 2100
rect 4295 2060 4344 2088
rect 4295 2057 4307 2060
rect 4249 2051 4307 2057
rect 4338 2048 4344 2060
rect 4396 2048 4402 2100
rect 3050 1980 3056 2032
rect 3108 1980 3114 2032
rect 5718 2020 5724 2032
rect 5644 1992 5724 2020
rect 3878 1912 3884 1964
rect 3936 1952 3942 1964
rect 5644 1961 5672 1992
rect 5718 1980 5724 1992
rect 5776 1980 5782 2032
rect 4065 1955 4123 1961
rect 4065 1952 4077 1955
rect 3936 1924 4077 1952
rect 3936 1912 3942 1924
rect 4065 1921 4077 1924
rect 4111 1921 4123 1955
rect 4065 1915 4123 1921
rect 5629 1955 5687 1961
rect 5629 1921 5641 1955
rect 5675 1921 5687 1955
rect 5810 1952 5816 1964
rect 5771 1924 5816 1952
rect 5629 1915 5687 1921
rect 5810 1912 5816 1924
rect 5868 1952 5874 1964
rect 6549 1955 6607 1961
rect 6549 1952 6561 1955
rect 5868 1924 6561 1952
rect 5868 1912 5874 1924
rect 6549 1921 6561 1924
rect 6595 1921 6607 1955
rect 6549 1915 6607 1921
rect 658 1844 664 1896
rect 716 1884 722 1896
rect 2225 1887 2283 1893
rect 2225 1884 2237 1887
rect 716 1856 2237 1884
rect 716 1844 722 1856
rect 2225 1853 2237 1856
rect 2271 1853 2283 1887
rect 2225 1847 2283 1853
rect 2593 1887 2651 1893
rect 2593 1853 2605 1887
rect 2639 1884 2651 1887
rect 2774 1884 2780 1896
rect 2639 1856 2780 1884
rect 2639 1853 2651 1856
rect 2593 1847 2651 1853
rect 2774 1844 2780 1856
rect 2832 1844 2838 1896
rect 5902 1884 5908 1896
rect 5863 1856 5908 1884
rect 5902 1844 5908 1856
rect 5960 1844 5966 1896
rect 1486 1708 1492 1760
rect 1544 1748 1550 1760
rect 1581 1751 1639 1757
rect 1581 1748 1593 1751
rect 1544 1720 1593 1748
rect 1544 1708 1550 1720
rect 1581 1717 1593 1720
rect 1627 1717 1639 1751
rect 1581 1711 1639 1717
rect 4525 1751 4583 1757
rect 4525 1717 4537 1751
rect 4571 1748 4583 1751
rect 6454 1748 6460 1760
rect 4571 1720 6460 1748
rect 4571 1717 4583 1720
rect 4525 1711 4583 1717
rect 6454 1708 6460 1720
rect 6512 1708 6518 1760
rect 1104 1658 7820 1680
rect 1104 1606 1150 1658
rect 1202 1606 1214 1658
rect 1266 1606 1278 1658
rect 1330 1606 1342 1658
rect 1394 1606 1406 1658
rect 1458 1606 5150 1658
rect 5202 1606 5214 1658
rect 5266 1606 5278 1658
rect 5330 1606 5342 1658
rect 5394 1606 5406 1658
rect 5458 1606 7820 1658
rect 1104 1584 7820 1606
rect 2774 1504 2780 1556
rect 2832 1544 2838 1556
rect 5261 1547 5319 1553
rect 5261 1544 5273 1547
rect 2832 1516 5273 1544
rect 2832 1504 2838 1516
rect 5261 1513 5273 1516
rect 5307 1544 5319 1547
rect 5994 1544 6000 1556
rect 5307 1516 6000 1544
rect 5307 1513 5319 1516
rect 5261 1507 5319 1513
rect 5994 1504 6000 1516
rect 6052 1504 6058 1556
rect 658 1368 664 1420
rect 716 1408 722 1420
rect 1581 1411 1639 1417
rect 1581 1408 1593 1411
rect 716 1380 1593 1408
rect 716 1368 722 1380
rect 1581 1377 1593 1380
rect 1627 1377 1639 1411
rect 1581 1371 1639 1377
rect 3050 1368 3056 1420
rect 3108 1408 3114 1420
rect 3237 1411 3295 1417
rect 3237 1408 3249 1411
rect 3108 1380 3249 1408
rect 3108 1368 3114 1380
rect 3237 1377 3249 1380
rect 3283 1377 3295 1411
rect 3237 1371 3295 1377
rect 3878 1368 3884 1420
rect 3936 1408 3942 1420
rect 3973 1411 4031 1417
rect 3973 1408 3985 1411
rect 3936 1380 3985 1408
rect 3936 1368 3942 1380
rect 3973 1377 3985 1380
rect 4019 1377 4031 1411
rect 3973 1371 4031 1377
rect 7006 1300 7012 1352
rect 7064 1340 7070 1352
rect 7101 1343 7159 1349
rect 7101 1340 7113 1343
rect 7064 1312 7113 1340
rect 7064 1300 7070 1312
rect 7101 1309 7113 1312
rect 7147 1309 7159 1343
rect 7101 1303 7159 1309
rect 7193 1207 7251 1213
rect 7193 1173 7205 1207
rect 7239 1204 7251 1207
rect 8386 1204 8392 1216
rect 7239 1176 8392 1204
rect 7239 1173 7251 1176
rect 7193 1167 7251 1173
rect 8386 1164 8392 1176
rect 8444 1164 8450 1216
rect 1104 1114 7820 1136
rect 1104 1062 3150 1114
rect 3202 1062 3214 1114
rect 3266 1062 3278 1114
rect 3330 1062 3342 1114
rect 3394 1062 3406 1114
rect 3458 1062 7150 1114
rect 7202 1062 7214 1114
rect 7266 1062 7278 1114
rect 7330 1062 7342 1114
rect 7394 1062 7406 1114
rect 7458 1062 7820 1114
rect 1104 1040 7820 1062
<< via1 >>
rect 2872 7896 2924 7948
rect 5724 7896 5776 7948
rect 3150 7590 3202 7642
rect 3214 7590 3266 7642
rect 3278 7590 3330 7642
rect 3342 7590 3394 7642
rect 3406 7590 3458 7642
rect 7150 7590 7202 7642
rect 7214 7590 7266 7642
rect 7278 7590 7330 7642
rect 7342 7590 7394 7642
rect 7406 7590 7458 7642
rect 2136 7395 2188 7404
rect 2136 7361 2145 7395
rect 2145 7361 2179 7395
rect 2179 7361 2188 7395
rect 2136 7352 2188 7361
rect 6828 7352 6880 7404
rect 7564 7352 7616 7404
rect 1150 7046 1202 7098
rect 1214 7046 1266 7098
rect 1278 7046 1330 7098
rect 1342 7046 1394 7098
rect 1406 7046 1458 7098
rect 5150 7046 5202 7098
rect 5214 7046 5266 7098
rect 5278 7046 5330 7098
rect 5342 7046 5394 7098
rect 5406 7046 5458 7098
rect 20 6944 72 6996
rect 1584 6851 1636 6860
rect 1584 6817 1593 6851
rect 1593 6817 1627 6851
rect 1627 6817 1636 6851
rect 1584 6808 1636 6817
rect 4252 6808 4304 6860
rect 6736 6808 6788 6860
rect 2136 6783 2188 6792
rect 2136 6749 2145 6783
rect 2145 6749 2179 6783
rect 2179 6749 2188 6783
rect 2136 6740 2188 6749
rect 2780 6740 2832 6792
rect 3056 6740 3108 6792
rect 8392 6740 8444 6792
rect 3150 6502 3202 6554
rect 3214 6502 3266 6554
rect 3278 6502 3330 6554
rect 3342 6502 3394 6554
rect 3406 6502 3458 6554
rect 7150 6502 7202 6554
rect 7214 6502 7266 6554
rect 7278 6502 7330 6554
rect 7342 6502 7394 6554
rect 7406 6502 7458 6554
rect 1584 6239 1636 6248
rect 1584 6205 1593 6239
rect 1593 6205 1627 6239
rect 1627 6205 1636 6239
rect 1584 6196 1636 6205
rect 3056 6264 3108 6316
rect 6736 6264 6788 6316
rect 4804 6196 4856 6248
rect 1584 6060 1636 6112
rect 7564 6060 7616 6112
rect 1150 5958 1202 6010
rect 1214 5958 1266 6010
rect 1278 5958 1330 6010
rect 1342 5958 1394 6010
rect 1406 5958 1458 6010
rect 5150 5958 5202 6010
rect 5214 5958 5266 6010
rect 5278 5958 5330 6010
rect 5342 5958 5394 6010
rect 5406 5958 5458 6010
rect 7012 5856 7064 5908
rect 6828 5763 6880 5772
rect 6828 5729 6837 5763
rect 6837 5729 6871 5763
rect 6871 5729 6880 5763
rect 6828 5720 6880 5729
rect 1584 5695 1636 5704
rect 1584 5661 1593 5695
rect 1593 5661 1627 5695
rect 1627 5661 1636 5695
rect 1584 5652 1636 5661
rect 6828 5584 6880 5636
rect 6552 5516 6604 5568
rect 3150 5414 3202 5466
rect 3214 5414 3266 5466
rect 3278 5414 3330 5466
rect 3342 5414 3394 5466
rect 3406 5414 3458 5466
rect 7150 5414 7202 5466
rect 7214 5414 7266 5466
rect 7278 5414 7330 5466
rect 7342 5414 7394 5466
rect 7406 5414 7458 5466
rect 6552 5015 6604 5024
rect 6552 4981 6561 5015
rect 6561 4981 6595 5015
rect 6595 4981 6604 5015
rect 6552 4972 6604 4981
rect 1150 4870 1202 4922
rect 1214 4870 1266 4922
rect 1278 4870 1330 4922
rect 1342 4870 1394 4922
rect 1406 4870 1458 4922
rect 5150 4870 5202 4922
rect 5214 4870 5266 4922
rect 5278 4870 5330 4922
rect 5342 4870 5394 4922
rect 5406 4870 5458 4922
rect 1952 4811 2004 4820
rect 1952 4777 1961 4811
rect 1961 4777 1995 4811
rect 1995 4777 2004 4811
rect 1952 4768 2004 4777
rect 6828 4768 6880 4820
rect 1492 4700 1544 4752
rect 7012 4700 7064 4752
rect 7748 4700 7800 4752
rect 3150 4326 3202 4378
rect 3214 4326 3266 4378
rect 3278 4326 3330 4378
rect 3342 4326 3394 4378
rect 3406 4326 3458 4378
rect 7150 4326 7202 4378
rect 7214 4326 7266 4378
rect 7278 4326 7330 4378
rect 7342 4326 7394 4378
rect 7406 4326 7458 4378
rect 1584 4156 1636 4208
rect 1952 4199 2004 4208
rect 1952 4165 1961 4199
rect 1961 4165 1995 4199
rect 1995 4165 2004 4199
rect 1952 4156 2004 4165
rect 4068 4156 4120 4208
rect 6460 4156 6512 4208
rect 1492 4088 1544 4140
rect 7012 4131 7064 4140
rect 7012 4097 7021 4131
rect 7021 4097 7055 4131
rect 7055 4097 7064 4131
rect 7012 4088 7064 4097
rect 7288 4131 7340 4140
rect 7288 4097 7297 4131
rect 7297 4097 7331 4131
rect 7331 4097 7340 4131
rect 7288 4088 7340 4097
rect 1032 4020 1084 4072
rect 4988 3952 5040 4004
rect 2780 3927 2832 3936
rect 2780 3893 2789 3927
rect 2789 3893 2823 3927
rect 2823 3893 2832 3927
rect 2780 3884 2832 3893
rect 1150 3782 1202 3834
rect 1214 3782 1266 3834
rect 1278 3782 1330 3834
rect 1342 3782 1394 3834
rect 1406 3782 1458 3834
rect 5150 3782 5202 3834
rect 5214 3782 5266 3834
rect 5278 3782 5330 3834
rect 5342 3782 5394 3834
rect 5406 3782 5458 3834
rect 6460 3723 6512 3732
rect 6460 3689 6469 3723
rect 6469 3689 6503 3723
rect 6503 3689 6512 3723
rect 6460 3680 6512 3689
rect 7012 3680 7064 3732
rect 7288 3723 7340 3732
rect 7288 3689 7297 3723
rect 7297 3689 7331 3723
rect 7331 3689 7340 3723
rect 7288 3680 7340 3689
rect 20 3612 72 3664
rect 6552 3612 6604 3664
rect 1584 3519 1636 3528
rect 1584 3485 1593 3519
rect 1593 3485 1627 3519
rect 1627 3485 1636 3519
rect 1584 3476 1636 3485
rect 3150 3238 3202 3290
rect 3214 3238 3266 3290
rect 3278 3238 3330 3290
rect 3342 3238 3394 3290
rect 3406 3238 3458 3290
rect 7150 3238 7202 3290
rect 7214 3238 7266 3290
rect 7278 3238 7330 3290
rect 7342 3238 7394 3290
rect 7406 3238 7458 3290
rect 4528 3136 4580 3188
rect 2596 3068 2648 3120
rect 1492 3000 1544 3052
rect 5080 3000 5132 3052
rect 7288 3043 7340 3052
rect 7288 3009 7297 3043
rect 7297 3009 7331 3043
rect 7331 3009 7340 3043
rect 7288 3000 7340 3009
rect 1952 2975 2004 2984
rect 1952 2941 1961 2975
rect 1961 2941 1995 2975
rect 1995 2941 2004 2975
rect 1952 2932 2004 2941
rect 4160 2796 4212 2848
rect 7840 2796 7892 2848
rect 1150 2694 1202 2746
rect 1214 2694 1266 2746
rect 1278 2694 1330 2746
rect 1342 2694 1394 2746
rect 1406 2694 1458 2746
rect 5150 2694 5202 2746
rect 5214 2694 5266 2746
rect 5278 2694 5330 2746
rect 5342 2694 5394 2746
rect 5406 2694 5458 2746
rect 5080 2592 5132 2644
rect 5724 2592 5776 2644
rect 1952 2499 2004 2508
rect 1952 2465 1961 2499
rect 1961 2465 1995 2499
rect 1995 2465 2004 2499
rect 1952 2456 2004 2465
rect 4252 2456 4304 2508
rect 2596 2431 2648 2440
rect 2596 2397 2605 2431
rect 2605 2397 2639 2431
rect 2639 2397 2648 2431
rect 2596 2388 2648 2397
rect 7288 2431 7340 2440
rect 7288 2397 7297 2431
rect 7297 2397 7331 2431
rect 7331 2397 7340 2431
rect 7288 2388 7340 2397
rect 7748 2388 7800 2440
rect 3150 2150 3202 2202
rect 3214 2150 3266 2202
rect 3278 2150 3330 2202
rect 3342 2150 3394 2202
rect 3406 2150 3458 2202
rect 7150 2150 7202 2202
rect 7214 2150 7266 2202
rect 7278 2150 7330 2202
rect 7342 2150 7394 2202
rect 7406 2150 7458 2202
rect 4344 2048 4396 2100
rect 3056 1980 3108 2032
rect 3884 1912 3936 1964
rect 5724 1980 5776 2032
rect 5816 1955 5868 1964
rect 5816 1921 5825 1955
rect 5825 1921 5859 1955
rect 5859 1921 5868 1955
rect 5816 1912 5868 1921
rect 664 1844 716 1896
rect 2780 1844 2832 1896
rect 5908 1887 5960 1896
rect 5908 1853 5917 1887
rect 5917 1853 5951 1887
rect 5951 1853 5960 1887
rect 5908 1844 5960 1853
rect 1492 1708 1544 1760
rect 6460 1708 6512 1760
rect 1150 1606 1202 1658
rect 1214 1606 1266 1658
rect 1278 1606 1330 1658
rect 1342 1606 1394 1658
rect 1406 1606 1458 1658
rect 5150 1606 5202 1658
rect 5214 1606 5266 1658
rect 5278 1606 5330 1658
rect 5342 1606 5394 1658
rect 5406 1606 5458 1658
rect 2780 1504 2832 1556
rect 6000 1504 6052 1556
rect 664 1368 716 1420
rect 3056 1368 3108 1420
rect 3884 1368 3936 1420
rect 7012 1300 7064 1352
rect 8392 1164 8444 1216
rect 3150 1062 3202 1114
rect 3214 1062 3266 1114
rect 3278 1062 3330 1114
rect 3342 1062 3394 1114
rect 3406 1062 3458 1114
rect 7150 1062 7202 1114
rect 7214 1062 7266 1114
rect 7278 1062 7330 1114
rect 7342 1062 7394 1114
rect 7406 1062 7458 1114
<< metal2 >>
rect 18 8200 74 9000
rect 662 8200 718 9000
rect 768 8214 1532 8242
rect 32 7002 60 8200
rect 676 8106 704 8200
rect 768 8106 796 8214
rect 676 8078 796 8106
rect 1150 7100 1458 7109
rect 1150 7098 1156 7100
rect 1212 7098 1236 7100
rect 1292 7098 1316 7100
rect 1372 7098 1396 7100
rect 1452 7098 1458 7100
rect 1212 7046 1214 7098
rect 1394 7046 1396 7098
rect 1150 7044 1156 7046
rect 1212 7044 1236 7046
rect 1292 7044 1316 7046
rect 1372 7044 1396 7046
rect 1452 7044 1458 7046
rect 1150 7035 1458 7044
rect 20 6996 72 7002
rect 20 6938 72 6944
rect 1150 6012 1458 6021
rect 1150 6010 1156 6012
rect 1212 6010 1236 6012
rect 1292 6010 1316 6012
rect 1372 6010 1396 6012
rect 1452 6010 1458 6012
rect 1212 5958 1214 6010
rect 1394 5958 1396 6010
rect 1150 5956 1156 5958
rect 1212 5956 1236 5958
rect 1292 5956 1316 5958
rect 1372 5956 1396 5958
rect 1452 5956 1458 5958
rect 1150 5947 1458 5956
rect 1150 4924 1458 4933
rect 1150 4922 1156 4924
rect 1212 4922 1236 4924
rect 1292 4922 1316 4924
rect 1372 4922 1396 4924
rect 1452 4922 1458 4924
rect 1212 4870 1214 4922
rect 1394 4870 1396 4922
rect 1150 4868 1156 4870
rect 1212 4868 1236 4870
rect 1292 4868 1316 4870
rect 1372 4868 1396 4870
rect 1452 4868 1458 4870
rect 1150 4859 1458 4868
rect 1504 4758 1532 8214
rect 1950 8200 2006 9000
rect 2148 8214 2544 8242
rect 1582 7576 1638 7585
rect 1582 7511 1638 7520
rect 1596 6866 1624 7511
rect 1584 6860 1636 6866
rect 1584 6802 1636 6808
rect 1584 6248 1636 6254
rect 1582 6216 1584 6225
rect 1636 6216 1638 6225
rect 1582 6151 1638 6160
rect 1584 6112 1636 6118
rect 1584 6054 1636 6060
rect 1596 5710 1624 6054
rect 1584 5704 1636 5710
rect 1584 5646 1636 5652
rect 1596 5137 1624 5646
rect 1582 5128 1638 5137
rect 1582 5063 1638 5072
rect 1964 4826 1992 8200
rect 2148 7410 2176 8214
rect 2516 8106 2544 8214
rect 2594 8200 2650 9000
rect 2870 8936 2926 8945
rect 2870 8871 2926 8880
rect 2608 8106 2636 8200
rect 2516 8078 2636 8106
rect 2884 7954 2912 8871
rect 3238 8200 3294 9000
rect 4526 8200 4582 9000
rect 4816 8214 5120 8242
rect 2872 7948 2924 7954
rect 2872 7890 2924 7896
rect 3252 7834 3280 8200
rect 3068 7806 3280 7834
rect 2136 7404 2188 7410
rect 2136 7346 2188 7352
rect 2148 6798 2176 7346
rect 3068 6798 3096 7806
rect 3150 7644 3458 7653
rect 3150 7642 3156 7644
rect 3212 7642 3236 7644
rect 3292 7642 3316 7644
rect 3372 7642 3396 7644
rect 3452 7642 3458 7644
rect 3212 7590 3214 7642
rect 3394 7590 3396 7642
rect 3150 7588 3156 7590
rect 3212 7588 3236 7590
rect 3292 7588 3316 7590
rect 3372 7588 3396 7590
rect 3452 7588 3458 7590
rect 3150 7579 3458 7588
rect 4250 6896 4306 6905
rect 4250 6831 4252 6840
rect 4304 6831 4306 6840
rect 4252 6802 4304 6808
rect 2136 6792 2188 6798
rect 2136 6734 2188 6740
rect 2780 6792 2832 6798
rect 2780 6734 2832 6740
rect 3056 6792 3108 6798
rect 3056 6734 3108 6740
rect 4342 6760 4398 6769
rect 1952 4820 2004 4826
rect 1952 4762 2004 4768
rect 1492 4752 1544 4758
rect 1492 4694 1544 4700
rect 1504 4146 1532 4694
rect 1964 4214 1992 4762
rect 1584 4208 1636 4214
rect 1584 4150 1636 4156
rect 1952 4208 2004 4214
rect 1952 4150 2004 4156
rect 1492 4140 1544 4146
rect 1492 4082 1544 4088
rect 1032 4072 1084 4078
rect 1032 4014 1084 4020
rect 20 3664 72 3670
rect 20 3606 72 3612
rect 32 800 60 3606
rect 664 1896 716 1902
rect 664 1838 716 1844
rect 676 1426 704 1838
rect 664 1420 716 1426
rect 664 1362 716 1368
rect 676 800 704 1362
rect 18 0 74 800
rect 662 0 718 800
rect 1044 762 1072 4014
rect 1150 3836 1458 3845
rect 1150 3834 1156 3836
rect 1212 3834 1236 3836
rect 1292 3834 1316 3836
rect 1372 3834 1396 3836
rect 1452 3834 1458 3836
rect 1212 3782 1214 3834
rect 1394 3782 1396 3834
rect 1150 3780 1156 3782
rect 1212 3780 1236 3782
rect 1292 3780 1316 3782
rect 1372 3780 1396 3782
rect 1452 3780 1458 3782
rect 1150 3771 1458 3780
rect 1596 3534 1624 4150
rect 2792 3942 2820 6734
rect 3068 6322 3096 6734
rect 4342 6695 4398 6704
rect 3150 6556 3458 6565
rect 3150 6554 3156 6556
rect 3212 6554 3236 6556
rect 3292 6554 3316 6556
rect 3372 6554 3396 6556
rect 3452 6554 3458 6556
rect 3212 6502 3214 6554
rect 3394 6502 3396 6554
rect 3150 6500 3156 6502
rect 3212 6500 3236 6502
rect 3292 6500 3316 6502
rect 3372 6500 3396 6502
rect 3452 6500 3458 6502
rect 3150 6491 3458 6500
rect 3056 6316 3108 6322
rect 3056 6258 3108 6264
rect 3150 5468 3458 5477
rect 3150 5466 3156 5468
rect 3212 5466 3236 5468
rect 3292 5466 3316 5468
rect 3372 5466 3396 5468
rect 3452 5466 3458 5468
rect 3212 5414 3214 5466
rect 3394 5414 3396 5466
rect 3150 5412 3156 5414
rect 3212 5412 3236 5414
rect 3292 5412 3316 5414
rect 3372 5412 3396 5414
rect 3452 5412 3458 5414
rect 3150 5403 3458 5412
rect 3150 4380 3458 4389
rect 3150 4378 3156 4380
rect 3212 4378 3236 4380
rect 3292 4378 3316 4380
rect 3372 4378 3396 4380
rect 3452 4378 3458 4380
rect 3212 4326 3214 4378
rect 3394 4326 3396 4378
rect 3150 4324 3156 4326
rect 3212 4324 3236 4326
rect 3292 4324 3316 4326
rect 3372 4324 3396 4326
rect 3452 4324 3458 4326
rect 3150 4315 3458 4324
rect 4068 4208 4120 4214
rect 4066 4176 4068 4185
rect 4120 4176 4122 4185
rect 4066 4111 4122 4120
rect 2780 3936 2832 3942
rect 2780 3878 2832 3884
rect 1584 3528 1636 3534
rect 2792 3505 2820 3878
rect 1584 3470 1636 3476
rect 2778 3496 2834 3505
rect 1492 3052 1544 3058
rect 1492 2994 1544 3000
rect 1150 2748 1458 2757
rect 1150 2746 1156 2748
rect 1212 2746 1236 2748
rect 1292 2746 1316 2748
rect 1372 2746 1396 2748
rect 1452 2746 1458 2748
rect 1212 2694 1214 2746
rect 1394 2694 1396 2746
rect 1150 2692 1156 2694
rect 1212 2692 1236 2694
rect 1292 2692 1316 2694
rect 1372 2692 1396 2694
rect 1452 2692 1458 2694
rect 1150 2683 1458 2692
rect 1504 1766 1532 2994
rect 1492 1760 1544 1766
rect 1492 1702 1544 1708
rect 1150 1660 1458 1669
rect 1150 1658 1156 1660
rect 1212 1658 1236 1660
rect 1292 1658 1316 1660
rect 1372 1658 1396 1660
rect 1452 1658 1458 1660
rect 1212 1606 1214 1658
rect 1394 1606 1396 1658
rect 1150 1604 1156 1606
rect 1212 1604 1236 1606
rect 1292 1604 1316 1606
rect 1372 1604 1396 1606
rect 1452 1604 1458 1606
rect 1150 1595 1458 1604
rect 1228 870 1348 898
rect 1228 762 1256 870
rect 1320 800 1348 870
rect 1044 734 1256 762
rect 1306 0 1362 800
rect 1504 785 1532 1702
rect 1596 1465 1624 3470
rect 2778 3431 2834 3440
rect 3150 3292 3458 3301
rect 3150 3290 3156 3292
rect 3212 3290 3236 3292
rect 3292 3290 3316 3292
rect 3372 3290 3396 3292
rect 3452 3290 3458 3292
rect 3212 3238 3214 3290
rect 3394 3238 3396 3290
rect 3150 3236 3156 3238
rect 3212 3236 3236 3238
rect 3292 3236 3316 3238
rect 3372 3236 3396 3238
rect 3452 3236 3458 3238
rect 3150 3227 3458 3236
rect 2596 3120 2648 3126
rect 2596 3062 2648 3068
rect 1952 2984 2004 2990
rect 1952 2926 2004 2932
rect 1964 2514 1992 2926
rect 1952 2508 2004 2514
rect 1952 2450 2004 2456
rect 2608 2446 2636 3062
rect 4160 2848 4212 2854
rect 4160 2790 4212 2796
rect 2596 2440 2648 2446
rect 2596 2382 2648 2388
rect 1582 1456 1638 1465
rect 1582 1391 1638 1400
rect 2608 800 2636 2382
rect 3150 2204 3458 2213
rect 3150 2202 3156 2204
rect 3212 2202 3236 2204
rect 3292 2202 3316 2204
rect 3372 2202 3396 2204
rect 3452 2202 3458 2204
rect 3212 2150 3214 2202
rect 3394 2150 3396 2202
rect 3150 2148 3156 2150
rect 3212 2148 3236 2150
rect 3292 2148 3316 2150
rect 3372 2148 3396 2150
rect 3452 2148 3458 2150
rect 3150 2139 3458 2148
rect 3056 2032 3108 2038
rect 3056 1974 3108 1980
rect 4066 2000 4122 2009
rect 2780 1896 2832 1902
rect 2780 1838 2832 1844
rect 2792 1562 2820 1838
rect 2780 1556 2832 1562
rect 2780 1498 2832 1504
rect 3068 1426 3096 1974
rect 3884 1964 3936 1970
rect 4172 1986 4200 2790
rect 4252 2508 4304 2514
rect 4252 2450 4304 2456
rect 4264 2417 4292 2450
rect 4250 2408 4306 2417
rect 4250 2343 4306 2352
rect 4356 2106 4384 6695
rect 4540 3194 4568 8200
rect 4816 6254 4844 8214
rect 5092 8106 5120 8214
rect 5170 8200 5226 9000
rect 5814 8200 5870 9000
rect 6734 8256 6790 8265
rect 7102 8200 7158 9000
rect 7746 8200 7802 9000
rect 8390 8200 8446 9000
rect 5184 8106 5212 8200
rect 5092 8078 5212 8106
rect 5724 7948 5776 7954
rect 5724 7890 5776 7896
rect 5150 7100 5458 7109
rect 5150 7098 5156 7100
rect 5212 7098 5236 7100
rect 5292 7098 5316 7100
rect 5372 7098 5396 7100
rect 5452 7098 5458 7100
rect 5212 7046 5214 7098
rect 5394 7046 5396 7098
rect 5150 7044 5156 7046
rect 5212 7044 5236 7046
rect 5292 7044 5316 7046
rect 5372 7044 5396 7046
rect 5452 7044 5458 7046
rect 5150 7035 5458 7044
rect 4804 6248 4856 6254
rect 4804 6190 4856 6196
rect 5150 6012 5458 6021
rect 5150 6010 5156 6012
rect 5212 6010 5236 6012
rect 5292 6010 5316 6012
rect 5372 6010 5396 6012
rect 5452 6010 5458 6012
rect 5212 5958 5214 6010
rect 5394 5958 5396 6010
rect 5150 5956 5156 5958
rect 5212 5956 5236 5958
rect 5292 5956 5316 5958
rect 5372 5956 5396 5958
rect 5452 5956 5458 5958
rect 5150 5947 5458 5956
rect 5150 4924 5458 4933
rect 5150 4922 5156 4924
rect 5212 4922 5236 4924
rect 5292 4922 5316 4924
rect 5372 4922 5396 4924
rect 5452 4922 5458 4924
rect 5212 4870 5214 4922
rect 5394 4870 5396 4922
rect 5150 4868 5156 4870
rect 5212 4868 5236 4870
rect 5292 4868 5316 4870
rect 5372 4868 5396 4870
rect 5452 4868 5458 4870
rect 5150 4859 5458 4868
rect 4988 4004 5040 4010
rect 4988 3946 5040 3952
rect 4528 3188 4580 3194
rect 4528 3130 4580 3136
rect 4344 2100 4396 2106
rect 4344 2042 4396 2048
rect 4122 1958 4200 1986
rect 4066 1935 4122 1944
rect 3884 1906 3936 1912
rect 3896 1426 3924 1906
rect 5000 1442 5028 3946
rect 5150 3836 5458 3845
rect 5150 3834 5156 3836
rect 5212 3834 5236 3836
rect 5292 3834 5316 3836
rect 5372 3834 5396 3836
rect 5452 3834 5458 3836
rect 5212 3782 5214 3834
rect 5394 3782 5396 3834
rect 5150 3780 5156 3782
rect 5212 3780 5236 3782
rect 5292 3780 5316 3782
rect 5372 3780 5396 3782
rect 5452 3780 5458 3782
rect 5150 3771 5458 3780
rect 5080 3052 5132 3058
rect 5080 2994 5132 3000
rect 5092 2961 5120 2994
rect 5078 2952 5134 2961
rect 5078 2887 5134 2896
rect 5092 2650 5120 2887
rect 5150 2748 5458 2757
rect 5150 2746 5156 2748
rect 5212 2746 5236 2748
rect 5292 2746 5316 2748
rect 5372 2746 5396 2748
rect 5452 2746 5458 2748
rect 5212 2694 5214 2746
rect 5394 2694 5396 2746
rect 5150 2692 5156 2694
rect 5212 2692 5236 2694
rect 5292 2692 5316 2694
rect 5372 2692 5396 2694
rect 5452 2692 5458 2694
rect 5150 2683 5458 2692
rect 5736 2650 5764 7890
rect 5828 6914 5856 8200
rect 6734 8191 6790 8200
rect 5828 6886 6040 6914
rect 5080 2644 5132 2650
rect 5080 2586 5132 2592
rect 5724 2644 5776 2650
rect 5724 2586 5776 2592
rect 5736 2038 5764 2586
rect 5724 2032 5776 2038
rect 5724 1974 5776 1980
rect 5816 1964 5868 1970
rect 5816 1906 5868 1912
rect 5150 1660 5458 1669
rect 5150 1658 5156 1660
rect 5212 1658 5236 1660
rect 5292 1658 5316 1660
rect 5372 1658 5396 1660
rect 5452 1658 5458 1660
rect 5212 1606 5214 1658
rect 5394 1606 5396 1658
rect 5150 1604 5156 1606
rect 5212 1604 5236 1606
rect 5292 1604 5316 1606
rect 5372 1604 5396 1606
rect 5452 1604 5458 1606
rect 5150 1595 5458 1604
rect 3056 1420 3108 1426
rect 3056 1362 3108 1368
rect 3884 1420 3936 1426
rect 5000 1414 5212 1442
rect 3884 1362 3936 1368
rect 3068 898 3096 1362
rect 3150 1116 3458 1125
rect 3150 1114 3156 1116
rect 3212 1114 3236 1116
rect 3292 1114 3316 1116
rect 3372 1114 3396 1116
rect 3452 1114 3458 1116
rect 3212 1062 3214 1114
rect 3394 1062 3396 1114
rect 3150 1060 3156 1062
rect 3212 1060 3236 1062
rect 3292 1060 3316 1062
rect 3372 1060 3396 1062
rect 3452 1060 3458 1062
rect 3150 1051 3458 1060
rect 3068 870 3280 898
rect 3252 800 3280 870
rect 3896 800 3924 1362
rect 5184 800 5212 1414
rect 5828 800 5856 1906
rect 5908 1896 5960 1902
rect 5908 1838 5960 1844
rect 5920 1465 5948 1838
rect 6012 1562 6040 6886
rect 6748 6866 6776 8191
rect 7116 7834 7144 8200
rect 7024 7806 7144 7834
rect 6828 7404 6880 7410
rect 6828 7346 6880 7352
rect 6736 6860 6788 6866
rect 6736 6802 6788 6808
rect 6748 6322 6776 6802
rect 6736 6316 6788 6322
rect 6736 6258 6788 6264
rect 6840 5778 6868 7346
rect 7024 5914 7052 7806
rect 7150 7644 7458 7653
rect 7150 7642 7156 7644
rect 7212 7642 7236 7644
rect 7292 7642 7316 7644
rect 7372 7642 7396 7644
rect 7452 7642 7458 7644
rect 7212 7590 7214 7642
rect 7394 7590 7396 7642
rect 7150 7588 7156 7590
rect 7212 7588 7236 7590
rect 7292 7588 7316 7590
rect 7372 7588 7396 7590
rect 7452 7588 7458 7590
rect 7150 7579 7458 7588
rect 7562 7576 7618 7585
rect 7562 7511 7618 7520
rect 7576 7410 7604 7511
rect 7564 7404 7616 7410
rect 7564 7346 7616 7352
rect 7150 6556 7458 6565
rect 7150 6554 7156 6556
rect 7212 6554 7236 6556
rect 7292 6554 7316 6556
rect 7372 6554 7396 6556
rect 7452 6554 7458 6556
rect 7212 6502 7214 6554
rect 7394 6502 7396 6554
rect 7150 6500 7156 6502
rect 7212 6500 7236 6502
rect 7292 6500 7316 6502
rect 7372 6500 7396 6502
rect 7452 6500 7458 6502
rect 7150 6491 7458 6500
rect 7564 6112 7616 6118
rect 7564 6054 7616 6060
rect 7012 5908 7064 5914
rect 7012 5850 7064 5856
rect 6828 5772 6880 5778
rect 6828 5714 6880 5720
rect 6828 5636 6880 5642
rect 6828 5578 6880 5584
rect 6552 5568 6604 5574
rect 6552 5510 6604 5516
rect 6564 5030 6592 5510
rect 6552 5024 6604 5030
rect 6552 4966 6604 4972
rect 6460 4208 6512 4214
rect 6460 4150 6512 4156
rect 6472 3738 6500 4150
rect 6460 3732 6512 3738
rect 6460 3674 6512 3680
rect 6564 3670 6592 4966
rect 6840 4865 6868 5578
rect 7576 5545 7604 6054
rect 7562 5536 7618 5545
rect 7150 5468 7458 5477
rect 7562 5471 7618 5480
rect 7150 5466 7156 5468
rect 7212 5466 7236 5468
rect 7292 5466 7316 5468
rect 7372 5466 7396 5468
rect 7452 5466 7458 5468
rect 7212 5414 7214 5466
rect 7394 5414 7396 5466
rect 7150 5412 7156 5414
rect 7212 5412 7236 5414
rect 7292 5412 7316 5414
rect 7372 5412 7396 5414
rect 7452 5412 7458 5414
rect 7150 5403 7458 5412
rect 6826 4856 6882 4865
rect 6826 4791 6828 4800
rect 6880 4791 6882 4800
rect 6828 4762 6880 4768
rect 6840 4731 6868 4762
rect 7760 4758 7788 8200
rect 8404 6798 8432 8200
rect 8392 6792 8444 6798
rect 8392 6734 8444 6740
rect 7012 4752 7064 4758
rect 7012 4694 7064 4700
rect 7748 4752 7800 4758
rect 7748 4694 7800 4700
rect 7024 4146 7052 4694
rect 7150 4380 7458 4389
rect 7150 4378 7156 4380
rect 7212 4378 7236 4380
rect 7292 4378 7316 4380
rect 7372 4378 7396 4380
rect 7452 4378 7458 4380
rect 7212 4326 7214 4378
rect 7394 4326 7396 4378
rect 7150 4324 7156 4326
rect 7212 4324 7236 4326
rect 7292 4324 7316 4326
rect 7372 4324 7396 4326
rect 7452 4324 7458 4326
rect 7150 4315 7458 4324
rect 7286 4176 7342 4185
rect 7012 4140 7064 4146
rect 7286 4111 7288 4120
rect 7012 4082 7064 4088
rect 7340 4111 7342 4120
rect 7288 4082 7340 4088
rect 7300 3738 7328 4082
rect 7012 3732 7064 3738
rect 7012 3674 7064 3680
rect 7288 3732 7340 3738
rect 7288 3674 7340 3680
rect 6552 3664 6604 3670
rect 6552 3606 6604 3612
rect 6460 1760 6512 1766
rect 6460 1702 6512 1708
rect 6000 1556 6052 1562
rect 6000 1498 6052 1504
rect 5906 1456 5962 1465
rect 5906 1391 5962 1400
rect 6472 800 6500 1702
rect 7024 1358 7052 3674
rect 7150 3292 7458 3301
rect 7150 3290 7156 3292
rect 7212 3290 7236 3292
rect 7292 3290 7316 3292
rect 7372 3290 7396 3292
rect 7452 3290 7458 3292
rect 7212 3238 7214 3290
rect 7394 3238 7396 3290
rect 7150 3236 7156 3238
rect 7212 3236 7236 3238
rect 7292 3236 7316 3238
rect 7372 3236 7396 3238
rect 7452 3236 7458 3238
rect 7150 3227 7458 3236
rect 7288 3052 7340 3058
rect 7288 2994 7340 3000
rect 7300 2446 7328 2994
rect 7840 2848 7892 2854
rect 7840 2790 7892 2796
rect 7288 2440 7340 2446
rect 7288 2382 7340 2388
rect 7748 2440 7800 2446
rect 7748 2382 7800 2388
rect 7150 2204 7458 2213
rect 7150 2202 7156 2204
rect 7212 2202 7236 2204
rect 7292 2202 7316 2204
rect 7372 2202 7396 2204
rect 7452 2202 7458 2204
rect 7212 2150 7214 2202
rect 7394 2150 7396 2202
rect 7150 2148 7156 2150
rect 7212 2148 7236 2150
rect 7292 2148 7316 2150
rect 7372 2148 7396 2150
rect 7452 2148 7458 2150
rect 7150 2139 7458 2148
rect 7012 1352 7064 1358
rect 7012 1294 7064 1300
rect 7150 1116 7458 1125
rect 7150 1114 7156 1116
rect 7212 1114 7236 1116
rect 7292 1114 7316 1116
rect 7372 1114 7396 1116
rect 7452 1114 7458 1116
rect 7212 1062 7214 1114
rect 7394 1062 7396 1114
rect 7150 1060 7156 1062
rect 7212 1060 7236 1062
rect 7292 1060 7316 1062
rect 7372 1060 7396 1062
rect 7452 1060 7458 1062
rect 7150 1051 7458 1060
rect 7760 800 7788 2382
rect 1490 776 1546 785
rect 1490 711 1546 720
rect 2594 0 2650 800
rect 3238 0 3294 800
rect 3882 0 3938 800
rect 5170 0 5226 800
rect 5814 0 5870 800
rect 6458 0 6514 800
rect 7746 0 7802 800
rect 7852 105 7880 2790
rect 8392 1216 8444 1222
rect 8392 1158 8444 1164
rect 8404 800 8432 1158
rect 7838 96 7894 105
rect 7838 31 7894 40
rect 8390 0 8446 800
<< via2 >>
rect 1156 7098 1212 7100
rect 1236 7098 1292 7100
rect 1316 7098 1372 7100
rect 1396 7098 1452 7100
rect 1156 7046 1202 7098
rect 1202 7046 1212 7098
rect 1236 7046 1266 7098
rect 1266 7046 1278 7098
rect 1278 7046 1292 7098
rect 1316 7046 1330 7098
rect 1330 7046 1342 7098
rect 1342 7046 1372 7098
rect 1396 7046 1406 7098
rect 1406 7046 1452 7098
rect 1156 7044 1212 7046
rect 1236 7044 1292 7046
rect 1316 7044 1372 7046
rect 1396 7044 1452 7046
rect 1156 6010 1212 6012
rect 1236 6010 1292 6012
rect 1316 6010 1372 6012
rect 1396 6010 1452 6012
rect 1156 5958 1202 6010
rect 1202 5958 1212 6010
rect 1236 5958 1266 6010
rect 1266 5958 1278 6010
rect 1278 5958 1292 6010
rect 1316 5958 1330 6010
rect 1330 5958 1342 6010
rect 1342 5958 1372 6010
rect 1396 5958 1406 6010
rect 1406 5958 1452 6010
rect 1156 5956 1212 5958
rect 1236 5956 1292 5958
rect 1316 5956 1372 5958
rect 1396 5956 1452 5958
rect 1156 4922 1212 4924
rect 1236 4922 1292 4924
rect 1316 4922 1372 4924
rect 1396 4922 1452 4924
rect 1156 4870 1202 4922
rect 1202 4870 1212 4922
rect 1236 4870 1266 4922
rect 1266 4870 1278 4922
rect 1278 4870 1292 4922
rect 1316 4870 1330 4922
rect 1330 4870 1342 4922
rect 1342 4870 1372 4922
rect 1396 4870 1406 4922
rect 1406 4870 1452 4922
rect 1156 4868 1212 4870
rect 1236 4868 1292 4870
rect 1316 4868 1372 4870
rect 1396 4868 1452 4870
rect 1582 7520 1638 7576
rect 1582 6196 1584 6216
rect 1584 6196 1636 6216
rect 1636 6196 1638 6216
rect 1582 6160 1638 6196
rect 1582 5072 1638 5128
rect 2870 8880 2926 8936
rect 3156 7642 3212 7644
rect 3236 7642 3292 7644
rect 3316 7642 3372 7644
rect 3396 7642 3452 7644
rect 3156 7590 3202 7642
rect 3202 7590 3212 7642
rect 3236 7590 3266 7642
rect 3266 7590 3278 7642
rect 3278 7590 3292 7642
rect 3316 7590 3330 7642
rect 3330 7590 3342 7642
rect 3342 7590 3372 7642
rect 3396 7590 3406 7642
rect 3406 7590 3452 7642
rect 3156 7588 3212 7590
rect 3236 7588 3292 7590
rect 3316 7588 3372 7590
rect 3396 7588 3452 7590
rect 4250 6860 4306 6896
rect 4250 6840 4252 6860
rect 4252 6840 4304 6860
rect 4304 6840 4306 6860
rect 1156 3834 1212 3836
rect 1236 3834 1292 3836
rect 1316 3834 1372 3836
rect 1396 3834 1452 3836
rect 1156 3782 1202 3834
rect 1202 3782 1212 3834
rect 1236 3782 1266 3834
rect 1266 3782 1278 3834
rect 1278 3782 1292 3834
rect 1316 3782 1330 3834
rect 1330 3782 1342 3834
rect 1342 3782 1372 3834
rect 1396 3782 1406 3834
rect 1406 3782 1452 3834
rect 1156 3780 1212 3782
rect 1236 3780 1292 3782
rect 1316 3780 1372 3782
rect 1396 3780 1452 3782
rect 4342 6704 4398 6760
rect 3156 6554 3212 6556
rect 3236 6554 3292 6556
rect 3316 6554 3372 6556
rect 3396 6554 3452 6556
rect 3156 6502 3202 6554
rect 3202 6502 3212 6554
rect 3236 6502 3266 6554
rect 3266 6502 3278 6554
rect 3278 6502 3292 6554
rect 3316 6502 3330 6554
rect 3330 6502 3342 6554
rect 3342 6502 3372 6554
rect 3396 6502 3406 6554
rect 3406 6502 3452 6554
rect 3156 6500 3212 6502
rect 3236 6500 3292 6502
rect 3316 6500 3372 6502
rect 3396 6500 3452 6502
rect 3156 5466 3212 5468
rect 3236 5466 3292 5468
rect 3316 5466 3372 5468
rect 3396 5466 3452 5468
rect 3156 5414 3202 5466
rect 3202 5414 3212 5466
rect 3236 5414 3266 5466
rect 3266 5414 3278 5466
rect 3278 5414 3292 5466
rect 3316 5414 3330 5466
rect 3330 5414 3342 5466
rect 3342 5414 3372 5466
rect 3396 5414 3406 5466
rect 3406 5414 3452 5466
rect 3156 5412 3212 5414
rect 3236 5412 3292 5414
rect 3316 5412 3372 5414
rect 3396 5412 3452 5414
rect 3156 4378 3212 4380
rect 3236 4378 3292 4380
rect 3316 4378 3372 4380
rect 3396 4378 3452 4380
rect 3156 4326 3202 4378
rect 3202 4326 3212 4378
rect 3236 4326 3266 4378
rect 3266 4326 3278 4378
rect 3278 4326 3292 4378
rect 3316 4326 3330 4378
rect 3330 4326 3342 4378
rect 3342 4326 3372 4378
rect 3396 4326 3406 4378
rect 3406 4326 3452 4378
rect 3156 4324 3212 4326
rect 3236 4324 3292 4326
rect 3316 4324 3372 4326
rect 3396 4324 3452 4326
rect 4066 4156 4068 4176
rect 4068 4156 4120 4176
rect 4120 4156 4122 4176
rect 4066 4120 4122 4156
rect 1156 2746 1212 2748
rect 1236 2746 1292 2748
rect 1316 2746 1372 2748
rect 1396 2746 1452 2748
rect 1156 2694 1202 2746
rect 1202 2694 1212 2746
rect 1236 2694 1266 2746
rect 1266 2694 1278 2746
rect 1278 2694 1292 2746
rect 1316 2694 1330 2746
rect 1330 2694 1342 2746
rect 1342 2694 1372 2746
rect 1396 2694 1406 2746
rect 1406 2694 1452 2746
rect 1156 2692 1212 2694
rect 1236 2692 1292 2694
rect 1316 2692 1372 2694
rect 1396 2692 1452 2694
rect 1156 1658 1212 1660
rect 1236 1658 1292 1660
rect 1316 1658 1372 1660
rect 1396 1658 1452 1660
rect 1156 1606 1202 1658
rect 1202 1606 1212 1658
rect 1236 1606 1266 1658
rect 1266 1606 1278 1658
rect 1278 1606 1292 1658
rect 1316 1606 1330 1658
rect 1330 1606 1342 1658
rect 1342 1606 1372 1658
rect 1396 1606 1406 1658
rect 1406 1606 1452 1658
rect 1156 1604 1212 1606
rect 1236 1604 1292 1606
rect 1316 1604 1372 1606
rect 1396 1604 1452 1606
rect 2778 3440 2834 3496
rect 3156 3290 3212 3292
rect 3236 3290 3292 3292
rect 3316 3290 3372 3292
rect 3396 3290 3452 3292
rect 3156 3238 3202 3290
rect 3202 3238 3212 3290
rect 3236 3238 3266 3290
rect 3266 3238 3278 3290
rect 3278 3238 3292 3290
rect 3316 3238 3330 3290
rect 3330 3238 3342 3290
rect 3342 3238 3372 3290
rect 3396 3238 3406 3290
rect 3406 3238 3452 3290
rect 3156 3236 3212 3238
rect 3236 3236 3292 3238
rect 3316 3236 3372 3238
rect 3396 3236 3452 3238
rect 1582 1400 1638 1456
rect 3156 2202 3212 2204
rect 3236 2202 3292 2204
rect 3316 2202 3372 2204
rect 3396 2202 3452 2204
rect 3156 2150 3202 2202
rect 3202 2150 3212 2202
rect 3236 2150 3266 2202
rect 3266 2150 3278 2202
rect 3278 2150 3292 2202
rect 3316 2150 3330 2202
rect 3330 2150 3342 2202
rect 3342 2150 3372 2202
rect 3396 2150 3406 2202
rect 3406 2150 3452 2202
rect 3156 2148 3212 2150
rect 3236 2148 3292 2150
rect 3316 2148 3372 2150
rect 3396 2148 3452 2150
rect 4066 1944 4122 2000
rect 4250 2352 4306 2408
rect 6734 8200 6790 8256
rect 5156 7098 5212 7100
rect 5236 7098 5292 7100
rect 5316 7098 5372 7100
rect 5396 7098 5452 7100
rect 5156 7046 5202 7098
rect 5202 7046 5212 7098
rect 5236 7046 5266 7098
rect 5266 7046 5278 7098
rect 5278 7046 5292 7098
rect 5316 7046 5330 7098
rect 5330 7046 5342 7098
rect 5342 7046 5372 7098
rect 5396 7046 5406 7098
rect 5406 7046 5452 7098
rect 5156 7044 5212 7046
rect 5236 7044 5292 7046
rect 5316 7044 5372 7046
rect 5396 7044 5452 7046
rect 5156 6010 5212 6012
rect 5236 6010 5292 6012
rect 5316 6010 5372 6012
rect 5396 6010 5452 6012
rect 5156 5958 5202 6010
rect 5202 5958 5212 6010
rect 5236 5958 5266 6010
rect 5266 5958 5278 6010
rect 5278 5958 5292 6010
rect 5316 5958 5330 6010
rect 5330 5958 5342 6010
rect 5342 5958 5372 6010
rect 5396 5958 5406 6010
rect 5406 5958 5452 6010
rect 5156 5956 5212 5958
rect 5236 5956 5292 5958
rect 5316 5956 5372 5958
rect 5396 5956 5452 5958
rect 5156 4922 5212 4924
rect 5236 4922 5292 4924
rect 5316 4922 5372 4924
rect 5396 4922 5452 4924
rect 5156 4870 5202 4922
rect 5202 4870 5212 4922
rect 5236 4870 5266 4922
rect 5266 4870 5278 4922
rect 5278 4870 5292 4922
rect 5316 4870 5330 4922
rect 5330 4870 5342 4922
rect 5342 4870 5372 4922
rect 5396 4870 5406 4922
rect 5406 4870 5452 4922
rect 5156 4868 5212 4870
rect 5236 4868 5292 4870
rect 5316 4868 5372 4870
rect 5396 4868 5452 4870
rect 5156 3834 5212 3836
rect 5236 3834 5292 3836
rect 5316 3834 5372 3836
rect 5396 3834 5452 3836
rect 5156 3782 5202 3834
rect 5202 3782 5212 3834
rect 5236 3782 5266 3834
rect 5266 3782 5278 3834
rect 5278 3782 5292 3834
rect 5316 3782 5330 3834
rect 5330 3782 5342 3834
rect 5342 3782 5372 3834
rect 5396 3782 5406 3834
rect 5406 3782 5452 3834
rect 5156 3780 5212 3782
rect 5236 3780 5292 3782
rect 5316 3780 5372 3782
rect 5396 3780 5452 3782
rect 5078 2896 5134 2952
rect 5156 2746 5212 2748
rect 5236 2746 5292 2748
rect 5316 2746 5372 2748
rect 5396 2746 5452 2748
rect 5156 2694 5202 2746
rect 5202 2694 5212 2746
rect 5236 2694 5266 2746
rect 5266 2694 5278 2746
rect 5278 2694 5292 2746
rect 5316 2694 5330 2746
rect 5330 2694 5342 2746
rect 5342 2694 5372 2746
rect 5396 2694 5406 2746
rect 5406 2694 5452 2746
rect 5156 2692 5212 2694
rect 5236 2692 5292 2694
rect 5316 2692 5372 2694
rect 5396 2692 5452 2694
rect 5156 1658 5212 1660
rect 5236 1658 5292 1660
rect 5316 1658 5372 1660
rect 5396 1658 5452 1660
rect 5156 1606 5202 1658
rect 5202 1606 5212 1658
rect 5236 1606 5266 1658
rect 5266 1606 5278 1658
rect 5278 1606 5292 1658
rect 5316 1606 5330 1658
rect 5330 1606 5342 1658
rect 5342 1606 5372 1658
rect 5396 1606 5406 1658
rect 5406 1606 5452 1658
rect 5156 1604 5212 1606
rect 5236 1604 5292 1606
rect 5316 1604 5372 1606
rect 5396 1604 5452 1606
rect 3156 1114 3212 1116
rect 3236 1114 3292 1116
rect 3316 1114 3372 1116
rect 3396 1114 3452 1116
rect 3156 1062 3202 1114
rect 3202 1062 3212 1114
rect 3236 1062 3266 1114
rect 3266 1062 3278 1114
rect 3278 1062 3292 1114
rect 3316 1062 3330 1114
rect 3330 1062 3342 1114
rect 3342 1062 3372 1114
rect 3396 1062 3406 1114
rect 3406 1062 3452 1114
rect 3156 1060 3212 1062
rect 3236 1060 3292 1062
rect 3316 1060 3372 1062
rect 3396 1060 3452 1062
rect 7156 7642 7212 7644
rect 7236 7642 7292 7644
rect 7316 7642 7372 7644
rect 7396 7642 7452 7644
rect 7156 7590 7202 7642
rect 7202 7590 7212 7642
rect 7236 7590 7266 7642
rect 7266 7590 7278 7642
rect 7278 7590 7292 7642
rect 7316 7590 7330 7642
rect 7330 7590 7342 7642
rect 7342 7590 7372 7642
rect 7396 7590 7406 7642
rect 7406 7590 7452 7642
rect 7156 7588 7212 7590
rect 7236 7588 7292 7590
rect 7316 7588 7372 7590
rect 7396 7588 7452 7590
rect 7562 7520 7618 7576
rect 7156 6554 7212 6556
rect 7236 6554 7292 6556
rect 7316 6554 7372 6556
rect 7396 6554 7452 6556
rect 7156 6502 7202 6554
rect 7202 6502 7212 6554
rect 7236 6502 7266 6554
rect 7266 6502 7278 6554
rect 7278 6502 7292 6554
rect 7316 6502 7330 6554
rect 7330 6502 7342 6554
rect 7342 6502 7372 6554
rect 7396 6502 7406 6554
rect 7406 6502 7452 6554
rect 7156 6500 7212 6502
rect 7236 6500 7292 6502
rect 7316 6500 7372 6502
rect 7396 6500 7452 6502
rect 7562 5480 7618 5536
rect 7156 5466 7212 5468
rect 7236 5466 7292 5468
rect 7316 5466 7372 5468
rect 7396 5466 7452 5468
rect 7156 5414 7202 5466
rect 7202 5414 7212 5466
rect 7236 5414 7266 5466
rect 7266 5414 7278 5466
rect 7278 5414 7292 5466
rect 7316 5414 7330 5466
rect 7330 5414 7342 5466
rect 7342 5414 7372 5466
rect 7396 5414 7406 5466
rect 7406 5414 7452 5466
rect 7156 5412 7212 5414
rect 7236 5412 7292 5414
rect 7316 5412 7372 5414
rect 7396 5412 7452 5414
rect 6826 4820 6882 4856
rect 6826 4800 6828 4820
rect 6828 4800 6880 4820
rect 6880 4800 6882 4820
rect 7156 4378 7212 4380
rect 7236 4378 7292 4380
rect 7316 4378 7372 4380
rect 7396 4378 7452 4380
rect 7156 4326 7202 4378
rect 7202 4326 7212 4378
rect 7236 4326 7266 4378
rect 7266 4326 7278 4378
rect 7278 4326 7292 4378
rect 7316 4326 7330 4378
rect 7330 4326 7342 4378
rect 7342 4326 7372 4378
rect 7396 4326 7406 4378
rect 7406 4326 7452 4378
rect 7156 4324 7212 4326
rect 7236 4324 7292 4326
rect 7316 4324 7372 4326
rect 7396 4324 7452 4326
rect 7286 4140 7342 4176
rect 7286 4120 7288 4140
rect 7288 4120 7340 4140
rect 7340 4120 7342 4140
rect 5906 1400 5962 1456
rect 7156 3290 7212 3292
rect 7236 3290 7292 3292
rect 7316 3290 7372 3292
rect 7396 3290 7452 3292
rect 7156 3238 7202 3290
rect 7202 3238 7212 3290
rect 7236 3238 7266 3290
rect 7266 3238 7278 3290
rect 7278 3238 7292 3290
rect 7316 3238 7330 3290
rect 7330 3238 7342 3290
rect 7342 3238 7372 3290
rect 7396 3238 7406 3290
rect 7406 3238 7452 3290
rect 7156 3236 7212 3238
rect 7236 3236 7292 3238
rect 7316 3236 7372 3238
rect 7396 3236 7452 3238
rect 7156 2202 7212 2204
rect 7236 2202 7292 2204
rect 7316 2202 7372 2204
rect 7396 2202 7452 2204
rect 7156 2150 7202 2202
rect 7202 2150 7212 2202
rect 7236 2150 7266 2202
rect 7266 2150 7278 2202
rect 7278 2150 7292 2202
rect 7316 2150 7330 2202
rect 7330 2150 7342 2202
rect 7342 2150 7372 2202
rect 7396 2150 7406 2202
rect 7406 2150 7452 2202
rect 7156 2148 7212 2150
rect 7236 2148 7292 2150
rect 7316 2148 7372 2150
rect 7396 2148 7452 2150
rect 7156 1114 7212 1116
rect 7236 1114 7292 1116
rect 7316 1114 7372 1116
rect 7396 1114 7452 1116
rect 7156 1062 7202 1114
rect 7202 1062 7212 1114
rect 7236 1062 7266 1114
rect 7266 1062 7278 1114
rect 7278 1062 7292 1114
rect 7316 1062 7330 1114
rect 7330 1062 7342 1114
rect 7342 1062 7372 1114
rect 7396 1062 7406 1114
rect 7406 1062 7452 1114
rect 7156 1060 7212 1062
rect 7236 1060 7292 1062
rect 7316 1060 7372 1062
rect 7396 1060 7452 1062
rect 1490 720 1546 776
rect 7838 40 7894 96
<< metal3 >>
rect 0 8938 800 8968
rect 2865 8938 2931 8941
rect 0 8936 2931 8938
rect 0 8880 2870 8936
rect 2926 8880 2931 8936
rect 0 8878 2931 8880
rect 0 8848 800 8878
rect 2865 8875 2931 8878
rect 6729 8258 6795 8261
rect 8200 8258 9000 8288
rect 6729 8256 9000 8258
rect 6729 8200 6734 8256
rect 6790 8200 9000 8256
rect 6729 8198 9000 8200
rect 6729 8195 6795 8198
rect 8200 8168 9000 8198
rect 3146 7648 3462 7649
rect 0 7578 800 7608
rect 3146 7584 3152 7648
rect 3216 7584 3232 7648
rect 3296 7584 3312 7648
rect 3376 7584 3392 7648
rect 3456 7584 3462 7648
rect 3146 7583 3462 7584
rect 7146 7648 7462 7649
rect 7146 7584 7152 7648
rect 7216 7584 7232 7648
rect 7296 7584 7312 7648
rect 7376 7584 7392 7648
rect 7456 7584 7462 7648
rect 7146 7583 7462 7584
rect 1577 7578 1643 7581
rect 0 7576 1643 7578
rect 0 7520 1582 7576
rect 1638 7520 1643 7576
rect 0 7518 1643 7520
rect 0 7488 800 7518
rect 1577 7515 1643 7518
rect 7557 7578 7623 7581
rect 8200 7578 9000 7608
rect 7557 7576 9000 7578
rect 7557 7520 7562 7576
rect 7618 7520 9000 7576
rect 7557 7518 9000 7520
rect 7557 7515 7623 7518
rect 8200 7488 9000 7518
rect 1146 7104 1462 7105
rect 1146 7040 1152 7104
rect 1216 7040 1232 7104
rect 1296 7040 1312 7104
rect 1376 7040 1392 7104
rect 1456 7040 1462 7104
rect 1146 7039 1462 7040
rect 5146 7104 5462 7105
rect 5146 7040 5152 7104
rect 5216 7040 5232 7104
rect 5296 7040 5312 7104
rect 5376 7040 5392 7104
rect 5456 7040 5462 7104
rect 5146 7039 5462 7040
rect 0 6898 800 6928
rect 4245 6898 4311 6901
rect 8200 6898 9000 6928
rect 0 6838 3986 6898
rect 0 6808 800 6838
rect 3926 6762 3986 6838
rect 4245 6896 9000 6898
rect 4245 6840 4250 6896
rect 4306 6840 9000 6896
rect 4245 6838 9000 6840
rect 4245 6835 4311 6838
rect 8200 6808 9000 6838
rect 4337 6762 4403 6765
rect 3926 6760 4403 6762
rect 3926 6704 4342 6760
rect 4398 6704 4403 6760
rect 3926 6702 4403 6704
rect 4337 6699 4403 6702
rect 3146 6560 3462 6561
rect 3146 6496 3152 6560
rect 3216 6496 3232 6560
rect 3296 6496 3312 6560
rect 3376 6496 3392 6560
rect 3456 6496 3462 6560
rect 3146 6495 3462 6496
rect 7146 6560 7462 6561
rect 7146 6496 7152 6560
rect 7216 6496 7232 6560
rect 7296 6496 7312 6560
rect 7376 6496 7392 6560
rect 7456 6496 7462 6560
rect 7146 6495 7462 6496
rect 0 6218 800 6248
rect 1577 6218 1643 6221
rect 0 6216 1643 6218
rect 0 6160 1582 6216
rect 1638 6160 1643 6216
rect 0 6158 1643 6160
rect 0 6128 800 6158
rect 1577 6155 1643 6158
rect 1146 6016 1462 6017
rect 1146 5952 1152 6016
rect 1216 5952 1232 6016
rect 1296 5952 1312 6016
rect 1376 5952 1392 6016
rect 1456 5952 1462 6016
rect 1146 5951 1462 5952
rect 5146 6016 5462 6017
rect 5146 5952 5152 6016
rect 5216 5952 5232 6016
rect 5296 5952 5312 6016
rect 5376 5952 5392 6016
rect 5456 5952 5462 6016
rect 5146 5951 5462 5952
rect 7557 5538 7623 5541
rect 8200 5538 9000 5568
rect 7557 5536 9000 5538
rect 7557 5480 7562 5536
rect 7618 5480 9000 5536
rect 7557 5478 9000 5480
rect 7557 5475 7623 5478
rect 3146 5472 3462 5473
rect 3146 5408 3152 5472
rect 3216 5408 3232 5472
rect 3296 5408 3312 5472
rect 3376 5408 3392 5472
rect 3456 5408 3462 5472
rect 3146 5407 3462 5408
rect 7146 5472 7462 5473
rect 7146 5408 7152 5472
rect 7216 5408 7232 5472
rect 7296 5408 7312 5472
rect 7376 5408 7392 5472
rect 7456 5408 7462 5472
rect 8200 5448 9000 5478
rect 7146 5407 7462 5408
rect 1577 5130 1643 5133
rect 982 5128 1643 5130
rect 982 5072 1582 5128
rect 1638 5072 1643 5128
rect 982 5070 1643 5072
rect 0 4858 800 4888
rect 982 4858 1042 5070
rect 1577 5067 1643 5070
rect 1146 4928 1462 4929
rect 1146 4864 1152 4928
rect 1216 4864 1232 4928
rect 1296 4864 1312 4928
rect 1376 4864 1392 4928
rect 1456 4864 1462 4928
rect 1146 4863 1462 4864
rect 5146 4928 5462 4929
rect 5146 4864 5152 4928
rect 5216 4864 5232 4928
rect 5296 4864 5312 4928
rect 5376 4864 5392 4928
rect 5456 4864 5462 4928
rect 5146 4863 5462 4864
rect 0 4798 1042 4858
rect 6821 4858 6887 4861
rect 8200 4858 9000 4888
rect 6821 4856 9000 4858
rect 6821 4800 6826 4856
rect 6882 4800 9000 4856
rect 6821 4798 9000 4800
rect 0 4768 800 4798
rect 6821 4795 6887 4798
rect 8200 4768 9000 4798
rect 3146 4384 3462 4385
rect 3146 4320 3152 4384
rect 3216 4320 3232 4384
rect 3296 4320 3312 4384
rect 3376 4320 3392 4384
rect 3456 4320 3462 4384
rect 3146 4319 3462 4320
rect 7146 4384 7462 4385
rect 7146 4320 7152 4384
rect 7216 4320 7232 4384
rect 7296 4320 7312 4384
rect 7376 4320 7392 4384
rect 7456 4320 7462 4384
rect 7146 4319 7462 4320
rect 0 4178 800 4208
rect 4061 4178 4127 4181
rect 0 4176 4127 4178
rect 0 4120 4066 4176
rect 4122 4120 4127 4176
rect 0 4118 4127 4120
rect 0 4088 800 4118
rect 4061 4115 4127 4118
rect 7281 4178 7347 4181
rect 8200 4178 9000 4208
rect 7281 4176 9000 4178
rect 7281 4120 7286 4176
rect 7342 4120 9000 4176
rect 7281 4118 9000 4120
rect 7281 4115 7347 4118
rect 8200 4088 9000 4118
rect 1146 3840 1462 3841
rect 1146 3776 1152 3840
rect 1216 3776 1232 3840
rect 1296 3776 1312 3840
rect 1376 3776 1392 3840
rect 1456 3776 1462 3840
rect 1146 3775 1462 3776
rect 5146 3840 5462 3841
rect 5146 3776 5152 3840
rect 5216 3776 5232 3840
rect 5296 3776 5312 3840
rect 5376 3776 5392 3840
rect 5456 3776 5462 3840
rect 5146 3775 5462 3776
rect 0 3498 800 3528
rect 2773 3498 2839 3501
rect 0 3496 2839 3498
rect 0 3440 2778 3496
rect 2834 3440 2839 3496
rect 0 3438 2839 3440
rect 0 3408 800 3438
rect 2773 3435 2839 3438
rect 3146 3296 3462 3297
rect 3146 3232 3152 3296
rect 3216 3232 3232 3296
rect 3296 3232 3312 3296
rect 3376 3232 3392 3296
rect 3456 3232 3462 3296
rect 3146 3231 3462 3232
rect 7146 3296 7462 3297
rect 7146 3232 7152 3296
rect 7216 3232 7232 3296
rect 7296 3232 7312 3296
rect 7376 3232 7392 3296
rect 7456 3232 7462 3296
rect 7146 3231 7462 3232
rect 5073 2954 5139 2957
rect 5073 2952 6930 2954
rect 5073 2896 5078 2952
rect 5134 2896 6930 2952
rect 5073 2894 6930 2896
rect 5073 2891 5139 2894
rect 6870 2818 6930 2894
rect 8200 2818 9000 2848
rect 6870 2758 9000 2818
rect 1146 2752 1462 2753
rect 1146 2688 1152 2752
rect 1216 2688 1232 2752
rect 1296 2688 1312 2752
rect 1376 2688 1392 2752
rect 1456 2688 1462 2752
rect 1146 2687 1462 2688
rect 5146 2752 5462 2753
rect 5146 2688 5152 2752
rect 5216 2688 5232 2752
rect 5296 2688 5312 2752
rect 5376 2688 5392 2752
rect 5456 2688 5462 2752
rect 8200 2728 9000 2758
rect 5146 2687 5462 2688
rect 4245 2410 4311 2413
rect 4245 2408 7666 2410
rect 4245 2352 4250 2408
rect 4306 2352 7666 2408
rect 4245 2350 7666 2352
rect 4245 2347 4311 2350
rect 3146 2208 3462 2209
rect 0 2138 800 2168
rect 3146 2144 3152 2208
rect 3216 2144 3232 2208
rect 3296 2144 3312 2208
rect 3376 2144 3392 2208
rect 3456 2144 3462 2208
rect 3146 2143 3462 2144
rect 7146 2208 7462 2209
rect 7146 2144 7152 2208
rect 7216 2144 7232 2208
rect 7296 2144 7312 2208
rect 7376 2144 7392 2208
rect 7456 2144 7462 2208
rect 7146 2143 7462 2144
rect 7606 2138 7666 2350
rect 8200 2138 9000 2168
rect 0 2078 2146 2138
rect 7606 2078 9000 2138
rect 0 2048 800 2078
rect 2086 2002 2146 2078
rect 8200 2048 9000 2078
rect 4061 2002 4127 2005
rect 2086 2000 4127 2002
rect 2086 1944 4066 2000
rect 4122 1944 4127 2000
rect 2086 1942 4127 1944
rect 4061 1939 4127 1942
rect 1146 1664 1462 1665
rect 1146 1600 1152 1664
rect 1216 1600 1232 1664
rect 1296 1600 1312 1664
rect 1376 1600 1392 1664
rect 1456 1600 1462 1664
rect 1146 1599 1462 1600
rect 5146 1664 5462 1665
rect 5146 1600 5152 1664
rect 5216 1600 5232 1664
rect 5296 1600 5312 1664
rect 5376 1600 5392 1664
rect 5456 1600 5462 1664
rect 5146 1599 5462 1600
rect 0 1458 800 1488
rect 1577 1458 1643 1461
rect 0 1456 1643 1458
rect 0 1400 1582 1456
rect 1638 1400 1643 1456
rect 0 1398 1643 1400
rect 0 1368 800 1398
rect 1577 1395 1643 1398
rect 5901 1458 5967 1461
rect 8200 1458 9000 1488
rect 5901 1456 9000 1458
rect 5901 1400 5906 1456
rect 5962 1400 9000 1456
rect 5901 1398 9000 1400
rect 5901 1395 5967 1398
rect 8200 1368 9000 1398
rect 3146 1120 3462 1121
rect 3146 1056 3152 1120
rect 3216 1056 3232 1120
rect 3296 1056 3312 1120
rect 3376 1056 3392 1120
rect 3456 1056 3462 1120
rect 3146 1055 3462 1056
rect 7146 1120 7462 1121
rect 7146 1056 7152 1120
rect 7216 1056 7232 1120
rect 7296 1056 7312 1120
rect 7376 1056 7392 1120
rect 7456 1056 7462 1120
rect 7146 1055 7462 1056
rect 0 778 800 808
rect 1485 778 1551 781
rect 0 776 1551 778
rect 0 720 1490 776
rect 1546 720 1551 776
rect 0 718 1551 720
rect 0 688 800 718
rect 1485 715 1551 718
rect 7833 98 7899 101
rect 8200 98 9000 128
rect 7833 96 9000 98
rect 7833 40 7838 96
rect 7894 40 9000 96
rect 7833 38 9000 40
rect 7833 35 7899 38
rect 8200 8 9000 38
<< via3 >>
rect 3152 7644 3216 7648
rect 3152 7588 3156 7644
rect 3156 7588 3212 7644
rect 3212 7588 3216 7644
rect 3152 7584 3216 7588
rect 3232 7644 3296 7648
rect 3232 7588 3236 7644
rect 3236 7588 3292 7644
rect 3292 7588 3296 7644
rect 3232 7584 3296 7588
rect 3312 7644 3376 7648
rect 3312 7588 3316 7644
rect 3316 7588 3372 7644
rect 3372 7588 3376 7644
rect 3312 7584 3376 7588
rect 3392 7644 3456 7648
rect 3392 7588 3396 7644
rect 3396 7588 3452 7644
rect 3452 7588 3456 7644
rect 3392 7584 3456 7588
rect 7152 7644 7216 7648
rect 7152 7588 7156 7644
rect 7156 7588 7212 7644
rect 7212 7588 7216 7644
rect 7152 7584 7216 7588
rect 7232 7644 7296 7648
rect 7232 7588 7236 7644
rect 7236 7588 7292 7644
rect 7292 7588 7296 7644
rect 7232 7584 7296 7588
rect 7312 7644 7376 7648
rect 7312 7588 7316 7644
rect 7316 7588 7372 7644
rect 7372 7588 7376 7644
rect 7312 7584 7376 7588
rect 7392 7644 7456 7648
rect 7392 7588 7396 7644
rect 7396 7588 7452 7644
rect 7452 7588 7456 7644
rect 7392 7584 7456 7588
rect 1152 7100 1216 7104
rect 1152 7044 1156 7100
rect 1156 7044 1212 7100
rect 1212 7044 1216 7100
rect 1152 7040 1216 7044
rect 1232 7100 1296 7104
rect 1232 7044 1236 7100
rect 1236 7044 1292 7100
rect 1292 7044 1296 7100
rect 1232 7040 1296 7044
rect 1312 7100 1376 7104
rect 1312 7044 1316 7100
rect 1316 7044 1372 7100
rect 1372 7044 1376 7100
rect 1312 7040 1376 7044
rect 1392 7100 1456 7104
rect 1392 7044 1396 7100
rect 1396 7044 1452 7100
rect 1452 7044 1456 7100
rect 1392 7040 1456 7044
rect 5152 7100 5216 7104
rect 5152 7044 5156 7100
rect 5156 7044 5212 7100
rect 5212 7044 5216 7100
rect 5152 7040 5216 7044
rect 5232 7100 5296 7104
rect 5232 7044 5236 7100
rect 5236 7044 5292 7100
rect 5292 7044 5296 7100
rect 5232 7040 5296 7044
rect 5312 7100 5376 7104
rect 5312 7044 5316 7100
rect 5316 7044 5372 7100
rect 5372 7044 5376 7100
rect 5312 7040 5376 7044
rect 5392 7100 5456 7104
rect 5392 7044 5396 7100
rect 5396 7044 5452 7100
rect 5452 7044 5456 7100
rect 5392 7040 5456 7044
rect 3152 6556 3216 6560
rect 3152 6500 3156 6556
rect 3156 6500 3212 6556
rect 3212 6500 3216 6556
rect 3152 6496 3216 6500
rect 3232 6556 3296 6560
rect 3232 6500 3236 6556
rect 3236 6500 3292 6556
rect 3292 6500 3296 6556
rect 3232 6496 3296 6500
rect 3312 6556 3376 6560
rect 3312 6500 3316 6556
rect 3316 6500 3372 6556
rect 3372 6500 3376 6556
rect 3312 6496 3376 6500
rect 3392 6556 3456 6560
rect 3392 6500 3396 6556
rect 3396 6500 3452 6556
rect 3452 6500 3456 6556
rect 3392 6496 3456 6500
rect 7152 6556 7216 6560
rect 7152 6500 7156 6556
rect 7156 6500 7212 6556
rect 7212 6500 7216 6556
rect 7152 6496 7216 6500
rect 7232 6556 7296 6560
rect 7232 6500 7236 6556
rect 7236 6500 7292 6556
rect 7292 6500 7296 6556
rect 7232 6496 7296 6500
rect 7312 6556 7376 6560
rect 7312 6500 7316 6556
rect 7316 6500 7372 6556
rect 7372 6500 7376 6556
rect 7312 6496 7376 6500
rect 7392 6556 7456 6560
rect 7392 6500 7396 6556
rect 7396 6500 7452 6556
rect 7452 6500 7456 6556
rect 7392 6496 7456 6500
rect 1152 6012 1216 6016
rect 1152 5956 1156 6012
rect 1156 5956 1212 6012
rect 1212 5956 1216 6012
rect 1152 5952 1216 5956
rect 1232 6012 1296 6016
rect 1232 5956 1236 6012
rect 1236 5956 1292 6012
rect 1292 5956 1296 6012
rect 1232 5952 1296 5956
rect 1312 6012 1376 6016
rect 1312 5956 1316 6012
rect 1316 5956 1372 6012
rect 1372 5956 1376 6012
rect 1312 5952 1376 5956
rect 1392 6012 1456 6016
rect 1392 5956 1396 6012
rect 1396 5956 1452 6012
rect 1452 5956 1456 6012
rect 1392 5952 1456 5956
rect 5152 6012 5216 6016
rect 5152 5956 5156 6012
rect 5156 5956 5212 6012
rect 5212 5956 5216 6012
rect 5152 5952 5216 5956
rect 5232 6012 5296 6016
rect 5232 5956 5236 6012
rect 5236 5956 5292 6012
rect 5292 5956 5296 6012
rect 5232 5952 5296 5956
rect 5312 6012 5376 6016
rect 5312 5956 5316 6012
rect 5316 5956 5372 6012
rect 5372 5956 5376 6012
rect 5312 5952 5376 5956
rect 5392 6012 5456 6016
rect 5392 5956 5396 6012
rect 5396 5956 5452 6012
rect 5452 5956 5456 6012
rect 5392 5952 5456 5956
rect 3152 5468 3216 5472
rect 3152 5412 3156 5468
rect 3156 5412 3212 5468
rect 3212 5412 3216 5468
rect 3152 5408 3216 5412
rect 3232 5468 3296 5472
rect 3232 5412 3236 5468
rect 3236 5412 3292 5468
rect 3292 5412 3296 5468
rect 3232 5408 3296 5412
rect 3312 5468 3376 5472
rect 3312 5412 3316 5468
rect 3316 5412 3372 5468
rect 3372 5412 3376 5468
rect 3312 5408 3376 5412
rect 3392 5468 3456 5472
rect 3392 5412 3396 5468
rect 3396 5412 3452 5468
rect 3452 5412 3456 5468
rect 3392 5408 3456 5412
rect 7152 5468 7216 5472
rect 7152 5412 7156 5468
rect 7156 5412 7212 5468
rect 7212 5412 7216 5468
rect 7152 5408 7216 5412
rect 7232 5468 7296 5472
rect 7232 5412 7236 5468
rect 7236 5412 7292 5468
rect 7292 5412 7296 5468
rect 7232 5408 7296 5412
rect 7312 5468 7376 5472
rect 7312 5412 7316 5468
rect 7316 5412 7372 5468
rect 7372 5412 7376 5468
rect 7312 5408 7376 5412
rect 7392 5468 7456 5472
rect 7392 5412 7396 5468
rect 7396 5412 7452 5468
rect 7452 5412 7456 5468
rect 7392 5408 7456 5412
rect 1152 4924 1216 4928
rect 1152 4868 1156 4924
rect 1156 4868 1212 4924
rect 1212 4868 1216 4924
rect 1152 4864 1216 4868
rect 1232 4924 1296 4928
rect 1232 4868 1236 4924
rect 1236 4868 1292 4924
rect 1292 4868 1296 4924
rect 1232 4864 1296 4868
rect 1312 4924 1376 4928
rect 1312 4868 1316 4924
rect 1316 4868 1372 4924
rect 1372 4868 1376 4924
rect 1312 4864 1376 4868
rect 1392 4924 1456 4928
rect 1392 4868 1396 4924
rect 1396 4868 1452 4924
rect 1452 4868 1456 4924
rect 1392 4864 1456 4868
rect 5152 4924 5216 4928
rect 5152 4868 5156 4924
rect 5156 4868 5212 4924
rect 5212 4868 5216 4924
rect 5152 4864 5216 4868
rect 5232 4924 5296 4928
rect 5232 4868 5236 4924
rect 5236 4868 5292 4924
rect 5292 4868 5296 4924
rect 5232 4864 5296 4868
rect 5312 4924 5376 4928
rect 5312 4868 5316 4924
rect 5316 4868 5372 4924
rect 5372 4868 5376 4924
rect 5312 4864 5376 4868
rect 5392 4924 5456 4928
rect 5392 4868 5396 4924
rect 5396 4868 5452 4924
rect 5452 4868 5456 4924
rect 5392 4864 5456 4868
rect 3152 4380 3216 4384
rect 3152 4324 3156 4380
rect 3156 4324 3212 4380
rect 3212 4324 3216 4380
rect 3152 4320 3216 4324
rect 3232 4380 3296 4384
rect 3232 4324 3236 4380
rect 3236 4324 3292 4380
rect 3292 4324 3296 4380
rect 3232 4320 3296 4324
rect 3312 4380 3376 4384
rect 3312 4324 3316 4380
rect 3316 4324 3372 4380
rect 3372 4324 3376 4380
rect 3312 4320 3376 4324
rect 3392 4380 3456 4384
rect 3392 4324 3396 4380
rect 3396 4324 3452 4380
rect 3452 4324 3456 4380
rect 3392 4320 3456 4324
rect 7152 4380 7216 4384
rect 7152 4324 7156 4380
rect 7156 4324 7212 4380
rect 7212 4324 7216 4380
rect 7152 4320 7216 4324
rect 7232 4380 7296 4384
rect 7232 4324 7236 4380
rect 7236 4324 7292 4380
rect 7292 4324 7296 4380
rect 7232 4320 7296 4324
rect 7312 4380 7376 4384
rect 7312 4324 7316 4380
rect 7316 4324 7372 4380
rect 7372 4324 7376 4380
rect 7312 4320 7376 4324
rect 7392 4380 7456 4384
rect 7392 4324 7396 4380
rect 7396 4324 7452 4380
rect 7452 4324 7456 4380
rect 7392 4320 7456 4324
rect 1152 3836 1216 3840
rect 1152 3780 1156 3836
rect 1156 3780 1212 3836
rect 1212 3780 1216 3836
rect 1152 3776 1216 3780
rect 1232 3836 1296 3840
rect 1232 3780 1236 3836
rect 1236 3780 1292 3836
rect 1292 3780 1296 3836
rect 1232 3776 1296 3780
rect 1312 3836 1376 3840
rect 1312 3780 1316 3836
rect 1316 3780 1372 3836
rect 1372 3780 1376 3836
rect 1312 3776 1376 3780
rect 1392 3836 1456 3840
rect 1392 3780 1396 3836
rect 1396 3780 1452 3836
rect 1452 3780 1456 3836
rect 1392 3776 1456 3780
rect 5152 3836 5216 3840
rect 5152 3780 5156 3836
rect 5156 3780 5212 3836
rect 5212 3780 5216 3836
rect 5152 3776 5216 3780
rect 5232 3836 5296 3840
rect 5232 3780 5236 3836
rect 5236 3780 5292 3836
rect 5292 3780 5296 3836
rect 5232 3776 5296 3780
rect 5312 3836 5376 3840
rect 5312 3780 5316 3836
rect 5316 3780 5372 3836
rect 5372 3780 5376 3836
rect 5312 3776 5376 3780
rect 5392 3836 5456 3840
rect 5392 3780 5396 3836
rect 5396 3780 5452 3836
rect 5452 3780 5456 3836
rect 5392 3776 5456 3780
rect 3152 3292 3216 3296
rect 3152 3236 3156 3292
rect 3156 3236 3212 3292
rect 3212 3236 3216 3292
rect 3152 3232 3216 3236
rect 3232 3292 3296 3296
rect 3232 3236 3236 3292
rect 3236 3236 3292 3292
rect 3292 3236 3296 3292
rect 3232 3232 3296 3236
rect 3312 3292 3376 3296
rect 3312 3236 3316 3292
rect 3316 3236 3372 3292
rect 3372 3236 3376 3292
rect 3312 3232 3376 3236
rect 3392 3292 3456 3296
rect 3392 3236 3396 3292
rect 3396 3236 3452 3292
rect 3452 3236 3456 3292
rect 3392 3232 3456 3236
rect 7152 3292 7216 3296
rect 7152 3236 7156 3292
rect 7156 3236 7212 3292
rect 7212 3236 7216 3292
rect 7152 3232 7216 3236
rect 7232 3292 7296 3296
rect 7232 3236 7236 3292
rect 7236 3236 7292 3292
rect 7292 3236 7296 3292
rect 7232 3232 7296 3236
rect 7312 3292 7376 3296
rect 7312 3236 7316 3292
rect 7316 3236 7372 3292
rect 7372 3236 7376 3292
rect 7312 3232 7376 3236
rect 7392 3292 7456 3296
rect 7392 3236 7396 3292
rect 7396 3236 7452 3292
rect 7452 3236 7456 3292
rect 7392 3232 7456 3236
rect 1152 2748 1216 2752
rect 1152 2692 1156 2748
rect 1156 2692 1212 2748
rect 1212 2692 1216 2748
rect 1152 2688 1216 2692
rect 1232 2748 1296 2752
rect 1232 2692 1236 2748
rect 1236 2692 1292 2748
rect 1292 2692 1296 2748
rect 1232 2688 1296 2692
rect 1312 2748 1376 2752
rect 1312 2692 1316 2748
rect 1316 2692 1372 2748
rect 1372 2692 1376 2748
rect 1312 2688 1376 2692
rect 1392 2748 1456 2752
rect 1392 2692 1396 2748
rect 1396 2692 1452 2748
rect 1452 2692 1456 2748
rect 1392 2688 1456 2692
rect 5152 2748 5216 2752
rect 5152 2692 5156 2748
rect 5156 2692 5212 2748
rect 5212 2692 5216 2748
rect 5152 2688 5216 2692
rect 5232 2748 5296 2752
rect 5232 2692 5236 2748
rect 5236 2692 5292 2748
rect 5292 2692 5296 2748
rect 5232 2688 5296 2692
rect 5312 2748 5376 2752
rect 5312 2692 5316 2748
rect 5316 2692 5372 2748
rect 5372 2692 5376 2748
rect 5312 2688 5376 2692
rect 5392 2748 5456 2752
rect 5392 2692 5396 2748
rect 5396 2692 5452 2748
rect 5452 2692 5456 2748
rect 5392 2688 5456 2692
rect 3152 2204 3216 2208
rect 3152 2148 3156 2204
rect 3156 2148 3212 2204
rect 3212 2148 3216 2204
rect 3152 2144 3216 2148
rect 3232 2204 3296 2208
rect 3232 2148 3236 2204
rect 3236 2148 3292 2204
rect 3292 2148 3296 2204
rect 3232 2144 3296 2148
rect 3312 2204 3376 2208
rect 3312 2148 3316 2204
rect 3316 2148 3372 2204
rect 3372 2148 3376 2204
rect 3312 2144 3376 2148
rect 3392 2204 3456 2208
rect 3392 2148 3396 2204
rect 3396 2148 3452 2204
rect 3452 2148 3456 2204
rect 3392 2144 3456 2148
rect 7152 2204 7216 2208
rect 7152 2148 7156 2204
rect 7156 2148 7212 2204
rect 7212 2148 7216 2204
rect 7152 2144 7216 2148
rect 7232 2204 7296 2208
rect 7232 2148 7236 2204
rect 7236 2148 7292 2204
rect 7292 2148 7296 2204
rect 7232 2144 7296 2148
rect 7312 2204 7376 2208
rect 7312 2148 7316 2204
rect 7316 2148 7372 2204
rect 7372 2148 7376 2204
rect 7312 2144 7376 2148
rect 7392 2204 7456 2208
rect 7392 2148 7396 2204
rect 7396 2148 7452 2204
rect 7452 2148 7456 2204
rect 7392 2144 7456 2148
rect 1152 1660 1216 1664
rect 1152 1604 1156 1660
rect 1156 1604 1212 1660
rect 1212 1604 1216 1660
rect 1152 1600 1216 1604
rect 1232 1660 1296 1664
rect 1232 1604 1236 1660
rect 1236 1604 1292 1660
rect 1292 1604 1296 1660
rect 1232 1600 1296 1604
rect 1312 1660 1376 1664
rect 1312 1604 1316 1660
rect 1316 1604 1372 1660
rect 1372 1604 1376 1660
rect 1312 1600 1376 1604
rect 1392 1660 1456 1664
rect 1392 1604 1396 1660
rect 1396 1604 1452 1660
rect 1452 1604 1456 1660
rect 1392 1600 1456 1604
rect 5152 1660 5216 1664
rect 5152 1604 5156 1660
rect 5156 1604 5212 1660
rect 5212 1604 5216 1660
rect 5152 1600 5216 1604
rect 5232 1660 5296 1664
rect 5232 1604 5236 1660
rect 5236 1604 5292 1660
rect 5292 1604 5296 1660
rect 5232 1600 5296 1604
rect 5312 1660 5376 1664
rect 5312 1604 5316 1660
rect 5316 1604 5372 1660
rect 5372 1604 5376 1660
rect 5312 1600 5376 1604
rect 5392 1660 5456 1664
rect 5392 1604 5396 1660
rect 5396 1604 5452 1660
rect 5452 1604 5456 1660
rect 5392 1600 5456 1604
rect 3152 1116 3216 1120
rect 3152 1060 3156 1116
rect 3156 1060 3212 1116
rect 3212 1060 3216 1116
rect 3152 1056 3216 1060
rect 3232 1116 3296 1120
rect 3232 1060 3236 1116
rect 3236 1060 3292 1116
rect 3292 1060 3296 1116
rect 3232 1056 3296 1060
rect 3312 1116 3376 1120
rect 3312 1060 3316 1116
rect 3316 1060 3372 1116
rect 3372 1060 3376 1116
rect 3312 1056 3376 1060
rect 3392 1116 3456 1120
rect 3392 1060 3396 1116
rect 3396 1060 3452 1116
rect 3452 1060 3456 1116
rect 3392 1056 3456 1060
rect 7152 1116 7216 1120
rect 7152 1060 7156 1116
rect 7156 1060 7212 1116
rect 7212 1060 7216 1116
rect 7152 1056 7216 1060
rect 7232 1116 7296 1120
rect 7232 1060 7236 1116
rect 7236 1060 7292 1116
rect 7292 1060 7296 1116
rect 7232 1056 7296 1060
rect 7312 1116 7376 1120
rect 7312 1060 7316 1116
rect 7316 1060 7372 1116
rect 7372 1060 7376 1116
rect 7312 1056 7376 1060
rect 7392 1116 7456 1120
rect 7392 1060 7396 1116
rect 7396 1060 7452 1116
rect 7452 1060 7456 1116
rect 7392 1056 7456 1060
<< metal4 >>
rect 1144 7104 1464 7664
rect 1144 7040 1152 7104
rect 1216 7040 1232 7104
rect 1296 7040 1312 7104
rect 1376 7040 1392 7104
rect 1456 7040 1464 7104
rect 1144 6016 1464 7040
rect 1144 5952 1152 6016
rect 1216 5952 1232 6016
rect 1296 5952 1312 6016
rect 1376 5952 1392 6016
rect 1456 5952 1464 6016
rect 1144 4928 1464 5952
rect 1144 4864 1152 4928
rect 1216 4864 1232 4928
rect 1296 4864 1312 4928
rect 1376 4864 1392 4928
rect 1456 4864 1464 4928
rect 1144 3840 1464 4864
rect 1144 3776 1152 3840
rect 1216 3776 1232 3840
rect 1296 3776 1312 3840
rect 1376 3776 1392 3840
rect 1456 3776 1464 3840
rect 1144 2752 1464 3776
rect 1144 2688 1152 2752
rect 1216 2688 1232 2752
rect 1296 2688 1312 2752
rect 1376 2688 1392 2752
rect 1456 2688 1464 2752
rect 1144 1664 1464 2688
rect 1144 1600 1152 1664
rect 1216 1600 1232 1664
rect 1296 1600 1312 1664
rect 1376 1600 1392 1664
rect 1456 1600 1464 1664
rect 1144 1040 1464 1600
rect 3144 7648 3464 7664
rect 3144 7584 3152 7648
rect 3216 7584 3232 7648
rect 3296 7584 3312 7648
rect 3376 7584 3392 7648
rect 3456 7584 3464 7648
rect 3144 6560 3464 7584
rect 3144 6496 3152 6560
rect 3216 6496 3232 6560
rect 3296 6496 3312 6560
rect 3376 6496 3392 6560
rect 3456 6496 3464 6560
rect 3144 5472 3464 6496
rect 3144 5408 3152 5472
rect 3216 5408 3232 5472
rect 3296 5408 3312 5472
rect 3376 5408 3392 5472
rect 3456 5408 3464 5472
rect 3144 4384 3464 5408
rect 3144 4320 3152 4384
rect 3216 4320 3232 4384
rect 3296 4320 3312 4384
rect 3376 4320 3392 4384
rect 3456 4320 3464 4384
rect 3144 3296 3464 4320
rect 3144 3232 3152 3296
rect 3216 3232 3232 3296
rect 3296 3232 3312 3296
rect 3376 3232 3392 3296
rect 3456 3232 3464 3296
rect 3144 2208 3464 3232
rect 3144 2144 3152 2208
rect 3216 2144 3232 2208
rect 3296 2144 3312 2208
rect 3376 2144 3392 2208
rect 3456 2144 3464 2208
rect 3144 1120 3464 2144
rect 3144 1056 3152 1120
rect 3216 1056 3232 1120
rect 3296 1056 3312 1120
rect 3376 1056 3392 1120
rect 3456 1056 3464 1120
rect 3144 1040 3464 1056
rect 5144 7104 5464 7664
rect 5144 7040 5152 7104
rect 5216 7040 5232 7104
rect 5296 7040 5312 7104
rect 5376 7040 5392 7104
rect 5456 7040 5464 7104
rect 5144 6016 5464 7040
rect 5144 5952 5152 6016
rect 5216 5952 5232 6016
rect 5296 5952 5312 6016
rect 5376 5952 5392 6016
rect 5456 5952 5464 6016
rect 5144 4928 5464 5952
rect 5144 4864 5152 4928
rect 5216 4864 5232 4928
rect 5296 4864 5312 4928
rect 5376 4864 5392 4928
rect 5456 4864 5464 4928
rect 5144 3840 5464 4864
rect 5144 3776 5152 3840
rect 5216 3776 5232 3840
rect 5296 3776 5312 3840
rect 5376 3776 5392 3840
rect 5456 3776 5464 3840
rect 5144 2752 5464 3776
rect 5144 2688 5152 2752
rect 5216 2688 5232 2752
rect 5296 2688 5312 2752
rect 5376 2688 5392 2752
rect 5456 2688 5464 2752
rect 5144 1664 5464 2688
rect 5144 1600 5152 1664
rect 5216 1600 5232 1664
rect 5296 1600 5312 1664
rect 5376 1600 5392 1664
rect 5456 1600 5464 1664
rect 5144 1040 5464 1600
rect 7144 7648 7464 7664
rect 7144 7584 7152 7648
rect 7216 7584 7232 7648
rect 7296 7584 7312 7648
rect 7376 7584 7392 7648
rect 7456 7584 7464 7648
rect 7144 6560 7464 7584
rect 7144 6496 7152 6560
rect 7216 6496 7232 6560
rect 7296 6496 7312 6560
rect 7376 6496 7392 6560
rect 7456 6496 7464 6560
rect 7144 5472 7464 6496
rect 7144 5408 7152 5472
rect 7216 5408 7232 5472
rect 7296 5408 7312 5472
rect 7376 5408 7392 5472
rect 7456 5408 7464 5472
rect 7144 4384 7464 5408
rect 7144 4320 7152 4384
rect 7216 4320 7232 4384
rect 7296 4320 7312 4384
rect 7376 4320 7392 4384
rect 7456 4320 7464 4384
rect 7144 3296 7464 4320
rect 7144 3232 7152 3296
rect 7216 3232 7232 3296
rect 7296 3232 7312 3296
rect 7376 3232 7392 3296
rect 7456 3232 7464 3296
rect 7144 2208 7464 3232
rect 7144 2144 7152 2208
rect 7216 2144 7232 2208
rect 7296 2144 7312 2208
rect 7376 2144 7392 2208
rect 7456 2144 7464 2208
rect 7144 1120 7464 2144
rect 7144 1056 7152 1120
rect 7216 1056 7232 1120
rect 7296 1056 7312 1120
rect 7376 1056 7392 1120
rect 7456 1056 7464 1120
rect 7144 1040 7464 1056
use sky130_fd_sc_hd__fill_2  FILLER_0_3 swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 1380 0 1 1088
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8 swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 1840 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20 swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 2944 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24 swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 3312 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1673029049
transform 1 0 3772 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34 swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 4232 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42 swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 4968 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48
timestamp 1673029049
transform 1 0 5520 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57
timestamp 1673029049
transform 1 0 6348 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68
timestamp 1673029049
transform 1 0 7360 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1673029049
transform 1 0 1380 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_8
timestamp 1673029049
transform 1 0 1840 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_38
timestamp 1673029049
transform 1 0 4600 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_46
timestamp 1673029049
transform 1 0 5336 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_53
timestamp 1673029049
transform 1 0 5980 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1673029049
transform 1 0 6348 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_62
timestamp 1673029049
transform 1 0 6808 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3 swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 1380 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_12
timestamp 1673029049
transform 1 0 2208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_19
timestamp 1673029049
transform 1 0 2852 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1673029049
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1673029049
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_41
timestamp 1673029049
transform 1 0 4876 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_47
timestamp 1673029049
transform 1 0 5428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_54
timestamp 1673029049
transform 1 0 6072 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_62
timestamp 1673029049
transform 1 0 6808 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_68
timestamp 1673029049
transform 1 0 7360 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3
timestamp 1673029049
transform 1 0 1380 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_35
timestamp 1673029049
transform 1 0 4324 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_47
timestamp 1673029049
transform 1 0 5428 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1673029049
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_57
timestamp 1673029049
transform 1 0 6348 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_68
timestamp 1673029049
transform 1 0 7360 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1673029049
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_8
timestamp 1673029049
transform 1 0 1840 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_20
timestamp 1673029049
transform 1 0 2944 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1673029049
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1673029049
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_53
timestamp 1673029049
transform 1 0 5980 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_57
timestamp 1673029049
transform 1 0 6348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_61
timestamp 1673029049
transform 1 0 6716 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_68
timestamp 1673029049
transform 1 0 7360 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1673029049
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_14
timestamp 1673029049
transform 1 0 2392 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_21
timestamp 1673029049
transform 1 0 3036 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_33
timestamp 1673029049
transform 1 0 4140 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_45
timestamp 1673029049
transform 1 0 5244 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_53
timestamp 1673029049
transform 1 0 5980 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_57
timestamp 1673029049
transform 1 0 6348 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_68
timestamp 1673029049
transform 1 0 7360 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_3
timestamp 1673029049
transform 1 0 1380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_10
timestamp 1673029049
transform 1 0 2024 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_17
timestamp 1673029049
transform 1 0 2668 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_25
timestamp 1673029049
transform 1 0 3404 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1673029049
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1673029049
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_53
timestamp 1673029049
transform 1 0 5980 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_57
timestamp 1673029049
transform 1 0 6348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_61
timestamp 1673029049
transform 1 0 6716 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_68
timestamp 1673029049
transform 1 0 7360 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1673029049
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1673029049
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1673029049
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1673029049
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1673029049
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1673029049
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_57
timestamp 1673029049
transform 1 0 6348 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_62
timestamp 1673029049
transform 1 0 6808 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1673029049
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_8
timestamp 1673029049
transform 1 0 1840 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_20
timestamp 1673029049
transform 1 0 2944 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1673029049
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1673029049
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_53
timestamp 1673029049
transform 1 0 5980 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_8_68
timestamp 1673029049
transform 1 0 7360 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1673029049
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_10
timestamp 1673029049
transform 1 0 2024 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_17
timestamp 1673029049
transform 1 0 2668 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_24
timestamp 1673029049
transform 1 0 3312 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_36
timestamp 1673029049
transform 1 0 4416 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_48
timestamp 1673029049
transform 1 0 5520 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_9_57
timestamp 1673029049
transform 1 0 6348 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_68
timestamp 1673029049
transform 1 0 7360 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1673029049
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_14
timestamp 1673029049
transform 1 0 2392 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_10_25
timestamp 1673029049
transform 1 0 3404 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1673029049
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_41
timestamp 1673029049
transform 1 0 4876 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_49
timestamp 1673029049
transform 1 0 5612 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_53
timestamp 1673029049
transform 1 0 5980 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_60
timestamp 1673029049
transform 1 0 6624 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_67
timestamp 1673029049
transform 1 0 7268 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_3
timestamp 1673029049
transform 1 0 1380 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_11_14
timestamp 1673029049
transform 1 0 2392 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_26
timestamp 1673029049
transform 1 0 3496 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_29
timestamp 1673029049
transform 1 0 3772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_41
timestamp 1673029049
transform 1 0 4876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_53
timestamp 1673029049
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_57
timestamp 1673029049
transform 1 0 6348 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_68
timestamp 1673029049
transform 1 0 7360 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1673029049
transform 1 0 1104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1673029049
transform -1 0 7820 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1673029049
transform 1 0 1104 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1673029049
transform -1 0 7820 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1673029049
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1673029049
transform -1 0 7820 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1673029049
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1673029049
transform -1 0 7820 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1673029049
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1673029049
transform -1 0 7820 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1673029049
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1673029049
transform -1 0 7820 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1673029049
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1673029049
transform -1 0 7820 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1673029049
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1673029049
transform -1 0 7820 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1673029049
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1673029049
transform -1 0 7820 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1673029049
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1673029049
transform -1 0 7820 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1673029049
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1673029049
transform -1 0 7820 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1673029049
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1673029049
transform -1 0 7820 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_24 swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 3680 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_25
timestamp 1673029049
transform 1 0 6256 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_26
timestamp 1673029049
transform 1 0 6256 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_27
timestamp 1673029049
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28
timestamp 1673029049
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1673029049
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1673029049
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 1673029049
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 1673029049
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 1673029049
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 1673029049
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1673029049
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1673029049
transform 1 0 3680 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1673029049
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  spare_logic_biginv swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 1564 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[0\] swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 6716 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[1\]
timestamp 1673029049
transform 1 0 7084 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[2\]
timestamp 1673029049
transform 1 0 5704 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[3\]
timestamp 1673029049
transform -1 0 7268 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[4\]
timestamp 1673029049
transform -1 0 2392 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[5\]
timestamp 1673029049
transform 1 0 3036 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[6\]
timestamp 1673029049
transform -1 0 6808 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[7\]
timestamp 1673029049
transform -1 0 3036 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[8\]
timestamp 1673029049
transform -1 0 6072 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[9\]
timestamp 1673029049
transform 1 0 7084 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[10\]
timestamp 1673029049
transform -1 0 2668 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[11\]
timestamp 1673029049
transform 1 0 6440 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[12\]
timestamp 1673029049
transform -1 0 1840 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[13\]
timestamp 1673029049
transform -1 0 7360 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[14\]
timestamp 1673029049
transform 1 0 1748 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[15\]
timestamp 1673029049
transform -1 0 6808 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[16\]
timestamp 1673029049
transform -1 0 1840 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[17\]
timestamp 1673029049
transform -1 0 7360 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[18\]
timestamp 1673029049
transform -1 0 2668 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[19\]
timestamp 1673029049
transform -1 0 1840 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[20\]
timestamp 1673029049
transform -1 0 5520 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[21\]
timestamp 1673029049
transform -1 0 2208 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[22\]
timestamp 1673029049
transform -1 0 1840 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[23\]
timestamp 1673029049
transform -1 0 2852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[24\]
timestamp 1673029049
transform 1 0 3036 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[25\]
timestamp 1673029049
transform -1 0 5428 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[26\]
timestamp 1673029049
transform -1 0 4232 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__dfbbp_1  spare_logic_flop\[0\] swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 1932 0 -1 3264
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbp_1  spare_logic_flop\[1\]
timestamp 1673029049
transform 1 0 2208 0 -1 2176
box -38 -48 2430 592
use sky130_fd_sc_hd__inv_2  spare_logic_inv\[0\] swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 7084 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  spare_logic_inv\[1\]
timestamp 1673029049
transform -1 0 7360 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  spare_logic_inv\[2\]
timestamp 1673029049
transform 1 0 7084 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  spare_logic_inv\[3\]
timestamp 1673029049
transform -1 0 6624 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  spare_logic_mux\[0\] swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 7360 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  spare_logic_mux\[1\]
timestamp 1673029049
transform -1 0 2392 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  spare_logic_nand\[0\] swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 2944 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  spare_logic_nand\[1\]
timestamp 1673029049
transform 1 0 5520 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  spare_logic_nor\[0\] swift/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 7360 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  spare_logic_nor\[1\]
timestamp 1673029049
transform -1 0 2024 0 -1 6528
box -38 -48 498 592
<< labels >>
flabel metal3 s 0 2048 800 2168 0 FreeSans 480 0 0 0 spare_xfq[0]
port 0 nsew signal tristate
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 spare_xfq[1]
port 1 nsew signal tristate
flabel metal2 s 4526 8200 4582 9000 0 FreeSans 224 90 0 0 spare_xfqn[0]
port 2 nsew signal tristate
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 spare_xfqn[1]
port 3 nsew signal tristate
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 spare_xi[0]
port 4 nsew signal tristate
flabel metal3 s 8200 8 9000 128 0 FreeSans 480 0 0 0 spare_xi[1]
port 5 nsew signal tristate
flabel metal3 s 8200 5448 9000 5568 0 FreeSans 480 0 0 0 spare_xi[2]
port 6 nsew signal tristate
flabel metal2 s 18 8200 74 9000 0 FreeSans 224 90 0 0 spare_xi[3]
port 7 nsew signal tristate
flabel metal3 s 0 7488 800 7608 0 FreeSans 480 0 0 0 spare_xib
port 8 nsew signal tristate
flabel metal2 s 7102 8200 7158 9000 0 FreeSans 224 90 0 0 spare_xmx[0]
port 9 nsew signal tristate
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 spare_xmx[1]
port 10 nsew signal tristate
flabel metal3 s 8200 6808 9000 6928 0 FreeSans 480 0 0 0 spare_xna[0]
port 11 nsew signal tristate
flabel metal3 s 8200 1368 9000 1488 0 FreeSans 480 0 0 0 spare_xna[1]
port 12 nsew signal tristate
flabel metal2 s 1306 0 1362 800 0 FreeSans 224 90 0 0 spare_xno[0]
port 13 nsew signal tristate
flabel metal3 s 0 6128 800 6248 0 FreeSans 480 0 0 0 spare_xno[1]
port 14 nsew signal tristate
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 spare_xz[0]
port 15 nsew signal tristate
flabel metal2 s 5170 8200 5226 9000 0 FreeSans 224 90 0 0 spare_xz[10]
port 16 nsew signal tristate
flabel metal2 s 7746 8200 7802 9000 0 FreeSans 224 90 0 0 spare_xz[11]
port 17 nsew signal tristate
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 spare_xz[12]
port 18 nsew signal tristate
flabel metal3 s 8200 7488 9000 7608 0 FreeSans 480 0 0 0 spare_xz[13]
port 19 nsew signal tristate
flabel metal2 s 1950 8200 2006 9000 0 FreeSans 224 90 0 0 spare_xz[14]
port 20 nsew signal tristate
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 spare_xz[15]
port 21 nsew signal tristate
flabel metal3 s 0 1368 800 1488 0 FreeSans 480 0 0 0 spare_xz[16]
port 22 nsew signal tristate
flabel metal3 s 8200 4768 9000 4888 0 FreeSans 480 0 0 0 spare_xz[17]
port 23 nsew signal tristate
flabel metal2 s 662 8200 718 9000 0 FreeSans 224 90 0 0 spare_xz[18]
port 24 nsew signal tristate
flabel metal3 s 0 688 800 808 0 FreeSans 480 0 0 0 spare_xz[19]
port 25 nsew signal tristate
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 spare_xz[1]
port 26 nsew signal tristate
flabel metal2 s 5814 8200 5870 9000 0 FreeSans 224 90 0 0 spare_xz[20]
port 27 nsew signal tristate
flabel metal3 s 8200 2048 9000 2168 0 FreeSans 480 0 0 0 spare_xz[21]
port 28 nsew signal tristate
flabel metal2 s 662 0 718 800 0 FreeSans 224 90 0 0 spare_xz[22]
port 29 nsew signal tristate
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 spare_xz[23]
port 30 nsew signal tristate
flabel metal2 s 3238 0 3294 800 0 FreeSans 224 90 0 0 spare_xz[24]
port 31 nsew signal tristate
flabel metal3 s 8200 2728 9000 2848 0 FreeSans 480 0 0 0 spare_xz[25]
port 32 nsew signal tristate
flabel metal2 s 3882 0 3938 800 0 FreeSans 224 90 0 0 spare_xz[26]
port 33 nsew signal tristate
flabel metal3 s 8200 8168 9000 8288 0 FreeSans 480 0 0 0 spare_xz[2]
port 34 nsew signal tristate
flabel metal2 s 8390 8200 8446 9000 0 FreeSans 224 90 0 0 spare_xz[3]
port 35 nsew signal tristate
flabel metal2 s 2594 8200 2650 9000 0 FreeSans 224 90 0 0 spare_xz[4]
port 36 nsew signal tristate
flabel metal2 s 3238 8200 3294 9000 0 FreeSans 224 90 0 0 spare_xz[5]
port 37 nsew signal tristate
flabel metal2 s 5814 0 5870 800 0 FreeSans 224 90 0 0 spare_xz[6]
port 38 nsew signal tristate
flabel metal3 s 0 3408 800 3528 0 FreeSans 480 0 0 0 spare_xz[7]
port 39 nsew signal tristate
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 spare_xz[8]
port 40 nsew signal tristate
flabel metal3 s 8200 4088 9000 4208 0 FreeSans 480 0 0 0 spare_xz[9]
port 41 nsew signal tristate
flabel metal4 s 1144 1040 1464 7664 0 FreeSans 1920 90 0 0 vccd
port 42 nsew power bidirectional
flabel metal4 s 5144 1040 5464 7664 0 FreeSans 1920 90 0 0 vccd
port 42 nsew power bidirectional
flabel metal4 s 3144 1040 3464 7664 0 FreeSans 1920 90 0 0 vssd
port 43 nsew ground bidirectional
flabel metal4 s 7144 1040 7464 7664 0 FreeSans 1920 90 0 0 vssd
port 43 nsew ground bidirectional
rlabel metal1 4462 7072 4462 7072 0 vccd
rlabel metal1 4462 7616 4462 7616 0 vssd
rlabel metal3 1395 2108 1395 2108 0 spare_xfq[0]
rlabel metal2 6486 1248 6486 1248 0 spare_xfq[1]
rlabel metal1 4278 3162 4278 3162 0 spare_xfqn[0]
rlabel metal1 4324 2074 4324 2074 0 spare_xfqn[1]
rlabel metal2 8418 976 8418 976 0 spare_xi[0]
rlabel metal1 7544 2822 7544 2822 0 spare_xi[1]
rlabel metal1 7406 6086 7406 6086 0 spare_xi[2]
rlabel metal1 3266 6970 3266 6970 0 spare_xi[3]
rlabel metal3 1142 7548 1142 7548 0 spare_xib
rlabel metal1 7130 5882 7130 5882 0 spare_xmx[0]
rlabel metal2 5198 1095 5198 1095 0 spare_xmx[1]
rlabel metal1 3818 6834 3818 6834 0 spare_xna[0]
rlabel metal2 5934 1649 5934 1649 0 spare_xna[1]
rlabel metal2 1334 823 1334 823 0 spare_xno[0]
rlabel metal3 1142 6188 1142 6188 0 spare_xno[1]
rlabel metal2 6486 3944 6486 3944 0 spare_xz[0]
rlabel metal1 3634 6222 3634 6222 0 spare_xz[10]
rlabel metal2 7038 4420 7038 4420 0 spare_xz[11]
rlabel metal2 1610 5389 1610 5389 0 spare_xz[12]
rlabel metal2 6854 6562 6854 6562 0 spare_xz[13]
rlabel metal2 1978 4488 1978 4488 0 spare_xz[14]
rlabel metal2 6578 4318 6578 4318 0 spare_xz[15]
rlabel metal2 1610 2465 1610 2465 0 spare_xz[16]
rlabel metal2 6854 5202 6854 5202 0 spare_xz[17]
rlabel metal1 1610 4114 1610 4114 0 spare_xz[18]
rlabel metal1 1564 1734 1564 1734 0 spare_xz[19]
rlabel metal1 7544 2414 7544 2414 0 spare_xz[1]
rlabel metal1 5658 1530 5658 1530 0 spare_xz[20]
rlabel metal1 3128 2482 3128 2482 0 spare_xz[21]
rlabel metal1 1150 1394 1150 1394 0 spare_xz[22]
rlabel metal2 2622 1588 2622 1588 0 spare_xz[23]
rlabel metal1 3174 1394 3174 1394 0 spare_xz[24]
rlabel metal1 5152 2618 5152 2618 0 spare_xz[25]
rlabel metal1 3956 1394 3956 1394 0 spare_xz[26]
rlabel metal1 6348 6834 6348 6834 0 spare_xz[2]
rlabel metal1 7498 6766 7498 6766 0 spare_xz[3]
rlabel metal2 2346 8228 2346 8228 0 spare_xz[4]
rlabel metal1 3128 6766 3128 6766 0 spare_xz[5]
rlabel metal2 5842 1350 5842 1350 0 spare_xz[6]
rlabel metal2 2806 3689 2806 3689 0 spare_xz[7]
rlabel metal1 5796 2618 5796 2618 0 spare_xz[8]
rlabel via2 7314 4131 7314 4131 0 spare_xz[9]
<< properties >>
string FIXED_BBOX 0 0 9000 9000
<< end >>
