magic
tech sky130A
magscale 1 2
timestamp 1637447660
<< error_p >>
rect 30970 218031 31724 218032
rect 30970 216955 30971 218031
rect 31723 216955 31724 218031
rect 30970 216954 31724 216955
rect 37508 216463 38270 216464
rect 37508 215381 37509 216463
rect 38269 215381 38270 216463
rect 37508 215380 38270 215381
<< metal3 >>
rect 6032 221346 43870 221382
rect 6032 221338 42656 221346
rect 6032 220224 6162 221338
rect 6862 220248 42656 221338
rect 43738 220248 43870 221346
rect 6862 220224 43870 220248
rect 6032 220182 43870 220224
rect 7246 219742 42226 219782
rect 7246 218628 7360 219742
rect 8060 219728 42226 219742
rect 8060 218630 41062 219728
rect 42144 218630 42226 219728
rect 8060 218628 42226 218630
rect 7246 218582 42226 218628
rect 17838 218068 31812 218100
rect 17838 216936 17896 218068
rect 18646 218032 31812 218068
rect 18646 216954 30970 218032
rect 31724 216954 31812 218032
rect 18646 216936 31812 216954
rect 17838 216900 31812 216936
rect 19032 216470 38402 216500
rect 19032 215338 19100 216470
rect 19850 216464 38402 216470
rect 19850 215380 37508 216464
rect 38270 215380 38402 216464
rect 19850 215338 38402 215380
rect 19032 215300 38402 215338
<< via3 >>
rect 6162 220224 6862 221338
rect 42656 220248 43738 221346
rect 7360 218628 8060 219742
rect 41062 218630 42144 219728
rect 17896 216936 18646 218068
rect 30970 216954 31724 218032
rect 19100 215338 19850 216470
rect 37508 215380 38270 216464
<< metal4 >>
rect 6116 221338 6916 221470
rect 6116 220224 6162 221338
rect 6862 220224 6916 221338
rect 6116 211888 6916 220224
rect 42594 221346 43800 221388
rect 42594 220248 42656 221346
rect 43738 220248 43800 221346
rect 42594 220174 43800 220248
rect 6116 211604 6134 211888
rect 6900 211604 6916 211888
rect 6116 208516 6916 211604
rect 6116 208236 6128 208516
rect 6902 208236 6916 208516
rect 6116 205138 6916 208236
rect 7316 219742 8116 219842
rect 7316 218628 7360 219742
rect 8060 218628 8116 219742
rect 7316 213578 8116 218628
rect 40990 219728 42196 219788
rect 40990 218630 41062 219728
rect 42144 218630 42196 219728
rect 40990 218574 42196 218630
rect 7316 213294 7332 213578
rect 8098 213294 8116 213578
rect 7316 210202 8116 213294
rect 7316 209918 7330 210202
rect 8096 209918 8116 210202
rect 7316 206826 8116 209918
rect 7316 206528 7326 206826
rect 8100 206528 8116 206826
rect 7316 206476 8116 206528
rect 17880 218068 18680 218110
rect 17880 216936 17896 218068
rect 18646 217338 18680 218068
rect 18656 217056 18680 217338
rect 18646 216936 18680 217056
rect 17880 212534 18680 216936
rect 17880 212246 17896 212534
rect 18668 212246 18680 212534
rect 17880 209152 18680 212246
rect 17880 208864 17890 209152
rect 18662 208864 18680 209152
rect 17880 205770 18680 208864
rect 17880 205482 17892 205770
rect 18664 205482 18680 205770
rect 17880 205422 18680 205482
rect 19080 216634 19880 216732
rect 19080 215338 19100 216634
rect 19856 216352 19880 216634
rect 19850 215338 19880 216352
rect 19080 210844 19880 215338
rect 19080 210556 19092 210844
rect 19864 210556 19880 210844
rect 19080 207464 19880 210556
rect 19080 207176 19096 207464
rect 19868 207176 19880 207464
rect 6116 204840 6132 205138
rect 6906 204840 6916 205138
rect 6116 204746 6916 204840
rect 19080 204084 19880 207176
rect 19080 203796 19096 204084
rect 19868 203796 19880 204084
rect 19080 203748 19880 203796
<< via4 >>
rect 6134 211604 6900 211888
rect 6128 208236 6902 208516
rect 7332 213294 8098 213578
rect 7330 209918 8096 210202
rect 7326 206528 8100 206826
rect 17900 217056 18646 217338
rect 18646 217056 18656 217338
rect 17896 212246 18668 212534
rect 17890 208864 18662 209152
rect 17892 205482 18664 205770
rect 19100 216470 19856 216634
rect 19100 216352 19850 216470
rect 19850 216352 19856 216470
rect 19092 210556 19864 210844
rect 19096 207176 19868 207464
rect 6132 204840 6906 205138
rect 19096 203796 19868 204084
<< metal5 >>
rect 17806 217350 18682 217372
rect 14320 217338 18682 217350
rect 14320 217056 17900 217338
rect 18656 217056 18682 217338
rect 14320 217030 18682 217056
rect 17806 217026 18682 217030
rect 19058 216650 19934 216670
rect 14320 216634 19934 216650
rect 14320 216352 19100 216634
rect 19856 216352 19934 216634
rect 14320 216330 19934 216352
rect 19058 216324 19934 216330
rect 7258 213598 8134 213614
rect 7258 213578 8592 213598
rect 7258 213294 7332 213578
rect 8098 213294 8592 213578
rect 7258 213278 8592 213294
rect 7258 213268 8134 213278
rect 17850 212550 18726 212568
rect 17434 212534 18726 212550
rect 17434 212246 17896 212534
rect 18668 212246 18726 212534
rect 17434 212230 18726 212246
rect 17850 212222 18726 212230
rect 6054 211908 6930 211912
rect 6054 211888 8592 211908
rect 6054 211604 6134 211888
rect 6900 211604 8592 211888
rect 6054 211588 8592 211604
rect 6054 211566 6930 211588
rect 19032 210860 19908 210870
rect 17434 210844 19910 210860
rect 17434 210556 19092 210844
rect 19864 210556 19910 210844
rect 17434 210540 19910 210556
rect 19032 210524 19908 210540
rect 7264 210218 8140 210226
rect 7264 210202 8592 210218
rect 7264 209918 7330 210202
rect 8096 209918 8592 210202
rect 7264 209898 8592 209918
rect 7264 209880 8140 209898
rect 17822 209170 18698 209180
rect 17434 209152 18698 209170
rect 17434 208864 17890 209152
rect 18662 208864 18698 209152
rect 17434 208850 18698 208864
rect 17822 208828 18698 208850
rect 6050 208528 6926 208548
rect 6050 208516 8592 208528
rect 6050 208236 6128 208516
rect 6902 208236 8592 208516
rect 6050 208208 8592 208236
rect 6050 208202 6926 208208
rect 19034 207480 19910 207494
rect 17434 207464 19910 207480
rect 17434 207176 19096 207464
rect 19868 207176 19910 207464
rect 17434 207160 19910 207176
rect 19034 207148 19910 207160
rect 7300 206838 8132 206852
rect 7300 206826 8624 206838
rect 7300 206528 7326 206826
rect 8100 206528 8624 206826
rect 7300 206518 8624 206528
rect 7300 206502 8132 206518
rect 17838 205790 18714 205802
rect 17434 205770 18714 205790
rect 17434 205482 17892 205770
rect 18664 205482 18714 205770
rect 17434 205470 18714 205482
rect 17838 205456 18714 205470
rect 6102 205148 6934 205162
rect 6102 205138 8624 205148
rect 6102 204840 6132 205138
rect 6906 204840 8624 205138
rect 6102 204828 8624 204840
rect 6102 204812 6934 204828
rect 19036 204100 19912 204114
rect 17434 204084 19912 204100
rect 17434 203796 19096 204084
rect 19868 203796 19912 204084
rect 17434 203780 19912 203796
rect 19036 203768 19912 203780
<< end >>
