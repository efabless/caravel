magic
tech sky130A
magscale 1 2
timestamp 1608587524
<< obsli1 >>
rect 480 797 3456 3273
<< obsm1 >>
rect 480 763 3456 3307
<< metal2 >>
rect 3284 2600 3340 3800
rect 596 -400 652 800
<< obsm2 >>
rect 598 2544 3228 3307
rect 598 856 3326 2544
rect 708 763 3326 856
<< obsm3 >>
rect 790 781 2270 3289
<< metal4 >>
rect 790 763 970 3307
rect 1670 814 1850 3256
rect 2090 763 2270 3307
rect 2970 814 3150 3256
<< labels >>
rlabel metal2 s 3284 2600 3340 3800 6 A
port 1 nsew signal input
rlabel metal2 s 596 -400 652 800 6 X
port 2 nsew signal output
rlabel metal4 s 790 763 970 3307 6 VPWR
port 3 nsew power bidirectional
rlabel metal4 s 2090 763 2270 3307 6 VGND
port 4 nsew ground bidirectional
rlabel metal4 s 1670 814 1850 3256 6 LVPWR
port 5 nsew power bidirectional
rlabel metal4 s 2970 814 3150 3256 6 LVGND
port 6 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 4000 3400
string LEFview TRUE
string GDS_FILE ../gds/xres_buf.gds
string GDS_END 48842
string GDS_START 40962
<< end >>
