magic
tech sky130A
magscale 1 2
timestamp 1636122974
<< locali >>
rect 2237 11543 2271 12257
rect 2421 11543 2455 12189
rect 6101 11747 6135 11917
<< viali >>
rect 2237 12257 2271 12291
rect 2237 11509 2271 11543
rect 2421 12189 2455 12223
rect 6101 11917 6135 11951
rect 6101 11713 6135 11747
rect 2421 11509 2455 11543
rect 1409 11305 1443 11339
rect 2053 11305 2087 11339
rect 2329 11305 2363 11339
rect 3157 11305 3191 11339
rect 3433 11305 3467 11339
rect 5641 11305 5675 11339
rect 6009 11305 6043 11339
rect 6285 11305 6319 11339
rect 6653 11305 6687 11339
rect 8033 11305 8067 11339
rect 2605 11237 2639 11271
rect 4077 11237 4111 11271
rect 4353 11237 4387 11271
rect 4537 11237 4571 11271
rect 5273 11237 5307 11271
rect 5549 11237 5583 11271
rect 7573 11237 7607 11271
rect 9045 11237 9079 11271
rect 1225 11101 1259 11135
rect 1501 11101 1535 11135
rect 1869 11101 1903 11135
rect 2145 11101 2179 11135
rect 2421 11101 2455 11135
rect 2697 11101 2731 11135
rect 2973 11101 3007 11135
rect 3249 11077 3283 11111
rect 3801 11101 3835 11135
rect 4261 11101 4295 11135
rect 4721 11101 4755 11135
rect 4997 11101 5031 11135
rect 5089 11101 5123 11135
rect 5365 11101 5399 11135
rect 5825 11101 5859 11135
rect 6745 11101 6779 11135
rect 6837 11101 6871 11135
rect 7113 11101 7147 11135
rect 7389 11101 7423 11135
rect 8125 11101 8159 11135
rect 8309 11101 8343 11135
rect 8861 11101 8895 11135
rect 9229 11101 9263 11135
rect 1685 10965 1719 10999
rect 2881 10965 2915 10999
rect 3709 10965 3743 10999
rect 3985 10965 4019 10999
rect 4813 10965 4847 10999
rect 7021 10965 7055 10999
rect 7297 10965 7331 10999
rect 7665 10965 7699 10999
rect 8493 10965 8527 10999
rect 9413 10965 9447 10999
rect 1409 10761 1443 10795
rect 4353 10761 4387 10795
rect 8953 10761 8987 10795
rect 8585 10693 8619 10727
rect 1225 10625 1259 10659
rect 1501 10625 1535 10659
rect 1777 10625 1811 10659
rect 2053 10625 2087 10659
rect 2329 10625 2363 10659
rect 2605 10625 2639 10659
rect 2881 10625 2915 10659
rect 3433 10625 3467 10659
rect 3617 10625 3651 10659
rect 3893 10625 3927 10659
rect 4445 10625 4479 10659
rect 4629 10625 4663 10659
rect 5089 10625 5123 10659
rect 5365 10625 5399 10659
rect 5641 10625 5675 10659
rect 5825 10625 5859 10659
rect 6009 10625 6043 10659
rect 6193 10625 6227 10659
rect 8033 10625 8067 10659
rect 8769 10625 8803 10659
rect 9229 10625 9263 10659
rect 3341 10557 3375 10591
rect 6561 10557 6595 10591
rect 1685 10489 1719 10523
rect 4813 10489 4847 10523
rect 9045 10489 9079 10523
rect 1961 10421 1995 10455
rect 2237 10421 2271 10455
rect 2513 10421 2547 10455
rect 2789 10421 2823 10455
rect 3157 10421 3191 10455
rect 3801 10421 3835 10455
rect 4077 10421 4111 10455
rect 4905 10421 4939 10455
rect 5273 10421 5307 10455
rect 5549 10421 5583 10455
rect 8493 10421 8527 10455
rect 9413 10421 9447 10455
rect 1317 10217 1351 10251
rect 1593 10217 1627 10251
rect 7585 10217 7619 10251
rect 7941 10217 7975 10251
rect 8217 10217 8251 10251
rect 6009 10149 6043 10183
rect 9045 10149 9079 10183
rect 3433 10081 3467 10115
rect 1409 10013 1443 10047
rect 3709 10013 3743 10047
rect 4077 10013 4111 10047
rect 5549 10013 5583 10047
rect 7849 10013 7883 10047
rect 8401 10013 8435 10047
rect 8861 10013 8895 10047
rect 9505 10013 9539 10047
rect 3157 9945 3191 9979
rect 1685 9877 1719 9911
rect 6101 9877 6135 9911
rect 8585 9877 8619 9911
rect 9321 9877 9355 9911
rect 1869 9673 1903 9707
rect 1317 9605 1351 9639
rect 6193 9605 6227 9639
rect 1409 9537 1443 9571
rect 1693 9541 1727 9575
rect 1961 9537 1995 9571
rect 2237 9537 2271 9571
rect 2697 9521 2731 9555
rect 3157 9537 3191 9571
rect 4629 9537 4663 9571
rect 5365 9537 5399 9571
rect 5641 9537 5675 9571
rect 6009 9537 6043 9571
rect 6837 9537 6871 9571
rect 6929 9537 6963 9571
rect 7205 9537 7239 9571
rect 9045 9537 9079 9571
rect 2789 9469 2823 9503
rect 7573 9469 7607 9503
rect 2145 9401 2179 9435
rect 2421 9401 2455 9435
rect 5181 9401 5215 9435
rect 5457 9401 5491 9435
rect 5825 9401 5859 9435
rect 7021 9401 7055 9435
rect 1593 9333 1627 9367
rect 2513 9333 2547 9367
rect 5089 9333 5123 9367
rect 9505 9333 9539 9367
rect 1225 9129 1259 9163
rect 1869 9129 1903 9163
rect 3433 9129 3467 9163
rect 3801 9129 3835 9163
rect 4629 9129 4663 9163
rect 9137 9129 9171 9163
rect 1593 9061 1627 9095
rect 4537 9061 4571 9095
rect 4077 8993 4111 9027
rect 5365 8993 5399 9027
rect 1409 8925 1443 8959
rect 1685 8925 1719 8959
rect 1961 8925 1995 8959
rect 2145 8925 2179 8959
rect 2421 8925 2455 8959
rect 2697 8925 2731 8959
rect 2973 8925 3007 8959
rect 3249 8925 3283 8959
rect 3617 8925 3651 8959
rect 4813 8925 4847 8959
rect 5273 8925 5307 8959
rect 8585 8925 8619 8959
rect 9229 8925 9263 8959
rect 4169 8857 4203 8891
rect 4353 8857 4387 8891
rect 5641 8857 5675 8891
rect 7665 8857 7699 8891
rect 8769 8857 8803 8891
rect 8953 8857 8987 8891
rect 2329 8789 2363 8823
rect 2605 8789 2639 8823
rect 2881 8789 2915 8823
rect 3157 8789 3191 8823
rect 5089 8789 5123 8823
rect 7113 8789 7147 8823
rect 9413 8789 9447 8823
rect 1225 8585 1259 8619
rect 1409 8585 1443 8619
rect 9505 8585 9539 8619
rect 2605 8517 2639 8551
rect 6193 8517 6227 8551
rect 6745 8517 6779 8551
rect 7113 8517 7147 8551
rect 1777 8449 1811 8483
rect 2053 8449 2087 8483
rect 4169 8449 4203 8483
rect 6377 8449 6411 8483
rect 6929 8449 6963 8483
rect 9045 8449 9079 8483
rect 1685 8381 1719 8415
rect 2329 8381 2363 8415
rect 4077 8381 4111 8415
rect 4445 8381 4479 8415
rect 7205 8381 7239 8415
rect 7573 8381 7607 8415
rect 1961 8313 1995 8347
rect 5917 8313 5951 8347
rect 2237 8245 2271 8279
rect 6561 8245 6595 8279
rect 3985 8041 4019 8075
rect 8769 8041 8803 8075
rect 1593 7973 1627 8007
rect 3433 7905 3467 7939
rect 5181 7905 5215 7939
rect 5549 7905 5583 7939
rect 7481 7905 7515 7939
rect 1409 7837 1443 7871
rect 3709 7837 3743 7871
rect 4261 7837 4295 7871
rect 4537 7837 4571 7871
rect 7021 7837 7055 7871
rect 8217 7837 8251 7871
rect 8585 7837 8619 7871
rect 8953 7837 8987 7871
rect 9045 7837 9079 7871
rect 9229 7837 9263 7871
rect 1317 7769 1351 7803
rect 3157 7769 3191 7803
rect 7573 7769 7607 7803
rect 7757 7769 7791 7803
rect 1685 7701 1719 7735
rect 4169 7701 4203 7735
rect 7941 7701 7975 7735
rect 8033 7701 8067 7735
rect 8401 7701 8435 7735
rect 9413 7701 9447 7735
rect 1317 7497 1351 7531
rect 1869 7497 1903 7531
rect 2329 7497 2363 7531
rect 4905 7497 4939 7531
rect 8217 7497 8251 7531
rect 9045 7497 9079 7531
rect 9413 7497 9447 7531
rect 2421 7429 2455 7463
rect 1409 7361 1443 7395
rect 1685 7361 1719 7395
rect 1961 7361 1995 7395
rect 2605 7361 2639 7395
rect 2973 7361 3007 7395
rect 4445 7361 4479 7395
rect 5917 7361 5951 7395
rect 6193 7361 6227 7395
rect 6469 7361 6503 7395
rect 8309 7361 8343 7395
rect 5641 7293 5675 7327
rect 6745 7293 6779 7327
rect 8769 7293 8803 7327
rect 8953 7293 8987 7327
rect 1593 7225 1627 7259
rect 2145 7157 2179 7191
rect 6377 7157 6411 7191
rect 8493 7157 8527 7191
rect 1225 6953 1259 6987
rect 6377 6953 6411 6987
rect 8321 6953 8355 6987
rect 8769 6953 8803 6987
rect 1685 6817 1719 6851
rect 3617 6817 3651 6851
rect 8585 6817 8619 6851
rect 9321 6817 9355 6851
rect 1409 6749 1443 6783
rect 3985 6749 4019 6783
rect 5457 6749 5491 6783
rect 6193 6749 6227 6783
rect 6285 6749 6319 6783
rect 1961 6681 1995 6715
rect 1593 6613 1627 6647
rect 3433 6613 3467 6647
rect 5917 6613 5951 6647
rect 6009 6613 6043 6647
rect 6745 6613 6779 6647
rect 6837 6613 6871 6647
rect 9137 6613 9171 6647
rect 9229 6613 9263 6647
rect 1777 6409 1811 6443
rect 4721 6409 4755 6443
rect 1961 6341 1995 6375
rect 2697 6341 2731 6375
rect 6009 6341 6043 6375
rect 2421 6273 2455 6307
rect 6285 6273 6319 6307
rect 8677 6273 8711 6307
rect 9229 6273 9263 6307
rect 6837 6205 6871 6239
rect 7205 6205 7239 6239
rect 4169 6069 4203 6103
rect 6377 6069 6411 6103
rect 6745 6069 6779 6103
rect 9137 6069 9171 6103
rect 9413 6069 9447 6103
rect 2973 5865 3007 5899
rect 3801 5865 3835 5899
rect 8033 5865 8067 5899
rect 9137 5865 9171 5899
rect 9321 5865 9355 5899
rect 3065 5797 3099 5831
rect 3617 5797 3651 5831
rect 4261 5729 4295 5763
rect 4537 5729 4571 5763
rect 6285 5729 6319 5763
rect 2513 5661 2547 5695
rect 2789 5661 2823 5695
rect 3433 5661 3467 5695
rect 4077 5661 4111 5695
rect 8309 5661 8343 5695
rect 9229 5661 9263 5695
rect 9505 5661 9539 5695
rect 3249 5593 3283 5627
rect 6561 5593 6595 5627
rect 8125 5593 8159 5627
rect 2697 5525 2731 5559
rect 6009 5525 6043 5559
rect 8493 5525 8527 5559
rect 8769 5525 8803 5559
rect 5089 5321 5123 5355
rect 5365 5321 5399 5355
rect 3341 5185 3375 5219
rect 5181 5185 5215 5219
rect 5641 5185 5675 5219
rect 6193 5185 6227 5219
rect 7665 5185 7699 5219
rect 8309 5185 8343 5219
rect 3617 5117 3651 5151
rect 5825 5117 5859 5151
rect 8125 5117 8159 5151
rect 8677 5117 8711 5151
rect 8861 5117 8895 5151
rect 8493 5049 8527 5083
rect 5457 4981 5491 5015
rect 9321 4981 9355 5015
rect 3801 4777 3835 4811
rect 4445 4777 4479 4811
rect 5549 4777 5583 4811
rect 7021 4777 7055 4811
rect 7297 4777 7331 4811
rect 9413 4777 9447 4811
rect 6745 4709 6779 4743
rect 8309 4709 8343 4743
rect 5273 4641 5307 4675
rect 8769 4641 8803 4675
rect 3617 4573 3651 4607
rect 3709 4573 3743 4607
rect 4353 4573 4387 4607
rect 4905 4573 4939 4607
rect 5089 4573 5123 4607
rect 5365 4573 5399 4607
rect 5733 4573 5767 4607
rect 6377 4573 6411 4607
rect 6561 4573 6595 4607
rect 6837 4573 6871 4607
rect 7113 4573 7147 4607
rect 7573 4573 7607 4607
rect 7757 4573 7791 4607
rect 7849 4573 7883 4607
rect 5917 4505 5951 4539
rect 7389 4505 7423 4539
rect 8401 4505 8435 4539
rect 3433 4437 3467 4471
rect 4169 4437 4203 4471
rect 4813 4437 4847 4471
rect 6101 4437 6135 4471
rect 6193 4437 6227 4471
rect 8493 4437 8527 4471
rect 8953 4437 8987 4471
rect 9045 4437 9079 4471
rect 8677 4233 8711 4267
rect 7297 4165 7331 4199
rect 9045 4165 9079 4199
rect 3341 4097 3375 4131
rect 3985 4097 4019 4131
rect 5457 4097 5491 4131
rect 6009 4097 6043 4131
rect 6285 4097 6319 4131
rect 6561 4097 6595 4131
rect 7113 4097 7147 4131
rect 7573 4097 7607 4131
rect 8125 4097 8159 4131
rect 8585 4097 8619 4131
rect 9137 4097 9171 4131
rect 3617 4029 3651 4063
rect 7021 4029 7055 4063
rect 9229 4029 9263 4063
rect 3525 3961 3559 3995
rect 6193 3961 6227 3995
rect 7941 3961 7975 3995
rect 5917 3893 5951 3927
rect 6469 3893 6503 3927
rect 6653 3893 6687 3927
rect 7481 3893 7515 3927
rect 7757 3893 7791 3927
rect 8401 3893 8435 3927
rect 4537 3689 4571 3723
rect 4905 3689 4939 3723
rect 8861 3689 8895 3723
rect 9229 3689 9263 3723
rect 6561 3553 6595 3587
rect 4353 3485 4387 3519
rect 4721 3485 4755 3519
rect 4997 3485 5031 3519
rect 6929 3485 6963 3519
rect 8401 3485 8435 3519
rect 8953 3485 8987 3519
rect 5181 3349 5215 3383
rect 8585 3349 8619 3383
rect 9413 3349 9447 3383
rect 7849 3145 7883 3179
rect 8125 3145 8159 3179
rect 8401 3145 8435 3179
rect 8769 3145 8803 3179
rect 4261 3009 4295 3043
rect 4629 3009 4663 3043
rect 6101 3009 6135 3043
rect 7665 3009 7699 3043
rect 7941 3009 7975 3043
rect 8309 3009 8343 3043
rect 8585 3009 8619 3043
rect 8861 3009 8895 3043
rect 9229 3009 9263 3043
rect 6561 2873 6595 2907
rect 9045 2873 9079 2907
rect 9413 2805 9447 2839
rect 8217 2601 8251 2635
rect 8953 2601 8987 2635
rect 9413 2601 9447 2635
rect 8861 2533 8895 2567
rect 8677 2397 8711 2431
rect 9137 2397 9171 2431
rect 9229 2397 9263 2431
rect 8585 2329 8619 2363
rect 9321 2057 9355 2091
rect 8861 1921 8895 1955
rect 9505 1921 9539 1955
rect 8953 1853 8987 1887
rect 9137 1717 9171 1751
<< metal1 >>
rect 2225 12291 2283 12297
rect 2225 12257 2237 12291
rect 2271 12288 2283 12291
rect 6178 12288 6184 12300
rect 2271 12260 6184 12288
rect 2271 12257 2283 12260
rect 2225 12251 2283 12257
rect 6178 12248 6184 12260
rect 6236 12248 6242 12300
rect 2409 12223 2467 12229
rect 2409 12189 2421 12223
rect 2455 12220 2467 12223
rect 6546 12220 6552 12232
rect 2455 12192 6552 12220
rect 2455 12189 2467 12192
rect 2409 12183 2467 12189
rect 6546 12180 6552 12192
rect 6604 12180 6610 12232
rect 1946 12112 1952 12164
rect 2004 12152 2010 12164
rect 8386 12152 8392 12164
rect 2004 12124 8392 12152
rect 2004 12112 2010 12124
rect 8386 12112 8392 12124
rect 8444 12112 8450 12164
rect 1762 12044 1768 12096
rect 1820 12084 1826 12096
rect 5994 12084 6000 12096
rect 1820 12056 6000 12084
rect 1820 12044 1826 12056
rect 5994 12044 6000 12056
rect 6052 12044 6058 12096
rect 3878 11976 3884 12028
rect 3936 12016 3942 12028
rect 6454 12016 6460 12028
rect 3936 11988 6460 12016
rect 3936 11976 3942 11988
rect 6454 11976 6460 11988
rect 6512 12016 6518 12028
rect 7834 12016 7840 12028
rect 6512 11988 7840 12016
rect 6512 11976 6518 11988
rect 7834 11976 7840 11988
rect 7892 11976 7898 12028
rect 1302 11908 1308 11960
rect 1360 11948 1366 11960
rect 4614 11948 4620 11960
rect 1360 11920 4620 11948
rect 1360 11908 1366 11920
rect 4614 11908 4620 11920
rect 4672 11908 4678 11960
rect 4706 11908 4712 11960
rect 4764 11948 4770 11960
rect 6089 11951 6147 11957
rect 6089 11948 6101 11951
rect 4764 11920 6101 11948
rect 4764 11908 4770 11920
rect 6089 11917 6101 11920
rect 6135 11917 6147 11951
rect 6089 11911 6147 11917
rect 5534 11880 5540 11892
rect 2746 11852 5540 11880
rect 2130 11772 2136 11824
rect 2188 11812 2194 11824
rect 2746 11812 2774 11852
rect 5534 11840 5540 11852
rect 5592 11880 5598 11892
rect 5994 11880 6000 11892
rect 5592 11852 6000 11880
rect 5592 11840 5598 11852
rect 5994 11840 6000 11852
rect 6052 11840 6058 11892
rect 2188 11784 2774 11812
rect 2188 11772 2194 11784
rect 3050 11772 3056 11824
rect 3108 11812 3114 11824
rect 9214 11812 9220 11824
rect 3108 11784 9220 11812
rect 3108 11772 3114 11784
rect 9214 11772 9220 11784
rect 9272 11772 9278 11824
rect 934 11704 940 11756
rect 992 11744 998 11756
rect 4338 11744 4344 11756
rect 992 11716 4344 11744
rect 992 11704 998 11716
rect 4338 11704 4344 11716
rect 4396 11704 4402 11756
rect 6086 11744 6092 11756
rect 5999 11716 6092 11744
rect 6086 11704 6092 11716
rect 6144 11744 6150 11756
rect 7650 11744 7656 11756
rect 6144 11716 7656 11744
rect 6144 11704 6150 11716
rect 7650 11704 7656 11716
rect 7708 11704 7714 11756
rect 3142 11636 3148 11688
rect 3200 11676 3206 11688
rect 7558 11676 7564 11688
rect 3200 11648 7564 11676
rect 3200 11636 3206 11648
rect 7558 11636 7564 11648
rect 7616 11636 7622 11688
rect 7742 11636 7748 11688
rect 7800 11676 7806 11688
rect 9122 11676 9128 11688
rect 7800 11648 9128 11676
rect 7800 11636 7806 11648
rect 9122 11636 9128 11648
rect 9180 11636 9186 11688
rect 1118 11568 1124 11620
rect 1176 11608 1182 11620
rect 2774 11608 2780 11620
rect 1176 11580 2780 11608
rect 1176 11568 1182 11580
rect 2774 11568 2780 11580
rect 2832 11568 2838 11620
rect 3234 11568 3240 11620
rect 3292 11608 3298 11620
rect 6270 11608 6276 11620
rect 3292 11580 6276 11608
rect 3292 11568 3298 11580
rect 6270 11568 6276 11580
rect 6328 11568 6334 11620
rect 7190 11568 7196 11620
rect 7248 11608 7254 11620
rect 9306 11608 9312 11620
rect 7248 11580 9312 11608
rect 7248 11568 7254 11580
rect 9306 11568 9312 11580
rect 9364 11568 9370 11620
rect 2038 11500 2044 11552
rect 2096 11540 2102 11552
rect 2225 11543 2283 11549
rect 2225 11540 2237 11543
rect 2096 11512 2237 11540
rect 2096 11500 2102 11512
rect 2225 11509 2237 11512
rect 2271 11509 2283 11543
rect 2225 11503 2283 11509
rect 2314 11500 2320 11552
rect 2372 11540 2378 11552
rect 2409 11543 2467 11549
rect 2409 11540 2421 11543
rect 2372 11512 2421 11540
rect 2372 11500 2378 11512
rect 2409 11509 2421 11512
rect 2455 11509 2467 11543
rect 2409 11503 2467 11509
rect 3602 11500 3608 11552
rect 3660 11540 3666 11552
rect 8662 11540 8668 11552
rect 3660 11512 8668 11540
rect 3660 11500 3666 11512
rect 8662 11500 8668 11512
rect 8720 11500 8726 11552
rect 920 11450 9844 11472
rect 920 11398 2566 11450
rect 2618 11398 2630 11450
rect 2682 11398 2694 11450
rect 2746 11398 2758 11450
rect 2810 11398 2822 11450
rect 2874 11398 5666 11450
rect 5718 11398 5730 11450
rect 5782 11398 5794 11450
rect 5846 11398 5858 11450
rect 5910 11398 5922 11450
rect 5974 11398 8766 11450
rect 8818 11398 8830 11450
rect 8882 11398 8894 11450
rect 8946 11398 8958 11450
rect 9010 11398 9022 11450
rect 9074 11398 9844 11450
rect 920 11376 9844 11398
rect 1397 11339 1455 11345
rect 1397 11305 1409 11339
rect 1443 11336 1455 11339
rect 1670 11336 1676 11348
rect 1443 11308 1676 11336
rect 1443 11305 1455 11308
rect 1397 11299 1455 11305
rect 1670 11296 1676 11308
rect 1728 11296 1734 11348
rect 2038 11336 2044 11348
rect 1999 11308 2044 11336
rect 2038 11296 2044 11308
rect 2096 11296 2102 11348
rect 2314 11336 2320 11348
rect 2275 11308 2320 11336
rect 2314 11296 2320 11308
rect 2372 11296 2378 11348
rect 3142 11336 3148 11348
rect 3103 11308 3148 11336
rect 3142 11296 3148 11308
rect 3200 11296 3206 11348
rect 3421 11339 3479 11345
rect 3421 11305 3433 11339
rect 3467 11336 3479 11339
rect 4430 11336 4436 11348
rect 3467 11308 4436 11336
rect 3467 11305 3479 11308
rect 3421 11299 3479 11305
rect 4430 11296 4436 11308
rect 4488 11296 4494 11348
rect 5629 11339 5687 11345
rect 5629 11336 5641 11339
rect 4632 11308 5641 11336
rect 2593 11271 2651 11277
rect 2593 11237 2605 11271
rect 2639 11268 2651 11271
rect 3602 11268 3608 11280
rect 2639 11240 3608 11268
rect 2639 11237 2651 11240
rect 2593 11231 2651 11237
rect 3602 11228 3608 11240
rect 3660 11228 3666 11280
rect 3694 11228 3700 11280
rect 3752 11268 3758 11280
rect 4065 11271 4123 11277
rect 4065 11268 4077 11271
rect 3752 11240 4077 11268
rect 3752 11228 3758 11240
rect 4065 11237 4077 11240
rect 4111 11237 4123 11271
rect 4338 11268 4344 11280
rect 4299 11240 4344 11268
rect 4065 11231 4123 11237
rect 4338 11228 4344 11240
rect 4396 11228 4402 11280
rect 4525 11271 4583 11277
rect 4525 11237 4537 11271
rect 4571 11237 4583 11271
rect 4525 11231 4583 11237
rect 1578 11160 1584 11212
rect 1636 11200 1642 11212
rect 3510 11200 3516 11212
rect 1636 11172 2452 11200
rect 1636 11160 1642 11172
rect 934 11092 940 11144
rect 992 11132 998 11144
rect 1213 11135 1271 11141
rect 1213 11132 1225 11135
rect 992 11104 1225 11132
rect 992 11092 998 11104
rect 1213 11101 1225 11104
rect 1259 11101 1271 11135
rect 1486 11132 1492 11144
rect 1447 11104 1492 11132
rect 1213 11095 1271 11101
rect 1486 11092 1492 11104
rect 1544 11092 1550 11144
rect 1762 11092 1768 11144
rect 1820 11132 1826 11144
rect 1857 11135 1915 11141
rect 1857 11132 1869 11135
rect 1820 11104 1869 11132
rect 1820 11092 1826 11104
rect 1857 11101 1869 11104
rect 1903 11101 1915 11135
rect 2130 11132 2136 11144
rect 2091 11104 2136 11132
rect 1857 11095 1915 11101
rect 2130 11092 2136 11104
rect 2188 11092 2194 11144
rect 2424 11141 2452 11172
rect 3160 11172 3516 11200
rect 2409 11135 2467 11141
rect 2409 11101 2421 11135
rect 2455 11132 2467 11135
rect 2590 11132 2596 11144
rect 2455 11104 2596 11132
rect 2455 11101 2467 11104
rect 2409 11095 2467 11101
rect 2590 11092 2596 11104
rect 2648 11092 2654 11144
rect 2685 11135 2743 11141
rect 2685 11101 2697 11135
rect 2731 11132 2743 11135
rect 2774 11132 2780 11144
rect 2731 11104 2780 11132
rect 2731 11101 2743 11104
rect 2685 11095 2743 11101
rect 2774 11092 2780 11104
rect 2832 11092 2838 11144
rect 2961 11135 3019 11141
rect 2961 11101 2973 11135
rect 3007 11132 3019 11135
rect 3160 11132 3188 11172
rect 3510 11160 3516 11172
rect 3568 11160 3574 11212
rect 4540 11200 4568 11231
rect 3804 11172 4568 11200
rect 3804 11141 3832 11172
rect 3007 11104 3188 11132
rect 3789 11135 3847 11141
rect 3007 11101 3019 11104
rect 2961 11095 3019 11101
rect 2314 11024 2320 11076
rect 2372 11064 2378 11076
rect 3234 11068 3240 11120
rect 3292 11108 3298 11120
rect 3292 11080 3337 11108
rect 3789 11101 3801 11135
rect 3835 11101 3847 11135
rect 3789 11095 3847 11101
rect 4249 11135 4307 11141
rect 4249 11101 4261 11135
rect 4295 11132 4307 11135
rect 4632 11132 4660 11308
rect 5629 11305 5641 11308
rect 5675 11305 5687 11339
rect 5994 11336 6000 11348
rect 5955 11308 6000 11336
rect 5629 11299 5687 11305
rect 5994 11296 6000 11308
rect 6052 11296 6058 11348
rect 6270 11336 6276 11348
rect 6231 11308 6276 11336
rect 6270 11296 6276 11308
rect 6328 11296 6334 11348
rect 6638 11336 6644 11348
rect 6599 11308 6644 11336
rect 6638 11296 6644 11308
rect 6696 11296 6702 11348
rect 7742 11336 7748 11348
rect 7484 11308 7748 11336
rect 5261 11271 5319 11277
rect 5261 11237 5273 11271
rect 5307 11237 5319 11271
rect 5261 11231 5319 11237
rect 5537 11271 5595 11277
rect 5537 11237 5549 11271
rect 5583 11268 5595 11271
rect 7484 11268 7512 11308
rect 7742 11296 7748 11308
rect 7800 11296 7806 11348
rect 8021 11339 8079 11345
rect 8021 11305 8033 11339
rect 8067 11336 8079 11339
rect 8202 11336 8208 11348
rect 8067 11308 8208 11336
rect 8067 11305 8079 11308
rect 8021 11299 8079 11305
rect 8202 11296 8208 11308
rect 8260 11296 8266 11348
rect 5583 11240 7512 11268
rect 7561 11271 7619 11277
rect 5583 11237 5595 11240
rect 5537 11231 5595 11237
rect 7561 11237 7573 11271
rect 7607 11268 7619 11271
rect 8478 11268 8484 11280
rect 7607 11240 8484 11268
rect 7607 11237 7619 11240
rect 7561 11231 7619 11237
rect 5276 11200 5304 11231
rect 8478 11228 8484 11240
rect 8536 11228 8542 11280
rect 9033 11271 9091 11277
rect 9033 11237 9045 11271
rect 9079 11268 9091 11271
rect 13814 11268 13820 11280
rect 9079 11240 13820 11268
rect 9079 11237 9091 11240
rect 9033 11231 9091 11237
rect 13814 11228 13820 11240
rect 13872 11228 13878 11280
rect 8386 11200 8392 11212
rect 5276 11172 6868 11200
rect 4295 11104 4660 11132
rect 4295 11101 4307 11104
rect 4249 11095 4307 11101
rect 4706 11092 4712 11144
rect 4764 11132 4770 11144
rect 4982 11132 4988 11144
rect 4764 11104 4809 11132
rect 4943 11104 4988 11132
rect 4764 11092 4770 11104
rect 4982 11092 4988 11104
rect 5040 11092 5046 11144
rect 5077 11135 5135 11141
rect 5077 11101 5089 11135
rect 5123 11132 5135 11135
rect 5258 11132 5264 11144
rect 5123 11104 5264 11132
rect 5123 11101 5135 11104
rect 5077 11095 5135 11101
rect 5258 11092 5264 11104
rect 5316 11092 5322 11144
rect 5353 11135 5411 11141
rect 5353 11101 5365 11135
rect 5399 11132 5411 11135
rect 5813 11135 5871 11141
rect 5399 11104 5764 11132
rect 5399 11101 5411 11104
rect 5353 11095 5411 11101
rect 3292 11068 3298 11080
rect 2372 11036 3188 11064
rect 2372 11024 2378 11036
rect 1673 10999 1731 11005
rect 1673 10965 1685 10999
rect 1719 10996 1731 10999
rect 2774 10996 2780 11008
rect 1719 10968 2780 10996
rect 1719 10965 1731 10968
rect 1673 10959 1731 10965
rect 2774 10956 2780 10968
rect 2832 10956 2838 11008
rect 2869 10999 2927 11005
rect 2869 10965 2881 10999
rect 2915 10996 2927 10999
rect 3050 10996 3056 11008
rect 2915 10968 3056 10996
rect 2915 10965 2927 10968
rect 2869 10959 2927 10965
rect 3050 10956 3056 10968
rect 3108 10956 3114 11008
rect 3160 10996 3188 11036
rect 4430 11024 4436 11076
rect 4488 11064 4494 11076
rect 5626 11064 5632 11076
rect 4488 11036 5632 11064
rect 4488 11024 4494 11036
rect 5626 11024 5632 11036
rect 5684 11024 5690 11076
rect 5736 11064 5764 11104
rect 5813 11101 5825 11135
rect 5859 11132 5871 11135
rect 5902 11132 5908 11144
rect 5859 11104 5908 11132
rect 5859 11101 5871 11104
rect 5813 11095 5871 11101
rect 5902 11092 5908 11104
rect 5960 11092 5966 11144
rect 6086 11092 6092 11144
rect 6144 11132 6150 11144
rect 6840 11141 6868 11172
rect 7300 11172 8064 11200
rect 6733 11135 6791 11141
rect 6733 11132 6745 11135
rect 6144 11104 6745 11132
rect 6144 11092 6150 11104
rect 6733 11101 6745 11104
rect 6779 11101 6791 11135
rect 6733 11095 6791 11101
rect 6825 11135 6883 11141
rect 6825 11101 6837 11135
rect 6871 11101 6883 11135
rect 7098 11132 7104 11144
rect 7059 11104 7104 11132
rect 6825 11095 6883 11101
rect 7098 11092 7104 11104
rect 7156 11092 7162 11144
rect 7190 11064 7196 11076
rect 5736 11036 7196 11064
rect 7190 11024 7196 11036
rect 7248 11024 7254 11076
rect 3697 10999 3755 11005
rect 3697 10996 3709 10999
rect 3160 10968 3709 10996
rect 3697 10965 3709 10968
rect 3743 10996 3755 10999
rect 3786 10996 3792 11008
rect 3743 10968 3792 10996
rect 3743 10965 3755 10968
rect 3697 10959 3755 10965
rect 3786 10956 3792 10968
rect 3844 10956 3850 11008
rect 3970 10996 3976 11008
rect 3931 10968 3976 10996
rect 3970 10956 3976 10968
rect 4028 10956 4034 11008
rect 4798 10996 4804 11008
rect 4759 10968 4804 10996
rect 4798 10956 4804 10968
rect 4856 10956 4862 11008
rect 4890 10956 4896 11008
rect 4948 10996 4954 11008
rect 5902 10996 5908 11008
rect 4948 10968 5908 10996
rect 4948 10956 4954 10968
rect 5902 10956 5908 10968
rect 5960 10996 5966 11008
rect 6638 10996 6644 11008
rect 5960 10968 6644 10996
rect 5960 10956 5966 10968
rect 6638 10956 6644 10968
rect 6696 10956 6702 11008
rect 7006 10996 7012 11008
rect 6967 10968 7012 10996
rect 7006 10956 7012 10968
rect 7064 10956 7070 11008
rect 7300 11005 7328 11172
rect 7377 11135 7435 11141
rect 7377 11101 7389 11135
rect 7423 11132 7435 11135
rect 7423 11104 7696 11132
rect 7423 11101 7435 11104
rect 7377 11095 7435 11101
rect 7668 11005 7696 11104
rect 8036 11064 8064 11172
rect 8128 11172 8392 11200
rect 8128 11141 8156 11172
rect 8386 11160 8392 11172
rect 8444 11160 8450 11212
rect 13722 11200 13728 11212
rect 8496 11172 13728 11200
rect 8113 11135 8171 11141
rect 8113 11101 8125 11135
rect 8159 11101 8171 11135
rect 8294 11132 8300 11144
rect 8255 11104 8300 11132
rect 8113 11095 8171 11101
rect 8294 11092 8300 11104
rect 8352 11092 8358 11144
rect 8386 11064 8392 11076
rect 8036 11036 8392 11064
rect 8386 11024 8392 11036
rect 8444 11024 8450 11076
rect 8496 11005 8524 11172
rect 13722 11160 13728 11172
rect 13780 11160 13786 11212
rect 8662 11092 8668 11144
rect 8720 11132 8726 11144
rect 8849 11135 8907 11141
rect 8849 11132 8861 11135
rect 8720 11104 8861 11132
rect 8720 11092 8726 11104
rect 8849 11101 8861 11104
rect 8895 11101 8907 11135
rect 9214 11132 9220 11144
rect 9175 11104 9220 11132
rect 8849 11095 8907 11101
rect 9214 11092 9220 11104
rect 9272 11092 9278 11144
rect 7285 10999 7343 11005
rect 7285 10965 7297 10999
rect 7331 10965 7343 10999
rect 7285 10959 7343 10965
rect 7653 10999 7711 11005
rect 7653 10965 7665 10999
rect 7699 10965 7711 10999
rect 7653 10959 7711 10965
rect 8481 10999 8539 11005
rect 8481 10965 8493 10999
rect 8527 10965 8539 10999
rect 9398 10996 9404 11008
rect 9359 10968 9404 10996
rect 8481 10959 8539 10965
rect 9398 10956 9404 10968
rect 9456 10956 9462 11008
rect 920 10906 9844 10928
rect 920 10854 4116 10906
rect 4168 10854 4180 10906
rect 4232 10854 4244 10906
rect 4296 10854 4308 10906
rect 4360 10854 4372 10906
rect 4424 10854 7216 10906
rect 7268 10854 7280 10906
rect 7332 10854 7344 10906
rect 7396 10854 7408 10906
rect 7460 10854 7472 10906
rect 7524 10854 9844 10906
rect 920 10832 9844 10854
rect 1397 10795 1455 10801
rect 1397 10761 1409 10795
rect 1443 10792 1455 10795
rect 1578 10792 1584 10804
rect 1443 10764 1584 10792
rect 1443 10761 1455 10764
rect 1397 10755 1455 10761
rect 1578 10752 1584 10764
rect 1636 10752 1642 10804
rect 3878 10792 3884 10804
rect 2608 10764 3884 10792
rect 1302 10684 1308 10736
rect 1360 10724 1366 10736
rect 1360 10696 1808 10724
rect 1360 10684 1366 10696
rect 1210 10656 1216 10668
rect 1171 10628 1216 10656
rect 1210 10616 1216 10628
rect 1268 10616 1274 10668
rect 1394 10616 1400 10668
rect 1452 10656 1458 10668
rect 1780 10665 1808 10696
rect 1489 10659 1547 10665
rect 1489 10656 1501 10659
rect 1452 10628 1501 10656
rect 1452 10616 1458 10628
rect 1489 10625 1501 10628
rect 1535 10625 1547 10659
rect 1489 10619 1547 10625
rect 1765 10659 1823 10665
rect 1765 10625 1777 10659
rect 1811 10625 1823 10659
rect 1765 10619 1823 10625
rect 2041 10659 2099 10665
rect 2041 10625 2053 10659
rect 2087 10656 2099 10659
rect 2130 10656 2136 10668
rect 2087 10628 2136 10656
rect 2087 10625 2099 10628
rect 2041 10619 2099 10625
rect 2130 10616 2136 10628
rect 2188 10616 2194 10668
rect 2314 10656 2320 10668
rect 2275 10628 2320 10656
rect 2314 10616 2320 10628
rect 2372 10616 2378 10668
rect 2608 10665 2636 10764
rect 3878 10752 3884 10764
rect 3936 10752 3942 10804
rect 4341 10795 4399 10801
rect 4341 10761 4353 10795
rect 4387 10792 4399 10795
rect 4982 10792 4988 10804
rect 4387 10764 4988 10792
rect 4387 10761 4399 10764
rect 4341 10755 4399 10761
rect 4982 10752 4988 10764
rect 5040 10752 5046 10804
rect 5626 10752 5632 10804
rect 5684 10792 5690 10804
rect 5684 10764 6960 10792
rect 5684 10752 5690 10764
rect 3068 10696 3556 10724
rect 2593 10659 2651 10665
rect 2593 10625 2605 10659
rect 2639 10625 2651 10659
rect 2593 10619 2651 10625
rect 2869 10659 2927 10665
rect 2869 10625 2881 10659
rect 2915 10656 2927 10659
rect 2958 10656 2964 10668
rect 2915 10628 2964 10656
rect 2915 10625 2927 10628
rect 2869 10619 2927 10625
rect 2958 10616 2964 10628
rect 3016 10616 3022 10668
rect 3068 10588 3096 10696
rect 3234 10616 3240 10668
rect 3292 10656 3298 10668
rect 3421 10659 3479 10665
rect 3421 10656 3433 10659
rect 3292 10628 3433 10656
rect 3292 10616 3298 10628
rect 3421 10625 3433 10628
rect 3467 10625 3479 10659
rect 3421 10619 3479 10625
rect 2884 10560 3096 10588
rect 1673 10523 1731 10529
rect 1673 10489 1685 10523
rect 1719 10520 1731 10523
rect 2130 10520 2136 10532
rect 1719 10492 2136 10520
rect 1719 10489 1731 10492
rect 1673 10483 1731 10489
rect 2130 10480 2136 10492
rect 2188 10480 2194 10532
rect 1946 10452 1952 10464
rect 1907 10424 1952 10452
rect 1946 10412 1952 10424
rect 2004 10412 2010 10464
rect 2225 10455 2283 10461
rect 2225 10421 2237 10455
rect 2271 10452 2283 10455
rect 2314 10452 2320 10464
rect 2271 10424 2320 10452
rect 2271 10421 2283 10424
rect 2225 10415 2283 10421
rect 2314 10412 2320 10424
rect 2372 10412 2378 10464
rect 2406 10412 2412 10464
rect 2464 10452 2470 10464
rect 2501 10455 2559 10461
rect 2501 10452 2513 10455
rect 2464 10424 2513 10452
rect 2464 10412 2470 10424
rect 2501 10421 2513 10424
rect 2547 10421 2559 10455
rect 2501 10415 2559 10421
rect 2777 10455 2835 10461
rect 2777 10421 2789 10455
rect 2823 10452 2835 10455
rect 2884 10452 2912 10560
rect 3142 10548 3148 10600
rect 3200 10588 3206 10600
rect 3329 10591 3387 10597
rect 3329 10588 3341 10591
rect 3200 10560 3341 10588
rect 3200 10548 3206 10560
rect 3329 10557 3341 10560
rect 3375 10557 3387 10591
rect 3329 10551 3387 10557
rect 3418 10480 3424 10532
rect 3476 10520 3482 10532
rect 3528 10520 3556 10696
rect 3970 10684 3976 10736
rect 4028 10724 4034 10736
rect 4028 10696 6224 10724
rect 6932 10710 6960 10764
rect 7098 10752 7104 10804
rect 7156 10792 7162 10804
rect 8941 10795 8999 10801
rect 8941 10792 8953 10795
rect 7156 10764 8953 10792
rect 7156 10752 7162 10764
rect 8941 10761 8953 10764
rect 8987 10761 8999 10795
rect 8941 10755 8999 10761
rect 8570 10724 8576 10736
rect 8531 10696 8576 10724
rect 4028 10684 4034 10696
rect 3605 10659 3663 10665
rect 3605 10625 3617 10659
rect 3651 10625 3663 10659
rect 3878 10656 3884 10668
rect 3839 10628 3884 10656
rect 3605 10619 3663 10625
rect 3476 10492 3556 10520
rect 3620 10588 3648 10619
rect 3878 10616 3884 10628
rect 3936 10656 3942 10668
rect 4433 10659 4491 10665
rect 4433 10656 4445 10659
rect 3936 10628 4445 10656
rect 3936 10616 3942 10628
rect 4433 10625 4445 10628
rect 4479 10625 4491 10659
rect 4433 10619 4491 10625
rect 4617 10659 4675 10665
rect 4617 10625 4629 10659
rect 4663 10656 4675 10659
rect 4890 10656 4896 10668
rect 4663 10628 4896 10656
rect 4663 10625 4675 10628
rect 4617 10619 4675 10625
rect 4632 10588 4660 10619
rect 4890 10616 4896 10628
rect 4948 10616 4954 10668
rect 5077 10659 5135 10665
rect 5077 10625 5089 10659
rect 5123 10656 5135 10659
rect 5350 10656 5356 10668
rect 5123 10628 5212 10656
rect 5311 10628 5356 10656
rect 5123 10625 5135 10628
rect 5077 10619 5135 10625
rect 3620 10560 4660 10588
rect 3476 10480 3482 10492
rect 3620 10464 3648 10560
rect 2823 10424 2912 10452
rect 3145 10455 3203 10461
rect 2823 10421 2835 10424
rect 2777 10415 2835 10421
rect 3145 10421 3157 10455
rect 3191 10452 3203 10455
rect 3602 10452 3608 10464
rect 3191 10424 3608 10452
rect 3191 10421 3203 10424
rect 3145 10415 3203 10421
rect 3602 10412 3608 10424
rect 3660 10412 3666 10464
rect 3786 10452 3792 10464
rect 3747 10424 3792 10452
rect 3786 10412 3792 10424
rect 3844 10412 3850 10464
rect 4080 10461 4108 10560
rect 4154 10480 4160 10532
rect 4212 10520 4218 10532
rect 4801 10523 4859 10529
rect 4801 10520 4813 10523
rect 4212 10492 4813 10520
rect 4212 10480 4218 10492
rect 4801 10489 4813 10492
rect 4847 10489 4859 10523
rect 5184 10520 5212 10628
rect 5350 10616 5356 10628
rect 5408 10616 5414 10668
rect 5534 10616 5540 10668
rect 5592 10656 5598 10668
rect 5629 10659 5687 10665
rect 5629 10656 5641 10659
rect 5592 10628 5641 10656
rect 5592 10616 5598 10628
rect 5629 10625 5641 10628
rect 5675 10625 5687 10659
rect 5629 10619 5687 10625
rect 5813 10659 5871 10665
rect 5813 10625 5825 10659
rect 5859 10625 5871 10659
rect 5813 10619 5871 10625
rect 5258 10548 5264 10600
rect 5316 10588 5322 10600
rect 5829 10588 5857 10619
rect 5902 10616 5908 10668
rect 5960 10656 5966 10668
rect 6196 10665 6224 10696
rect 8570 10684 8576 10696
rect 8628 10684 8634 10736
rect 5997 10659 6055 10665
rect 5997 10656 6009 10659
rect 5960 10628 6009 10656
rect 5960 10616 5966 10628
rect 5997 10625 6009 10628
rect 6043 10625 6055 10659
rect 5997 10619 6055 10625
rect 6181 10659 6239 10665
rect 6181 10625 6193 10659
rect 6227 10625 6239 10659
rect 6181 10619 6239 10625
rect 7558 10616 7564 10668
rect 7616 10656 7622 10668
rect 8021 10659 8079 10665
rect 8021 10656 8033 10659
rect 7616 10628 8033 10656
rect 7616 10616 7622 10628
rect 8021 10625 8033 10628
rect 8067 10625 8079 10659
rect 8021 10619 8079 10625
rect 8202 10616 8208 10668
rect 8260 10656 8266 10668
rect 8757 10659 8815 10665
rect 8757 10656 8769 10659
rect 8260 10628 8769 10656
rect 8260 10616 8266 10628
rect 8757 10625 8769 10628
rect 8803 10625 8815 10659
rect 8757 10619 8815 10625
rect 9217 10659 9275 10665
rect 9217 10625 9229 10659
rect 9263 10625 9275 10659
rect 9217 10619 9275 10625
rect 6086 10588 6092 10600
rect 5316 10560 6092 10588
rect 5316 10548 5322 10560
rect 6086 10548 6092 10560
rect 6144 10548 6150 10600
rect 6549 10591 6607 10597
rect 6549 10557 6561 10591
rect 6595 10588 6607 10591
rect 6822 10588 6828 10600
rect 6595 10560 6828 10588
rect 6595 10557 6607 10560
rect 6549 10551 6607 10557
rect 6822 10548 6828 10560
rect 6880 10548 6886 10600
rect 8110 10548 8116 10600
rect 8168 10588 8174 10600
rect 9232 10588 9260 10619
rect 8168 10560 9260 10588
rect 8168 10548 8174 10560
rect 5184 10492 6316 10520
rect 4801 10483 4859 10489
rect 4065 10455 4123 10461
rect 4065 10421 4077 10455
rect 4111 10421 4123 10455
rect 4065 10415 4123 10421
rect 4522 10412 4528 10464
rect 4580 10452 4586 10464
rect 4893 10455 4951 10461
rect 4893 10452 4905 10455
rect 4580 10424 4905 10452
rect 4580 10412 4586 10424
rect 4893 10421 4905 10424
rect 4939 10421 4951 10455
rect 5258 10452 5264 10464
rect 5219 10424 5264 10452
rect 4893 10415 4951 10421
rect 5258 10412 5264 10424
rect 5316 10412 5322 10464
rect 5534 10452 5540 10464
rect 5495 10424 5540 10452
rect 5534 10412 5540 10424
rect 5592 10412 5598 10464
rect 6288 10452 6316 10492
rect 7834 10480 7840 10532
rect 7892 10520 7898 10532
rect 9033 10523 9091 10529
rect 9033 10520 9045 10523
rect 7892 10492 9045 10520
rect 7892 10480 7898 10492
rect 9033 10489 9045 10492
rect 9079 10489 9091 10523
rect 9033 10483 9091 10489
rect 7926 10452 7932 10464
rect 6288 10424 7932 10452
rect 7926 10412 7932 10424
rect 7984 10412 7990 10464
rect 8481 10455 8539 10461
rect 8481 10421 8493 10455
rect 8527 10452 8539 10455
rect 8662 10452 8668 10464
rect 8527 10424 8668 10452
rect 8527 10421 8539 10424
rect 8481 10415 8539 10421
rect 8662 10412 8668 10424
rect 8720 10412 8726 10464
rect 9401 10455 9459 10461
rect 9401 10421 9413 10455
rect 9447 10452 9459 10455
rect 16574 10452 16580 10464
rect 9447 10424 16580 10452
rect 9447 10421 9459 10424
rect 9401 10415 9459 10421
rect 16574 10412 16580 10424
rect 16632 10412 16638 10464
rect 920 10362 9844 10384
rect 920 10310 2566 10362
rect 2618 10310 2630 10362
rect 2682 10310 2694 10362
rect 2746 10310 2758 10362
rect 2810 10310 2822 10362
rect 2874 10310 5666 10362
rect 5718 10310 5730 10362
rect 5782 10310 5794 10362
rect 5846 10310 5858 10362
rect 5910 10310 5922 10362
rect 5974 10310 8766 10362
rect 8818 10310 8830 10362
rect 8882 10310 8894 10362
rect 8946 10310 8958 10362
rect 9010 10310 9022 10362
rect 9074 10310 9844 10362
rect 920 10288 9844 10310
rect 1302 10248 1308 10260
rect 1263 10220 1308 10248
rect 1302 10208 1308 10220
rect 1360 10208 1366 10260
rect 1581 10251 1639 10257
rect 1581 10217 1593 10251
rect 1627 10248 1639 10251
rect 7573 10251 7631 10257
rect 7573 10248 7585 10251
rect 1627 10220 7585 10248
rect 1627 10217 1639 10220
rect 1581 10211 1639 10217
rect 7573 10217 7585 10220
rect 7619 10217 7631 10251
rect 7926 10248 7932 10260
rect 7887 10220 7932 10248
rect 7573 10211 7631 10217
rect 7926 10208 7932 10220
rect 7984 10208 7990 10260
rect 8202 10248 8208 10260
rect 8163 10220 8208 10248
rect 8202 10208 8208 10220
rect 8260 10208 8266 10260
rect 3602 10180 3608 10192
rect 3344 10152 3608 10180
rect 2498 10112 2504 10124
rect 2056 10084 2504 10112
rect 1394 10044 1400 10056
rect 1355 10016 1400 10044
rect 1394 10004 1400 10016
rect 1452 10004 1458 10056
rect 2056 10030 2084 10084
rect 2498 10072 2504 10084
rect 2556 10112 2562 10124
rect 3344 10112 3372 10152
rect 3602 10140 3608 10152
rect 3660 10140 3666 10192
rect 5534 10140 5540 10192
rect 5592 10140 5598 10192
rect 5997 10183 6055 10189
rect 5997 10149 6009 10183
rect 6043 10180 6055 10183
rect 6454 10180 6460 10192
rect 6043 10152 6460 10180
rect 6043 10149 6055 10152
rect 5997 10143 6055 10149
rect 6454 10140 6460 10152
rect 6512 10140 6518 10192
rect 7834 10140 7840 10192
rect 7892 10180 7898 10192
rect 9033 10183 9091 10189
rect 9033 10180 9045 10183
rect 7892 10152 9045 10180
rect 7892 10140 7898 10152
rect 9033 10149 9045 10152
rect 9079 10149 9091 10183
rect 9033 10143 9091 10149
rect 2556 10084 3372 10112
rect 3421 10115 3479 10121
rect 2556 10072 2562 10084
rect 3421 10081 3433 10115
rect 3467 10112 3479 10115
rect 4522 10112 4528 10124
rect 3467 10084 4528 10112
rect 3467 10081 3479 10084
rect 3421 10075 3479 10081
rect 4522 10072 4528 10084
rect 4580 10072 4586 10124
rect 5552 10112 5580 10140
rect 6914 10112 6920 10124
rect 5552 10084 6920 10112
rect 6914 10072 6920 10084
rect 6972 10072 6978 10124
rect 7098 10072 7104 10124
rect 7156 10112 7162 10124
rect 7156 10084 8892 10112
rect 7156 10072 7162 10084
rect 3694 10044 3700 10056
rect 3655 10016 3700 10044
rect 3694 10004 3700 10016
rect 3752 10004 3758 10056
rect 3970 10004 3976 10056
rect 4028 10044 4034 10056
rect 4065 10047 4123 10053
rect 4065 10044 4077 10047
rect 4028 10016 4077 10044
rect 4028 10004 4034 10016
rect 4065 10013 4077 10016
rect 4111 10013 4123 10047
rect 4065 10007 4123 10013
rect 4982 10004 4988 10056
rect 5040 10044 5046 10056
rect 7852 10053 7880 10084
rect 8864 10053 8892 10084
rect 5537 10047 5595 10053
rect 5537 10044 5549 10047
rect 5040 10016 5549 10044
rect 5040 10004 5046 10016
rect 5537 10013 5549 10016
rect 5583 10013 5595 10047
rect 5537 10007 5595 10013
rect 7837 10047 7895 10053
rect 7837 10013 7849 10047
rect 7883 10013 7895 10047
rect 7837 10007 7895 10013
rect 8389 10047 8447 10053
rect 8389 10013 8401 10047
rect 8435 10013 8447 10047
rect 8389 10007 8447 10013
rect 8849 10047 8907 10053
rect 8849 10013 8861 10047
rect 8895 10013 8907 10047
rect 9490 10044 9496 10056
rect 9451 10016 9496 10044
rect 8849 10007 8907 10013
rect 3142 9976 3148 9988
rect 3103 9948 3148 9976
rect 3142 9936 3148 9948
rect 3200 9936 3206 9988
rect 3418 9936 3424 9988
rect 3476 9976 3482 9988
rect 3602 9976 3608 9988
rect 3476 9948 3608 9976
rect 3476 9936 3482 9948
rect 3602 9936 3608 9948
rect 3660 9936 3666 9988
rect 4798 9936 4804 9988
rect 4856 9936 4862 9988
rect 1673 9911 1731 9917
rect 1673 9877 1685 9911
rect 1719 9908 1731 9911
rect 2222 9908 2228 9920
rect 1719 9880 2228 9908
rect 1719 9877 1731 9880
rect 1673 9871 1731 9877
rect 2222 9868 2228 9880
rect 2280 9908 2286 9920
rect 2498 9908 2504 9920
rect 2280 9880 2504 9908
rect 2280 9868 2286 9880
rect 2498 9868 2504 9880
rect 2556 9868 2562 9920
rect 6089 9911 6147 9917
rect 6089 9877 6101 9911
rect 6135 9908 6147 9911
rect 6822 9908 6828 9920
rect 6135 9880 6828 9908
rect 6135 9877 6147 9880
rect 6089 9871 6147 9877
rect 6822 9868 6828 9880
rect 6880 9868 6886 9920
rect 7116 9908 7144 9962
rect 7466 9936 7472 9988
rect 7524 9976 7530 9988
rect 8404 9976 8432 10007
rect 9490 10004 9496 10016
rect 9548 10004 9554 10056
rect 7524 9948 8892 9976
rect 7524 9936 7530 9948
rect 8864 9920 8892 9948
rect 8202 9908 8208 9920
rect 7116 9880 8208 9908
rect 8202 9868 8208 9880
rect 8260 9868 8266 9920
rect 8570 9908 8576 9920
rect 8531 9880 8576 9908
rect 8570 9868 8576 9880
rect 8628 9868 8634 9920
rect 8846 9868 8852 9920
rect 8904 9868 8910 9920
rect 9309 9911 9367 9917
rect 9309 9877 9321 9911
rect 9355 9908 9367 9911
rect 10870 9908 10876 9920
rect 9355 9880 10876 9908
rect 9355 9877 9367 9880
rect 9309 9871 9367 9877
rect 10870 9868 10876 9880
rect 10928 9868 10934 9920
rect 920 9818 9844 9840
rect 920 9766 4116 9818
rect 4168 9766 4180 9818
rect 4232 9766 4244 9818
rect 4296 9766 4308 9818
rect 4360 9766 4372 9818
rect 4424 9766 7216 9818
rect 7268 9766 7280 9818
rect 7332 9766 7344 9818
rect 7396 9766 7408 9818
rect 7460 9766 7472 9818
rect 7524 9766 9844 9818
rect 920 9744 9844 9766
rect 1857 9707 1915 9713
rect 1857 9673 1869 9707
rect 1903 9704 1915 9707
rect 2958 9704 2964 9716
rect 1903 9676 1937 9704
rect 2608 9676 2964 9704
rect 1903 9673 1915 9676
rect 1857 9667 1915 9673
rect 1302 9636 1308 9648
rect 1263 9608 1308 9636
rect 1302 9596 1308 9608
rect 1360 9596 1366 9648
rect 1872 9636 1900 9667
rect 2608 9636 2636 9676
rect 2958 9664 2964 9676
rect 3016 9664 3022 9716
rect 3142 9664 3148 9716
rect 3200 9704 3206 9716
rect 3200 9676 4384 9704
rect 3200 9664 3206 9676
rect 1872 9608 2636 9636
rect 2682 9596 2688 9648
rect 2740 9636 2746 9648
rect 2740 9608 2820 9636
rect 2740 9596 2746 9608
rect 1026 9528 1032 9580
rect 1084 9568 1090 9580
rect 1397 9571 1455 9577
rect 1397 9568 1409 9571
rect 1084 9540 1409 9568
rect 1084 9528 1090 9540
rect 1397 9537 1409 9540
rect 1443 9568 1455 9571
rect 1681 9575 1739 9581
rect 1443 9540 1624 9568
rect 1443 9537 1455 9540
rect 1397 9531 1455 9537
rect 1596 9500 1624 9540
rect 1681 9541 1693 9575
rect 1727 9572 1739 9575
rect 1727 9568 1808 9572
rect 1854 9568 1860 9580
rect 1727 9544 1860 9568
rect 1727 9541 1739 9544
rect 1681 9535 1739 9541
rect 1780 9540 1860 9544
rect 1854 9528 1860 9540
rect 1912 9528 1918 9580
rect 1949 9571 2007 9577
rect 1949 9537 1961 9571
rect 1995 9568 2007 9571
rect 2038 9568 2044 9580
rect 1995 9540 2044 9568
rect 1995 9537 2007 9540
rect 1949 9531 2007 9537
rect 2038 9528 2044 9540
rect 2096 9528 2102 9580
rect 2130 9528 2136 9580
rect 2188 9528 2194 9580
rect 2225 9571 2283 9577
rect 2225 9537 2237 9571
rect 2271 9537 2283 9571
rect 2225 9531 2283 9537
rect 2148 9500 2176 9528
rect 1596 9472 2176 9500
rect 1670 9392 1676 9444
rect 1728 9432 1734 9444
rect 2133 9435 2191 9441
rect 2133 9432 2145 9435
rect 1728 9404 2145 9432
rect 1728 9392 1734 9404
rect 2133 9401 2145 9404
rect 2179 9401 2191 9435
rect 2133 9395 2191 9401
rect 1581 9367 1639 9373
rect 1581 9333 1593 9367
rect 1627 9364 1639 9367
rect 2038 9364 2044 9376
rect 1627 9336 2044 9364
rect 1627 9333 1639 9336
rect 1581 9327 1639 9333
rect 2038 9324 2044 9336
rect 2096 9324 2102 9376
rect 2240 9364 2268 9531
rect 2590 9528 2596 9580
rect 2648 9568 2654 9580
rect 2792 9568 2820 9608
rect 3418 9596 3424 9648
rect 3476 9636 3482 9648
rect 4356 9636 4384 9676
rect 5258 9664 5264 9716
rect 5316 9704 5322 9716
rect 8018 9704 8024 9716
rect 5316 9676 8024 9704
rect 5316 9664 5322 9676
rect 8018 9664 8024 9676
rect 8076 9664 8082 9716
rect 6181 9639 6239 9645
rect 6181 9636 6193 9639
rect 3476 9608 3542 9636
rect 4356 9608 6193 9636
rect 3476 9596 3482 9608
rect 6181 9605 6193 9608
rect 6227 9605 6239 9639
rect 6181 9599 6239 9605
rect 8478 9596 8484 9648
rect 8536 9596 8542 9648
rect 8846 9596 8852 9648
rect 8904 9636 8910 9648
rect 9398 9636 9404 9648
rect 8904 9608 9404 9636
rect 8904 9596 8910 9608
rect 9398 9596 9404 9608
rect 9456 9596 9462 9648
rect 3145 9571 3203 9577
rect 3145 9568 3157 9571
rect 2648 9561 2728 9568
rect 2648 9555 2743 9561
rect 2648 9540 2697 9555
rect 2648 9528 2654 9540
rect 2685 9521 2697 9540
rect 2731 9521 2743 9555
rect 2792 9540 3157 9568
rect 3145 9537 3157 9540
rect 3191 9537 3203 9571
rect 4614 9568 4620 9580
rect 4575 9540 4620 9568
rect 3145 9531 3203 9537
rect 4614 9528 4620 9540
rect 4672 9528 4678 9580
rect 4890 9528 4896 9580
rect 4948 9568 4954 9580
rect 5353 9571 5411 9577
rect 5353 9568 5365 9571
rect 4948 9540 5365 9568
rect 4948 9528 4954 9540
rect 5353 9537 5365 9540
rect 5399 9537 5411 9571
rect 5629 9571 5687 9577
rect 5629 9568 5641 9571
rect 5353 9531 5411 9537
rect 5460 9540 5641 9568
rect 2685 9515 2743 9521
rect 2777 9503 2835 9509
rect 2777 9469 2789 9503
rect 2823 9469 2835 9503
rect 2777 9463 2835 9469
rect 2409 9435 2467 9441
rect 2409 9401 2421 9435
rect 2455 9432 2467 9435
rect 2792 9432 2820 9463
rect 4706 9460 4712 9512
rect 4764 9500 4770 9512
rect 5460 9500 5488 9540
rect 5629 9537 5641 9540
rect 5675 9537 5687 9571
rect 5994 9568 6000 9580
rect 5955 9540 6000 9568
rect 5629 9531 5687 9537
rect 5994 9528 6000 9540
rect 6052 9528 6058 9580
rect 6822 9568 6828 9580
rect 6783 9540 6828 9568
rect 6822 9528 6828 9540
rect 6880 9528 6886 9580
rect 6917 9571 6975 9577
rect 6917 9537 6929 9571
rect 6963 9537 6975 9571
rect 6917 9531 6975 9537
rect 4764 9472 5488 9500
rect 4764 9460 4770 9472
rect 5718 9460 5724 9512
rect 5776 9500 5782 9512
rect 6932 9500 6960 9531
rect 7006 9528 7012 9580
rect 7064 9568 7070 9580
rect 7193 9571 7251 9577
rect 7193 9568 7205 9571
rect 7064 9540 7205 9568
rect 7064 9528 7070 9540
rect 7193 9537 7205 9540
rect 7239 9537 7251 9571
rect 7650 9568 7656 9580
rect 7193 9531 7251 9537
rect 7300 9540 7656 9568
rect 5776 9472 6960 9500
rect 5776 9460 5782 9472
rect 5169 9435 5227 9441
rect 5169 9432 5181 9435
rect 2455 9404 2820 9432
rect 4080 9404 5181 9432
rect 2455 9401 2467 9404
rect 2409 9395 2467 9401
rect 2501 9367 2559 9373
rect 2501 9364 2513 9367
rect 2240 9336 2513 9364
rect 2501 9333 2513 9336
rect 2547 9333 2559 9367
rect 2501 9327 2559 9333
rect 3878 9324 3884 9376
rect 3936 9364 3942 9376
rect 4080 9364 4108 9404
rect 5169 9401 5181 9404
rect 5215 9401 5227 9435
rect 5169 9395 5227 9401
rect 5258 9392 5264 9444
rect 5316 9432 5322 9444
rect 5445 9435 5503 9441
rect 5445 9432 5457 9435
rect 5316 9404 5457 9432
rect 5316 9392 5322 9404
rect 5445 9401 5457 9404
rect 5491 9401 5503 9435
rect 5445 9395 5503 9401
rect 5534 9392 5540 9444
rect 5592 9432 5598 9444
rect 5813 9435 5871 9441
rect 5813 9432 5825 9435
rect 5592 9404 5825 9432
rect 5592 9392 5598 9404
rect 5813 9401 5825 9404
rect 5859 9401 5871 9435
rect 5813 9395 5871 9401
rect 7009 9435 7067 9441
rect 7009 9401 7021 9435
rect 7055 9432 7067 9435
rect 7300 9432 7328 9540
rect 7650 9528 7656 9540
rect 7708 9528 7714 9580
rect 9033 9571 9091 9577
rect 9033 9537 9045 9571
rect 9079 9537 9091 9571
rect 9033 9531 9091 9537
rect 7558 9500 7564 9512
rect 7519 9472 7564 9500
rect 7558 9460 7564 9472
rect 7616 9460 7622 9512
rect 7055 9404 7328 9432
rect 7055 9401 7067 9404
rect 7009 9395 7067 9401
rect 8478 9392 8484 9444
rect 8536 9432 8542 9444
rect 9048 9432 9076 9531
rect 8536 9404 9076 9432
rect 8536 9392 8542 9404
rect 3936 9336 4108 9364
rect 5077 9367 5135 9373
rect 3936 9324 3942 9336
rect 5077 9333 5089 9367
rect 5123 9364 5135 9367
rect 6362 9364 6368 9376
rect 5123 9336 6368 9364
rect 5123 9333 5135 9336
rect 5077 9327 5135 9333
rect 6362 9324 6368 9336
rect 6420 9324 6426 9376
rect 7190 9324 7196 9376
rect 7248 9364 7254 9376
rect 9493 9367 9551 9373
rect 9493 9364 9505 9367
rect 7248 9336 9505 9364
rect 7248 9324 7254 9336
rect 9493 9333 9505 9336
rect 9539 9333 9551 9367
rect 9493 9327 9551 9333
rect 920 9274 9844 9296
rect 920 9222 2566 9274
rect 2618 9222 2630 9274
rect 2682 9222 2694 9274
rect 2746 9222 2758 9274
rect 2810 9222 2822 9274
rect 2874 9222 5666 9274
rect 5718 9222 5730 9274
rect 5782 9222 5794 9274
rect 5846 9222 5858 9274
rect 5910 9222 5922 9274
rect 5974 9222 8766 9274
rect 8818 9222 8830 9274
rect 8882 9222 8894 9274
rect 8946 9222 8958 9274
rect 9010 9222 9022 9274
rect 9074 9222 9844 9274
rect 920 9200 9844 9222
rect 1210 9160 1216 9172
rect 1171 9132 1216 9160
rect 1210 9120 1216 9132
rect 1268 9120 1274 9172
rect 1857 9163 1915 9169
rect 1857 9129 1869 9163
rect 1903 9160 1915 9163
rect 3142 9160 3148 9172
rect 1903 9132 3148 9160
rect 1903 9129 1915 9132
rect 1857 9123 1915 9129
rect 3142 9120 3148 9132
rect 3200 9120 3206 9172
rect 3418 9160 3424 9172
rect 3379 9132 3424 9160
rect 3418 9120 3424 9132
rect 3476 9120 3482 9172
rect 3789 9163 3847 9169
rect 3789 9129 3801 9163
rect 3835 9160 3847 9163
rect 4338 9160 4344 9172
rect 3835 9132 4344 9160
rect 3835 9129 3847 9132
rect 3789 9123 3847 9129
rect 4338 9120 4344 9132
rect 4396 9120 4402 9172
rect 4614 9160 4620 9172
rect 4575 9132 4620 9160
rect 4614 9120 4620 9132
rect 4672 9120 4678 9172
rect 7190 9160 7196 9172
rect 5276 9132 7196 9160
rect 1581 9095 1639 9101
rect 1581 9061 1593 9095
rect 1627 9092 1639 9095
rect 3602 9092 3608 9104
rect 1627 9064 3608 9092
rect 1627 9061 1639 9064
rect 1581 9055 1639 9061
rect 3602 9052 3608 9064
rect 3660 9052 3666 9104
rect 4430 9092 4436 9104
rect 3988 9064 4436 9092
rect 2314 9024 2320 9036
rect 1412 8996 2320 9024
rect 1412 8965 1440 8996
rect 2314 8984 2320 8996
rect 2372 8984 2378 9036
rect 3988 9024 4016 9064
rect 4430 9052 4436 9064
rect 4488 9052 4494 9104
rect 4525 9095 4583 9101
rect 4525 9061 4537 9095
rect 4571 9092 4583 9095
rect 4706 9092 4712 9104
rect 4571 9064 4712 9092
rect 4571 9061 4583 9064
rect 4525 9055 4583 9061
rect 4706 9052 4712 9064
rect 4764 9052 4770 9104
rect 2884 8996 4016 9024
rect 4065 9027 4123 9033
rect 1397 8959 1455 8965
rect 1397 8925 1409 8959
rect 1443 8925 1455 8959
rect 1673 8959 1731 8965
rect 1673 8956 1685 8959
rect 1397 8919 1455 8925
rect 1504 8928 1685 8956
rect 1118 8848 1124 8900
rect 1176 8888 1182 8900
rect 1504 8888 1532 8928
rect 1673 8925 1685 8928
rect 1719 8925 1731 8959
rect 1946 8956 1952 8968
rect 1907 8928 1952 8956
rect 1673 8919 1731 8925
rect 1946 8916 1952 8928
rect 2004 8916 2010 8968
rect 2130 8956 2136 8968
rect 2091 8928 2136 8956
rect 2130 8916 2136 8928
rect 2188 8916 2194 8968
rect 2406 8956 2412 8968
rect 2367 8928 2412 8956
rect 2406 8916 2412 8928
rect 2464 8916 2470 8968
rect 2685 8959 2743 8965
rect 2685 8956 2697 8959
rect 2516 8928 2697 8956
rect 1176 8860 1532 8888
rect 1176 8848 1182 8860
rect 1578 8848 1584 8900
rect 1636 8888 1642 8900
rect 2516 8888 2544 8928
rect 2685 8925 2697 8928
rect 2731 8925 2743 8959
rect 2884 8956 2912 8996
rect 4065 8993 4077 9027
rect 4111 9024 4123 9027
rect 4890 9024 4896 9036
rect 4111 8996 4896 9024
rect 4111 8993 4123 8996
rect 4065 8987 4123 8993
rect 4890 8984 4896 8996
rect 4948 8984 4954 9036
rect 2685 8919 2743 8925
rect 2792 8928 2912 8956
rect 2961 8959 3019 8965
rect 1636 8860 2544 8888
rect 1636 8848 1642 8860
rect 2317 8823 2375 8829
rect 2317 8789 2329 8823
rect 2363 8820 2375 8823
rect 2406 8820 2412 8832
rect 2363 8792 2412 8820
rect 2363 8789 2375 8792
rect 2317 8783 2375 8789
rect 2406 8780 2412 8792
rect 2464 8780 2470 8832
rect 2593 8823 2651 8829
rect 2593 8789 2605 8823
rect 2639 8820 2651 8823
rect 2792 8820 2820 8928
rect 2961 8925 2973 8959
rect 3007 8956 3019 8959
rect 3050 8956 3056 8968
rect 3007 8928 3056 8956
rect 3007 8925 3019 8928
rect 2961 8919 3019 8925
rect 3050 8916 3056 8928
rect 3108 8916 3114 8968
rect 3234 8956 3240 8968
rect 3195 8928 3240 8956
rect 3234 8916 3240 8928
rect 3292 8916 3298 8968
rect 3418 8916 3424 8968
rect 3476 8956 3482 8968
rect 3605 8959 3663 8965
rect 3605 8956 3617 8959
rect 3476 8928 3617 8956
rect 3476 8916 3482 8928
rect 3605 8925 3617 8928
rect 3651 8925 3663 8959
rect 3605 8919 3663 8925
rect 3620 8888 3648 8919
rect 3786 8916 3792 8968
rect 3844 8956 3850 8968
rect 5276 8965 5304 9132
rect 7190 9120 7196 9132
rect 7248 9120 7254 9172
rect 9125 9163 9183 9169
rect 9125 9129 9137 9163
rect 9171 9160 9183 9163
rect 9306 9160 9312 9172
rect 9171 9132 9312 9160
rect 9171 9129 9183 9132
rect 9125 9123 9183 9129
rect 9306 9120 9312 9132
rect 9364 9120 9370 9172
rect 13814 9120 13820 9172
rect 13872 9160 13878 9172
rect 16666 9160 16672 9172
rect 13872 9132 16672 9160
rect 13872 9120 13878 9132
rect 16666 9120 16672 9132
rect 16724 9120 16730 9172
rect 8754 9052 8760 9104
rect 8812 9092 8818 9104
rect 9398 9092 9404 9104
rect 8812 9064 9404 9092
rect 8812 9052 8818 9064
rect 9398 9052 9404 9064
rect 9456 9052 9462 9104
rect 5353 9027 5411 9033
rect 5353 8993 5365 9027
rect 5399 9024 5411 9027
rect 6822 9024 6828 9036
rect 5399 8996 6828 9024
rect 5399 8993 5411 8996
rect 5353 8987 5411 8993
rect 6822 8984 6828 8996
rect 6880 9024 6886 9036
rect 7098 9024 7104 9036
rect 6880 8996 7104 9024
rect 6880 8984 6886 8996
rect 7098 8984 7104 8996
rect 7156 8984 7162 9036
rect 4801 8959 4859 8965
rect 4801 8956 4813 8959
rect 3844 8928 4813 8956
rect 3844 8916 3850 8928
rect 4801 8925 4813 8928
rect 4847 8925 4859 8959
rect 4801 8919 4859 8925
rect 5261 8959 5319 8965
rect 5261 8925 5273 8959
rect 5307 8925 5319 8959
rect 8110 8956 8116 8968
rect 5261 8919 5319 8925
rect 7024 8928 8116 8956
rect 4157 8891 4215 8897
rect 4157 8888 4169 8891
rect 3620 8860 4169 8888
rect 4157 8857 4169 8860
rect 4203 8857 4215 8891
rect 4338 8888 4344 8900
rect 4299 8860 4344 8888
rect 4157 8851 4215 8857
rect 4338 8848 4344 8860
rect 4396 8848 4402 8900
rect 4430 8848 4436 8900
rect 4488 8888 4494 8900
rect 5629 8891 5687 8897
rect 4488 8860 5396 8888
rect 4488 8848 4494 8860
rect 2639 8792 2820 8820
rect 2869 8823 2927 8829
rect 2639 8789 2651 8792
rect 2593 8783 2651 8789
rect 2869 8789 2881 8823
rect 2915 8820 2927 8823
rect 3050 8820 3056 8832
rect 2915 8792 3056 8820
rect 2915 8789 2927 8792
rect 2869 8783 2927 8789
rect 3050 8780 3056 8792
rect 3108 8780 3114 8832
rect 3145 8823 3203 8829
rect 3145 8789 3157 8823
rect 3191 8820 3203 8823
rect 4982 8820 4988 8832
rect 3191 8792 4988 8820
rect 3191 8789 3203 8792
rect 3145 8783 3203 8789
rect 4982 8780 4988 8792
rect 5040 8780 5046 8832
rect 5074 8780 5080 8832
rect 5132 8820 5138 8832
rect 5368 8820 5396 8860
rect 5629 8857 5641 8891
rect 5675 8888 5687 8891
rect 5902 8888 5908 8900
rect 5675 8860 5908 8888
rect 5675 8857 5687 8860
rect 5629 8851 5687 8857
rect 5902 8848 5908 8860
rect 5960 8848 5966 8900
rect 6638 8848 6644 8900
rect 6696 8848 6702 8900
rect 7024 8820 7052 8928
rect 8110 8916 8116 8928
rect 8168 8916 8174 8968
rect 8570 8956 8576 8968
rect 8483 8928 8576 8956
rect 8570 8916 8576 8928
rect 8628 8956 8634 8968
rect 9214 8956 9220 8968
rect 8628 8928 9076 8956
rect 9175 8928 9220 8956
rect 8628 8916 8634 8928
rect 7190 8888 7196 8900
rect 7116 8860 7196 8888
rect 7116 8829 7144 8860
rect 7190 8848 7196 8860
rect 7248 8888 7254 8900
rect 7558 8888 7564 8900
rect 7248 8860 7564 8888
rect 7248 8848 7254 8860
rect 7558 8848 7564 8860
rect 7616 8848 7622 8900
rect 7653 8891 7711 8897
rect 7653 8857 7665 8891
rect 7699 8888 7711 8891
rect 7742 8888 7748 8900
rect 7699 8860 7748 8888
rect 7699 8857 7711 8860
rect 7653 8851 7711 8857
rect 7742 8848 7748 8860
rect 7800 8888 7806 8900
rect 8754 8888 8760 8900
rect 7800 8860 8294 8888
rect 8715 8860 8760 8888
rect 7800 8848 7806 8860
rect 5132 8792 5177 8820
rect 5368 8792 7052 8820
rect 7101 8823 7159 8829
rect 5132 8780 5138 8792
rect 7101 8789 7113 8823
rect 7147 8789 7159 8823
rect 8266 8820 8294 8860
rect 8754 8848 8760 8860
rect 8812 8848 8818 8900
rect 8941 8891 8999 8897
rect 8941 8857 8953 8891
rect 8987 8857 8999 8891
rect 9048 8888 9076 8928
rect 9214 8916 9220 8928
rect 9272 8916 9278 8968
rect 9306 8888 9312 8900
rect 9048 8860 9312 8888
rect 8941 8851 8999 8857
rect 8956 8820 8984 8851
rect 9306 8848 9312 8860
rect 9364 8848 9370 8900
rect 9398 8820 9404 8832
rect 8266 8792 8984 8820
rect 9359 8792 9404 8820
rect 7101 8783 7159 8789
rect 9398 8780 9404 8792
rect 9456 8780 9462 8832
rect 920 8730 9844 8752
rect 920 8678 4116 8730
rect 4168 8678 4180 8730
rect 4232 8678 4244 8730
rect 4296 8678 4308 8730
rect 4360 8678 4372 8730
rect 4424 8678 7216 8730
rect 7268 8678 7280 8730
rect 7332 8678 7344 8730
rect 7396 8678 7408 8730
rect 7460 8678 7472 8730
rect 7524 8678 9844 8730
rect 920 8656 9844 8678
rect 1210 8616 1216 8628
rect 1171 8588 1216 8616
rect 1210 8576 1216 8588
rect 1268 8576 1274 8628
rect 1302 8576 1308 8628
rect 1360 8616 1366 8628
rect 1397 8619 1455 8625
rect 1397 8616 1409 8619
rect 1360 8588 1409 8616
rect 1360 8576 1366 8588
rect 1397 8585 1409 8588
rect 1443 8585 1455 8619
rect 7834 8616 7840 8628
rect 1397 8579 1455 8585
rect 1780 8588 7840 8616
rect 1780 8489 1808 8588
rect 7834 8576 7840 8588
rect 7892 8576 7898 8628
rect 9490 8616 9496 8628
rect 9451 8588 9496 8616
rect 9490 8576 9496 8588
rect 9548 8576 9554 8628
rect 2222 8508 2228 8560
rect 2280 8548 2286 8560
rect 2593 8551 2651 8557
rect 2593 8548 2605 8551
rect 2280 8520 2605 8548
rect 2280 8508 2286 8520
rect 2593 8517 2605 8520
rect 2639 8517 2651 8551
rect 4522 8548 4528 8560
rect 2593 8511 2651 8517
rect 4172 8520 4528 8548
rect 4172 8492 4200 8520
rect 4522 8508 4528 8520
rect 4580 8508 4586 8560
rect 5718 8508 5724 8560
rect 5776 8548 5782 8560
rect 6181 8551 6239 8557
rect 6181 8548 6193 8551
rect 5776 8520 6193 8548
rect 5776 8508 5782 8520
rect 6181 8517 6193 8520
rect 6227 8517 6239 8551
rect 6730 8548 6736 8560
rect 6691 8520 6736 8548
rect 6181 8511 6239 8517
rect 6730 8508 6736 8520
rect 6788 8508 6794 8560
rect 6822 8508 6828 8560
rect 6880 8548 6886 8560
rect 7101 8551 7159 8557
rect 7101 8548 7113 8551
rect 6880 8520 7113 8548
rect 6880 8508 6886 8520
rect 7101 8517 7113 8520
rect 7147 8517 7159 8551
rect 7101 8511 7159 8517
rect 8018 8508 8024 8560
rect 8076 8508 8082 8560
rect 1765 8483 1823 8489
rect 1765 8449 1777 8483
rect 1811 8449 1823 8483
rect 2038 8480 2044 8492
rect 1999 8452 2044 8480
rect 1765 8443 1823 8449
rect 2038 8440 2044 8452
rect 2096 8440 2102 8492
rect 4154 8480 4160 8492
rect 3726 8452 3832 8480
rect 4067 8452 4160 8480
rect 3804 8424 3832 8452
rect 4154 8440 4160 8452
rect 4212 8440 4218 8492
rect 5534 8440 5540 8492
rect 5592 8480 5598 8492
rect 6365 8483 6423 8489
rect 6365 8480 6377 8483
rect 5592 8452 6377 8480
rect 5592 8440 5598 8452
rect 6365 8449 6377 8452
rect 6411 8480 6423 8483
rect 6638 8480 6644 8492
rect 6411 8452 6644 8480
rect 6411 8449 6423 8452
rect 6365 8443 6423 8449
rect 6638 8440 6644 8452
rect 6696 8440 6702 8492
rect 6917 8483 6975 8489
rect 6917 8449 6929 8483
rect 6963 8449 6975 8483
rect 6917 8443 6975 8449
rect 9033 8483 9091 8489
rect 9033 8449 9045 8483
rect 9079 8480 9091 8483
rect 9122 8480 9128 8492
rect 9079 8452 9128 8480
rect 9079 8449 9091 8452
rect 9033 8443 9091 8449
rect 1673 8415 1731 8421
rect 1673 8381 1685 8415
rect 1719 8412 1731 8415
rect 2130 8412 2136 8424
rect 1719 8384 2136 8412
rect 1719 8381 1731 8384
rect 1673 8375 1731 8381
rect 2130 8372 2136 8384
rect 2188 8372 2194 8424
rect 2314 8412 2320 8424
rect 2275 8384 2320 8412
rect 2314 8372 2320 8384
rect 2372 8372 2378 8424
rect 3786 8372 3792 8424
rect 3844 8372 3850 8424
rect 3970 8372 3976 8424
rect 4028 8412 4034 8424
rect 4065 8415 4123 8421
rect 4065 8412 4077 8415
rect 4028 8384 4077 8412
rect 4028 8372 4034 8384
rect 4065 8381 4077 8384
rect 4111 8381 4123 8415
rect 4065 8375 4123 8381
rect 4433 8415 4491 8421
rect 4433 8381 4445 8415
rect 4479 8412 4491 8415
rect 4522 8412 4528 8424
rect 4479 8384 4528 8412
rect 4479 8381 4491 8384
rect 4433 8375 4491 8381
rect 4522 8372 4528 8384
rect 4580 8372 4586 8424
rect 4798 8372 4804 8424
rect 4856 8412 4862 8424
rect 6932 8412 6960 8443
rect 9122 8440 9128 8452
rect 9180 8440 9186 8492
rect 4856 8384 6960 8412
rect 7193 8415 7251 8421
rect 4856 8372 4862 8384
rect 7193 8381 7205 8415
rect 7239 8381 7251 8415
rect 7558 8412 7564 8424
rect 7519 8384 7564 8412
rect 7193 8375 7251 8381
rect 1946 8344 1952 8356
rect 1907 8316 1952 8344
rect 1946 8304 1952 8316
rect 2004 8304 2010 8356
rect 5534 8304 5540 8356
rect 5592 8344 5598 8356
rect 5902 8344 5908 8356
rect 5592 8316 5908 8344
rect 5592 8304 5598 8316
rect 5902 8304 5908 8316
rect 5960 8304 5966 8356
rect 6380 8316 6684 8344
rect 1302 8236 1308 8288
rect 1360 8276 1366 8288
rect 1854 8276 1860 8288
rect 1360 8248 1860 8276
rect 1360 8236 1366 8248
rect 1854 8236 1860 8248
rect 1912 8236 1918 8288
rect 2222 8276 2228 8288
rect 2183 8248 2228 8276
rect 2222 8236 2228 8248
rect 2280 8236 2286 8288
rect 2406 8236 2412 8288
rect 2464 8276 2470 8288
rect 6380 8276 6408 8316
rect 6546 8276 6552 8288
rect 2464 8248 6408 8276
rect 6507 8248 6552 8276
rect 2464 8236 2470 8248
rect 6546 8236 6552 8248
rect 6604 8236 6610 8288
rect 6656 8276 6684 8316
rect 6914 8304 6920 8356
rect 6972 8344 6978 8356
rect 7208 8344 7236 8375
rect 7558 8372 7564 8384
rect 7616 8372 7622 8424
rect 6972 8316 7236 8344
rect 6972 8304 6978 8316
rect 9122 8276 9128 8288
rect 6656 8248 9128 8276
rect 9122 8236 9128 8248
rect 9180 8236 9186 8288
rect 920 8186 9844 8208
rect 920 8134 2566 8186
rect 2618 8134 2630 8186
rect 2682 8134 2694 8186
rect 2746 8134 2758 8186
rect 2810 8134 2822 8186
rect 2874 8134 5666 8186
rect 5718 8134 5730 8186
rect 5782 8134 5794 8186
rect 5846 8134 5858 8186
rect 5910 8134 5922 8186
rect 5974 8134 8766 8186
rect 8818 8134 8830 8186
rect 8882 8134 8894 8186
rect 8946 8134 8958 8186
rect 9010 8134 9022 8186
rect 9074 8134 9844 8186
rect 920 8112 9844 8134
rect 1412 8044 3372 8072
rect 1412 7877 1440 8044
rect 1578 8004 1584 8016
rect 1539 7976 1584 8004
rect 1578 7964 1584 7976
rect 1636 7964 1642 8016
rect 3344 8004 3372 8044
rect 3418 8032 3424 8084
rect 3476 8072 3482 8084
rect 3973 8075 4031 8081
rect 3476 8044 3924 8072
rect 3476 8032 3482 8044
rect 3786 8004 3792 8016
rect 3344 7976 3792 8004
rect 3786 7964 3792 7976
rect 3844 7964 3850 8016
rect 3896 8004 3924 8044
rect 3973 8041 3985 8075
rect 4019 8072 4031 8075
rect 4062 8072 4068 8084
rect 4019 8044 4068 8072
rect 4019 8041 4031 8044
rect 3973 8035 4031 8041
rect 4062 8032 4068 8044
rect 4120 8032 4126 8084
rect 5166 8032 5172 8084
rect 5224 8072 5230 8084
rect 8757 8075 8815 8081
rect 8757 8072 8769 8075
rect 5224 8044 8769 8072
rect 5224 8032 5230 8044
rect 8757 8041 8769 8044
rect 8803 8041 8815 8075
rect 8757 8035 8815 8041
rect 3896 7976 5212 8004
rect 2406 7896 2412 7948
rect 2464 7936 2470 7948
rect 3421 7939 3479 7945
rect 3421 7936 3433 7939
rect 2464 7908 3433 7936
rect 2464 7896 2470 7908
rect 3421 7905 3433 7908
rect 3467 7936 3479 7939
rect 4154 7936 4160 7948
rect 3467 7908 4160 7936
rect 3467 7905 3479 7908
rect 3421 7899 3479 7905
rect 4154 7896 4160 7908
rect 4212 7896 4218 7948
rect 5184 7945 5212 7976
rect 6546 7964 6552 8016
rect 6604 8004 6610 8016
rect 8110 8004 8116 8016
rect 6604 7976 8116 8004
rect 6604 7964 6610 7976
rect 8110 7964 8116 7976
rect 8168 7964 8174 8016
rect 9582 8004 9588 8016
rect 8220 7976 9588 8004
rect 5169 7939 5227 7945
rect 5169 7905 5181 7939
rect 5215 7905 5227 7939
rect 5534 7936 5540 7948
rect 5495 7908 5540 7936
rect 5169 7899 5227 7905
rect 5534 7896 5540 7908
rect 5592 7896 5598 7948
rect 5994 7936 6000 7948
rect 5644 7908 6000 7936
rect 1397 7871 1455 7877
rect 1397 7837 1409 7871
rect 1443 7837 1455 7871
rect 1397 7831 1455 7837
rect 3510 7828 3516 7880
rect 3568 7868 3574 7880
rect 3697 7871 3755 7877
rect 3697 7868 3709 7871
rect 3568 7840 3709 7868
rect 3568 7828 3574 7840
rect 3697 7837 3709 7840
rect 3743 7837 3755 7871
rect 3697 7831 3755 7837
rect 3786 7828 3792 7880
rect 3844 7868 3850 7880
rect 4249 7871 4307 7877
rect 4249 7868 4261 7871
rect 3844 7840 4261 7868
rect 3844 7828 3850 7840
rect 4249 7837 4261 7840
rect 4295 7837 4307 7871
rect 4249 7831 4307 7837
rect 4525 7871 4583 7877
rect 4525 7837 4537 7871
rect 4571 7868 4583 7871
rect 5644 7868 5672 7908
rect 5994 7896 6000 7908
rect 6052 7896 6058 7948
rect 7469 7939 7527 7945
rect 7469 7905 7481 7939
rect 7515 7936 7527 7939
rect 8220 7936 8248 7976
rect 9582 7964 9588 7976
rect 9640 7964 9646 8016
rect 7515 7908 8248 7936
rect 8312 7908 9260 7936
rect 7515 7905 7527 7908
rect 7469 7899 7527 7905
rect 4571 7840 5672 7868
rect 7009 7871 7067 7877
rect 4571 7837 4583 7840
rect 4525 7831 4583 7837
rect 7009 7837 7021 7871
rect 7055 7868 7067 7871
rect 8202 7868 8208 7880
rect 7055 7840 8064 7868
rect 8163 7840 8208 7868
rect 7055 7837 7067 7840
rect 7009 7831 7067 7837
rect 1305 7803 1363 7809
rect 1305 7769 1317 7803
rect 1351 7800 1363 7803
rect 1486 7800 1492 7812
rect 1351 7772 1492 7800
rect 1351 7769 1363 7772
rect 1305 7763 1363 7769
rect 1486 7760 1492 7772
rect 1544 7760 1550 7812
rect 2682 7760 2688 7812
rect 2740 7760 2746 7812
rect 3145 7803 3203 7809
rect 3145 7769 3157 7803
rect 3191 7800 3203 7803
rect 3970 7800 3976 7812
rect 3191 7772 3976 7800
rect 3191 7769 3203 7772
rect 3145 7763 3203 7769
rect 3970 7760 3976 7772
rect 4028 7760 4034 7812
rect 5166 7800 5172 7812
rect 4080 7772 5172 7800
rect 1670 7732 1676 7744
rect 1631 7704 1676 7732
rect 1670 7692 1676 7704
rect 1728 7692 1734 7744
rect 1854 7692 1860 7744
rect 1912 7732 1918 7744
rect 4080 7732 4108 7772
rect 5166 7760 5172 7772
rect 5224 7760 5230 7812
rect 6270 7760 6276 7812
rect 6328 7760 6334 7812
rect 6914 7760 6920 7812
rect 6972 7800 6978 7812
rect 7561 7803 7619 7809
rect 7561 7800 7573 7803
rect 6972 7772 7573 7800
rect 6972 7760 6978 7772
rect 7561 7769 7573 7772
rect 7607 7769 7619 7803
rect 7742 7800 7748 7812
rect 7703 7772 7748 7800
rect 7561 7763 7619 7769
rect 7742 7760 7748 7772
rect 7800 7760 7806 7812
rect 1912 7704 4108 7732
rect 4157 7735 4215 7741
rect 1912 7692 1918 7704
rect 4157 7701 4169 7735
rect 4203 7732 4215 7735
rect 6178 7732 6184 7744
rect 4203 7704 6184 7732
rect 4203 7701 4215 7704
rect 4157 7695 4215 7701
rect 6178 7692 6184 7704
rect 6236 7692 6242 7744
rect 6362 7692 6368 7744
rect 6420 7732 6426 7744
rect 7650 7732 7656 7744
rect 6420 7704 7656 7732
rect 6420 7692 6426 7704
rect 7650 7692 7656 7704
rect 7708 7692 7714 7744
rect 7926 7732 7932 7744
rect 7887 7704 7932 7732
rect 7926 7692 7932 7704
rect 7984 7692 7990 7744
rect 8036 7741 8064 7840
rect 8202 7828 8208 7840
rect 8260 7828 8266 7880
rect 8110 7760 8116 7812
rect 8168 7800 8174 7812
rect 8312 7800 8340 7908
rect 8570 7868 8576 7880
rect 8531 7840 8576 7868
rect 8570 7828 8576 7840
rect 8628 7828 8634 7880
rect 8941 7871 8999 7877
rect 8941 7837 8953 7871
rect 8987 7837 8999 7871
rect 8941 7831 8999 7837
rect 8168 7772 8340 7800
rect 8168 7760 8174 7772
rect 8478 7760 8484 7812
rect 8536 7800 8542 7812
rect 8956 7800 8984 7831
rect 9030 7828 9036 7880
rect 9088 7868 9094 7880
rect 9232 7877 9260 7908
rect 9217 7871 9275 7877
rect 9088 7840 9133 7868
rect 9088 7828 9094 7840
rect 9217 7837 9229 7871
rect 9263 7837 9275 7871
rect 9217 7831 9275 7837
rect 8536 7772 8984 7800
rect 8536 7760 8542 7772
rect 8021 7735 8079 7741
rect 8021 7701 8033 7735
rect 8067 7701 8079 7735
rect 8386 7732 8392 7744
rect 8347 7704 8392 7732
rect 8021 7695 8079 7701
rect 8386 7692 8392 7704
rect 8444 7692 8450 7744
rect 9401 7735 9459 7741
rect 9401 7701 9413 7735
rect 9447 7732 9459 7735
rect 12250 7732 12256 7744
rect 9447 7704 12256 7732
rect 9447 7701 9459 7704
rect 9401 7695 9459 7701
rect 12250 7692 12256 7704
rect 12308 7692 12314 7744
rect 920 7642 9844 7664
rect 920 7590 4116 7642
rect 4168 7590 4180 7642
rect 4232 7590 4244 7642
rect 4296 7590 4308 7642
rect 4360 7590 4372 7642
rect 4424 7590 7216 7642
rect 7268 7590 7280 7642
rect 7332 7590 7344 7642
rect 7396 7590 7408 7642
rect 7460 7590 7472 7642
rect 7524 7590 9844 7642
rect 920 7568 9844 7590
rect 1302 7528 1308 7540
rect 1263 7500 1308 7528
rect 1302 7488 1308 7500
rect 1360 7488 1366 7540
rect 1857 7531 1915 7537
rect 1857 7497 1869 7531
rect 1903 7528 1915 7531
rect 2038 7528 2044 7540
rect 1903 7500 2044 7528
rect 1903 7497 1915 7500
rect 1857 7491 1915 7497
rect 2038 7488 2044 7500
rect 2096 7488 2102 7540
rect 2314 7528 2320 7540
rect 2275 7500 2320 7528
rect 2314 7488 2320 7500
rect 2372 7488 2378 7540
rect 4798 7528 4804 7540
rect 2424 7500 4804 7528
rect 2424 7469 2452 7500
rect 4798 7488 4804 7500
rect 4856 7488 4862 7540
rect 4893 7531 4951 7537
rect 4893 7497 4905 7531
rect 4939 7497 4951 7531
rect 7098 7528 7104 7540
rect 4893 7491 4951 7497
rect 6380 7500 7104 7528
rect 2409 7463 2467 7469
rect 2409 7429 2421 7463
rect 2455 7429 2467 7463
rect 2409 7423 2467 7429
rect 3878 7420 3884 7472
rect 3936 7420 3942 7472
rect 4908 7460 4936 7491
rect 6380 7460 6408 7500
rect 7098 7488 7104 7500
rect 7156 7488 7162 7540
rect 7558 7488 7564 7540
rect 7616 7528 7622 7540
rect 8202 7528 8208 7540
rect 7616 7500 8208 7528
rect 7616 7488 7622 7500
rect 8202 7488 8208 7500
rect 8260 7488 8266 7540
rect 9033 7531 9091 7537
rect 9033 7497 9045 7531
rect 9079 7528 9091 7531
rect 9122 7528 9128 7540
rect 9079 7500 9128 7528
rect 9079 7497 9091 7500
rect 9033 7491 9091 7497
rect 9122 7488 9128 7500
rect 9180 7488 9186 7540
rect 9214 7488 9220 7540
rect 9272 7528 9278 7540
rect 9401 7531 9459 7537
rect 9401 7528 9413 7531
rect 9272 7500 9413 7528
rect 9272 7488 9278 7500
rect 9401 7497 9413 7500
rect 9447 7497 9459 7531
rect 9401 7491 9459 7497
rect 6822 7460 6828 7472
rect 4908 7432 6408 7460
rect 6472 7432 6828 7460
rect 1397 7395 1455 7401
rect 1397 7361 1409 7395
rect 1443 7361 1455 7395
rect 1397 7355 1455 7361
rect 1673 7395 1731 7401
rect 1673 7361 1685 7395
rect 1719 7392 1731 7395
rect 1762 7392 1768 7404
rect 1719 7364 1768 7392
rect 1719 7361 1731 7364
rect 1673 7355 1731 7361
rect 1412 7324 1440 7355
rect 1762 7352 1768 7364
rect 1820 7392 1826 7404
rect 1949 7395 2007 7401
rect 1949 7392 1961 7395
rect 1820 7364 1961 7392
rect 1820 7352 1826 7364
rect 1949 7361 1961 7364
rect 1995 7361 2007 7395
rect 1949 7355 2007 7361
rect 2222 7352 2228 7404
rect 2280 7392 2286 7404
rect 2593 7395 2651 7401
rect 2593 7392 2605 7395
rect 2280 7364 2605 7392
rect 2280 7352 2286 7364
rect 2593 7361 2605 7364
rect 2639 7361 2651 7395
rect 2593 7355 2651 7361
rect 2774 7352 2780 7404
rect 2832 7392 2838 7404
rect 2961 7395 3019 7401
rect 2961 7392 2973 7395
rect 2832 7364 2973 7392
rect 2832 7352 2838 7364
rect 2961 7361 2973 7364
rect 3007 7361 3019 7395
rect 2961 7355 3019 7361
rect 4433 7395 4491 7401
rect 4433 7361 4445 7395
rect 4479 7392 4491 7395
rect 5258 7392 5264 7404
rect 4479 7364 5264 7392
rect 4479 7361 4491 7364
rect 4433 7355 4491 7361
rect 5258 7352 5264 7364
rect 5316 7352 5322 7404
rect 5905 7395 5963 7401
rect 5905 7392 5917 7395
rect 5368 7364 5917 7392
rect 1854 7324 1860 7336
rect 1412 7296 1860 7324
rect 1854 7284 1860 7296
rect 1912 7284 1918 7336
rect 5368 7324 5396 7364
rect 5905 7361 5917 7364
rect 5951 7361 5963 7395
rect 6178 7392 6184 7404
rect 6139 7364 6184 7392
rect 5905 7355 5963 7361
rect 4724 7296 5396 7324
rect 5629 7327 5687 7333
rect 1581 7259 1639 7265
rect 1581 7225 1593 7259
rect 1627 7256 1639 7259
rect 1627 7228 2636 7256
rect 1627 7225 1639 7228
rect 1581 7219 1639 7225
rect 2130 7188 2136 7200
rect 2091 7160 2136 7188
rect 2130 7148 2136 7160
rect 2188 7148 2194 7200
rect 2608 7188 2636 7228
rect 3878 7216 3884 7268
rect 3936 7256 3942 7268
rect 4724 7256 4752 7296
rect 5629 7293 5641 7327
rect 5675 7293 5687 7327
rect 5920 7324 5948 7355
rect 6178 7352 6184 7364
rect 6236 7352 6242 7404
rect 6472 7401 6500 7432
rect 6822 7420 6828 7432
rect 6880 7420 6886 7472
rect 7282 7420 7288 7472
rect 7340 7420 7346 7472
rect 6457 7395 6515 7401
rect 6457 7361 6469 7395
rect 6503 7361 6515 7395
rect 6457 7355 6515 7361
rect 8297 7395 8355 7401
rect 8297 7361 8309 7395
rect 8343 7392 8355 7395
rect 9490 7392 9496 7404
rect 8343 7364 9496 7392
rect 8343 7361 8355 7364
rect 8297 7355 8355 7361
rect 6362 7324 6368 7336
rect 5920 7296 6368 7324
rect 5629 7287 5687 7293
rect 3936 7228 4752 7256
rect 5644 7256 5672 7287
rect 6362 7284 6368 7296
rect 6420 7284 6426 7336
rect 6733 7327 6791 7333
rect 6733 7293 6745 7327
rect 6779 7324 6791 7327
rect 7098 7324 7104 7336
rect 6779 7296 7104 7324
rect 6779 7293 6791 7296
rect 6733 7287 6791 7293
rect 7098 7284 7104 7296
rect 7156 7284 7162 7336
rect 7190 7284 7196 7336
rect 7248 7324 7254 7336
rect 8312 7324 8340 7355
rect 9490 7352 9496 7364
rect 9548 7352 9554 7404
rect 7248 7296 8340 7324
rect 7248 7284 7254 7296
rect 8662 7284 8668 7336
rect 8720 7324 8726 7336
rect 8757 7327 8815 7333
rect 8757 7324 8769 7327
rect 8720 7296 8769 7324
rect 8720 7284 8726 7296
rect 8757 7293 8769 7296
rect 8803 7293 8815 7327
rect 8757 7287 8815 7293
rect 8941 7327 8999 7333
rect 8941 7293 8953 7327
rect 8987 7293 8999 7327
rect 8941 7287 8999 7293
rect 6086 7256 6092 7268
rect 5644 7228 6092 7256
rect 3936 7216 3942 7228
rect 6086 7216 6092 7228
rect 6144 7216 6150 7268
rect 6270 7216 6276 7268
rect 6328 7256 6334 7268
rect 8956 7256 8984 7287
rect 6328 7228 6408 7256
rect 6328 7216 6334 7228
rect 6178 7188 6184 7200
rect 2608 7160 6184 7188
rect 6178 7148 6184 7160
rect 6236 7148 6242 7200
rect 6380 7197 6408 7228
rect 7760 7228 8984 7256
rect 6365 7191 6423 7197
rect 6365 7157 6377 7191
rect 6411 7157 6423 7191
rect 6365 7151 6423 7157
rect 6454 7148 6460 7200
rect 6512 7188 6518 7200
rect 7760 7188 7788 7228
rect 6512 7160 7788 7188
rect 8481 7191 8539 7197
rect 6512 7148 6518 7160
rect 8481 7157 8493 7191
rect 8527 7188 8539 7191
rect 11054 7188 11060 7200
rect 8527 7160 11060 7188
rect 8527 7157 8539 7160
rect 8481 7151 8539 7157
rect 11054 7148 11060 7160
rect 11112 7148 11118 7200
rect 920 7098 9844 7120
rect 920 7046 2566 7098
rect 2618 7046 2630 7098
rect 2682 7046 2694 7098
rect 2746 7046 2758 7098
rect 2810 7046 2822 7098
rect 2874 7046 5666 7098
rect 5718 7046 5730 7098
rect 5782 7046 5794 7098
rect 5846 7046 5858 7098
rect 5910 7046 5922 7098
rect 5974 7046 8766 7098
rect 8818 7046 8830 7098
rect 8882 7046 8894 7098
rect 8946 7046 8958 7098
rect 9010 7046 9022 7098
rect 9074 7046 9844 7098
rect 920 7024 9844 7046
rect 1026 6944 1032 6996
rect 1084 6984 1090 6996
rect 1213 6987 1271 6993
rect 1213 6984 1225 6987
rect 1084 6956 1225 6984
rect 1084 6944 1090 6956
rect 1213 6953 1225 6956
rect 1259 6953 1271 6987
rect 1213 6947 1271 6953
rect 2314 6944 2320 6996
rect 2372 6984 2378 6996
rect 3326 6984 3332 6996
rect 2372 6956 3332 6984
rect 2372 6944 2378 6956
rect 3326 6944 3332 6956
rect 3384 6944 3390 6996
rect 3694 6944 3700 6996
rect 3752 6984 3758 6996
rect 6362 6984 6368 6996
rect 3752 6956 5212 6984
rect 6323 6956 6368 6984
rect 3752 6944 3758 6956
rect 5184 6916 5212 6956
rect 6362 6944 6368 6956
rect 6420 6984 6426 6996
rect 7190 6984 7196 6996
rect 6420 6956 7196 6984
rect 6420 6944 6426 6956
rect 7190 6944 7196 6956
rect 7248 6984 7254 6996
rect 7742 6984 7748 6996
rect 7248 6956 7748 6984
rect 7248 6944 7254 6956
rect 7742 6944 7748 6956
rect 7800 6944 7806 6996
rect 8202 6944 8208 6996
rect 8260 6984 8266 6996
rect 8309 6987 8367 6993
rect 8309 6984 8321 6987
rect 8260 6956 8321 6984
rect 8260 6944 8266 6956
rect 8309 6953 8321 6956
rect 8355 6953 8367 6987
rect 8309 6947 8367 6953
rect 8570 6944 8576 6996
rect 8628 6984 8634 6996
rect 8757 6987 8815 6993
rect 8757 6984 8769 6987
rect 8628 6956 8769 6984
rect 8628 6944 8634 6956
rect 8757 6953 8769 6956
rect 8803 6953 8815 6987
rect 8757 6947 8815 6953
rect 5184 6888 5580 6916
rect 1673 6851 1731 6857
rect 1673 6817 1685 6851
rect 1719 6848 1731 6851
rect 2314 6848 2320 6860
rect 1719 6820 2320 6848
rect 1719 6817 1731 6820
rect 1673 6811 1731 6817
rect 2314 6808 2320 6820
rect 2372 6808 2378 6860
rect 2590 6808 2596 6860
rect 2648 6848 2654 6860
rect 3605 6851 3663 6857
rect 2648 6820 3372 6848
rect 2648 6808 2654 6820
rect 1394 6780 1400 6792
rect 1355 6752 1400 6780
rect 1394 6740 1400 6752
rect 1452 6740 1458 6792
rect 3050 6740 3056 6792
rect 3108 6740 3114 6792
rect 1670 6672 1676 6724
rect 1728 6712 1734 6724
rect 1949 6715 2007 6721
rect 1949 6712 1961 6715
rect 1728 6684 1961 6712
rect 1728 6672 1734 6684
rect 1949 6681 1961 6684
rect 1995 6681 2007 6715
rect 3344 6712 3372 6820
rect 3605 6817 3617 6851
rect 3651 6848 3663 6851
rect 3694 6848 3700 6860
rect 3651 6820 3700 6848
rect 3651 6817 3663 6820
rect 3605 6811 3663 6817
rect 3694 6808 3700 6820
rect 3752 6808 3758 6860
rect 5552 6848 5580 6888
rect 6270 6876 6276 6928
rect 6328 6916 6334 6928
rect 6638 6916 6644 6928
rect 6328 6888 6644 6916
rect 6328 6876 6334 6888
rect 6638 6876 6644 6888
rect 6696 6876 6702 6928
rect 5552 6820 6316 6848
rect 3418 6740 3424 6792
rect 3476 6780 3482 6792
rect 3973 6783 4031 6789
rect 3973 6780 3985 6783
rect 3476 6752 3985 6780
rect 3476 6740 3482 6752
rect 3973 6749 3985 6752
rect 4019 6749 4031 6783
rect 3973 6743 4031 6749
rect 5445 6783 5503 6789
rect 5445 6749 5457 6783
rect 5491 6749 5503 6783
rect 5445 6743 5503 6749
rect 3344 6684 3556 6712
rect 1949 6675 2007 6681
rect 1581 6647 1639 6653
rect 1581 6613 1593 6647
rect 1627 6644 1639 6647
rect 2590 6644 2596 6656
rect 1627 6616 2596 6644
rect 1627 6613 1639 6616
rect 1581 6607 1639 6613
rect 2590 6604 2596 6616
rect 2648 6604 2654 6656
rect 2682 6604 2688 6656
rect 2740 6644 2746 6656
rect 3418 6644 3424 6656
rect 2740 6616 3424 6644
rect 2740 6604 2746 6616
rect 3418 6604 3424 6616
rect 3476 6604 3482 6656
rect 3528 6644 3556 6684
rect 4706 6672 4712 6724
rect 4764 6672 4770 6724
rect 5460 6644 5488 6743
rect 6086 6740 6092 6792
rect 6144 6780 6150 6792
rect 6288 6789 6316 6820
rect 6546 6808 6552 6860
rect 6604 6848 6610 6860
rect 6822 6848 6828 6860
rect 6604 6820 6828 6848
rect 6604 6808 6610 6820
rect 6822 6808 6828 6820
rect 6880 6848 6886 6860
rect 8573 6851 8631 6857
rect 8573 6848 8585 6851
rect 6880 6820 8585 6848
rect 6880 6808 6886 6820
rect 8573 6817 8585 6820
rect 8619 6817 8631 6851
rect 8573 6811 8631 6817
rect 8662 6808 8668 6860
rect 8720 6848 8726 6860
rect 9309 6851 9367 6857
rect 9309 6848 9321 6851
rect 8720 6820 9321 6848
rect 8720 6808 8726 6820
rect 9309 6817 9321 6820
rect 9355 6817 9367 6851
rect 9309 6811 9367 6817
rect 6181 6783 6239 6789
rect 6181 6780 6193 6783
rect 6144 6752 6193 6780
rect 6144 6740 6150 6752
rect 6181 6749 6193 6752
rect 6227 6749 6239 6783
rect 6181 6743 6239 6749
rect 6273 6783 6331 6789
rect 6273 6749 6285 6783
rect 6319 6780 6331 6783
rect 6914 6780 6920 6792
rect 6319 6752 6920 6780
rect 6319 6749 6331 6752
rect 6273 6743 6331 6749
rect 6914 6740 6920 6752
rect 6972 6740 6978 6792
rect 7190 6740 7196 6792
rect 7248 6740 7254 6792
rect 9122 6780 9128 6792
rect 8680 6752 9128 6780
rect 8680 6724 8708 6752
rect 9122 6740 9128 6752
rect 9180 6740 9186 6792
rect 5920 6684 7052 6712
rect 5920 6653 5948 6684
rect 3528 6616 5488 6644
rect 5905 6647 5963 6653
rect 5905 6613 5917 6647
rect 5951 6613 5963 6647
rect 5905 6607 5963 6613
rect 5994 6604 6000 6656
rect 6052 6644 6058 6656
rect 6052 6616 6097 6644
rect 6052 6604 6058 6616
rect 6638 6604 6644 6656
rect 6696 6644 6702 6656
rect 6733 6647 6791 6653
rect 6733 6644 6745 6647
rect 6696 6616 6745 6644
rect 6696 6604 6702 6616
rect 6733 6613 6745 6616
rect 6779 6613 6791 6647
rect 6733 6607 6791 6613
rect 6825 6647 6883 6653
rect 6825 6613 6837 6647
rect 6871 6644 6883 6647
rect 6914 6644 6920 6656
rect 6871 6616 6920 6644
rect 6871 6613 6883 6616
rect 6825 6607 6883 6613
rect 6914 6604 6920 6616
rect 6972 6604 6978 6656
rect 7024 6644 7052 6684
rect 8662 6672 8668 6724
rect 8720 6672 8726 6724
rect 8110 6644 8116 6656
rect 7024 6616 8116 6644
rect 8110 6604 8116 6616
rect 8168 6604 8174 6656
rect 9122 6644 9128 6656
rect 9083 6616 9128 6644
rect 9122 6604 9128 6616
rect 9180 6604 9186 6656
rect 9214 6604 9220 6656
rect 9272 6644 9278 6656
rect 9272 6616 9317 6644
rect 9272 6604 9278 6616
rect 920 6554 9844 6576
rect 920 6502 4116 6554
rect 4168 6502 4180 6554
rect 4232 6502 4244 6554
rect 4296 6502 4308 6554
rect 4360 6502 4372 6554
rect 4424 6502 7216 6554
rect 7268 6502 7280 6554
rect 7332 6502 7344 6554
rect 7396 6502 7408 6554
rect 7460 6502 7472 6554
rect 7524 6502 9844 6554
rect 920 6480 9844 6502
rect 1765 6443 1823 6449
rect 1765 6409 1777 6443
rect 1811 6440 1823 6443
rect 2406 6440 2412 6452
rect 1811 6412 2412 6440
rect 1811 6409 1823 6412
rect 1765 6403 1823 6409
rect 2406 6400 2412 6412
rect 2464 6400 2470 6452
rect 3050 6400 3056 6452
rect 3108 6400 3114 6452
rect 4709 6443 4767 6449
rect 4709 6409 4721 6443
rect 4755 6440 4767 6443
rect 4798 6440 4804 6452
rect 4755 6412 4804 6440
rect 4755 6409 4767 6412
rect 4709 6403 4767 6409
rect 4798 6400 4804 6412
rect 4856 6400 4862 6452
rect 9122 6440 9128 6452
rect 5460 6412 9128 6440
rect 1118 6332 1124 6384
rect 1176 6372 1182 6384
rect 1949 6375 2007 6381
rect 1949 6372 1961 6375
rect 1176 6344 1961 6372
rect 1176 6332 1182 6344
rect 1949 6341 1961 6344
rect 1995 6341 2007 6375
rect 2682 6372 2688 6384
rect 2643 6344 2688 6372
rect 1949 6335 2007 6341
rect 2682 6332 2688 6344
rect 2740 6332 2746 6384
rect 3068 6372 3096 6400
rect 3068 6344 3174 6372
rect 2314 6264 2320 6316
rect 2372 6304 2378 6316
rect 2409 6307 2467 6313
rect 2409 6304 2421 6307
rect 2372 6276 2421 6304
rect 2372 6264 2378 6276
rect 2409 6273 2421 6276
rect 2455 6273 2467 6307
rect 2409 6267 2467 6273
rect 1578 6196 1584 6248
rect 1636 6236 1642 6248
rect 5460 6236 5488 6412
rect 9122 6400 9128 6412
rect 9180 6400 9186 6452
rect 5997 6375 6055 6381
rect 5997 6341 6009 6375
rect 6043 6372 6055 6375
rect 6730 6372 6736 6384
rect 6043 6344 6736 6372
rect 6043 6341 6055 6344
rect 5997 6335 6055 6341
rect 6730 6332 6736 6344
rect 6788 6332 6794 6384
rect 6822 6332 6828 6384
rect 6880 6332 6886 6384
rect 9306 6372 9312 6384
rect 8326 6344 9312 6372
rect 9306 6332 9312 6344
rect 9364 6332 9370 6384
rect 5902 6264 5908 6316
rect 5960 6304 5966 6316
rect 6273 6307 6331 6313
rect 6273 6304 6285 6307
rect 5960 6276 6285 6304
rect 5960 6264 5966 6276
rect 6273 6273 6285 6276
rect 6319 6304 6331 6307
rect 6840 6304 6868 6332
rect 6319 6276 6868 6304
rect 6319 6273 6331 6276
rect 6273 6267 6331 6273
rect 8478 6264 8484 6316
rect 8536 6304 8542 6316
rect 8665 6307 8723 6313
rect 8665 6304 8677 6307
rect 8536 6276 8677 6304
rect 8536 6264 8542 6276
rect 8665 6273 8677 6276
rect 8711 6273 8723 6307
rect 9217 6307 9275 6313
rect 9217 6304 9229 6307
rect 8665 6267 8723 6273
rect 8772 6276 9229 6304
rect 1636 6208 5488 6236
rect 1636 6196 1642 6208
rect 5534 6196 5540 6248
rect 5592 6236 5598 6248
rect 6825 6239 6883 6245
rect 6825 6236 6837 6239
rect 5592 6208 6837 6236
rect 5592 6196 5598 6208
rect 6825 6205 6837 6208
rect 6871 6205 6883 6239
rect 7190 6236 7196 6248
rect 7151 6208 7196 6236
rect 6825 6199 6883 6205
rect 7190 6196 7196 6208
rect 7248 6196 7254 6248
rect 6454 6128 6460 6180
rect 6512 6168 6518 6180
rect 6512 6140 6960 6168
rect 6512 6128 6518 6140
rect 3970 6060 3976 6112
rect 4028 6100 4034 6112
rect 4157 6103 4215 6109
rect 4157 6100 4169 6103
rect 4028 6072 4169 6100
rect 4028 6060 4034 6072
rect 4157 6069 4169 6072
rect 4203 6069 4215 6103
rect 4157 6063 4215 6069
rect 4982 6060 4988 6112
rect 5040 6100 5046 6112
rect 6362 6100 6368 6112
rect 5040 6072 6368 6100
rect 5040 6060 5046 6072
rect 6362 6060 6368 6072
rect 6420 6060 6426 6112
rect 6733 6103 6791 6109
rect 6733 6069 6745 6103
rect 6779 6100 6791 6103
rect 6822 6100 6828 6112
rect 6779 6072 6828 6100
rect 6779 6069 6791 6072
rect 6733 6063 6791 6069
rect 6822 6060 6828 6072
rect 6880 6060 6886 6112
rect 6932 6100 6960 6140
rect 8772 6100 8800 6276
rect 9217 6273 9229 6276
rect 9263 6273 9275 6307
rect 9217 6267 9275 6273
rect 9122 6100 9128 6112
rect 6932 6072 8800 6100
rect 9083 6072 9128 6100
rect 9122 6060 9128 6072
rect 9180 6060 9186 6112
rect 9398 6100 9404 6112
rect 9359 6072 9404 6100
rect 9398 6060 9404 6072
rect 9456 6060 9462 6112
rect 920 6010 9844 6032
rect 920 5958 2566 6010
rect 2618 5958 2630 6010
rect 2682 5958 2694 6010
rect 2746 5958 2758 6010
rect 2810 5958 2822 6010
rect 2874 5958 5666 6010
rect 5718 5958 5730 6010
rect 5782 5958 5794 6010
rect 5846 5958 5858 6010
rect 5910 5958 5922 6010
rect 5974 5958 8766 6010
rect 8818 5958 8830 6010
rect 8882 5958 8894 6010
rect 8946 5958 8958 6010
rect 9010 5958 9022 6010
rect 9074 5958 9844 6010
rect 920 5936 9844 5958
rect 2961 5899 3019 5905
rect 2961 5865 2973 5899
rect 3007 5896 3019 5899
rect 3694 5896 3700 5908
rect 3007 5868 3700 5896
rect 3007 5865 3019 5868
rect 2961 5859 3019 5865
rect 3694 5856 3700 5868
rect 3752 5856 3758 5908
rect 3786 5856 3792 5908
rect 3844 5896 3850 5908
rect 7006 5896 7012 5908
rect 3844 5868 3889 5896
rect 5552 5868 7012 5896
rect 3844 5856 3850 5868
rect 1394 5788 1400 5840
rect 1452 5828 1458 5840
rect 3053 5831 3111 5837
rect 3053 5828 3065 5831
rect 1452 5800 3065 5828
rect 1452 5788 1458 5800
rect 3053 5797 3065 5800
rect 3099 5797 3111 5831
rect 3605 5831 3663 5837
rect 3605 5828 3617 5831
rect 3053 5791 3111 5797
rect 3160 5800 3617 5828
rect 3160 5760 3188 5800
rect 3605 5797 3617 5800
rect 3651 5797 3663 5831
rect 3605 5791 3663 5797
rect 2516 5732 3188 5760
rect 2516 5701 2544 5732
rect 3326 5720 3332 5772
rect 3384 5760 3390 5772
rect 4249 5763 4307 5769
rect 4249 5760 4261 5763
rect 3384 5732 4261 5760
rect 3384 5720 3390 5732
rect 4249 5729 4261 5732
rect 4295 5729 4307 5763
rect 4249 5723 4307 5729
rect 4525 5763 4583 5769
rect 4525 5729 4537 5763
rect 4571 5760 4583 5763
rect 5552 5760 5580 5868
rect 7006 5856 7012 5868
rect 7064 5856 7070 5908
rect 7190 5856 7196 5908
rect 7248 5896 7254 5908
rect 7558 5896 7564 5908
rect 7248 5868 7564 5896
rect 7248 5856 7254 5868
rect 7558 5856 7564 5868
rect 7616 5896 7622 5908
rect 8021 5899 8079 5905
rect 8021 5896 8033 5899
rect 7616 5868 8033 5896
rect 7616 5856 7622 5868
rect 8021 5865 8033 5868
rect 8067 5865 8079 5899
rect 8021 5859 8079 5865
rect 9125 5899 9183 5905
rect 9125 5865 9137 5899
rect 9171 5865 9183 5899
rect 9306 5896 9312 5908
rect 9267 5868 9312 5896
rect 9125 5859 9183 5865
rect 9140 5828 9168 5859
rect 9306 5856 9312 5868
rect 9364 5856 9370 5908
rect 9490 5828 9496 5840
rect 9140 5800 9496 5828
rect 9490 5788 9496 5800
rect 9548 5788 9554 5840
rect 4571 5732 5580 5760
rect 6273 5763 6331 5769
rect 4571 5729 4583 5732
rect 4525 5723 4583 5729
rect 6273 5729 6285 5763
rect 6319 5760 6331 5763
rect 6546 5760 6552 5772
rect 6319 5732 6552 5760
rect 6319 5729 6331 5732
rect 6273 5723 6331 5729
rect 6546 5720 6552 5732
rect 6604 5720 6610 5772
rect 6638 5720 6644 5772
rect 6696 5760 6702 5772
rect 6696 5732 9536 5760
rect 6696 5720 6702 5732
rect 2501 5695 2559 5701
rect 2501 5661 2513 5695
rect 2547 5661 2559 5695
rect 2501 5655 2559 5661
rect 2777 5695 2835 5701
rect 2777 5661 2789 5695
rect 2823 5661 2835 5695
rect 2777 5655 2835 5661
rect 2130 5584 2136 5636
rect 2188 5624 2194 5636
rect 2792 5624 2820 5655
rect 3142 5652 3148 5704
rect 3200 5692 3206 5704
rect 3421 5695 3479 5701
rect 3421 5692 3433 5695
rect 3200 5664 3433 5692
rect 3200 5652 3206 5664
rect 3421 5661 3433 5664
rect 3467 5692 3479 5695
rect 4065 5695 4123 5701
rect 4065 5692 4077 5695
rect 3467 5664 4077 5692
rect 3467 5661 3479 5664
rect 3421 5655 3479 5661
rect 4065 5661 4077 5664
rect 4111 5661 4123 5695
rect 4065 5655 4123 5661
rect 7650 5652 7656 5704
rect 7708 5692 7714 5704
rect 8297 5695 8355 5701
rect 8297 5692 8309 5695
rect 7708 5664 8309 5692
rect 7708 5652 7714 5664
rect 8297 5661 8309 5664
rect 8343 5661 8355 5695
rect 8297 5655 8355 5661
rect 8662 5652 8668 5704
rect 8720 5692 8726 5704
rect 9508 5701 9536 5732
rect 9217 5695 9275 5701
rect 9217 5692 9229 5695
rect 8720 5664 9229 5692
rect 8720 5652 8726 5664
rect 9217 5661 9229 5664
rect 9263 5661 9275 5695
rect 9217 5655 9275 5661
rect 9493 5695 9551 5701
rect 9493 5661 9505 5695
rect 9539 5661 9551 5695
rect 9493 5655 9551 5661
rect 2188 5596 2820 5624
rect 2188 5584 2194 5596
rect 3050 5584 3056 5636
rect 3108 5624 3114 5636
rect 3237 5627 3295 5633
rect 3237 5624 3249 5627
rect 3108 5596 3249 5624
rect 3108 5584 3114 5596
rect 3237 5593 3249 5596
rect 3283 5624 3295 5627
rect 3786 5624 3792 5636
rect 3283 5596 3792 5624
rect 3283 5593 3295 5596
rect 3237 5587 3295 5593
rect 3786 5584 3792 5596
rect 3844 5624 3850 5636
rect 4982 5624 4988 5636
rect 3844 5596 4988 5624
rect 3844 5584 3850 5596
rect 4982 5584 4988 5596
rect 5040 5584 5046 5636
rect 6178 5624 6184 5636
rect 6012 5596 6184 5624
rect 2685 5559 2743 5565
rect 2685 5525 2697 5559
rect 2731 5556 2743 5559
rect 4706 5556 4712 5568
rect 2731 5528 4712 5556
rect 2731 5525 2743 5528
rect 2685 5519 2743 5525
rect 4706 5516 4712 5528
rect 4764 5516 4770 5568
rect 6012 5565 6040 5596
rect 6178 5584 6184 5596
rect 6236 5624 6242 5636
rect 6549 5627 6607 5633
rect 6549 5624 6561 5627
rect 6236 5596 6561 5624
rect 6236 5584 6242 5596
rect 6549 5593 6561 5596
rect 6595 5593 6607 5627
rect 8113 5627 8171 5633
rect 8113 5624 8125 5627
rect 6549 5587 6607 5593
rect 7852 5596 8125 5624
rect 5997 5559 6055 5565
rect 5997 5525 6009 5559
rect 6043 5525 6055 5559
rect 5997 5519 6055 5525
rect 6730 5516 6736 5568
rect 6788 5556 6794 5568
rect 7852 5556 7880 5596
rect 8113 5593 8125 5596
rect 8159 5593 8171 5627
rect 8113 5587 8171 5593
rect 9030 5584 9036 5636
rect 9088 5624 9094 5636
rect 9306 5624 9312 5636
rect 9088 5596 9312 5624
rect 9088 5584 9094 5596
rect 9306 5584 9312 5596
rect 9364 5584 9370 5636
rect 6788 5528 7880 5556
rect 6788 5516 6794 5528
rect 8018 5516 8024 5568
rect 8076 5556 8082 5568
rect 8481 5559 8539 5565
rect 8481 5556 8493 5559
rect 8076 5528 8493 5556
rect 8076 5516 8082 5528
rect 8481 5525 8493 5528
rect 8527 5525 8539 5559
rect 8481 5519 8539 5525
rect 8757 5559 8815 5565
rect 8757 5525 8769 5559
rect 8803 5556 8815 5559
rect 9122 5556 9128 5568
rect 8803 5528 9128 5556
rect 8803 5525 8815 5528
rect 8757 5519 8815 5525
rect 9122 5516 9128 5528
rect 9180 5516 9186 5568
rect 920 5466 9844 5488
rect 920 5414 4116 5466
rect 4168 5414 4180 5466
rect 4232 5414 4244 5466
rect 4296 5414 4308 5466
rect 4360 5414 4372 5466
rect 4424 5414 7216 5466
rect 7268 5414 7280 5466
rect 7332 5414 7344 5466
rect 7396 5414 7408 5466
rect 7460 5414 7472 5466
rect 7524 5414 9844 5466
rect 920 5392 9844 5414
rect 3786 5312 3792 5364
rect 3844 5312 3850 5364
rect 4614 5312 4620 5364
rect 4672 5352 4678 5364
rect 5077 5355 5135 5361
rect 5077 5352 5089 5355
rect 4672 5324 5089 5352
rect 4672 5312 4678 5324
rect 5077 5321 5089 5324
rect 5123 5321 5135 5355
rect 5077 5315 5135 5321
rect 5353 5355 5411 5361
rect 5353 5321 5365 5355
rect 5399 5352 5411 5355
rect 5442 5352 5448 5364
rect 5399 5324 5448 5352
rect 5399 5321 5411 5324
rect 5353 5315 5411 5321
rect 5442 5312 5448 5324
rect 5500 5312 5506 5364
rect 5994 5352 6000 5364
rect 5552 5324 6000 5352
rect 3804 5284 3832 5312
rect 3804 5256 4094 5284
rect 3326 5216 3332 5228
rect 3287 5188 3332 5216
rect 3326 5176 3332 5188
rect 3384 5176 3390 5228
rect 5169 5219 5227 5225
rect 5169 5185 5181 5219
rect 5215 5216 5227 5219
rect 5552 5216 5580 5324
rect 5994 5312 6000 5324
rect 6052 5312 6058 5364
rect 6914 5244 6920 5296
rect 6972 5244 6978 5296
rect 5215 5188 5580 5216
rect 5629 5219 5687 5225
rect 5215 5185 5227 5188
rect 5169 5179 5227 5185
rect 5629 5185 5641 5219
rect 5675 5216 5687 5219
rect 5994 5216 6000 5228
rect 5675 5188 6000 5216
rect 5675 5185 5687 5188
rect 5629 5179 5687 5185
rect 3605 5151 3663 5157
rect 3605 5117 3617 5151
rect 3651 5148 3663 5151
rect 3970 5148 3976 5160
rect 3651 5120 3976 5148
rect 3651 5117 3663 5120
rect 3605 5111 3663 5117
rect 3970 5108 3976 5120
rect 4028 5108 4034 5160
rect 5534 5108 5540 5160
rect 5592 5148 5598 5160
rect 5644 5148 5672 5179
rect 5994 5176 6000 5188
rect 6052 5176 6058 5228
rect 6178 5216 6184 5228
rect 6139 5188 6184 5216
rect 6178 5176 6184 5188
rect 6236 5176 6242 5228
rect 7650 5216 7656 5228
rect 7611 5188 7656 5216
rect 7650 5176 7656 5188
rect 7708 5176 7714 5228
rect 8297 5219 8355 5225
rect 8297 5216 8309 5219
rect 8128 5188 8309 5216
rect 5592 5120 5672 5148
rect 5813 5151 5871 5157
rect 5592 5108 5598 5120
rect 5813 5117 5825 5151
rect 5859 5148 5871 5151
rect 6086 5148 6092 5160
rect 5859 5120 6092 5148
rect 5859 5117 5871 5120
rect 5813 5111 5871 5117
rect 6086 5108 6092 5120
rect 6144 5108 6150 5160
rect 8128 5157 8156 5188
rect 8297 5185 8309 5188
rect 8343 5216 8355 5219
rect 9490 5216 9496 5228
rect 8343 5188 9496 5216
rect 8343 5185 8355 5188
rect 8297 5179 8355 5185
rect 9490 5176 9496 5188
rect 9548 5176 9554 5228
rect 8113 5151 8171 5157
rect 8113 5117 8125 5151
rect 8159 5117 8171 5151
rect 8113 5111 8171 5117
rect 8570 5108 8576 5160
rect 8628 5148 8634 5160
rect 8665 5151 8723 5157
rect 8665 5148 8677 5151
rect 8628 5120 8677 5148
rect 8628 5108 8634 5120
rect 8665 5117 8677 5120
rect 8711 5117 8723 5151
rect 8665 5111 8723 5117
rect 8754 5108 8760 5160
rect 8812 5148 8818 5160
rect 8849 5151 8907 5157
rect 8849 5148 8861 5151
rect 8812 5120 8861 5148
rect 8812 5108 8818 5120
rect 8849 5117 8861 5120
rect 8895 5117 8907 5151
rect 8849 5111 8907 5117
rect 8481 5083 8539 5089
rect 8481 5049 8493 5083
rect 8527 5080 8539 5083
rect 16574 5080 16580 5092
rect 8527 5052 16580 5080
rect 8527 5049 8539 5052
rect 8481 5043 8539 5049
rect 16574 5040 16580 5052
rect 16632 5040 16638 5092
rect 5442 4972 5448 5024
rect 5500 5012 5506 5024
rect 5500 4984 5545 5012
rect 5500 4972 5506 4984
rect 7190 4972 7196 5024
rect 7248 5012 7254 5024
rect 8018 5012 8024 5024
rect 7248 4984 8024 5012
rect 7248 4972 7254 4984
rect 8018 4972 8024 4984
rect 8076 4972 8082 5024
rect 9309 5015 9367 5021
rect 9309 4981 9321 5015
rect 9355 5012 9367 5015
rect 9582 5012 9588 5024
rect 9355 4984 9588 5012
rect 9355 4981 9367 4984
rect 9309 4975 9367 4981
rect 9582 4972 9588 4984
rect 9640 4972 9646 5024
rect 3036 4922 9844 4944
rect 3036 4870 5666 4922
rect 5718 4870 5730 4922
rect 5782 4870 5794 4922
rect 5846 4870 5858 4922
rect 5910 4870 5922 4922
rect 5974 4870 8766 4922
rect 8818 4870 8830 4922
rect 8882 4870 8894 4922
rect 8946 4870 8958 4922
rect 9010 4870 9022 4922
rect 9074 4870 9844 4922
rect 3036 4848 9844 4870
rect 3786 4808 3792 4820
rect 3747 4780 3792 4808
rect 3786 4768 3792 4780
rect 3844 4808 3850 4820
rect 4433 4811 4491 4817
rect 4433 4808 4445 4811
rect 3844 4780 4445 4808
rect 3844 4768 3850 4780
rect 4433 4777 4445 4780
rect 4479 4777 4491 4811
rect 4433 4771 4491 4777
rect 5537 4811 5595 4817
rect 5537 4777 5549 4811
rect 5583 4808 5595 4811
rect 6086 4808 6092 4820
rect 5583 4780 6092 4808
rect 5583 4777 5595 4780
rect 5537 4771 5595 4777
rect 4448 4672 4476 4771
rect 6086 4768 6092 4780
rect 6144 4768 6150 4820
rect 6914 4768 6920 4820
rect 6972 4808 6978 4820
rect 7009 4811 7067 4817
rect 7009 4808 7021 4811
rect 6972 4780 7021 4808
rect 6972 4768 6978 4780
rect 7009 4777 7021 4780
rect 7055 4777 7067 4811
rect 7009 4771 7067 4777
rect 7285 4811 7343 4817
rect 7285 4777 7297 4811
rect 7331 4808 7343 4811
rect 8478 4808 8484 4820
rect 7331 4780 8484 4808
rect 7331 4777 7343 4780
rect 7285 4771 7343 4777
rect 8478 4768 8484 4780
rect 8536 4768 8542 4820
rect 9214 4768 9220 4820
rect 9272 4808 9278 4820
rect 9401 4811 9459 4817
rect 9401 4808 9413 4811
rect 9272 4780 9413 4808
rect 9272 4768 9278 4780
rect 9401 4777 9413 4780
rect 9447 4777 9459 4811
rect 9401 4771 9459 4777
rect 6733 4743 6791 4749
rect 6733 4709 6745 4743
rect 6779 4740 6791 4743
rect 7650 4740 7656 4752
rect 6779 4712 7656 4740
rect 6779 4709 6791 4712
rect 6733 4703 6791 4709
rect 7650 4700 7656 4712
rect 7708 4700 7714 4752
rect 8294 4740 8300 4752
rect 8255 4712 8300 4740
rect 8294 4700 8300 4712
rect 8352 4700 8358 4752
rect 5261 4675 5319 4681
rect 2746 4644 4384 4672
rect 4448 4644 5120 4672
rect 1486 4564 1492 4616
rect 1544 4604 1550 4616
rect 2746 4604 2774 4644
rect 1544 4576 2774 4604
rect 3605 4607 3663 4613
rect 1544 4564 1550 4576
rect 3605 4573 3617 4607
rect 3651 4573 3663 4607
rect 3605 4567 3663 4573
rect 3620 4536 3648 4567
rect 3694 4564 3700 4616
rect 3752 4604 3758 4616
rect 4356 4613 4384 4644
rect 5092 4613 5120 4644
rect 5261 4641 5273 4675
rect 5307 4672 5319 4675
rect 7926 4672 7932 4684
rect 5307 4644 6408 4672
rect 5307 4641 5319 4644
rect 5261 4635 5319 4641
rect 4341 4607 4399 4613
rect 3752 4576 3797 4604
rect 3752 4564 3758 4576
rect 4341 4573 4353 4607
rect 4387 4604 4399 4607
rect 4893 4607 4951 4613
rect 4893 4604 4905 4607
rect 4387 4576 4905 4604
rect 4387 4573 4399 4576
rect 4341 4567 4399 4573
rect 4893 4573 4905 4576
rect 4939 4573 4951 4607
rect 4893 4567 4951 4573
rect 5077 4607 5135 4613
rect 5077 4573 5089 4607
rect 5123 4573 5135 4607
rect 5077 4567 5135 4573
rect 5353 4607 5411 4613
rect 5353 4573 5365 4607
rect 5399 4604 5411 4607
rect 5442 4604 5448 4616
rect 5399 4576 5448 4604
rect 5399 4573 5411 4576
rect 5353 4567 5411 4573
rect 3970 4536 3976 4548
rect 3620 4508 3976 4536
rect 3970 4496 3976 4508
rect 4028 4496 4034 4548
rect 5092 4536 5120 4567
rect 5442 4564 5448 4576
rect 5500 4564 5506 4616
rect 5718 4604 5724 4616
rect 5679 4576 5724 4604
rect 5718 4564 5724 4576
rect 5776 4564 5782 4616
rect 6380 4613 6408 4644
rect 7116 4644 7932 4672
rect 6365 4607 6423 4613
rect 6365 4573 6377 4607
rect 6411 4573 6423 4607
rect 6365 4567 6423 4573
rect 6549 4607 6607 4613
rect 6549 4573 6561 4607
rect 6595 4573 6607 4607
rect 6822 4604 6828 4616
rect 6783 4576 6828 4604
rect 6549 4567 6607 4573
rect 5905 4539 5963 4545
rect 5905 4536 5917 4539
rect 5092 4508 5917 4536
rect 5905 4505 5917 4508
rect 5951 4536 5963 4539
rect 6454 4536 6460 4548
rect 5951 4508 6460 4536
rect 5951 4505 5963 4508
rect 5905 4499 5963 4505
rect 6454 4496 6460 4508
rect 6512 4496 6518 4548
rect 6564 4536 6592 4567
rect 6822 4564 6828 4576
rect 6880 4564 6886 4616
rect 7116 4613 7144 4644
rect 7926 4632 7932 4644
rect 7984 4632 7990 4684
rect 8202 4632 8208 4684
rect 8260 4672 8266 4684
rect 8386 4672 8392 4684
rect 8260 4644 8392 4672
rect 8260 4632 8266 4644
rect 8386 4632 8392 4644
rect 8444 4672 8450 4684
rect 8757 4675 8815 4681
rect 8757 4672 8769 4675
rect 8444 4644 8769 4672
rect 8444 4632 8450 4644
rect 8757 4641 8769 4644
rect 8803 4641 8815 4675
rect 8757 4635 8815 4641
rect 7101 4607 7159 4613
rect 7101 4573 7113 4607
rect 7147 4573 7159 4607
rect 7558 4604 7564 4616
rect 7519 4576 7564 4604
rect 7101 4567 7159 4573
rect 7558 4564 7564 4576
rect 7616 4564 7622 4616
rect 7745 4607 7803 4613
rect 7745 4573 7757 4607
rect 7791 4573 7803 4607
rect 7745 4567 7803 4573
rect 7190 4536 7196 4548
rect 6564 4508 7196 4536
rect 7190 4496 7196 4508
rect 7248 4496 7254 4548
rect 7377 4539 7435 4545
rect 7377 4505 7389 4539
rect 7423 4536 7435 4539
rect 7650 4536 7656 4548
rect 7423 4508 7656 4536
rect 7423 4505 7435 4508
rect 7377 4499 7435 4505
rect 7650 4496 7656 4508
rect 7708 4496 7714 4548
rect 7760 4536 7788 4567
rect 7834 4564 7840 4616
rect 7892 4604 7898 4616
rect 7892 4576 7937 4604
rect 7892 4564 7898 4576
rect 7760 4508 8064 4536
rect 8036 4480 8064 4508
rect 8386 4496 8392 4548
rect 8444 4536 8450 4548
rect 8444 4508 8489 4536
rect 8444 4496 8450 4508
rect 3326 4428 3332 4480
rect 3384 4468 3390 4480
rect 3421 4471 3479 4477
rect 3421 4468 3433 4471
rect 3384 4440 3433 4468
rect 3384 4428 3390 4440
rect 3421 4437 3433 4440
rect 3467 4437 3479 4471
rect 3421 4431 3479 4437
rect 4157 4471 4215 4477
rect 4157 4437 4169 4471
rect 4203 4468 4215 4471
rect 4614 4468 4620 4480
rect 4203 4440 4620 4468
rect 4203 4437 4215 4440
rect 4157 4431 4215 4437
rect 4614 4428 4620 4440
rect 4672 4428 4678 4480
rect 4801 4471 4859 4477
rect 4801 4437 4813 4471
rect 4847 4468 4859 4471
rect 4982 4468 4988 4480
rect 4847 4440 4988 4468
rect 4847 4437 4859 4440
rect 4801 4431 4859 4437
rect 4982 4428 4988 4440
rect 5040 4428 5046 4480
rect 6086 4468 6092 4480
rect 6047 4440 6092 4468
rect 6086 4428 6092 4440
rect 6144 4428 6150 4480
rect 6178 4428 6184 4480
rect 6236 4468 6242 4480
rect 6236 4440 6281 4468
rect 6236 4428 6242 4440
rect 8018 4428 8024 4480
rect 8076 4468 8082 4480
rect 8481 4471 8539 4477
rect 8481 4468 8493 4471
rect 8076 4440 8493 4468
rect 8076 4428 8082 4440
rect 8481 4437 8493 4440
rect 8527 4437 8539 4471
rect 8938 4468 8944 4480
rect 8899 4440 8944 4468
rect 8481 4431 8539 4437
rect 8938 4428 8944 4440
rect 8996 4428 9002 4480
rect 9033 4471 9091 4477
rect 9033 4437 9045 4471
rect 9079 4468 9091 4471
rect 9306 4468 9312 4480
rect 9079 4440 9312 4468
rect 9079 4437 9091 4440
rect 9033 4431 9091 4437
rect 9306 4428 9312 4440
rect 9364 4428 9370 4480
rect 3036 4378 9844 4400
rect 3036 4326 4116 4378
rect 4168 4326 4180 4378
rect 4232 4326 4244 4378
rect 4296 4326 4308 4378
rect 4360 4326 4372 4378
rect 4424 4326 7216 4378
rect 7268 4326 7280 4378
rect 7332 4326 7344 4378
rect 7396 4326 7408 4378
rect 7460 4326 7472 4378
rect 7524 4326 9844 4378
rect 3036 4304 9844 4326
rect 3970 4224 3976 4276
rect 4028 4264 4034 4276
rect 5534 4264 5540 4276
rect 4028 4236 5540 4264
rect 4028 4224 4034 4236
rect 5534 4224 5540 4236
rect 5592 4264 5598 4276
rect 5592 4236 6040 4264
rect 5592 4224 5598 4236
rect 4522 4156 4528 4208
rect 4580 4156 4586 4208
rect 3326 4128 3332 4140
rect 3287 4100 3332 4128
rect 3326 4088 3332 4100
rect 3384 4088 3390 4140
rect 3878 4088 3884 4140
rect 3936 4128 3942 4140
rect 3973 4131 4031 4137
rect 3973 4128 3985 4131
rect 3936 4100 3985 4128
rect 3936 4088 3942 4100
rect 3973 4097 3985 4100
rect 4019 4097 4031 4131
rect 3973 4091 4031 4097
rect 4890 4088 4896 4140
rect 4948 4128 4954 4140
rect 6012 4137 6040 4236
rect 8294 4224 8300 4276
rect 8352 4264 8358 4276
rect 8570 4264 8576 4276
rect 8352 4236 8576 4264
rect 8352 4224 8358 4236
rect 8570 4224 8576 4236
rect 8628 4224 8634 4276
rect 8665 4267 8723 4273
rect 8665 4233 8677 4267
rect 8711 4264 8723 4267
rect 8938 4264 8944 4276
rect 8711 4236 8944 4264
rect 8711 4233 8723 4236
rect 8665 4227 8723 4233
rect 8938 4224 8944 4236
rect 8996 4224 9002 4276
rect 6454 4156 6460 4208
rect 6512 4196 6518 4208
rect 6638 4196 6644 4208
rect 6512 4168 6644 4196
rect 6512 4156 6518 4168
rect 6638 4156 6644 4168
rect 6696 4196 6702 4208
rect 7285 4199 7343 4205
rect 7285 4196 7297 4199
rect 6696 4168 7297 4196
rect 6696 4156 6702 4168
rect 7285 4165 7297 4168
rect 7331 4165 7343 4199
rect 7285 4159 7343 4165
rect 8478 4156 8484 4208
rect 8536 4196 8542 4208
rect 9033 4199 9091 4205
rect 9033 4196 9045 4199
rect 8536 4168 9045 4196
rect 8536 4156 8542 4168
rect 9033 4165 9045 4168
rect 9079 4165 9091 4199
rect 9033 4159 9091 4165
rect 5445 4131 5503 4137
rect 5445 4128 5457 4131
rect 4948 4100 5457 4128
rect 4948 4088 4954 4100
rect 5445 4097 5457 4100
rect 5491 4097 5503 4131
rect 5445 4091 5503 4097
rect 5997 4131 6055 4137
rect 5997 4097 6009 4131
rect 6043 4097 6055 4131
rect 6273 4131 6331 4137
rect 6273 4128 6285 4131
rect 5997 4091 6055 4097
rect 6196 4100 6285 4128
rect 3605 4063 3663 4069
rect 3605 4029 3617 4063
rect 3651 4029 3663 4063
rect 3605 4023 3663 4029
rect 3513 3995 3571 4001
rect 3513 3961 3525 3995
rect 3559 3992 3571 3995
rect 3620 3992 3648 4023
rect 6196 4001 6224 4100
rect 6273 4097 6285 4100
rect 6319 4097 6331 4131
rect 6273 4091 6331 4097
rect 6362 4088 6368 4140
rect 6420 4128 6426 4140
rect 6549 4131 6607 4137
rect 6549 4128 6561 4131
rect 6420 4100 6561 4128
rect 6420 4088 6426 4100
rect 6549 4097 6561 4100
rect 6595 4128 6607 4131
rect 7101 4131 7159 4137
rect 7101 4128 7113 4131
rect 6595 4100 7113 4128
rect 6595 4097 6607 4100
rect 6549 4091 6607 4097
rect 7101 4097 7113 4100
rect 7147 4097 7159 4131
rect 7101 4091 7159 4097
rect 7561 4131 7619 4137
rect 7561 4097 7573 4131
rect 7607 4097 7619 4131
rect 7561 4091 7619 4097
rect 8113 4131 8171 4137
rect 8113 4097 8125 4131
rect 8159 4097 8171 4131
rect 8570 4128 8576 4140
rect 8531 4100 8576 4128
rect 8113 4091 8171 4097
rect 7009 4063 7067 4069
rect 7009 4029 7021 4063
rect 7055 4060 7067 4063
rect 7576 4060 7604 4091
rect 7055 4032 7604 4060
rect 7055 4029 7067 4032
rect 7009 4023 7067 4029
rect 3559 3964 3648 3992
rect 6181 3995 6239 4001
rect 3559 3961 3571 3964
rect 3513 3955 3571 3961
rect 6181 3961 6193 3995
rect 6227 3961 6239 3995
rect 7926 3992 7932 4004
rect 7887 3964 7932 3992
rect 6181 3955 6239 3961
rect 7926 3952 7932 3964
rect 7984 3952 7990 4004
rect 8128 3992 8156 4091
rect 8570 4088 8576 4100
rect 8628 4088 8634 4140
rect 9125 4131 9183 4137
rect 9125 4097 9137 4131
rect 9171 4128 9183 4131
rect 9306 4128 9312 4140
rect 9171 4100 9312 4128
rect 9171 4097 9183 4100
rect 9125 4091 9183 4097
rect 9306 4088 9312 4100
rect 9364 4088 9370 4140
rect 9214 4020 9220 4072
rect 9272 4060 9278 4072
rect 9272 4032 9317 4060
rect 9272 4020 9278 4032
rect 9398 3992 9404 4004
rect 8128 3964 9404 3992
rect 9398 3952 9404 3964
rect 9456 3952 9462 4004
rect 5905 3927 5963 3933
rect 5905 3893 5917 3927
rect 5951 3924 5963 3927
rect 6362 3924 6368 3936
rect 5951 3896 6368 3924
rect 5951 3893 5963 3896
rect 5905 3887 5963 3893
rect 6362 3884 6368 3896
rect 6420 3884 6426 3936
rect 6457 3927 6515 3933
rect 6457 3893 6469 3927
rect 6503 3924 6515 3927
rect 6546 3924 6552 3936
rect 6503 3896 6552 3924
rect 6503 3893 6515 3896
rect 6457 3887 6515 3893
rect 6546 3884 6552 3896
rect 6604 3884 6610 3936
rect 6638 3884 6644 3936
rect 6696 3924 6702 3936
rect 7469 3927 7527 3933
rect 6696 3896 6741 3924
rect 6696 3884 6702 3896
rect 7469 3893 7481 3927
rect 7515 3924 7527 3927
rect 7650 3924 7656 3936
rect 7515 3896 7656 3924
rect 7515 3893 7527 3896
rect 7469 3887 7527 3893
rect 7650 3884 7656 3896
rect 7708 3884 7714 3936
rect 7745 3927 7803 3933
rect 7745 3893 7757 3927
rect 7791 3924 7803 3927
rect 7834 3924 7840 3936
rect 7791 3896 7840 3924
rect 7791 3893 7803 3896
rect 7745 3887 7803 3893
rect 7834 3884 7840 3896
rect 7892 3884 7898 3936
rect 8389 3927 8447 3933
rect 8389 3893 8401 3927
rect 8435 3924 8447 3927
rect 16574 3924 16580 3936
rect 8435 3896 16580 3924
rect 8435 3893 8447 3896
rect 8389 3887 8447 3893
rect 16574 3884 16580 3896
rect 16632 3884 16638 3936
rect 3036 3834 9844 3856
rect 3036 3782 5666 3834
rect 5718 3782 5730 3834
rect 5782 3782 5794 3834
rect 5846 3782 5858 3834
rect 5910 3782 5922 3834
rect 5974 3782 8766 3834
rect 8818 3782 8830 3834
rect 8882 3782 8894 3834
rect 8946 3782 8958 3834
rect 9010 3782 9022 3834
rect 9074 3782 9844 3834
rect 3036 3760 9844 3782
rect 4522 3720 4528 3732
rect 4483 3692 4528 3720
rect 4522 3680 4528 3692
rect 4580 3680 4586 3732
rect 4890 3720 4896 3732
rect 4851 3692 4896 3720
rect 4890 3680 4896 3692
rect 4948 3680 4954 3732
rect 8570 3680 8576 3732
rect 8628 3720 8634 3732
rect 8849 3723 8907 3729
rect 8849 3720 8861 3723
rect 8628 3692 8861 3720
rect 8628 3680 8634 3692
rect 8849 3689 8861 3692
rect 8895 3689 8907 3723
rect 8849 3683 8907 3689
rect 9217 3723 9275 3729
rect 9217 3689 9229 3723
rect 9263 3720 9275 3723
rect 9398 3720 9404 3732
rect 9263 3692 9404 3720
rect 9263 3689 9275 3692
rect 9217 3683 9275 3689
rect 9398 3680 9404 3692
rect 9456 3680 9462 3732
rect 6086 3584 6092 3596
rect 4724 3556 6092 3584
rect 4341 3519 4399 3525
rect 4341 3485 4353 3519
rect 4387 3516 4399 3519
rect 4614 3516 4620 3528
rect 4387 3488 4620 3516
rect 4387 3485 4399 3488
rect 4341 3479 4399 3485
rect 4614 3476 4620 3488
rect 4672 3476 4678 3528
rect 4724 3525 4752 3556
rect 6086 3544 6092 3556
rect 6144 3544 6150 3596
rect 6546 3584 6552 3596
rect 6507 3556 6552 3584
rect 6546 3544 6552 3556
rect 6604 3544 6610 3596
rect 4709 3519 4767 3525
rect 4709 3485 4721 3519
rect 4755 3485 4767 3519
rect 4982 3516 4988 3528
rect 4943 3488 4988 3516
rect 4709 3479 4767 3485
rect 4982 3476 4988 3488
rect 5040 3476 5046 3528
rect 6917 3519 6975 3525
rect 6917 3485 6929 3519
rect 6963 3516 6975 3519
rect 7006 3516 7012 3528
rect 6963 3488 7012 3516
rect 6963 3485 6975 3488
rect 6917 3479 6975 3485
rect 7006 3476 7012 3488
rect 7064 3476 7070 3528
rect 7926 3476 7932 3528
rect 7984 3516 7990 3528
rect 8389 3519 8447 3525
rect 8389 3516 8401 3519
rect 7984 3488 8401 3516
rect 7984 3476 7990 3488
rect 8389 3485 8401 3488
rect 8435 3485 8447 3519
rect 8389 3479 8447 3485
rect 8941 3519 8999 3525
rect 8941 3485 8953 3519
rect 8987 3516 8999 3519
rect 9490 3516 9496 3528
rect 8987 3488 9496 3516
rect 8987 3485 8999 3488
rect 8941 3479 8999 3485
rect 9490 3476 9496 3488
rect 9548 3476 9554 3528
rect 2682 3408 2688 3460
rect 2740 3448 2746 3460
rect 2740 3420 5304 3448
rect 2740 3408 2746 3420
rect 5166 3380 5172 3392
rect 5127 3352 5172 3380
rect 5166 3340 5172 3352
rect 5224 3340 5230 3392
rect 5276 3380 5304 3420
rect 7834 3408 7840 3460
rect 7892 3408 7898 3460
rect 7742 3380 7748 3392
rect 5276 3352 7748 3380
rect 7742 3340 7748 3352
rect 7800 3340 7806 3392
rect 8478 3340 8484 3392
rect 8536 3380 8542 3392
rect 8573 3383 8631 3389
rect 8573 3380 8585 3383
rect 8536 3352 8585 3380
rect 8536 3340 8542 3352
rect 8573 3349 8585 3352
rect 8619 3349 8631 3383
rect 8573 3343 8631 3349
rect 9122 3340 9128 3392
rect 9180 3380 9186 3392
rect 9401 3383 9459 3389
rect 9401 3380 9413 3383
rect 9180 3352 9413 3380
rect 9180 3340 9186 3352
rect 9401 3349 9413 3352
rect 9447 3349 9459 3383
rect 9401 3343 9459 3349
rect 3036 3290 9844 3312
rect 3036 3238 4116 3290
rect 4168 3238 4180 3290
rect 4232 3238 4244 3290
rect 4296 3238 4308 3290
rect 4360 3238 4372 3290
rect 4424 3238 7216 3290
rect 7268 3238 7280 3290
rect 7332 3238 7344 3290
rect 7396 3238 7408 3290
rect 7460 3238 7472 3290
rect 7524 3238 9844 3290
rect 3036 3216 9844 3238
rect 7837 3179 7895 3185
rect 7837 3145 7849 3179
rect 7883 3176 7895 3179
rect 7926 3176 7932 3188
rect 7883 3148 7932 3176
rect 7883 3145 7895 3148
rect 7837 3139 7895 3145
rect 7926 3136 7932 3148
rect 7984 3136 7990 3188
rect 8113 3179 8171 3185
rect 8113 3145 8125 3179
rect 8159 3145 8171 3179
rect 8386 3176 8392 3188
rect 8347 3148 8392 3176
rect 8113 3139 8171 3145
rect 5166 3068 5172 3120
rect 5224 3068 5230 3120
rect 8128 3108 8156 3139
rect 8386 3136 8392 3148
rect 8444 3136 8450 3188
rect 8662 3136 8668 3188
rect 8720 3176 8726 3188
rect 8757 3179 8815 3185
rect 8757 3176 8769 3179
rect 8720 3148 8769 3176
rect 8720 3136 8726 3148
rect 8757 3145 8769 3148
rect 8803 3145 8815 3179
rect 8757 3139 8815 3145
rect 9030 3108 9036 3120
rect 8128 3080 8340 3108
rect 8312 3052 8340 3080
rect 8588 3080 9036 3108
rect 3970 3000 3976 3052
rect 4028 3040 4034 3052
rect 4249 3043 4307 3049
rect 4249 3040 4261 3043
rect 4028 3012 4261 3040
rect 4028 3000 4034 3012
rect 4249 3009 4261 3012
rect 4295 3009 4307 3043
rect 4249 3003 4307 3009
rect 4617 3043 4675 3049
rect 4617 3009 4629 3043
rect 4663 3040 4675 3043
rect 4706 3040 4712 3052
rect 4663 3012 4712 3040
rect 4663 3009 4675 3012
rect 4617 3003 4675 3009
rect 4706 3000 4712 3012
rect 4764 3000 4770 3052
rect 6089 3043 6147 3049
rect 6089 3009 6101 3043
rect 6135 3040 6147 3043
rect 6178 3040 6184 3052
rect 6135 3012 6184 3040
rect 6135 3009 6147 3012
rect 6089 3003 6147 3009
rect 6178 3000 6184 3012
rect 6236 3000 6242 3052
rect 7650 3040 7656 3052
rect 7611 3012 7656 3040
rect 7650 3000 7656 3012
rect 7708 3000 7714 3052
rect 7929 3043 7987 3049
rect 7929 3009 7941 3043
rect 7975 3040 7987 3043
rect 8110 3040 8116 3052
rect 7975 3012 8116 3040
rect 7975 3009 7987 3012
rect 7929 3003 7987 3009
rect 8110 3000 8116 3012
rect 8168 3000 8174 3052
rect 8294 3040 8300 3052
rect 8255 3012 8300 3040
rect 8294 3000 8300 3012
rect 8352 3000 8358 3052
rect 8588 3049 8616 3080
rect 9030 3068 9036 3080
rect 9088 3068 9094 3120
rect 9674 3108 9680 3120
rect 9140 3080 9680 3108
rect 8573 3043 8631 3049
rect 8573 3009 8585 3043
rect 8619 3009 8631 3043
rect 8573 3003 8631 3009
rect 8849 3043 8907 3049
rect 8849 3009 8861 3043
rect 8895 3040 8907 3043
rect 9140 3040 9168 3080
rect 9674 3068 9680 3080
rect 9732 3068 9738 3120
rect 8895 3012 9168 3040
rect 9217 3043 9275 3049
rect 8895 3009 8907 3012
rect 8849 3003 8907 3009
rect 9217 3009 9229 3043
rect 9263 3009 9275 3043
rect 9217 3003 9275 3009
rect 6362 2932 6368 2984
rect 6420 2972 6426 2984
rect 9232 2972 9260 3003
rect 16574 2972 16580 2984
rect 6420 2944 9260 2972
rect 6420 2932 6426 2944
rect 16546 2932 16580 2972
rect 16632 2932 16638 2984
rect 6549 2907 6607 2913
rect 6549 2873 6561 2907
rect 6595 2904 6607 2907
rect 8294 2904 8300 2916
rect 6595 2876 8300 2904
rect 6595 2873 6607 2876
rect 6549 2867 6607 2873
rect 8294 2864 8300 2876
rect 8352 2864 8358 2916
rect 9033 2907 9091 2913
rect 9033 2873 9045 2907
rect 9079 2904 9091 2907
rect 16546 2904 16574 2932
rect 9079 2876 16574 2904
rect 9079 2873 9091 2876
rect 9033 2867 9091 2873
rect 9398 2836 9404 2848
rect 9359 2808 9404 2836
rect 9398 2796 9404 2808
rect 9456 2796 9462 2848
rect 3036 2746 9844 2768
rect 3036 2694 5666 2746
rect 5718 2694 5730 2746
rect 5782 2694 5794 2746
rect 5846 2694 5858 2746
rect 5910 2694 5922 2746
rect 5974 2694 8766 2746
rect 8818 2694 8830 2746
rect 8882 2694 8894 2746
rect 8946 2694 8958 2746
rect 9010 2694 9022 2746
rect 9074 2694 9844 2746
rect 3036 2672 9844 2694
rect 7926 2592 7932 2644
rect 7984 2632 7990 2644
rect 8205 2635 8263 2641
rect 8205 2632 8217 2635
rect 7984 2604 8217 2632
rect 7984 2592 7990 2604
rect 8205 2601 8217 2604
rect 8251 2601 8263 2635
rect 8205 2595 8263 2601
rect 8941 2635 8999 2641
rect 8941 2601 8953 2635
rect 8987 2632 8999 2635
rect 9214 2632 9220 2644
rect 8987 2604 9220 2632
rect 8987 2601 8999 2604
rect 8941 2595 8999 2601
rect 9214 2592 9220 2604
rect 9272 2592 9278 2644
rect 9401 2635 9459 2641
rect 9401 2601 9413 2635
rect 9447 2632 9459 2635
rect 9490 2632 9496 2644
rect 9447 2604 9496 2632
rect 9447 2601 9459 2604
rect 9401 2595 9459 2601
rect 9490 2592 9496 2604
rect 9548 2592 9554 2644
rect 8849 2567 8907 2573
rect 8849 2533 8861 2567
rect 8895 2564 8907 2567
rect 9306 2564 9312 2576
rect 8895 2536 9312 2564
rect 8895 2533 8907 2536
rect 8849 2527 8907 2533
rect 9306 2524 9312 2536
rect 9364 2524 9370 2576
rect 8294 2456 8300 2508
rect 8352 2496 8358 2508
rect 8352 2468 9260 2496
rect 8352 2456 8358 2468
rect 8665 2431 8723 2437
rect 8665 2397 8677 2431
rect 8711 2397 8723 2431
rect 9122 2428 9128 2440
rect 9083 2400 9128 2428
rect 8665 2391 8723 2397
rect 8573 2363 8631 2369
rect 8573 2329 8585 2363
rect 8619 2360 8631 2363
rect 8680 2360 8708 2391
rect 9122 2388 9128 2400
rect 9180 2388 9186 2440
rect 9232 2437 9260 2468
rect 9217 2431 9275 2437
rect 9217 2397 9229 2431
rect 9263 2397 9275 2431
rect 9217 2391 9275 2397
rect 16574 2360 16580 2372
rect 8619 2332 16580 2360
rect 8619 2329 8631 2332
rect 8573 2323 8631 2329
rect 16574 2320 16580 2332
rect 16632 2320 16638 2372
rect 3036 2202 9844 2224
rect 3036 2150 4116 2202
rect 4168 2150 4180 2202
rect 4232 2150 4244 2202
rect 4296 2150 4308 2202
rect 4360 2150 4372 2202
rect 4424 2150 7216 2202
rect 7268 2150 7280 2202
rect 7332 2150 7344 2202
rect 7396 2150 7408 2202
rect 7460 2150 7472 2202
rect 7524 2150 9844 2202
rect 3036 2128 9844 2150
rect 8202 2048 8208 2100
rect 8260 2088 8266 2100
rect 9309 2091 9367 2097
rect 9309 2088 9321 2091
rect 8260 2060 9321 2088
rect 8260 2048 8266 2060
rect 9309 2057 9321 2060
rect 9355 2057 9367 2091
rect 9309 2051 9367 2057
rect 8849 1955 8907 1961
rect 8849 1921 8861 1955
rect 8895 1952 8907 1955
rect 9493 1955 9551 1961
rect 9493 1952 9505 1955
rect 8895 1924 9505 1952
rect 8895 1921 8907 1924
rect 8849 1915 8907 1921
rect 9493 1921 9505 1924
rect 9539 1952 9551 1955
rect 9539 1924 16574 1952
rect 9539 1921 9551 1924
rect 9493 1915 9551 1921
rect 7834 1844 7840 1896
rect 7892 1884 7898 1896
rect 8941 1887 8999 1893
rect 8941 1884 8953 1887
rect 7892 1856 8953 1884
rect 7892 1844 7898 1856
rect 8941 1853 8953 1856
rect 8987 1884 8999 1887
rect 9214 1884 9220 1896
rect 8987 1856 9220 1884
rect 8987 1853 8999 1856
rect 8941 1847 8999 1853
rect 9214 1844 9220 1856
rect 9272 1844 9278 1896
rect 16546 1828 16574 1924
rect 16546 1788 16580 1828
rect 16574 1776 16580 1788
rect 16632 1776 16638 1828
rect 9122 1748 9128 1760
rect 9083 1720 9128 1748
rect 9122 1708 9128 1720
rect 9180 1708 9186 1760
rect 3036 1658 9844 1680
rect 3036 1606 5666 1658
rect 5718 1606 5730 1658
rect 5782 1606 5794 1658
rect 5846 1606 5858 1658
rect 5910 1606 5922 1658
rect 5974 1606 8766 1658
rect 8818 1606 8830 1658
rect 8882 1606 8894 1658
rect 8946 1606 8958 1658
rect 9010 1606 9022 1658
rect 9074 1606 9844 1658
rect 3036 1584 9844 1606
rect 3036 1114 9844 1136
rect 3036 1062 4116 1114
rect 4168 1062 4180 1114
rect 4232 1062 4244 1114
rect 4296 1062 4308 1114
rect 4360 1062 4372 1114
rect 4424 1062 7216 1114
rect 7268 1062 7280 1114
rect 7332 1062 7344 1114
rect 7396 1062 7408 1114
rect 7460 1062 7472 1114
rect 7524 1062 9844 1114
rect 3036 1040 9844 1062
<< via1 >>
rect 6184 12248 6236 12300
rect 6552 12180 6604 12232
rect 1952 12112 2004 12164
rect 8392 12112 8444 12164
rect 1768 12044 1820 12096
rect 6000 12044 6052 12096
rect 3884 11976 3936 12028
rect 6460 11976 6512 12028
rect 7840 11976 7892 12028
rect 1308 11908 1360 11960
rect 4620 11908 4672 11960
rect 4712 11908 4764 11960
rect 2136 11772 2188 11824
rect 5540 11840 5592 11892
rect 6000 11840 6052 11892
rect 3056 11772 3108 11824
rect 9220 11772 9272 11824
rect 940 11704 992 11756
rect 4344 11704 4396 11756
rect 6092 11747 6144 11756
rect 6092 11713 6101 11747
rect 6101 11713 6135 11747
rect 6135 11713 6144 11747
rect 6092 11704 6144 11713
rect 7656 11704 7708 11756
rect 3148 11636 3200 11688
rect 7564 11636 7616 11688
rect 7748 11636 7800 11688
rect 9128 11636 9180 11688
rect 1124 11568 1176 11620
rect 2780 11568 2832 11620
rect 3240 11568 3292 11620
rect 6276 11568 6328 11620
rect 7196 11568 7248 11620
rect 9312 11568 9364 11620
rect 2044 11500 2096 11552
rect 2320 11500 2372 11552
rect 3608 11500 3660 11552
rect 8668 11500 8720 11552
rect 2566 11398 2618 11450
rect 2630 11398 2682 11450
rect 2694 11398 2746 11450
rect 2758 11398 2810 11450
rect 2822 11398 2874 11450
rect 5666 11398 5718 11450
rect 5730 11398 5782 11450
rect 5794 11398 5846 11450
rect 5858 11398 5910 11450
rect 5922 11398 5974 11450
rect 8766 11398 8818 11450
rect 8830 11398 8882 11450
rect 8894 11398 8946 11450
rect 8958 11398 9010 11450
rect 9022 11398 9074 11450
rect 1676 11296 1728 11348
rect 2044 11339 2096 11348
rect 2044 11305 2053 11339
rect 2053 11305 2087 11339
rect 2087 11305 2096 11339
rect 2044 11296 2096 11305
rect 2320 11339 2372 11348
rect 2320 11305 2329 11339
rect 2329 11305 2363 11339
rect 2363 11305 2372 11339
rect 2320 11296 2372 11305
rect 3148 11339 3200 11348
rect 3148 11305 3157 11339
rect 3157 11305 3191 11339
rect 3191 11305 3200 11339
rect 3148 11296 3200 11305
rect 4436 11296 4488 11348
rect 3608 11228 3660 11280
rect 3700 11228 3752 11280
rect 4344 11271 4396 11280
rect 4344 11237 4353 11271
rect 4353 11237 4387 11271
rect 4387 11237 4396 11271
rect 4344 11228 4396 11237
rect 1584 11160 1636 11212
rect 940 11092 992 11144
rect 1492 11135 1544 11144
rect 1492 11101 1501 11135
rect 1501 11101 1535 11135
rect 1535 11101 1544 11135
rect 1492 11092 1544 11101
rect 1768 11092 1820 11144
rect 2136 11135 2188 11144
rect 2136 11101 2145 11135
rect 2145 11101 2179 11135
rect 2179 11101 2188 11135
rect 2136 11092 2188 11101
rect 2596 11092 2648 11144
rect 2780 11092 2832 11144
rect 3516 11160 3568 11212
rect 2320 11024 2372 11076
rect 3240 11111 3292 11120
rect 3240 11077 3249 11111
rect 3249 11077 3283 11111
rect 3283 11077 3292 11111
rect 6000 11339 6052 11348
rect 6000 11305 6009 11339
rect 6009 11305 6043 11339
rect 6043 11305 6052 11339
rect 6000 11296 6052 11305
rect 6276 11339 6328 11348
rect 6276 11305 6285 11339
rect 6285 11305 6319 11339
rect 6319 11305 6328 11339
rect 6276 11296 6328 11305
rect 6644 11339 6696 11348
rect 6644 11305 6653 11339
rect 6653 11305 6687 11339
rect 6687 11305 6696 11339
rect 6644 11296 6696 11305
rect 7748 11296 7800 11348
rect 8208 11296 8260 11348
rect 8484 11228 8536 11280
rect 13820 11228 13872 11280
rect 4712 11135 4764 11144
rect 4712 11101 4721 11135
rect 4721 11101 4755 11135
rect 4755 11101 4764 11135
rect 4988 11135 5040 11144
rect 4712 11092 4764 11101
rect 4988 11101 4997 11135
rect 4997 11101 5031 11135
rect 5031 11101 5040 11135
rect 4988 11092 5040 11101
rect 5264 11092 5316 11144
rect 3240 11068 3292 11077
rect 2780 10956 2832 11008
rect 3056 10956 3108 11008
rect 4436 11024 4488 11076
rect 5632 11024 5684 11076
rect 5908 11092 5960 11144
rect 6092 11092 6144 11144
rect 7104 11135 7156 11144
rect 7104 11101 7113 11135
rect 7113 11101 7147 11135
rect 7147 11101 7156 11135
rect 7104 11092 7156 11101
rect 7196 11024 7248 11076
rect 3792 10956 3844 11008
rect 3976 10999 4028 11008
rect 3976 10965 3985 10999
rect 3985 10965 4019 10999
rect 4019 10965 4028 10999
rect 3976 10956 4028 10965
rect 4804 10999 4856 11008
rect 4804 10965 4813 10999
rect 4813 10965 4847 10999
rect 4847 10965 4856 10999
rect 4804 10956 4856 10965
rect 4896 10956 4948 11008
rect 5908 10956 5960 11008
rect 6644 10956 6696 11008
rect 7012 10999 7064 11008
rect 7012 10965 7021 10999
rect 7021 10965 7055 10999
rect 7055 10965 7064 10999
rect 7012 10956 7064 10965
rect 8392 11160 8444 11212
rect 8300 11135 8352 11144
rect 8300 11101 8309 11135
rect 8309 11101 8343 11135
rect 8343 11101 8352 11135
rect 8300 11092 8352 11101
rect 8392 11024 8444 11076
rect 13728 11160 13780 11212
rect 8668 11092 8720 11144
rect 9220 11135 9272 11144
rect 9220 11101 9229 11135
rect 9229 11101 9263 11135
rect 9263 11101 9272 11135
rect 9220 11092 9272 11101
rect 9404 10999 9456 11008
rect 9404 10965 9413 10999
rect 9413 10965 9447 10999
rect 9447 10965 9456 10999
rect 9404 10956 9456 10965
rect 4116 10854 4168 10906
rect 4180 10854 4232 10906
rect 4244 10854 4296 10906
rect 4308 10854 4360 10906
rect 4372 10854 4424 10906
rect 7216 10854 7268 10906
rect 7280 10854 7332 10906
rect 7344 10854 7396 10906
rect 7408 10854 7460 10906
rect 7472 10854 7524 10906
rect 1584 10752 1636 10804
rect 1308 10684 1360 10736
rect 1216 10659 1268 10668
rect 1216 10625 1225 10659
rect 1225 10625 1259 10659
rect 1259 10625 1268 10659
rect 1216 10616 1268 10625
rect 1400 10616 1452 10668
rect 2136 10616 2188 10668
rect 2320 10659 2372 10668
rect 2320 10625 2329 10659
rect 2329 10625 2363 10659
rect 2363 10625 2372 10659
rect 2320 10616 2372 10625
rect 3884 10752 3936 10804
rect 4988 10752 5040 10804
rect 5632 10752 5684 10804
rect 2964 10616 3016 10668
rect 3240 10616 3292 10668
rect 2136 10480 2188 10532
rect 1952 10455 2004 10464
rect 1952 10421 1961 10455
rect 1961 10421 1995 10455
rect 1995 10421 2004 10455
rect 1952 10412 2004 10421
rect 2320 10412 2372 10464
rect 2412 10412 2464 10464
rect 3148 10548 3200 10600
rect 3424 10480 3476 10532
rect 3976 10684 4028 10736
rect 7104 10752 7156 10804
rect 8576 10727 8628 10736
rect 3884 10659 3936 10668
rect 3884 10625 3893 10659
rect 3893 10625 3927 10659
rect 3927 10625 3936 10659
rect 3884 10616 3936 10625
rect 4896 10616 4948 10668
rect 5356 10659 5408 10668
rect 3608 10412 3660 10464
rect 3792 10455 3844 10464
rect 3792 10421 3801 10455
rect 3801 10421 3835 10455
rect 3835 10421 3844 10455
rect 3792 10412 3844 10421
rect 4160 10480 4212 10532
rect 5356 10625 5365 10659
rect 5365 10625 5399 10659
rect 5399 10625 5408 10659
rect 5356 10616 5408 10625
rect 5540 10616 5592 10668
rect 5264 10548 5316 10600
rect 5908 10616 5960 10668
rect 8576 10693 8585 10727
rect 8585 10693 8619 10727
rect 8619 10693 8628 10727
rect 8576 10684 8628 10693
rect 7564 10616 7616 10668
rect 8208 10616 8260 10668
rect 6092 10548 6144 10600
rect 6828 10548 6880 10600
rect 8116 10548 8168 10600
rect 4528 10412 4580 10464
rect 5264 10455 5316 10464
rect 5264 10421 5273 10455
rect 5273 10421 5307 10455
rect 5307 10421 5316 10455
rect 5264 10412 5316 10421
rect 5540 10455 5592 10464
rect 5540 10421 5549 10455
rect 5549 10421 5583 10455
rect 5583 10421 5592 10455
rect 5540 10412 5592 10421
rect 7840 10480 7892 10532
rect 7932 10412 7984 10464
rect 8668 10412 8720 10464
rect 16580 10412 16632 10464
rect 2566 10310 2618 10362
rect 2630 10310 2682 10362
rect 2694 10310 2746 10362
rect 2758 10310 2810 10362
rect 2822 10310 2874 10362
rect 5666 10310 5718 10362
rect 5730 10310 5782 10362
rect 5794 10310 5846 10362
rect 5858 10310 5910 10362
rect 5922 10310 5974 10362
rect 8766 10310 8818 10362
rect 8830 10310 8882 10362
rect 8894 10310 8946 10362
rect 8958 10310 9010 10362
rect 9022 10310 9074 10362
rect 1308 10251 1360 10260
rect 1308 10217 1317 10251
rect 1317 10217 1351 10251
rect 1351 10217 1360 10251
rect 1308 10208 1360 10217
rect 7932 10251 7984 10260
rect 7932 10217 7941 10251
rect 7941 10217 7975 10251
rect 7975 10217 7984 10251
rect 7932 10208 7984 10217
rect 8208 10251 8260 10260
rect 8208 10217 8217 10251
rect 8217 10217 8251 10251
rect 8251 10217 8260 10251
rect 8208 10208 8260 10217
rect 1400 10047 1452 10056
rect 1400 10013 1409 10047
rect 1409 10013 1443 10047
rect 1443 10013 1452 10047
rect 1400 10004 1452 10013
rect 2504 10072 2556 10124
rect 3608 10140 3660 10192
rect 5540 10140 5592 10192
rect 6460 10140 6512 10192
rect 7840 10140 7892 10192
rect 4528 10072 4580 10124
rect 6920 10072 6972 10124
rect 7104 10072 7156 10124
rect 3700 10047 3752 10056
rect 3700 10013 3709 10047
rect 3709 10013 3743 10047
rect 3743 10013 3752 10047
rect 3700 10004 3752 10013
rect 3976 10004 4028 10056
rect 4988 10004 5040 10056
rect 9496 10047 9548 10056
rect 3148 9979 3200 9988
rect 3148 9945 3157 9979
rect 3157 9945 3191 9979
rect 3191 9945 3200 9979
rect 3148 9936 3200 9945
rect 3424 9936 3476 9988
rect 3608 9936 3660 9988
rect 4804 9936 4856 9988
rect 2228 9868 2280 9920
rect 2504 9868 2556 9920
rect 6828 9868 6880 9920
rect 7472 9936 7524 9988
rect 9496 10013 9505 10047
rect 9505 10013 9539 10047
rect 9539 10013 9548 10047
rect 9496 10004 9548 10013
rect 8208 9868 8260 9920
rect 8576 9911 8628 9920
rect 8576 9877 8585 9911
rect 8585 9877 8619 9911
rect 8619 9877 8628 9911
rect 8576 9868 8628 9877
rect 8852 9868 8904 9920
rect 10876 9868 10928 9920
rect 4116 9766 4168 9818
rect 4180 9766 4232 9818
rect 4244 9766 4296 9818
rect 4308 9766 4360 9818
rect 4372 9766 4424 9818
rect 7216 9766 7268 9818
rect 7280 9766 7332 9818
rect 7344 9766 7396 9818
rect 7408 9766 7460 9818
rect 7472 9766 7524 9818
rect 1308 9639 1360 9648
rect 1308 9605 1317 9639
rect 1317 9605 1351 9639
rect 1351 9605 1360 9639
rect 1308 9596 1360 9605
rect 2964 9664 3016 9716
rect 3148 9664 3200 9716
rect 2688 9596 2740 9648
rect 1032 9528 1084 9580
rect 1860 9528 1912 9580
rect 2044 9528 2096 9580
rect 2136 9528 2188 9580
rect 1676 9392 1728 9444
rect 2044 9324 2096 9376
rect 2596 9528 2648 9580
rect 3424 9596 3476 9648
rect 5264 9664 5316 9716
rect 8024 9664 8076 9716
rect 8484 9596 8536 9648
rect 8852 9596 8904 9648
rect 9404 9596 9456 9648
rect 4620 9571 4672 9580
rect 4620 9537 4629 9571
rect 4629 9537 4663 9571
rect 4663 9537 4672 9571
rect 4620 9528 4672 9537
rect 4896 9528 4948 9580
rect 4712 9460 4764 9512
rect 6000 9571 6052 9580
rect 6000 9537 6009 9571
rect 6009 9537 6043 9571
rect 6043 9537 6052 9571
rect 6000 9528 6052 9537
rect 6828 9571 6880 9580
rect 6828 9537 6837 9571
rect 6837 9537 6871 9571
rect 6871 9537 6880 9571
rect 6828 9528 6880 9537
rect 5724 9460 5776 9512
rect 7012 9528 7064 9580
rect 3884 9324 3936 9376
rect 5264 9392 5316 9444
rect 5540 9392 5592 9444
rect 7656 9528 7708 9580
rect 7564 9503 7616 9512
rect 7564 9469 7573 9503
rect 7573 9469 7607 9503
rect 7607 9469 7616 9503
rect 7564 9460 7616 9469
rect 8484 9392 8536 9444
rect 6368 9324 6420 9376
rect 7196 9324 7248 9376
rect 2566 9222 2618 9274
rect 2630 9222 2682 9274
rect 2694 9222 2746 9274
rect 2758 9222 2810 9274
rect 2822 9222 2874 9274
rect 5666 9222 5718 9274
rect 5730 9222 5782 9274
rect 5794 9222 5846 9274
rect 5858 9222 5910 9274
rect 5922 9222 5974 9274
rect 8766 9222 8818 9274
rect 8830 9222 8882 9274
rect 8894 9222 8946 9274
rect 8958 9222 9010 9274
rect 9022 9222 9074 9274
rect 1216 9163 1268 9172
rect 1216 9129 1225 9163
rect 1225 9129 1259 9163
rect 1259 9129 1268 9163
rect 1216 9120 1268 9129
rect 3148 9120 3200 9172
rect 3424 9163 3476 9172
rect 3424 9129 3433 9163
rect 3433 9129 3467 9163
rect 3467 9129 3476 9163
rect 3424 9120 3476 9129
rect 4344 9120 4396 9172
rect 4620 9163 4672 9172
rect 4620 9129 4629 9163
rect 4629 9129 4663 9163
rect 4663 9129 4672 9163
rect 4620 9120 4672 9129
rect 3608 9052 3660 9104
rect 2320 8984 2372 9036
rect 4436 9052 4488 9104
rect 4712 9052 4764 9104
rect 1124 8848 1176 8900
rect 1952 8959 2004 8968
rect 1952 8925 1961 8959
rect 1961 8925 1995 8959
rect 1995 8925 2004 8959
rect 1952 8916 2004 8925
rect 2136 8959 2188 8968
rect 2136 8925 2145 8959
rect 2145 8925 2179 8959
rect 2179 8925 2188 8959
rect 2136 8916 2188 8925
rect 2412 8959 2464 8968
rect 2412 8925 2421 8959
rect 2421 8925 2455 8959
rect 2455 8925 2464 8959
rect 2412 8916 2464 8925
rect 1584 8848 1636 8900
rect 4896 8984 4948 9036
rect 2412 8780 2464 8832
rect 3056 8916 3108 8968
rect 3240 8959 3292 8968
rect 3240 8925 3249 8959
rect 3249 8925 3283 8959
rect 3283 8925 3292 8959
rect 3240 8916 3292 8925
rect 3424 8916 3476 8968
rect 3792 8916 3844 8968
rect 7196 9120 7248 9172
rect 9312 9120 9364 9172
rect 13820 9120 13872 9172
rect 16672 9120 16724 9172
rect 8760 9052 8812 9104
rect 9404 9052 9456 9104
rect 6828 8984 6880 9036
rect 7104 8984 7156 9036
rect 4344 8891 4396 8900
rect 4344 8857 4353 8891
rect 4353 8857 4387 8891
rect 4387 8857 4396 8891
rect 4344 8848 4396 8857
rect 4436 8848 4488 8900
rect 3056 8780 3108 8832
rect 4988 8780 5040 8832
rect 5080 8823 5132 8832
rect 5080 8789 5089 8823
rect 5089 8789 5123 8823
rect 5123 8789 5132 8823
rect 5908 8848 5960 8900
rect 6644 8848 6696 8900
rect 8116 8916 8168 8968
rect 8576 8959 8628 8968
rect 8576 8925 8585 8959
rect 8585 8925 8619 8959
rect 8619 8925 8628 8959
rect 9220 8959 9272 8968
rect 8576 8916 8628 8925
rect 7196 8848 7248 8900
rect 7564 8848 7616 8900
rect 7748 8848 7800 8900
rect 8760 8891 8812 8900
rect 5080 8780 5132 8789
rect 8760 8857 8769 8891
rect 8769 8857 8803 8891
rect 8803 8857 8812 8891
rect 8760 8848 8812 8857
rect 9220 8925 9229 8959
rect 9229 8925 9263 8959
rect 9263 8925 9272 8959
rect 9220 8916 9272 8925
rect 9312 8848 9364 8900
rect 9404 8823 9456 8832
rect 9404 8789 9413 8823
rect 9413 8789 9447 8823
rect 9447 8789 9456 8823
rect 9404 8780 9456 8789
rect 4116 8678 4168 8730
rect 4180 8678 4232 8730
rect 4244 8678 4296 8730
rect 4308 8678 4360 8730
rect 4372 8678 4424 8730
rect 7216 8678 7268 8730
rect 7280 8678 7332 8730
rect 7344 8678 7396 8730
rect 7408 8678 7460 8730
rect 7472 8678 7524 8730
rect 1216 8619 1268 8628
rect 1216 8585 1225 8619
rect 1225 8585 1259 8619
rect 1259 8585 1268 8619
rect 1216 8576 1268 8585
rect 1308 8576 1360 8628
rect 7840 8576 7892 8628
rect 9496 8619 9548 8628
rect 9496 8585 9505 8619
rect 9505 8585 9539 8619
rect 9539 8585 9548 8619
rect 9496 8576 9548 8585
rect 2228 8508 2280 8560
rect 4528 8508 4580 8560
rect 5724 8508 5776 8560
rect 6736 8551 6788 8560
rect 6736 8517 6745 8551
rect 6745 8517 6779 8551
rect 6779 8517 6788 8551
rect 6736 8508 6788 8517
rect 6828 8508 6880 8560
rect 8024 8508 8076 8560
rect 2044 8483 2096 8492
rect 2044 8449 2053 8483
rect 2053 8449 2087 8483
rect 2087 8449 2096 8483
rect 2044 8440 2096 8449
rect 4160 8483 4212 8492
rect 4160 8449 4169 8483
rect 4169 8449 4203 8483
rect 4203 8449 4212 8483
rect 4160 8440 4212 8449
rect 5540 8440 5592 8492
rect 6644 8440 6696 8492
rect 2136 8372 2188 8424
rect 2320 8415 2372 8424
rect 2320 8381 2329 8415
rect 2329 8381 2363 8415
rect 2363 8381 2372 8415
rect 2320 8372 2372 8381
rect 3792 8372 3844 8424
rect 3976 8372 4028 8424
rect 4528 8372 4580 8424
rect 4804 8372 4856 8424
rect 9128 8440 9180 8492
rect 7564 8415 7616 8424
rect 1952 8347 2004 8356
rect 1952 8313 1961 8347
rect 1961 8313 1995 8347
rect 1995 8313 2004 8347
rect 1952 8304 2004 8313
rect 5540 8304 5592 8356
rect 5908 8347 5960 8356
rect 5908 8313 5917 8347
rect 5917 8313 5951 8347
rect 5951 8313 5960 8347
rect 5908 8304 5960 8313
rect 1308 8236 1360 8288
rect 1860 8236 1912 8288
rect 2228 8279 2280 8288
rect 2228 8245 2237 8279
rect 2237 8245 2271 8279
rect 2271 8245 2280 8279
rect 2228 8236 2280 8245
rect 2412 8236 2464 8288
rect 6552 8279 6604 8288
rect 6552 8245 6561 8279
rect 6561 8245 6595 8279
rect 6595 8245 6604 8279
rect 6552 8236 6604 8245
rect 6920 8304 6972 8356
rect 7564 8381 7573 8415
rect 7573 8381 7607 8415
rect 7607 8381 7616 8415
rect 7564 8372 7616 8381
rect 9128 8236 9180 8288
rect 2566 8134 2618 8186
rect 2630 8134 2682 8186
rect 2694 8134 2746 8186
rect 2758 8134 2810 8186
rect 2822 8134 2874 8186
rect 5666 8134 5718 8186
rect 5730 8134 5782 8186
rect 5794 8134 5846 8186
rect 5858 8134 5910 8186
rect 5922 8134 5974 8186
rect 8766 8134 8818 8186
rect 8830 8134 8882 8186
rect 8894 8134 8946 8186
rect 8958 8134 9010 8186
rect 9022 8134 9074 8186
rect 1584 8007 1636 8016
rect 1584 7973 1593 8007
rect 1593 7973 1627 8007
rect 1627 7973 1636 8007
rect 1584 7964 1636 7973
rect 3424 8032 3476 8084
rect 3792 7964 3844 8016
rect 4068 8032 4120 8084
rect 5172 8032 5224 8084
rect 2412 7896 2464 7948
rect 4160 7896 4212 7948
rect 6552 7964 6604 8016
rect 8116 7964 8168 8016
rect 5540 7939 5592 7948
rect 5540 7905 5549 7939
rect 5549 7905 5583 7939
rect 5583 7905 5592 7939
rect 5540 7896 5592 7905
rect 3516 7828 3568 7880
rect 3792 7828 3844 7880
rect 6000 7896 6052 7948
rect 9588 7964 9640 8016
rect 8208 7871 8260 7880
rect 1492 7760 1544 7812
rect 2688 7760 2740 7812
rect 3976 7760 4028 7812
rect 1676 7735 1728 7744
rect 1676 7701 1685 7735
rect 1685 7701 1719 7735
rect 1719 7701 1728 7735
rect 1676 7692 1728 7701
rect 1860 7692 1912 7744
rect 5172 7760 5224 7812
rect 6276 7760 6328 7812
rect 6920 7760 6972 7812
rect 7748 7803 7800 7812
rect 7748 7769 7757 7803
rect 7757 7769 7791 7803
rect 7791 7769 7800 7803
rect 7748 7760 7800 7769
rect 6184 7692 6236 7744
rect 6368 7692 6420 7744
rect 7656 7692 7708 7744
rect 7932 7735 7984 7744
rect 7932 7701 7941 7735
rect 7941 7701 7975 7735
rect 7975 7701 7984 7735
rect 7932 7692 7984 7701
rect 8208 7837 8217 7871
rect 8217 7837 8251 7871
rect 8251 7837 8260 7871
rect 8208 7828 8260 7837
rect 8116 7760 8168 7812
rect 8576 7871 8628 7880
rect 8576 7837 8585 7871
rect 8585 7837 8619 7871
rect 8619 7837 8628 7871
rect 8576 7828 8628 7837
rect 8484 7760 8536 7812
rect 9036 7871 9088 7880
rect 9036 7837 9045 7871
rect 9045 7837 9079 7871
rect 9079 7837 9088 7871
rect 9036 7828 9088 7837
rect 8392 7735 8444 7744
rect 8392 7701 8401 7735
rect 8401 7701 8435 7735
rect 8435 7701 8444 7735
rect 8392 7692 8444 7701
rect 12256 7692 12308 7744
rect 4116 7590 4168 7642
rect 4180 7590 4232 7642
rect 4244 7590 4296 7642
rect 4308 7590 4360 7642
rect 4372 7590 4424 7642
rect 7216 7590 7268 7642
rect 7280 7590 7332 7642
rect 7344 7590 7396 7642
rect 7408 7590 7460 7642
rect 7472 7590 7524 7642
rect 1308 7531 1360 7540
rect 1308 7497 1317 7531
rect 1317 7497 1351 7531
rect 1351 7497 1360 7531
rect 1308 7488 1360 7497
rect 2044 7488 2096 7540
rect 2320 7531 2372 7540
rect 2320 7497 2329 7531
rect 2329 7497 2363 7531
rect 2363 7497 2372 7531
rect 2320 7488 2372 7497
rect 4804 7488 4856 7540
rect 3884 7420 3936 7472
rect 7104 7488 7156 7540
rect 7564 7488 7616 7540
rect 8208 7531 8260 7540
rect 8208 7497 8217 7531
rect 8217 7497 8251 7531
rect 8251 7497 8260 7531
rect 8208 7488 8260 7497
rect 9128 7488 9180 7540
rect 9220 7488 9272 7540
rect 1768 7352 1820 7404
rect 2228 7352 2280 7404
rect 2780 7352 2832 7404
rect 5264 7352 5316 7404
rect 1860 7284 1912 7336
rect 6184 7395 6236 7404
rect 2136 7191 2188 7200
rect 2136 7157 2145 7191
rect 2145 7157 2179 7191
rect 2179 7157 2188 7191
rect 2136 7148 2188 7157
rect 3884 7216 3936 7268
rect 6184 7361 6193 7395
rect 6193 7361 6227 7395
rect 6227 7361 6236 7395
rect 6184 7352 6236 7361
rect 6828 7420 6880 7472
rect 7288 7420 7340 7472
rect 6368 7284 6420 7336
rect 7104 7284 7156 7336
rect 7196 7284 7248 7336
rect 9496 7352 9548 7404
rect 8668 7284 8720 7336
rect 6092 7216 6144 7268
rect 6276 7216 6328 7268
rect 6184 7148 6236 7200
rect 6460 7148 6512 7200
rect 11060 7148 11112 7200
rect 2566 7046 2618 7098
rect 2630 7046 2682 7098
rect 2694 7046 2746 7098
rect 2758 7046 2810 7098
rect 2822 7046 2874 7098
rect 5666 7046 5718 7098
rect 5730 7046 5782 7098
rect 5794 7046 5846 7098
rect 5858 7046 5910 7098
rect 5922 7046 5974 7098
rect 8766 7046 8818 7098
rect 8830 7046 8882 7098
rect 8894 7046 8946 7098
rect 8958 7046 9010 7098
rect 9022 7046 9074 7098
rect 1032 6944 1084 6996
rect 2320 6944 2372 6996
rect 3332 6944 3384 6996
rect 3700 6944 3752 6996
rect 6368 6987 6420 6996
rect 6368 6953 6377 6987
rect 6377 6953 6411 6987
rect 6411 6953 6420 6987
rect 6368 6944 6420 6953
rect 7196 6944 7248 6996
rect 7748 6944 7800 6996
rect 8208 6944 8260 6996
rect 8576 6944 8628 6996
rect 2320 6808 2372 6860
rect 2596 6808 2648 6860
rect 1400 6783 1452 6792
rect 1400 6749 1409 6783
rect 1409 6749 1443 6783
rect 1443 6749 1452 6783
rect 1400 6740 1452 6749
rect 3056 6740 3108 6792
rect 1676 6672 1728 6724
rect 3700 6808 3752 6860
rect 6276 6876 6328 6928
rect 6644 6876 6696 6928
rect 3424 6740 3476 6792
rect 2596 6604 2648 6656
rect 2688 6604 2740 6656
rect 3424 6647 3476 6656
rect 3424 6613 3433 6647
rect 3433 6613 3467 6647
rect 3467 6613 3476 6647
rect 3424 6604 3476 6613
rect 4712 6672 4764 6724
rect 6092 6740 6144 6792
rect 6552 6808 6604 6860
rect 6828 6808 6880 6860
rect 8668 6808 8720 6860
rect 6920 6740 6972 6792
rect 7196 6740 7248 6792
rect 9128 6740 9180 6792
rect 6000 6647 6052 6656
rect 6000 6613 6009 6647
rect 6009 6613 6043 6647
rect 6043 6613 6052 6647
rect 6000 6604 6052 6613
rect 6644 6604 6696 6656
rect 6920 6604 6972 6656
rect 8668 6672 8720 6724
rect 8116 6604 8168 6656
rect 9128 6647 9180 6656
rect 9128 6613 9137 6647
rect 9137 6613 9171 6647
rect 9171 6613 9180 6647
rect 9128 6604 9180 6613
rect 9220 6647 9272 6656
rect 9220 6613 9229 6647
rect 9229 6613 9263 6647
rect 9263 6613 9272 6647
rect 9220 6604 9272 6613
rect 4116 6502 4168 6554
rect 4180 6502 4232 6554
rect 4244 6502 4296 6554
rect 4308 6502 4360 6554
rect 4372 6502 4424 6554
rect 7216 6502 7268 6554
rect 7280 6502 7332 6554
rect 7344 6502 7396 6554
rect 7408 6502 7460 6554
rect 7472 6502 7524 6554
rect 2412 6400 2464 6452
rect 3056 6400 3108 6452
rect 4804 6400 4856 6452
rect 1124 6332 1176 6384
rect 2688 6375 2740 6384
rect 2688 6341 2697 6375
rect 2697 6341 2731 6375
rect 2731 6341 2740 6375
rect 2688 6332 2740 6341
rect 2320 6264 2372 6316
rect 1584 6196 1636 6248
rect 9128 6400 9180 6452
rect 6736 6332 6788 6384
rect 6828 6332 6880 6384
rect 9312 6332 9364 6384
rect 5908 6264 5960 6316
rect 8484 6264 8536 6316
rect 5540 6196 5592 6248
rect 7196 6239 7248 6248
rect 7196 6205 7205 6239
rect 7205 6205 7239 6239
rect 7239 6205 7248 6239
rect 7196 6196 7248 6205
rect 6460 6128 6512 6180
rect 3976 6060 4028 6112
rect 4988 6060 5040 6112
rect 6368 6103 6420 6112
rect 6368 6069 6377 6103
rect 6377 6069 6411 6103
rect 6411 6069 6420 6103
rect 6368 6060 6420 6069
rect 6828 6060 6880 6112
rect 9128 6103 9180 6112
rect 9128 6069 9137 6103
rect 9137 6069 9171 6103
rect 9171 6069 9180 6103
rect 9128 6060 9180 6069
rect 9404 6103 9456 6112
rect 9404 6069 9413 6103
rect 9413 6069 9447 6103
rect 9447 6069 9456 6103
rect 9404 6060 9456 6069
rect 2566 5958 2618 6010
rect 2630 5958 2682 6010
rect 2694 5958 2746 6010
rect 2758 5958 2810 6010
rect 2822 5958 2874 6010
rect 5666 5958 5718 6010
rect 5730 5958 5782 6010
rect 5794 5958 5846 6010
rect 5858 5958 5910 6010
rect 5922 5958 5974 6010
rect 8766 5958 8818 6010
rect 8830 5958 8882 6010
rect 8894 5958 8946 6010
rect 8958 5958 9010 6010
rect 9022 5958 9074 6010
rect 3700 5856 3752 5908
rect 3792 5899 3844 5908
rect 3792 5865 3801 5899
rect 3801 5865 3835 5899
rect 3835 5865 3844 5899
rect 3792 5856 3844 5865
rect 1400 5788 1452 5840
rect 3332 5720 3384 5772
rect 7012 5856 7064 5908
rect 7196 5856 7248 5908
rect 7564 5856 7616 5908
rect 9312 5899 9364 5908
rect 9312 5865 9321 5899
rect 9321 5865 9355 5899
rect 9355 5865 9364 5899
rect 9312 5856 9364 5865
rect 9496 5788 9548 5840
rect 6552 5720 6604 5772
rect 6644 5720 6696 5772
rect 2136 5584 2188 5636
rect 3148 5652 3200 5704
rect 7656 5652 7708 5704
rect 8668 5652 8720 5704
rect 3056 5584 3108 5636
rect 3792 5584 3844 5636
rect 4988 5584 5040 5636
rect 4712 5516 4764 5568
rect 6184 5584 6236 5636
rect 6736 5516 6788 5568
rect 9036 5584 9088 5636
rect 9312 5584 9364 5636
rect 8024 5516 8076 5568
rect 9128 5516 9180 5568
rect 4116 5414 4168 5466
rect 4180 5414 4232 5466
rect 4244 5414 4296 5466
rect 4308 5414 4360 5466
rect 4372 5414 4424 5466
rect 7216 5414 7268 5466
rect 7280 5414 7332 5466
rect 7344 5414 7396 5466
rect 7408 5414 7460 5466
rect 7472 5414 7524 5466
rect 3792 5312 3844 5364
rect 4620 5312 4672 5364
rect 5448 5312 5500 5364
rect 3332 5219 3384 5228
rect 3332 5185 3341 5219
rect 3341 5185 3375 5219
rect 3375 5185 3384 5219
rect 3332 5176 3384 5185
rect 6000 5312 6052 5364
rect 6920 5244 6972 5296
rect 3976 5108 4028 5160
rect 5540 5108 5592 5160
rect 6000 5176 6052 5228
rect 6184 5219 6236 5228
rect 6184 5185 6193 5219
rect 6193 5185 6227 5219
rect 6227 5185 6236 5219
rect 6184 5176 6236 5185
rect 7656 5219 7708 5228
rect 7656 5185 7665 5219
rect 7665 5185 7699 5219
rect 7699 5185 7708 5219
rect 7656 5176 7708 5185
rect 6092 5108 6144 5160
rect 9496 5176 9548 5228
rect 8576 5108 8628 5160
rect 8760 5108 8812 5160
rect 16580 5040 16632 5092
rect 5448 5015 5500 5024
rect 5448 4981 5457 5015
rect 5457 4981 5491 5015
rect 5491 4981 5500 5015
rect 5448 4972 5500 4981
rect 7196 4972 7248 5024
rect 8024 4972 8076 5024
rect 9588 4972 9640 5024
rect 5666 4870 5718 4922
rect 5730 4870 5782 4922
rect 5794 4870 5846 4922
rect 5858 4870 5910 4922
rect 5922 4870 5974 4922
rect 8766 4870 8818 4922
rect 8830 4870 8882 4922
rect 8894 4870 8946 4922
rect 8958 4870 9010 4922
rect 9022 4870 9074 4922
rect 3792 4811 3844 4820
rect 3792 4777 3801 4811
rect 3801 4777 3835 4811
rect 3835 4777 3844 4811
rect 3792 4768 3844 4777
rect 6092 4768 6144 4820
rect 6920 4768 6972 4820
rect 8484 4768 8536 4820
rect 9220 4768 9272 4820
rect 7656 4700 7708 4752
rect 8300 4743 8352 4752
rect 8300 4709 8309 4743
rect 8309 4709 8343 4743
rect 8343 4709 8352 4743
rect 8300 4700 8352 4709
rect 1492 4564 1544 4616
rect 3700 4607 3752 4616
rect 3700 4573 3709 4607
rect 3709 4573 3743 4607
rect 3743 4573 3752 4607
rect 3700 4564 3752 4573
rect 3976 4496 4028 4548
rect 5448 4564 5500 4616
rect 5724 4607 5776 4616
rect 5724 4573 5733 4607
rect 5733 4573 5767 4607
rect 5767 4573 5776 4607
rect 5724 4564 5776 4573
rect 6828 4607 6880 4616
rect 6460 4496 6512 4548
rect 6828 4573 6837 4607
rect 6837 4573 6871 4607
rect 6871 4573 6880 4607
rect 6828 4564 6880 4573
rect 7932 4632 7984 4684
rect 8208 4632 8260 4684
rect 8392 4632 8444 4684
rect 7564 4607 7616 4616
rect 7564 4573 7573 4607
rect 7573 4573 7607 4607
rect 7607 4573 7616 4607
rect 7564 4564 7616 4573
rect 7196 4496 7248 4548
rect 7656 4496 7708 4548
rect 7840 4607 7892 4616
rect 7840 4573 7849 4607
rect 7849 4573 7883 4607
rect 7883 4573 7892 4607
rect 7840 4564 7892 4573
rect 8392 4539 8444 4548
rect 8392 4505 8401 4539
rect 8401 4505 8435 4539
rect 8435 4505 8444 4539
rect 8392 4496 8444 4505
rect 3332 4428 3384 4480
rect 4620 4428 4672 4480
rect 4988 4428 5040 4480
rect 6092 4471 6144 4480
rect 6092 4437 6101 4471
rect 6101 4437 6135 4471
rect 6135 4437 6144 4471
rect 6092 4428 6144 4437
rect 6184 4471 6236 4480
rect 6184 4437 6193 4471
rect 6193 4437 6227 4471
rect 6227 4437 6236 4471
rect 6184 4428 6236 4437
rect 8024 4428 8076 4480
rect 8944 4471 8996 4480
rect 8944 4437 8953 4471
rect 8953 4437 8987 4471
rect 8987 4437 8996 4471
rect 8944 4428 8996 4437
rect 9312 4428 9364 4480
rect 4116 4326 4168 4378
rect 4180 4326 4232 4378
rect 4244 4326 4296 4378
rect 4308 4326 4360 4378
rect 4372 4326 4424 4378
rect 7216 4326 7268 4378
rect 7280 4326 7332 4378
rect 7344 4326 7396 4378
rect 7408 4326 7460 4378
rect 7472 4326 7524 4378
rect 3976 4224 4028 4276
rect 5540 4224 5592 4276
rect 4528 4156 4580 4208
rect 3332 4131 3384 4140
rect 3332 4097 3341 4131
rect 3341 4097 3375 4131
rect 3375 4097 3384 4131
rect 3332 4088 3384 4097
rect 3884 4088 3936 4140
rect 4896 4088 4948 4140
rect 8300 4224 8352 4276
rect 8576 4224 8628 4276
rect 8944 4224 8996 4276
rect 6460 4156 6512 4208
rect 6644 4156 6696 4208
rect 8484 4156 8536 4208
rect 6368 4088 6420 4140
rect 8576 4131 8628 4140
rect 7932 3995 7984 4004
rect 7932 3961 7941 3995
rect 7941 3961 7975 3995
rect 7975 3961 7984 3995
rect 7932 3952 7984 3961
rect 8576 4097 8585 4131
rect 8585 4097 8619 4131
rect 8619 4097 8628 4131
rect 8576 4088 8628 4097
rect 9312 4088 9364 4140
rect 9220 4063 9272 4072
rect 9220 4029 9229 4063
rect 9229 4029 9263 4063
rect 9263 4029 9272 4063
rect 9220 4020 9272 4029
rect 9404 3952 9456 4004
rect 6368 3884 6420 3936
rect 6552 3884 6604 3936
rect 6644 3927 6696 3936
rect 6644 3893 6653 3927
rect 6653 3893 6687 3927
rect 6687 3893 6696 3927
rect 6644 3884 6696 3893
rect 7656 3884 7708 3936
rect 7840 3884 7892 3936
rect 16580 3884 16632 3936
rect 5666 3782 5718 3834
rect 5730 3782 5782 3834
rect 5794 3782 5846 3834
rect 5858 3782 5910 3834
rect 5922 3782 5974 3834
rect 8766 3782 8818 3834
rect 8830 3782 8882 3834
rect 8894 3782 8946 3834
rect 8958 3782 9010 3834
rect 9022 3782 9074 3834
rect 4528 3723 4580 3732
rect 4528 3689 4537 3723
rect 4537 3689 4571 3723
rect 4571 3689 4580 3723
rect 4528 3680 4580 3689
rect 4896 3723 4948 3732
rect 4896 3689 4905 3723
rect 4905 3689 4939 3723
rect 4939 3689 4948 3723
rect 4896 3680 4948 3689
rect 8576 3680 8628 3732
rect 9404 3680 9456 3732
rect 4620 3476 4672 3528
rect 6092 3544 6144 3596
rect 6552 3587 6604 3596
rect 6552 3553 6561 3587
rect 6561 3553 6595 3587
rect 6595 3553 6604 3587
rect 6552 3544 6604 3553
rect 4988 3519 5040 3528
rect 4988 3485 4997 3519
rect 4997 3485 5031 3519
rect 5031 3485 5040 3519
rect 4988 3476 5040 3485
rect 7012 3476 7064 3528
rect 7932 3476 7984 3528
rect 9496 3476 9548 3528
rect 2688 3408 2740 3460
rect 5172 3383 5224 3392
rect 5172 3349 5181 3383
rect 5181 3349 5215 3383
rect 5215 3349 5224 3383
rect 5172 3340 5224 3349
rect 7840 3408 7892 3460
rect 7748 3340 7800 3392
rect 8484 3340 8536 3392
rect 9128 3340 9180 3392
rect 4116 3238 4168 3290
rect 4180 3238 4232 3290
rect 4244 3238 4296 3290
rect 4308 3238 4360 3290
rect 4372 3238 4424 3290
rect 7216 3238 7268 3290
rect 7280 3238 7332 3290
rect 7344 3238 7396 3290
rect 7408 3238 7460 3290
rect 7472 3238 7524 3290
rect 7932 3136 7984 3188
rect 8392 3179 8444 3188
rect 5172 3068 5224 3120
rect 8392 3145 8401 3179
rect 8401 3145 8435 3179
rect 8435 3145 8444 3179
rect 8392 3136 8444 3145
rect 8668 3136 8720 3188
rect 3976 3000 4028 3052
rect 4712 3000 4764 3052
rect 6184 3000 6236 3052
rect 7656 3043 7708 3052
rect 7656 3009 7665 3043
rect 7665 3009 7699 3043
rect 7699 3009 7708 3043
rect 7656 3000 7708 3009
rect 8116 3000 8168 3052
rect 8300 3043 8352 3052
rect 8300 3009 8309 3043
rect 8309 3009 8343 3043
rect 8343 3009 8352 3043
rect 8300 3000 8352 3009
rect 9036 3068 9088 3120
rect 9680 3068 9732 3120
rect 6368 2932 6420 2984
rect 16580 2932 16632 2984
rect 8300 2864 8352 2916
rect 9404 2839 9456 2848
rect 9404 2805 9413 2839
rect 9413 2805 9447 2839
rect 9447 2805 9456 2839
rect 9404 2796 9456 2805
rect 5666 2694 5718 2746
rect 5730 2694 5782 2746
rect 5794 2694 5846 2746
rect 5858 2694 5910 2746
rect 5922 2694 5974 2746
rect 8766 2694 8818 2746
rect 8830 2694 8882 2746
rect 8894 2694 8946 2746
rect 8958 2694 9010 2746
rect 9022 2694 9074 2746
rect 7932 2592 7984 2644
rect 9220 2592 9272 2644
rect 9496 2592 9548 2644
rect 9312 2524 9364 2576
rect 8300 2456 8352 2508
rect 9128 2431 9180 2440
rect 9128 2397 9137 2431
rect 9137 2397 9171 2431
rect 9171 2397 9180 2431
rect 9128 2388 9180 2397
rect 16580 2320 16632 2372
rect 4116 2150 4168 2202
rect 4180 2150 4232 2202
rect 4244 2150 4296 2202
rect 4308 2150 4360 2202
rect 4372 2150 4424 2202
rect 7216 2150 7268 2202
rect 7280 2150 7332 2202
rect 7344 2150 7396 2202
rect 7408 2150 7460 2202
rect 7472 2150 7524 2202
rect 8208 2048 8260 2100
rect 7840 1844 7892 1896
rect 9220 1844 9272 1896
rect 16580 1776 16632 1828
rect 9128 1751 9180 1760
rect 9128 1717 9137 1751
rect 9137 1717 9171 1751
rect 9171 1717 9180 1751
rect 9128 1708 9180 1717
rect 5666 1606 5718 1658
rect 5730 1606 5782 1658
rect 5794 1606 5846 1658
rect 5858 1606 5910 1658
rect 5922 1606 5974 1658
rect 8766 1606 8818 1658
rect 8830 1606 8882 1658
rect 8894 1606 8946 1658
rect 8958 1606 9010 1658
rect 9022 1606 9074 1658
rect 4116 1062 4168 1114
rect 4180 1062 4232 1114
rect 4244 1062 4296 1114
rect 4308 1062 4360 1114
rect 4372 1062 4424 1114
rect 7216 1062 7268 1114
rect 7280 1062 7332 1114
rect 7344 1062 7396 1114
rect 7408 1062 7460 1114
rect 7472 1062 7524 1114
<< metal2 >>
rect 938 12200 994 13000
rect 1398 12200 1454 13000
rect 1858 12200 1914 13000
rect 2318 12200 2374 13000
rect 2410 12200 2466 12209
rect 2778 12200 2834 13000
rect 3238 12200 3294 13000
rect 3698 12200 3754 13000
rect 4158 12200 4214 13000
rect 4264 12294 4568 12322
rect 952 11762 980 12200
rect 1308 11960 1360 11966
rect 1308 11902 1360 11908
rect 940 11756 992 11762
rect 940 11698 992 11704
rect 952 11150 980 11698
rect 1124 11620 1176 11626
rect 1124 11562 1176 11568
rect 940 11144 992 11150
rect 940 11086 992 11092
rect 1032 9580 1084 9586
rect 1032 9522 1084 9528
rect 1044 7002 1072 9522
rect 1136 8906 1164 11562
rect 1320 10742 1348 11902
rect 1412 11234 1440 12200
rect 1768 12096 1820 12102
rect 1768 12038 1820 12044
rect 1674 11656 1730 11665
rect 1674 11591 1730 11600
rect 1688 11354 1716 11591
rect 1676 11348 1728 11354
rect 1676 11290 1728 11296
rect 1412 11206 1532 11234
rect 1504 11150 1532 11206
rect 1584 11212 1636 11218
rect 1584 11154 1636 11160
rect 1492 11144 1544 11150
rect 1492 11086 1544 11092
rect 1398 10976 1454 10985
rect 1398 10911 1454 10920
rect 1308 10736 1360 10742
rect 1308 10678 1360 10684
rect 1216 10668 1268 10674
rect 1216 10610 1268 10616
rect 1228 10169 1256 10610
rect 1320 10266 1348 10678
rect 1412 10674 1440 10911
rect 1400 10668 1452 10674
rect 1400 10610 1452 10616
rect 1308 10260 1360 10266
rect 1308 10202 1360 10208
rect 1214 10160 1270 10169
rect 1412 10146 1440 10610
rect 1214 10095 1270 10104
rect 1320 10118 1440 10146
rect 1228 9178 1256 10095
rect 1320 9654 1348 10118
rect 1400 10056 1452 10062
rect 1398 10024 1400 10033
rect 1452 10024 1454 10033
rect 1398 9959 1454 9968
rect 1398 9888 1454 9897
rect 1398 9823 1454 9832
rect 1308 9648 1360 9654
rect 1308 9590 1360 9596
rect 1306 9480 1362 9489
rect 1306 9415 1362 9424
rect 1216 9172 1268 9178
rect 1216 9114 1268 9120
rect 1214 9072 1270 9081
rect 1214 9007 1270 9016
rect 1124 8900 1176 8906
rect 1124 8842 1176 8848
rect 1032 6996 1084 7002
rect 1032 6938 1084 6944
rect 1136 6390 1164 8842
rect 1228 8634 1256 9007
rect 1320 8634 1348 9415
rect 1216 8628 1268 8634
rect 1216 8570 1268 8576
rect 1308 8628 1360 8634
rect 1308 8570 1360 8576
rect 1308 8288 1360 8294
rect 1308 8230 1360 8236
rect 1320 7546 1348 8230
rect 1308 7540 1360 7546
rect 1308 7482 1360 7488
rect 1412 6882 1440 9823
rect 1504 7818 1532 11086
rect 1596 10810 1624 11154
rect 1780 11150 1808 12038
rect 1768 11144 1820 11150
rect 1688 11104 1768 11132
rect 1584 10804 1636 10810
rect 1584 10746 1636 10752
rect 1688 9674 1716 11104
rect 1768 11086 1820 11092
rect 1596 9646 1716 9674
rect 1596 9081 1624 9646
rect 1766 9616 1822 9625
rect 1872 9586 1900 12200
rect 1952 12164 2004 12170
rect 1952 12106 2004 12112
rect 1964 10470 1992 12106
rect 2136 11824 2188 11830
rect 2136 11766 2188 11772
rect 2044 11552 2096 11558
rect 2044 11494 2096 11500
rect 2056 11354 2084 11494
rect 2044 11348 2096 11354
rect 2044 11290 2096 11296
rect 2148 11150 2176 11766
rect 2332 11642 2360 12200
rect 2410 12135 2466 12144
rect 2240 11614 2360 11642
rect 2136 11144 2188 11150
rect 2042 11112 2098 11121
rect 2136 11086 2188 11092
rect 2042 11047 2098 11056
rect 1952 10464 2004 10470
rect 1952 10406 2004 10412
rect 1950 10024 2006 10033
rect 1950 9959 2006 9968
rect 1766 9551 1822 9560
rect 1860 9580 1912 9586
rect 1676 9444 1728 9450
rect 1676 9386 1728 9392
rect 1582 9072 1638 9081
rect 1582 9007 1638 9016
rect 1584 8900 1636 8906
rect 1584 8842 1636 8848
rect 1596 8022 1624 8842
rect 1584 8016 1636 8022
rect 1584 7958 1636 7964
rect 1688 7834 1716 9386
rect 1492 7812 1544 7818
rect 1492 7754 1544 7760
rect 1596 7806 1716 7834
rect 1412 6854 1532 6882
rect 1400 6792 1452 6798
rect 1400 6734 1452 6740
rect 1124 6384 1176 6390
rect 1124 6326 1176 6332
rect 1412 5846 1440 6734
rect 1400 5840 1452 5846
rect 1400 5782 1452 5788
rect 1504 4622 1532 6854
rect 1596 6254 1624 7806
rect 1676 7744 1728 7750
rect 1676 7686 1728 7692
rect 1688 7585 1716 7686
rect 1674 7576 1730 7585
rect 1674 7511 1730 7520
rect 1688 6730 1716 7511
rect 1780 7410 1808 9551
rect 1860 9522 1912 9528
rect 1872 8294 1900 9522
rect 1964 8974 1992 9959
rect 2056 9586 2084 11047
rect 2134 10704 2190 10713
rect 2134 10639 2136 10648
rect 2188 10639 2190 10648
rect 2136 10610 2188 10616
rect 2134 10568 2190 10577
rect 2134 10503 2136 10512
rect 2188 10503 2190 10512
rect 2136 10474 2188 10480
rect 2240 10010 2268 11614
rect 2320 11552 2372 11558
rect 2320 11494 2372 11500
rect 2332 11354 2360 11494
rect 2320 11348 2372 11354
rect 2320 11290 2372 11296
rect 2424 11121 2452 12135
rect 2792 11626 2820 12200
rect 3056 11824 3108 11830
rect 2870 11792 2926 11801
rect 3056 11766 3108 11772
rect 3252 11778 3280 12200
rect 2870 11727 2926 11736
rect 2780 11620 2832 11626
rect 2780 11562 2832 11568
rect 2884 11540 2912 11727
rect 2884 11512 3004 11540
rect 2566 11452 2874 11472
rect 2566 11450 2572 11452
rect 2628 11450 2652 11452
rect 2708 11450 2732 11452
rect 2788 11450 2812 11452
rect 2868 11450 2874 11452
rect 2628 11398 2630 11450
rect 2810 11398 2812 11450
rect 2566 11396 2572 11398
rect 2628 11396 2652 11398
rect 2708 11396 2732 11398
rect 2788 11396 2812 11398
rect 2868 11396 2874 11398
rect 2566 11376 2874 11396
rect 2976 11336 3004 11512
rect 2792 11308 3004 11336
rect 2594 11248 2650 11257
rect 2594 11183 2650 11192
rect 2608 11150 2636 11183
rect 2792 11150 2820 11308
rect 2596 11144 2648 11150
rect 2410 11112 2466 11121
rect 2320 11076 2372 11082
rect 2596 11086 2648 11092
rect 2780 11144 2832 11150
rect 2780 11086 2832 11092
rect 2410 11047 2466 11056
rect 2320 11018 2372 11024
rect 2332 10674 2360 11018
rect 3068 11014 3096 11766
rect 3252 11750 3372 11778
rect 3148 11688 3200 11694
rect 3148 11630 3200 11636
rect 3160 11354 3188 11630
rect 3240 11620 3292 11626
rect 3240 11562 3292 11568
rect 3148 11348 3200 11354
rect 3148 11290 3200 11296
rect 3252 11126 3280 11562
rect 3240 11120 3292 11126
rect 3240 11062 3292 11068
rect 2780 11008 2832 11014
rect 3056 11008 3108 11014
rect 2832 10968 3004 10996
rect 2780 10950 2832 10956
rect 2778 10840 2834 10849
rect 2700 10784 2778 10792
rect 2700 10775 2834 10784
rect 2700 10764 2820 10775
rect 2320 10668 2372 10674
rect 2320 10610 2372 10616
rect 2700 10554 2728 10764
rect 2976 10690 3004 10968
rect 3056 10950 3108 10956
rect 2976 10674 3280 10690
rect 2964 10668 3292 10674
rect 3016 10662 3240 10668
rect 2964 10610 3016 10616
rect 3240 10610 3292 10616
rect 2332 10526 2728 10554
rect 3148 10600 3200 10606
rect 3148 10542 3200 10548
rect 2332 10470 2360 10526
rect 2320 10464 2372 10470
rect 2320 10406 2372 10412
rect 2412 10464 2464 10470
rect 2412 10406 2464 10412
rect 3054 10432 3110 10441
rect 2424 10112 2452 10406
rect 2566 10364 2874 10384
rect 3054 10367 3110 10376
rect 2566 10362 2572 10364
rect 2628 10362 2652 10364
rect 2708 10362 2732 10364
rect 2788 10362 2812 10364
rect 2868 10362 2874 10364
rect 2628 10310 2630 10362
rect 2810 10310 2812 10362
rect 2566 10308 2572 10310
rect 2628 10308 2652 10310
rect 2708 10308 2732 10310
rect 2788 10308 2812 10310
rect 2868 10308 2874 10310
rect 2566 10288 2874 10308
rect 2962 10296 3018 10305
rect 2962 10231 3018 10240
rect 2148 9982 2268 10010
rect 2332 10084 2452 10112
rect 2504 10124 2556 10130
rect 2148 9586 2176 9982
rect 2228 9920 2280 9926
rect 2332 9897 2360 10084
rect 2504 10066 2556 10072
rect 2516 10010 2544 10066
rect 2424 9982 2544 10010
rect 2228 9862 2280 9868
rect 2318 9888 2374 9897
rect 2044 9580 2096 9586
rect 2044 9522 2096 9528
rect 2136 9580 2188 9586
rect 2136 9522 2188 9528
rect 2056 9489 2084 9522
rect 2042 9480 2098 9489
rect 2042 9415 2098 9424
rect 2044 9376 2096 9382
rect 2044 9318 2096 9324
rect 1952 8968 2004 8974
rect 2056 8945 2084 9318
rect 2134 9072 2190 9081
rect 2134 9007 2190 9016
rect 2148 8974 2176 9007
rect 2136 8968 2188 8974
rect 1952 8910 2004 8916
rect 2042 8936 2098 8945
rect 2136 8910 2188 8916
rect 2042 8871 2098 8880
rect 2044 8492 2096 8498
rect 2044 8434 2096 8440
rect 1950 8392 2006 8401
rect 1950 8327 1952 8336
rect 2004 8327 2006 8336
rect 1952 8298 2004 8304
rect 1860 8288 1912 8294
rect 1860 8230 1912 8236
rect 1860 7744 1912 7750
rect 1860 7686 1912 7692
rect 1768 7404 1820 7410
rect 1768 7346 1820 7352
rect 1872 7342 1900 7686
rect 2056 7546 2084 8434
rect 2148 8430 2176 8910
rect 2240 8566 2268 9862
rect 2318 9823 2374 9832
rect 2318 9480 2374 9489
rect 2318 9415 2374 9424
rect 2332 9042 2360 9415
rect 2320 9036 2372 9042
rect 2320 8978 2372 8984
rect 2424 8974 2452 9982
rect 2504 9920 2556 9926
rect 2504 9862 2556 9868
rect 2516 9738 2544 9862
rect 2516 9710 2728 9738
rect 2976 9722 3004 10231
rect 2700 9654 2728 9710
rect 2964 9716 3016 9722
rect 2964 9658 3016 9664
rect 2688 9648 2740 9654
rect 2594 9616 2650 9625
rect 2688 9590 2740 9596
rect 2594 9551 2596 9560
rect 2648 9551 2650 9560
rect 2596 9522 2648 9528
rect 2962 9480 3018 9489
rect 2962 9415 3018 9424
rect 2566 9276 2874 9296
rect 2566 9274 2572 9276
rect 2628 9274 2652 9276
rect 2708 9274 2732 9276
rect 2788 9274 2812 9276
rect 2868 9274 2874 9276
rect 2628 9222 2630 9274
rect 2810 9222 2812 9274
rect 2566 9220 2572 9222
rect 2628 9220 2652 9222
rect 2708 9220 2732 9222
rect 2788 9220 2812 9222
rect 2868 9220 2874 9222
rect 2566 9200 2874 9220
rect 2412 8968 2464 8974
rect 2412 8910 2464 8916
rect 2412 8832 2464 8838
rect 2412 8774 2464 8780
rect 2228 8560 2280 8566
rect 2228 8502 2280 8508
rect 2136 8424 2188 8430
rect 2136 8366 2188 8372
rect 2320 8424 2372 8430
rect 2320 8366 2372 8372
rect 2228 8288 2280 8294
rect 2228 8230 2280 8236
rect 2044 7540 2096 7546
rect 2044 7482 2096 7488
rect 2240 7410 2268 8230
rect 2332 7970 2360 8366
rect 2424 8294 2452 8774
rect 2412 8288 2464 8294
rect 2412 8230 2464 8236
rect 2566 8188 2874 8208
rect 2566 8186 2572 8188
rect 2628 8186 2652 8188
rect 2708 8186 2732 8188
rect 2788 8186 2812 8188
rect 2868 8186 2874 8188
rect 2628 8134 2630 8186
rect 2810 8134 2812 8186
rect 2566 8132 2572 8134
rect 2628 8132 2652 8134
rect 2708 8132 2732 8134
rect 2788 8132 2812 8134
rect 2868 8132 2874 8134
rect 2566 8112 2874 8132
rect 2686 7984 2742 7993
rect 2332 7954 2452 7970
rect 2332 7948 2464 7954
rect 2332 7942 2412 7948
rect 2332 7546 2360 7942
rect 2686 7919 2742 7928
rect 2412 7890 2464 7896
rect 2700 7818 2728 7919
rect 2688 7812 2740 7818
rect 2688 7754 2740 7760
rect 2778 7576 2834 7585
rect 2320 7540 2372 7546
rect 2778 7511 2834 7520
rect 2320 7482 2372 7488
rect 2228 7404 2280 7410
rect 2228 7346 2280 7352
rect 1860 7336 1912 7342
rect 1860 7278 1912 7284
rect 2136 7200 2188 7206
rect 2136 7142 2188 7148
rect 1676 6724 1728 6730
rect 1676 6666 1728 6672
rect 1584 6248 1636 6254
rect 1584 6190 1636 6196
rect 2148 5642 2176 7142
rect 2332 7002 2360 7482
rect 2792 7410 2820 7511
rect 2780 7404 2832 7410
rect 2780 7346 2832 7352
rect 2976 7313 3004 9415
rect 3068 8974 3096 10367
rect 3160 10112 3188 10542
rect 3160 10084 3280 10112
rect 3148 9988 3200 9994
rect 3148 9930 3200 9936
rect 3160 9722 3188 9930
rect 3148 9716 3200 9722
rect 3148 9658 3200 9664
rect 3148 9172 3200 9178
rect 3148 9114 3200 9120
rect 3056 8968 3108 8974
rect 3056 8910 3108 8916
rect 3056 8832 3108 8838
rect 3056 8774 3108 8780
rect 3068 8129 3096 8774
rect 3054 8120 3110 8129
rect 3054 8055 3110 8064
rect 3054 7984 3110 7993
rect 3054 7919 3110 7928
rect 2410 7304 2466 7313
rect 2410 7239 2466 7248
rect 2962 7304 3018 7313
rect 2962 7239 3018 7248
rect 2320 6996 2372 7002
rect 2320 6938 2372 6944
rect 2332 6866 2360 6938
rect 2320 6860 2372 6866
rect 2320 6802 2372 6808
rect 2332 6322 2360 6802
rect 2424 6458 2452 7239
rect 2566 7100 2874 7120
rect 2566 7098 2572 7100
rect 2628 7098 2652 7100
rect 2708 7098 2732 7100
rect 2788 7098 2812 7100
rect 2868 7098 2874 7100
rect 2628 7046 2630 7098
rect 2810 7046 2812 7098
rect 2566 7044 2572 7046
rect 2628 7044 2652 7046
rect 2708 7044 2732 7046
rect 2788 7044 2812 7046
rect 2868 7044 2874 7046
rect 2566 7024 2874 7044
rect 2596 6860 2648 6866
rect 2596 6802 2648 6808
rect 2608 6662 2636 6802
rect 3068 6798 3096 7919
rect 3056 6792 3108 6798
rect 3056 6734 3108 6740
rect 2596 6656 2648 6662
rect 2596 6598 2648 6604
rect 2688 6656 2740 6662
rect 2688 6598 2740 6604
rect 2412 6452 2464 6458
rect 2412 6394 2464 6400
rect 2700 6390 2728 6598
rect 3068 6458 3096 6734
rect 3056 6452 3108 6458
rect 3056 6394 3108 6400
rect 2688 6384 2740 6390
rect 2688 6326 2740 6332
rect 2320 6316 2372 6322
rect 2320 6258 2372 6264
rect 2566 6012 2874 6032
rect 2566 6010 2572 6012
rect 2628 6010 2652 6012
rect 2708 6010 2732 6012
rect 2788 6010 2812 6012
rect 2868 6010 2874 6012
rect 2628 5958 2630 6010
rect 2810 5958 2812 6010
rect 2566 5956 2572 5958
rect 2628 5956 2652 5958
rect 2708 5956 2732 5958
rect 2788 5956 2812 5958
rect 2868 5956 2874 5958
rect 2566 5936 2874 5956
rect 3068 5642 3096 6394
rect 3160 5710 3188 9114
rect 3252 8974 3280 10084
rect 3344 9489 3372 11750
rect 3608 11552 3660 11558
rect 3608 11494 3660 11500
rect 3514 11384 3570 11393
rect 3514 11319 3570 11328
rect 3528 11218 3556 11319
rect 3620 11286 3648 11494
rect 3712 11370 3740 12200
rect 4172 12152 4200 12200
rect 4264 12152 4292 12294
rect 4172 12124 4292 12152
rect 3884 12028 3936 12034
rect 3884 11970 3936 11976
rect 3712 11342 3832 11370
rect 3608 11280 3660 11286
rect 3608 11222 3660 11228
rect 3700 11280 3752 11286
rect 3700 11222 3752 11228
rect 3516 11212 3568 11218
rect 3516 11154 3568 11160
rect 3514 10840 3570 10849
rect 3514 10775 3570 10784
rect 3424 10532 3476 10538
rect 3424 10474 3476 10480
rect 3436 9994 3464 10474
rect 3424 9988 3476 9994
rect 3424 9930 3476 9936
rect 3424 9648 3476 9654
rect 3424 9590 3476 9596
rect 3330 9480 3386 9489
rect 3330 9415 3386 9424
rect 3436 9178 3464 9590
rect 3424 9172 3476 9178
rect 3424 9114 3476 9120
rect 3240 8968 3292 8974
rect 3424 8968 3476 8974
rect 3240 8910 3292 8916
rect 3422 8936 3424 8945
rect 3476 8936 3478 8945
rect 3422 8871 3478 8880
rect 3528 8537 3556 10775
rect 3608 10464 3660 10470
rect 3608 10406 3660 10412
rect 3620 10198 3648 10406
rect 3608 10192 3660 10198
rect 3608 10134 3660 10140
rect 3712 10062 3740 11222
rect 3804 11014 3832 11342
rect 3792 11008 3844 11014
rect 3792 10950 3844 10956
rect 3896 10810 3924 11970
rect 4344 11756 4396 11762
rect 4344 11698 4396 11704
rect 4356 11286 4384 11698
rect 4436 11348 4488 11354
rect 4436 11290 4488 11296
rect 4344 11280 4396 11286
rect 4344 11222 4396 11228
rect 4448 11082 4476 11290
rect 4436 11076 4488 11082
rect 4436 11018 4488 11024
rect 3976 11008 4028 11014
rect 3976 10950 4028 10956
rect 3884 10804 3936 10810
rect 3884 10746 3936 10752
rect 3988 10742 4016 10950
rect 4116 10908 4424 10928
rect 4116 10906 4122 10908
rect 4178 10906 4202 10908
rect 4258 10906 4282 10908
rect 4338 10906 4362 10908
rect 4418 10906 4424 10908
rect 4178 10854 4180 10906
rect 4360 10854 4362 10906
rect 4116 10852 4122 10854
rect 4178 10852 4202 10854
rect 4258 10852 4282 10854
rect 4338 10852 4362 10854
rect 4418 10852 4424 10854
rect 4116 10832 4424 10852
rect 3976 10736 4028 10742
rect 4540 10713 4568 12294
rect 4618 12200 4674 13000
rect 5078 12200 5134 13000
rect 5538 12200 5594 13000
rect 5998 12200 6054 13000
rect 6184 12300 6236 12306
rect 6184 12242 6236 12248
rect 4632 11966 4660 12200
rect 4620 11960 4672 11966
rect 4620 11902 4672 11908
rect 4712 11960 4764 11966
rect 4712 11902 4764 11908
rect 4724 11150 4752 11902
rect 4712 11144 4764 11150
rect 4712 11086 4764 11092
rect 4988 11144 5040 11150
rect 5092 11121 5120 12200
rect 5552 11898 5580 12200
rect 6012 12102 6040 12200
rect 6000 12096 6052 12102
rect 6000 12038 6052 12044
rect 5540 11892 5592 11898
rect 5540 11834 5592 11840
rect 6000 11892 6052 11898
rect 6000 11834 6052 11840
rect 5170 11656 5226 11665
rect 5170 11591 5226 11600
rect 4988 11086 5040 11092
rect 5078 11112 5134 11121
rect 4804 11008 4856 11014
rect 4804 10950 4856 10956
rect 4896 11008 4948 11014
rect 4896 10950 4948 10956
rect 3976 10678 4028 10684
rect 4526 10704 4582 10713
rect 3884 10668 3936 10674
rect 4526 10639 4582 10648
rect 3884 10610 3936 10616
rect 3792 10464 3844 10470
rect 3792 10406 3844 10412
rect 3700 10056 3752 10062
rect 3700 9998 3752 10004
rect 3608 9988 3660 9994
rect 3608 9930 3660 9936
rect 3620 9194 3648 9930
rect 3620 9166 3740 9194
rect 3608 9104 3660 9110
rect 3608 9046 3660 9052
rect 3514 8528 3570 8537
rect 3514 8463 3570 8472
rect 3422 8120 3478 8129
rect 3422 8055 3424 8064
rect 3476 8055 3478 8064
rect 3424 8026 3476 8032
rect 3528 7886 3556 8463
rect 3516 7880 3568 7886
rect 3516 7822 3568 7828
rect 3332 6996 3384 7002
rect 3332 6938 3384 6944
rect 3344 5778 3372 6938
rect 3424 6792 3476 6798
rect 3424 6734 3476 6740
rect 3436 6662 3464 6734
rect 3424 6656 3476 6662
rect 3424 6598 3476 6604
rect 3332 5772 3384 5778
rect 3332 5714 3384 5720
rect 3148 5704 3200 5710
rect 3148 5646 3200 5652
rect 2136 5636 2188 5642
rect 2136 5578 2188 5584
rect 3056 5636 3108 5642
rect 3056 5578 3108 5584
rect 3344 5234 3372 5714
rect 3332 5228 3384 5234
rect 3332 5170 3384 5176
rect 1492 4616 1544 4622
rect 3620 4604 3648 9046
rect 3712 7002 3740 9166
rect 3804 8974 3832 10406
rect 3896 10305 3924 10610
rect 4160 10532 4212 10538
rect 4160 10474 4212 10480
rect 4172 10441 4200 10474
rect 4540 10470 4568 10639
rect 4528 10464 4580 10470
rect 4158 10432 4214 10441
rect 4528 10406 4580 10412
rect 4158 10367 4214 10376
rect 3882 10296 3938 10305
rect 3882 10231 3938 10240
rect 4528 10124 4580 10130
rect 4528 10066 4580 10072
rect 3976 10056 4028 10062
rect 3976 9998 4028 10004
rect 3884 9376 3936 9382
rect 3884 9318 3936 9324
rect 3792 8968 3844 8974
rect 3792 8910 3844 8916
rect 3790 8800 3846 8809
rect 3790 8735 3846 8744
rect 3804 8430 3832 8735
rect 3792 8424 3844 8430
rect 3792 8366 3844 8372
rect 3804 8129 3832 8366
rect 3790 8120 3846 8129
rect 3790 8055 3846 8064
rect 3792 8016 3844 8022
rect 3792 7958 3844 7964
rect 3804 7886 3832 7958
rect 3792 7880 3844 7886
rect 3792 7822 3844 7828
rect 3804 7290 3832 7822
rect 3896 7478 3924 9318
rect 3988 8430 4016 9998
rect 4116 9820 4424 9840
rect 4116 9818 4122 9820
rect 4178 9818 4202 9820
rect 4258 9818 4282 9820
rect 4338 9818 4362 9820
rect 4418 9818 4424 9820
rect 4178 9766 4180 9818
rect 4360 9766 4362 9818
rect 4116 9764 4122 9766
rect 4178 9764 4202 9766
rect 4258 9764 4282 9766
rect 4338 9764 4362 9766
rect 4418 9764 4424 9766
rect 4116 9744 4424 9764
rect 4344 9172 4396 9178
rect 4344 9114 4396 9120
rect 4356 8945 4384 9114
rect 4436 9104 4488 9110
rect 4436 9046 4488 9052
rect 4342 8936 4398 8945
rect 4448 8906 4476 9046
rect 4342 8871 4344 8880
rect 4396 8871 4398 8880
rect 4436 8900 4488 8906
rect 4344 8842 4396 8848
rect 4436 8842 4488 8848
rect 4116 8732 4424 8752
rect 4116 8730 4122 8732
rect 4178 8730 4202 8732
rect 4258 8730 4282 8732
rect 4338 8730 4362 8732
rect 4418 8730 4424 8732
rect 4178 8678 4180 8730
rect 4360 8678 4362 8730
rect 4116 8676 4122 8678
rect 4178 8676 4202 8678
rect 4258 8676 4282 8678
rect 4338 8676 4362 8678
rect 4418 8676 4424 8678
rect 4116 8656 4424 8676
rect 4540 8566 4568 10066
rect 4816 9994 4844 10950
rect 4908 10674 4936 10950
rect 5000 10810 5028 11086
rect 5078 11047 5134 11056
rect 4988 10804 5040 10810
rect 4988 10746 5040 10752
rect 4896 10668 4948 10674
rect 4896 10610 4948 10616
rect 5184 10588 5212 11591
rect 5666 11452 5974 11472
rect 5666 11450 5672 11452
rect 5728 11450 5752 11452
rect 5808 11450 5832 11452
rect 5888 11450 5912 11452
rect 5968 11450 5974 11452
rect 5728 11398 5730 11450
rect 5910 11398 5912 11450
rect 5666 11396 5672 11398
rect 5728 11396 5752 11398
rect 5808 11396 5832 11398
rect 5888 11396 5912 11398
rect 5968 11396 5974 11398
rect 5538 11384 5594 11393
rect 5666 11376 5974 11396
rect 6012 11354 6040 11834
rect 6092 11756 6144 11762
rect 6092 11698 6144 11704
rect 5538 11319 5594 11328
rect 6000 11348 6052 11354
rect 5446 11248 5502 11257
rect 5446 11183 5502 11192
rect 5264 11144 5316 11150
rect 5262 11112 5264 11121
rect 5316 11112 5318 11121
rect 5262 11047 5318 11056
rect 5356 10668 5408 10674
rect 5356 10610 5408 10616
rect 5264 10600 5316 10606
rect 5184 10560 5264 10588
rect 5264 10542 5316 10548
rect 5264 10464 5316 10470
rect 5264 10406 5316 10412
rect 4988 10056 5040 10062
rect 4988 9998 5040 10004
rect 4804 9988 4856 9994
rect 4804 9930 4856 9936
rect 4620 9580 4672 9586
rect 4620 9522 4672 9528
rect 4896 9580 4948 9586
rect 4896 9522 4948 9528
rect 4632 9178 4660 9522
rect 4712 9512 4764 9518
rect 4712 9454 4764 9460
rect 4620 9172 4672 9178
rect 4620 9114 4672 9120
rect 4724 9110 4752 9454
rect 4712 9104 4764 9110
rect 4712 9046 4764 9052
rect 4908 9042 4936 9522
rect 4896 9036 4948 9042
rect 4896 8978 4948 8984
rect 5000 8838 5028 9998
rect 5276 9722 5304 10406
rect 5264 9716 5316 9722
rect 5264 9658 5316 9664
rect 5368 9466 5396 10610
rect 5460 9602 5488 11183
rect 5552 10674 5580 11319
rect 6000 11290 6052 11296
rect 6104 11234 6132 11698
rect 5920 11206 6132 11234
rect 5920 11150 5948 11206
rect 5908 11144 5960 11150
rect 6092 11144 6144 11150
rect 5908 11086 5960 11092
rect 5998 11112 6054 11121
rect 5632 11076 5684 11082
rect 6092 11086 6144 11092
rect 5998 11047 6054 11056
rect 5632 11018 5684 11024
rect 5644 10810 5672 11018
rect 5908 11008 5960 11014
rect 5908 10950 5960 10956
rect 5632 10804 5684 10810
rect 5632 10746 5684 10752
rect 5920 10674 5948 10950
rect 5540 10668 5592 10674
rect 5540 10610 5592 10616
rect 5908 10668 5960 10674
rect 5908 10610 5960 10616
rect 5540 10464 5592 10470
rect 5540 10406 5592 10412
rect 5552 10198 5580 10406
rect 5666 10364 5974 10384
rect 5666 10362 5672 10364
rect 5728 10362 5752 10364
rect 5808 10362 5832 10364
rect 5888 10362 5912 10364
rect 5968 10362 5974 10364
rect 5728 10310 5730 10362
rect 5910 10310 5912 10362
rect 5666 10308 5672 10310
rect 5728 10308 5752 10310
rect 5808 10308 5832 10310
rect 5888 10308 5912 10310
rect 5968 10308 5974 10310
rect 5666 10288 5974 10308
rect 5540 10192 5592 10198
rect 5540 10134 5592 10140
rect 6012 9625 6040 11047
rect 6104 10606 6132 11086
rect 6092 10600 6144 10606
rect 6092 10542 6144 10548
rect 5998 9616 6054 9625
rect 5460 9574 5764 9602
rect 5736 9518 5764 9574
rect 5998 9551 6000 9560
rect 6052 9551 6054 9560
rect 6000 9522 6052 9528
rect 5724 9512 5776 9518
rect 5368 9450 5580 9466
rect 5724 9454 5776 9460
rect 5264 9444 5316 9450
rect 5368 9444 5592 9450
rect 5368 9438 5540 9444
rect 5264 9386 5316 9392
rect 5540 9386 5592 9392
rect 4988 8832 5040 8838
rect 4988 8774 5040 8780
rect 5080 8832 5132 8838
rect 5080 8774 5132 8780
rect 4528 8560 4580 8566
rect 4528 8502 4580 8508
rect 4160 8492 4212 8498
rect 4160 8434 4212 8440
rect 3976 8424 4028 8430
rect 3976 8366 4028 8372
rect 3988 7818 4016 8366
rect 4066 8120 4122 8129
rect 4066 8055 4068 8064
rect 4120 8055 4122 8064
rect 4068 8026 4120 8032
rect 4172 7954 4200 8434
rect 4528 8424 4580 8430
rect 4804 8424 4856 8430
rect 4580 8384 4660 8412
rect 4528 8366 4580 8372
rect 4160 7948 4212 7954
rect 4160 7890 4212 7896
rect 3976 7812 4028 7818
rect 3976 7754 4028 7760
rect 4116 7644 4424 7664
rect 4116 7642 4122 7644
rect 4178 7642 4202 7644
rect 4258 7642 4282 7644
rect 4338 7642 4362 7644
rect 4418 7642 4424 7644
rect 4178 7590 4180 7642
rect 4360 7590 4362 7642
rect 4116 7588 4122 7590
rect 4178 7588 4202 7590
rect 4258 7588 4282 7590
rect 4338 7588 4362 7590
rect 4418 7588 4424 7590
rect 4116 7568 4424 7588
rect 3884 7472 3936 7478
rect 3884 7414 3936 7420
rect 3804 7274 3924 7290
rect 3804 7268 3936 7274
rect 3804 7262 3884 7268
rect 3884 7210 3936 7216
rect 3700 6996 3752 7002
rect 3700 6938 3752 6944
rect 3700 6860 3752 6866
rect 3700 6802 3752 6808
rect 3712 5914 3740 6802
rect 4116 6556 4424 6576
rect 4116 6554 4122 6556
rect 4178 6554 4202 6556
rect 4258 6554 4282 6556
rect 4338 6554 4362 6556
rect 4418 6554 4424 6556
rect 4178 6502 4180 6554
rect 4360 6502 4362 6554
rect 4116 6500 4122 6502
rect 4178 6500 4202 6502
rect 4258 6500 4282 6502
rect 4338 6500 4362 6502
rect 4418 6500 4424 6502
rect 4116 6480 4424 6500
rect 3976 6112 4028 6118
rect 3976 6054 4028 6060
rect 3700 5908 3752 5914
rect 3700 5850 3752 5856
rect 3792 5908 3844 5914
rect 3792 5850 3844 5856
rect 3804 5642 3832 5850
rect 3792 5636 3844 5642
rect 3792 5578 3844 5584
rect 3804 5370 3832 5578
rect 3792 5364 3844 5370
rect 3792 5306 3844 5312
rect 3804 4826 3832 5306
rect 3988 5166 4016 6054
rect 4116 5468 4424 5488
rect 4116 5466 4122 5468
rect 4178 5466 4202 5468
rect 4258 5466 4282 5468
rect 4338 5466 4362 5468
rect 4418 5466 4424 5468
rect 4178 5414 4180 5466
rect 4360 5414 4362 5466
rect 4116 5412 4122 5414
rect 4178 5412 4202 5414
rect 4258 5412 4282 5414
rect 4338 5412 4362 5414
rect 4418 5412 4424 5414
rect 4116 5392 4424 5412
rect 4632 5370 4660 8384
rect 4804 8366 4856 8372
rect 4816 7546 4844 8366
rect 4804 7540 4856 7546
rect 4804 7482 4856 7488
rect 4712 6724 4764 6730
rect 4712 6666 4764 6672
rect 4724 5574 4752 6666
rect 4816 6458 4844 7482
rect 5092 7449 5120 8774
rect 5172 8084 5224 8090
rect 5172 8026 5224 8032
rect 5184 7818 5212 8026
rect 5172 7812 5224 7818
rect 5172 7754 5224 7760
rect 5078 7440 5134 7449
rect 5276 7410 5304 9386
rect 5666 9276 5974 9296
rect 5666 9274 5672 9276
rect 5728 9274 5752 9276
rect 5808 9274 5832 9276
rect 5888 9274 5912 9276
rect 5968 9274 5974 9276
rect 5728 9222 5730 9274
rect 5910 9222 5912 9274
rect 5666 9220 5672 9222
rect 5728 9220 5752 9222
rect 5808 9220 5832 9222
rect 5888 9220 5912 9222
rect 5968 9220 5974 9222
rect 5666 9200 5974 9220
rect 5538 8936 5594 8945
rect 5538 8871 5594 8880
rect 5908 8900 5960 8906
rect 5552 8498 5580 8871
rect 5908 8842 5960 8848
rect 5724 8560 5776 8566
rect 5722 8528 5724 8537
rect 5776 8528 5778 8537
rect 5540 8492 5592 8498
rect 5722 8463 5778 8472
rect 5540 8434 5592 8440
rect 5920 8362 5948 8842
rect 5540 8356 5592 8362
rect 5540 8298 5592 8304
rect 5908 8356 5960 8362
rect 5908 8298 5960 8304
rect 5552 7954 5580 8298
rect 5666 8188 5974 8208
rect 5666 8186 5672 8188
rect 5728 8186 5752 8188
rect 5808 8186 5832 8188
rect 5888 8186 5912 8188
rect 5968 8186 5974 8188
rect 5728 8134 5730 8186
rect 5910 8134 5912 8186
rect 5666 8132 5672 8134
rect 5728 8132 5752 8134
rect 5808 8132 5832 8134
rect 5888 8132 5912 8134
rect 5968 8132 5974 8134
rect 5666 8112 5974 8132
rect 6012 7954 6040 9522
rect 5540 7948 5592 7954
rect 5540 7890 5592 7896
rect 6000 7948 6052 7954
rect 6000 7890 6052 7896
rect 6196 7834 6224 12242
rect 6458 12200 6514 13000
rect 6552 12232 6604 12238
rect 6472 12034 6500 12200
rect 6552 12174 6604 12180
rect 6460 12028 6512 12034
rect 6460 11970 6512 11976
rect 6276 11620 6328 11626
rect 6276 11562 6328 11568
rect 6288 11354 6316 11562
rect 6276 11348 6328 11354
rect 6276 11290 6328 11296
rect 6460 10192 6512 10198
rect 6460 10134 6512 10140
rect 6368 9376 6420 9382
rect 6368 9318 6420 9324
rect 6380 7993 6408 9318
rect 6366 7984 6422 7993
rect 6366 7919 6422 7928
rect 6012 7806 6224 7834
rect 6276 7812 6328 7818
rect 5078 7375 5134 7384
rect 5264 7404 5316 7410
rect 5264 7346 5316 7352
rect 5666 7100 5974 7120
rect 5666 7098 5672 7100
rect 5728 7098 5752 7100
rect 5808 7098 5832 7100
rect 5888 7098 5912 7100
rect 5968 7098 5974 7100
rect 5728 7046 5730 7098
rect 5910 7046 5912 7098
rect 5666 7044 5672 7046
rect 5728 7044 5752 7046
rect 5808 7044 5832 7046
rect 5888 7044 5912 7046
rect 5968 7044 5974 7046
rect 5666 7024 5974 7044
rect 6012 6746 6040 7806
rect 6276 7754 6328 7760
rect 6184 7744 6236 7750
rect 6184 7686 6236 7692
rect 6196 7410 6224 7686
rect 6184 7404 6236 7410
rect 6184 7346 6236 7352
rect 6288 7274 6316 7754
rect 6368 7744 6420 7750
rect 6368 7686 6420 7692
rect 6380 7342 6408 7686
rect 6368 7336 6420 7342
rect 6368 7278 6420 7284
rect 6472 7290 6500 10134
rect 6564 8378 6592 12174
rect 8392 12164 8444 12170
rect 8392 12106 8444 12112
rect 7840 12028 7892 12034
rect 7840 11970 7892 11976
rect 7656 11756 7708 11762
rect 7656 11698 7708 11704
rect 7564 11688 7616 11694
rect 7564 11630 7616 11636
rect 7196 11620 7248 11626
rect 7196 11562 7248 11568
rect 6642 11384 6698 11393
rect 6642 11319 6644 11328
rect 6696 11319 6698 11328
rect 6644 11290 6696 11296
rect 6656 11014 6684 11290
rect 7104 11144 7156 11150
rect 7104 11086 7156 11092
rect 6644 11008 6696 11014
rect 6644 10950 6696 10956
rect 7012 11008 7064 11014
rect 7012 10950 7064 10956
rect 6656 8906 6684 10950
rect 6828 10600 6880 10606
rect 6828 10542 6880 10548
rect 6840 9926 6868 10542
rect 6920 10124 6972 10130
rect 6920 10066 6972 10072
rect 6828 9920 6880 9926
rect 6828 9862 6880 9868
rect 6840 9586 6868 9862
rect 6828 9580 6880 9586
rect 6828 9522 6880 9528
rect 6734 9072 6790 9081
rect 6734 9007 6790 9016
rect 6828 9036 6880 9042
rect 6644 8900 6696 8906
rect 6644 8842 6696 8848
rect 6656 8498 6684 8842
rect 6748 8566 6776 9007
rect 6828 8978 6880 8984
rect 6840 8566 6868 8978
rect 6736 8560 6788 8566
rect 6736 8502 6788 8508
rect 6828 8560 6880 8566
rect 6828 8502 6880 8508
rect 6644 8492 6696 8498
rect 6644 8434 6696 8440
rect 6564 8350 6684 8378
rect 6552 8288 6604 8294
rect 6552 8230 6604 8236
rect 6564 8022 6592 8230
rect 6552 8016 6604 8022
rect 6552 7958 6604 7964
rect 6092 7268 6144 7274
rect 6092 7210 6144 7216
rect 6276 7268 6328 7274
rect 6472 7262 6592 7290
rect 6276 7210 6328 7216
rect 6104 6798 6132 7210
rect 6184 7200 6236 7206
rect 6460 7200 6512 7206
rect 6236 7148 6460 7154
rect 6184 7142 6512 7148
rect 6196 7126 6500 7142
rect 6368 6996 6420 7002
rect 6564 6984 6592 7262
rect 6368 6938 6420 6944
rect 6472 6956 6592 6984
rect 6276 6928 6328 6934
rect 6276 6870 6328 6876
rect 5920 6718 6040 6746
rect 6092 6792 6144 6798
rect 6092 6734 6144 6740
rect 4804 6452 4856 6458
rect 4804 6394 4856 6400
rect 5920 6322 5948 6718
rect 6000 6656 6052 6662
rect 6000 6598 6052 6604
rect 5908 6316 5960 6322
rect 5908 6258 5960 6264
rect 5540 6248 5592 6254
rect 5540 6190 5592 6196
rect 4988 6112 5040 6118
rect 4988 6054 5040 6060
rect 5000 5642 5028 6054
rect 4988 5636 5040 5642
rect 4988 5578 5040 5584
rect 4712 5568 4764 5574
rect 4712 5510 4764 5516
rect 5552 5386 5580 6190
rect 5666 6012 5974 6032
rect 5666 6010 5672 6012
rect 5728 6010 5752 6012
rect 5808 6010 5832 6012
rect 5888 6010 5912 6012
rect 5968 6010 5974 6012
rect 5728 5958 5730 6010
rect 5910 5958 5912 6010
rect 5666 5956 5672 5958
rect 5728 5956 5752 5958
rect 5808 5956 5832 5958
rect 5888 5956 5912 5958
rect 5968 5956 5974 5958
rect 5666 5936 5974 5956
rect 5460 5370 5580 5386
rect 6012 5370 6040 6598
rect 4620 5364 4672 5370
rect 4620 5306 4672 5312
rect 5448 5364 5580 5370
rect 5500 5358 5580 5364
rect 6000 5364 6052 5370
rect 5448 5306 5500 5312
rect 6000 5306 6052 5312
rect 3976 5160 4028 5166
rect 3976 5102 4028 5108
rect 3792 4820 3844 4826
rect 3792 4762 3844 4768
rect 3988 4672 4016 5102
rect 3896 4644 4016 4672
rect 3700 4616 3752 4622
rect 3620 4584 3700 4604
rect 3752 4584 3754 4593
rect 3620 4576 3698 4584
rect 1492 4558 1544 4564
rect 3698 4519 3754 4528
rect 3332 4480 3384 4486
rect 3332 4422 3384 4428
rect 3344 4146 3372 4422
rect 3896 4146 3924 4644
rect 4632 4570 4660 5306
rect 6104 5250 6132 6734
rect 6184 5636 6236 5642
rect 6184 5578 6236 5584
rect 6012 5234 6132 5250
rect 6196 5234 6224 5578
rect 6000 5228 6132 5234
rect 6052 5222 6132 5228
rect 6184 5228 6236 5234
rect 6000 5170 6052 5176
rect 6184 5170 6236 5176
rect 5540 5160 5592 5166
rect 5540 5102 5592 5108
rect 6092 5160 6144 5166
rect 6092 5102 6144 5108
rect 5448 5024 5500 5030
rect 5448 4966 5500 4972
rect 5460 4622 5488 4966
rect 5448 4616 5500 4622
rect 3976 4548 4028 4554
rect 4632 4542 4752 4570
rect 5448 4558 5500 4564
rect 3976 4490 4028 4496
rect 3988 4282 4016 4490
rect 4620 4480 4672 4486
rect 4620 4422 4672 4428
rect 4116 4380 4424 4400
rect 4116 4378 4122 4380
rect 4178 4378 4202 4380
rect 4258 4378 4282 4380
rect 4338 4378 4362 4380
rect 4418 4378 4424 4380
rect 4178 4326 4180 4378
rect 4360 4326 4362 4378
rect 4116 4324 4122 4326
rect 4178 4324 4202 4326
rect 4258 4324 4282 4326
rect 4338 4324 4362 4326
rect 4418 4324 4424 4326
rect 4116 4304 4424 4324
rect 3976 4276 4028 4282
rect 3976 4218 4028 4224
rect 3332 4140 3384 4146
rect 3332 4082 3384 4088
rect 3884 4140 3936 4146
rect 3884 4082 3936 4088
rect 2688 3460 2740 3466
rect 2688 3402 2740 3408
rect 2700 3369 2728 3402
rect 2686 3360 2742 3369
rect 2686 3295 2742 3304
rect 3988 3058 4016 4218
rect 4528 4208 4580 4214
rect 4528 4150 4580 4156
rect 4540 3738 4568 4150
rect 4528 3732 4580 3738
rect 4528 3674 4580 3680
rect 4632 3534 4660 4422
rect 4620 3528 4672 3534
rect 4620 3470 4672 3476
rect 4116 3292 4424 3312
rect 4116 3290 4122 3292
rect 4178 3290 4202 3292
rect 4258 3290 4282 3292
rect 4338 3290 4362 3292
rect 4418 3290 4424 3292
rect 4178 3238 4180 3290
rect 4360 3238 4362 3290
rect 4116 3236 4122 3238
rect 4178 3236 4202 3238
rect 4258 3236 4282 3238
rect 4338 3236 4362 3238
rect 4418 3236 4424 3238
rect 4116 3216 4424 3236
rect 4724 3058 4752 4542
rect 4988 4480 5040 4486
rect 4988 4422 5040 4428
rect 4896 4140 4948 4146
rect 4896 4082 4948 4088
rect 4908 3738 4936 4082
rect 4896 3732 4948 3738
rect 4896 3674 4948 3680
rect 5000 3534 5028 4422
rect 5552 4282 5580 5102
rect 5666 4924 5974 4944
rect 5666 4922 5672 4924
rect 5728 4922 5752 4924
rect 5808 4922 5832 4924
rect 5888 4922 5912 4924
rect 5968 4922 5974 4924
rect 5728 4870 5730 4922
rect 5910 4870 5912 4922
rect 5666 4868 5672 4870
rect 5728 4868 5752 4870
rect 5808 4868 5832 4870
rect 5888 4868 5912 4870
rect 5968 4868 5974 4870
rect 5666 4848 5974 4868
rect 6104 4826 6132 5102
rect 6092 4820 6144 4826
rect 6092 4762 6144 4768
rect 5724 4616 5776 4622
rect 5722 4584 5724 4593
rect 5776 4584 5778 4593
rect 5722 4519 5778 4528
rect 6092 4480 6144 4486
rect 6092 4422 6144 4428
rect 6184 4480 6236 4486
rect 6184 4422 6236 4428
rect 5540 4276 5592 4282
rect 5540 4218 5592 4224
rect 5666 3836 5974 3856
rect 5666 3834 5672 3836
rect 5728 3834 5752 3836
rect 5808 3834 5832 3836
rect 5888 3834 5912 3836
rect 5968 3834 5974 3836
rect 5728 3782 5730 3834
rect 5910 3782 5912 3834
rect 5666 3780 5672 3782
rect 5728 3780 5752 3782
rect 5808 3780 5832 3782
rect 5888 3780 5912 3782
rect 5968 3780 5974 3782
rect 5666 3760 5974 3780
rect 6104 3602 6132 4422
rect 6092 3596 6144 3602
rect 6092 3538 6144 3544
rect 4988 3528 5040 3534
rect 4988 3470 5040 3476
rect 5172 3392 5224 3398
rect 5172 3334 5224 3340
rect 5184 3126 5212 3334
rect 5172 3120 5224 3126
rect 5172 3062 5224 3068
rect 6196 3058 6224 4422
rect 6288 4162 6316 6870
rect 6380 6118 6408 6938
rect 6472 6186 6500 6956
rect 6656 6934 6684 8350
rect 6644 6928 6696 6934
rect 6644 6870 6696 6876
rect 6552 6860 6604 6866
rect 6552 6802 6604 6808
rect 6460 6180 6512 6186
rect 6460 6122 6512 6128
rect 6368 6112 6420 6118
rect 6368 6054 6420 6060
rect 6564 5778 6592 6802
rect 6644 6656 6696 6662
rect 6644 6598 6696 6604
rect 6656 5778 6684 6598
rect 6748 6390 6776 8502
rect 6840 7478 6868 8502
rect 6932 8362 6960 10066
rect 7024 9586 7052 10950
rect 7116 10810 7144 11086
rect 7208 11082 7236 11562
rect 7196 11076 7248 11082
rect 7196 11018 7248 11024
rect 7216 10908 7524 10928
rect 7216 10906 7222 10908
rect 7278 10906 7302 10908
rect 7358 10906 7382 10908
rect 7438 10906 7462 10908
rect 7518 10906 7524 10908
rect 7278 10854 7280 10906
rect 7460 10854 7462 10906
rect 7216 10852 7222 10854
rect 7278 10852 7302 10854
rect 7358 10852 7382 10854
rect 7438 10852 7462 10854
rect 7518 10852 7524 10854
rect 7216 10832 7524 10852
rect 7104 10804 7156 10810
rect 7104 10746 7156 10752
rect 7576 10674 7604 11630
rect 7564 10668 7616 10674
rect 7564 10610 7616 10616
rect 7470 10568 7526 10577
rect 7470 10503 7526 10512
rect 7104 10124 7156 10130
rect 7104 10066 7156 10072
rect 7012 9580 7064 9586
rect 7012 9522 7064 9528
rect 7116 9042 7144 10066
rect 7484 9994 7512 10503
rect 7472 9988 7524 9994
rect 7472 9930 7524 9936
rect 7216 9820 7524 9840
rect 7216 9818 7222 9820
rect 7278 9818 7302 9820
rect 7358 9818 7382 9820
rect 7438 9818 7462 9820
rect 7518 9818 7524 9820
rect 7278 9766 7280 9818
rect 7460 9766 7462 9818
rect 7216 9764 7222 9766
rect 7278 9764 7302 9766
rect 7358 9764 7382 9766
rect 7438 9764 7462 9766
rect 7518 9764 7524 9766
rect 7216 9744 7524 9764
rect 7668 9586 7696 11698
rect 7748 11688 7800 11694
rect 7748 11630 7800 11636
rect 7760 11354 7788 11630
rect 7748 11348 7800 11354
rect 7748 11290 7800 11296
rect 7852 10538 7880 11970
rect 8022 11792 8078 11801
rect 8022 11727 8078 11736
rect 7840 10532 7892 10538
rect 7840 10474 7892 10480
rect 7932 10464 7984 10470
rect 7932 10406 7984 10412
rect 7944 10266 7972 10406
rect 7932 10260 7984 10266
rect 7932 10202 7984 10208
rect 7840 10192 7892 10198
rect 8036 10146 8064 11727
rect 8206 11384 8262 11393
rect 8206 11319 8208 11328
rect 8260 11319 8262 11328
rect 8404 11370 8432 12106
rect 16670 11928 16726 11937
rect 16670 11863 16726 11872
rect 9220 11824 9272 11830
rect 9220 11766 9272 11772
rect 9128 11688 9180 11694
rect 9128 11630 9180 11636
rect 8668 11552 8720 11558
rect 8668 11494 8720 11500
rect 8404 11342 8616 11370
rect 8208 11290 8260 11296
rect 8220 10674 8248 11290
rect 8404 11218 8432 11342
rect 8484 11280 8536 11286
rect 8484 11222 8536 11228
rect 8392 11212 8444 11218
rect 8392 11154 8444 11160
rect 8300 11144 8352 11150
rect 8300 11086 8352 11092
rect 8208 10668 8260 10674
rect 8208 10610 8260 10616
rect 8116 10600 8168 10606
rect 8116 10542 8168 10548
rect 7840 10134 7892 10140
rect 7656 9580 7708 9586
rect 7656 9522 7708 9528
rect 7564 9512 7616 9518
rect 7564 9454 7616 9460
rect 7196 9376 7248 9382
rect 7196 9318 7248 9324
rect 7208 9178 7236 9318
rect 7196 9172 7248 9178
rect 7196 9114 7248 9120
rect 7104 9036 7156 9042
rect 7104 8978 7156 8984
rect 7576 8906 7604 9454
rect 7196 8900 7248 8906
rect 7024 8860 7196 8888
rect 6920 8356 6972 8362
rect 6920 8298 6972 8304
rect 6920 7812 6972 7818
rect 6920 7754 6972 7760
rect 6828 7472 6880 7478
rect 6828 7414 6880 7420
rect 6840 6866 6868 7414
rect 6828 6860 6880 6866
rect 6828 6802 6880 6808
rect 6932 6798 6960 7754
rect 7024 7324 7052 8860
rect 7196 8842 7248 8848
rect 7564 8900 7616 8906
rect 7564 8842 7616 8848
rect 7216 8732 7524 8752
rect 7216 8730 7222 8732
rect 7278 8730 7302 8732
rect 7358 8730 7382 8732
rect 7438 8730 7462 8732
rect 7518 8730 7524 8732
rect 7278 8678 7280 8730
rect 7460 8678 7462 8730
rect 7216 8676 7222 8678
rect 7278 8676 7302 8678
rect 7358 8676 7382 8678
rect 7438 8676 7462 8678
rect 7518 8676 7524 8678
rect 7216 8656 7524 8676
rect 7564 8424 7616 8430
rect 7564 8366 7616 8372
rect 7216 7644 7524 7664
rect 7216 7642 7222 7644
rect 7278 7642 7302 7644
rect 7358 7642 7382 7644
rect 7438 7642 7462 7644
rect 7518 7642 7524 7644
rect 7278 7590 7280 7642
rect 7460 7590 7462 7642
rect 7216 7588 7222 7590
rect 7278 7588 7302 7590
rect 7358 7588 7382 7590
rect 7438 7588 7462 7590
rect 7518 7588 7524 7590
rect 7216 7568 7524 7588
rect 7576 7546 7604 8366
rect 7668 7750 7696 9522
rect 7748 8900 7800 8906
rect 7748 8842 7800 8848
rect 7760 7818 7788 8842
rect 7852 8634 7880 10134
rect 7944 10118 8064 10146
rect 7840 8628 7892 8634
rect 7840 8570 7892 8576
rect 7944 7834 7972 10118
rect 8024 9716 8076 9722
rect 8024 9658 8076 9664
rect 8036 8566 8064 9658
rect 8128 8974 8156 10542
rect 8220 10266 8248 10610
rect 8208 10260 8260 10266
rect 8208 10202 8260 10208
rect 8220 9926 8248 10202
rect 8208 9920 8260 9926
rect 8208 9862 8260 9868
rect 8206 9480 8262 9489
rect 8206 9415 8262 9424
rect 8116 8968 8168 8974
rect 8116 8910 8168 8916
rect 8024 8560 8076 8566
rect 8024 8502 8076 8508
rect 8220 8401 8248 9415
rect 8206 8392 8262 8401
rect 8206 8327 8262 8336
rect 8116 8016 8168 8022
rect 8168 7964 8248 7970
rect 8116 7958 8248 7964
rect 8128 7942 8248 7958
rect 8220 7886 8248 7942
rect 7748 7812 7800 7818
rect 7748 7754 7800 7760
rect 7852 7806 7972 7834
rect 8208 7880 8260 7886
rect 8208 7822 8260 7828
rect 8116 7812 8168 7818
rect 7656 7744 7708 7750
rect 7656 7686 7708 7692
rect 7104 7540 7156 7546
rect 7564 7540 7616 7546
rect 7156 7500 7236 7528
rect 7104 7482 7156 7488
rect 7208 7342 7236 7500
rect 7564 7482 7616 7488
rect 7288 7472 7340 7478
rect 7288 7414 7340 7420
rect 7104 7336 7156 7342
rect 7024 7296 7104 7324
rect 7104 7278 7156 7284
rect 7196 7336 7248 7342
rect 7196 7278 7248 7284
rect 7196 6996 7248 7002
rect 7300 6984 7328 7414
rect 7760 7002 7788 7754
rect 7248 6956 7328 6984
rect 7748 6996 7800 7002
rect 7196 6938 7248 6944
rect 7748 6938 7800 6944
rect 7208 6798 7236 6938
rect 6920 6792 6972 6798
rect 6920 6734 6972 6740
rect 7196 6792 7248 6798
rect 7196 6734 7248 6740
rect 6920 6656 6972 6662
rect 6972 6616 7052 6644
rect 6920 6598 6972 6604
rect 6736 6384 6788 6390
rect 6736 6326 6788 6332
rect 6828 6384 6880 6390
rect 6828 6326 6880 6332
rect 6840 6202 6868 6326
rect 6748 6174 6868 6202
rect 6552 5772 6604 5778
rect 6552 5714 6604 5720
rect 6644 5772 6696 5778
rect 6644 5714 6696 5720
rect 6748 5574 6776 6174
rect 6828 6112 6880 6118
rect 6828 6054 6880 6060
rect 6736 5568 6788 5574
rect 6736 5510 6788 5516
rect 6840 4622 6868 6054
rect 7024 5914 7052 6616
rect 7216 6556 7524 6576
rect 7216 6554 7222 6556
rect 7278 6554 7302 6556
rect 7358 6554 7382 6556
rect 7438 6554 7462 6556
rect 7518 6554 7524 6556
rect 7278 6502 7280 6554
rect 7460 6502 7462 6554
rect 7216 6500 7222 6502
rect 7278 6500 7302 6502
rect 7358 6500 7382 6502
rect 7438 6500 7462 6502
rect 7518 6500 7524 6502
rect 7216 6480 7524 6500
rect 7196 6248 7248 6254
rect 7196 6190 7248 6196
rect 7208 5914 7236 6190
rect 7012 5908 7064 5914
rect 7012 5850 7064 5856
rect 7196 5908 7248 5914
rect 7196 5850 7248 5856
rect 7564 5908 7616 5914
rect 7564 5850 7616 5856
rect 6920 5296 6972 5302
rect 6920 5238 6972 5244
rect 6932 4826 6960 5238
rect 6920 4820 6972 4826
rect 6920 4762 6972 4768
rect 6828 4616 6880 4622
rect 6828 4558 6880 4564
rect 6460 4548 6512 4554
rect 6460 4490 6512 4496
rect 6472 4214 6500 4490
rect 6460 4208 6512 4214
rect 6288 4146 6408 4162
rect 6460 4150 6512 4156
rect 6644 4208 6696 4214
rect 6644 4150 6696 4156
rect 6288 4140 6420 4146
rect 6288 4134 6368 4140
rect 6368 4082 6420 4088
rect 6656 3942 6684 4150
rect 6368 3936 6420 3942
rect 6368 3878 6420 3884
rect 6552 3936 6604 3942
rect 6552 3878 6604 3884
rect 6644 3936 6696 3942
rect 6644 3878 6696 3884
rect 3976 3052 4028 3058
rect 3976 2994 4028 3000
rect 4712 3052 4764 3058
rect 4712 2994 4764 3000
rect 6184 3052 6236 3058
rect 6184 2994 6236 3000
rect 6380 2990 6408 3878
rect 6564 3602 6592 3878
rect 6552 3596 6604 3602
rect 6552 3538 6604 3544
rect 7024 3534 7052 5850
rect 7216 5468 7524 5488
rect 7216 5466 7222 5468
rect 7278 5466 7302 5468
rect 7358 5466 7382 5468
rect 7438 5466 7462 5468
rect 7518 5466 7524 5468
rect 7278 5414 7280 5466
rect 7460 5414 7462 5466
rect 7216 5412 7222 5414
rect 7278 5412 7302 5414
rect 7358 5412 7382 5414
rect 7438 5412 7462 5414
rect 7518 5412 7524 5414
rect 7216 5392 7524 5412
rect 7196 5024 7248 5030
rect 7196 4966 7248 4972
rect 7208 4554 7236 4966
rect 7576 4622 7604 5850
rect 7656 5704 7708 5710
rect 7760 5692 7788 6938
rect 7708 5664 7788 5692
rect 7656 5646 7708 5652
rect 7656 5228 7708 5234
rect 7656 5170 7708 5176
rect 7668 4758 7696 5170
rect 7656 4752 7708 4758
rect 7852 4706 7880 7806
rect 8116 7754 8168 7760
rect 7932 7744 7984 7750
rect 7932 7686 7984 7692
rect 7656 4694 7708 4700
rect 7760 4678 7880 4706
rect 7944 4690 7972 7686
rect 8128 6662 8156 7754
rect 8208 7540 8260 7546
rect 8208 7482 8260 7488
rect 8220 7002 8248 7482
rect 8208 6996 8260 7002
rect 8208 6938 8260 6944
rect 8116 6656 8168 6662
rect 8116 6598 8168 6604
rect 8114 5808 8170 5817
rect 8114 5743 8170 5752
rect 8024 5568 8076 5574
rect 8024 5510 8076 5516
rect 8036 5030 8064 5510
rect 8024 5024 8076 5030
rect 8024 4966 8076 4972
rect 7932 4684 7984 4690
rect 7564 4616 7616 4622
rect 7760 4570 7788 4678
rect 7932 4626 7984 4632
rect 7564 4558 7616 4564
rect 7668 4554 7788 4570
rect 7840 4616 7892 4622
rect 7840 4558 7892 4564
rect 7930 4584 7986 4593
rect 7196 4548 7248 4554
rect 7196 4490 7248 4496
rect 7656 4548 7788 4554
rect 7708 4542 7788 4548
rect 7656 4490 7708 4496
rect 7216 4380 7524 4400
rect 7216 4378 7222 4380
rect 7278 4378 7302 4380
rect 7358 4378 7382 4380
rect 7438 4378 7462 4380
rect 7518 4378 7524 4380
rect 7278 4326 7280 4378
rect 7460 4326 7462 4378
rect 7216 4324 7222 4326
rect 7278 4324 7302 4326
rect 7358 4324 7382 4326
rect 7438 4324 7462 4326
rect 7518 4324 7524 4326
rect 7216 4304 7524 4324
rect 7852 4026 7880 4558
rect 7930 4519 7986 4528
rect 7760 3998 7880 4026
rect 7944 4010 7972 4519
rect 8024 4480 8076 4486
rect 8024 4422 8076 4428
rect 7932 4004 7984 4010
rect 7656 3936 7708 3942
rect 7656 3878 7708 3884
rect 7012 3528 7064 3534
rect 7012 3470 7064 3476
rect 7216 3292 7524 3312
rect 7216 3290 7222 3292
rect 7278 3290 7302 3292
rect 7358 3290 7382 3292
rect 7438 3290 7462 3292
rect 7518 3290 7524 3292
rect 7278 3238 7280 3290
rect 7460 3238 7462 3290
rect 7216 3236 7222 3238
rect 7278 3236 7302 3238
rect 7358 3236 7382 3238
rect 7438 3236 7462 3238
rect 7518 3236 7524 3238
rect 7216 3216 7524 3236
rect 7668 3058 7696 3878
rect 7760 3398 7788 3998
rect 7932 3946 7984 3952
rect 7840 3936 7892 3942
rect 7840 3878 7892 3884
rect 7852 3466 7880 3878
rect 7932 3528 7984 3534
rect 7932 3470 7984 3476
rect 7840 3460 7892 3466
rect 7840 3402 7892 3408
rect 7748 3392 7800 3398
rect 7748 3334 7800 3340
rect 7944 3194 7972 3470
rect 7932 3188 7984 3194
rect 7932 3130 7984 3136
rect 8036 3074 8064 4422
rect 7656 3052 7708 3058
rect 7656 2994 7708 3000
rect 7852 3046 8064 3074
rect 8128 3058 8156 5743
rect 8312 4758 8340 11086
rect 8392 11076 8444 11082
rect 8392 11018 8444 11024
rect 8404 9466 8432 11018
rect 8496 9654 8524 11222
rect 8588 10742 8616 11342
rect 8680 11150 8708 11494
rect 8766 11452 9074 11472
rect 8766 11450 8772 11452
rect 8828 11450 8852 11452
rect 8908 11450 8932 11452
rect 8988 11450 9012 11452
rect 9068 11450 9074 11452
rect 8828 11398 8830 11450
rect 9010 11398 9012 11450
rect 8766 11396 8772 11398
rect 8828 11396 8852 11398
rect 8908 11396 8932 11398
rect 8988 11396 9012 11398
rect 9068 11396 9074 11398
rect 8766 11376 9074 11396
rect 8668 11144 8720 11150
rect 8668 11086 8720 11092
rect 8576 10736 8628 10742
rect 8576 10678 8628 10684
rect 8668 10464 8720 10470
rect 8668 10406 8720 10412
rect 8576 9920 8628 9926
rect 8576 9862 8628 9868
rect 8484 9648 8536 9654
rect 8484 9590 8536 9596
rect 8404 9450 8524 9466
rect 8404 9444 8536 9450
rect 8404 9438 8484 9444
rect 8484 9386 8536 9392
rect 8588 8974 8616 9862
rect 8576 8968 8628 8974
rect 8576 8910 8628 8916
rect 8576 7880 8628 7886
rect 8576 7822 8628 7828
rect 8484 7812 8536 7818
rect 8484 7754 8536 7760
rect 8392 7744 8444 7750
rect 8392 7686 8444 7692
rect 8404 6633 8432 7686
rect 8390 6624 8446 6633
rect 8390 6559 8446 6568
rect 8496 6474 8524 7754
rect 8588 7002 8616 7822
rect 8680 7342 8708 10406
rect 8766 10364 9074 10384
rect 8766 10362 8772 10364
rect 8828 10362 8852 10364
rect 8908 10362 8932 10364
rect 8988 10362 9012 10364
rect 9068 10362 9074 10364
rect 8828 10310 8830 10362
rect 9010 10310 9012 10362
rect 8766 10308 8772 10310
rect 8828 10308 8852 10310
rect 8908 10308 8932 10310
rect 8988 10308 9012 10310
rect 9068 10308 9074 10310
rect 8766 10288 9074 10308
rect 8852 9920 8904 9926
rect 8852 9862 8904 9868
rect 8864 9654 8892 9862
rect 8852 9648 8904 9654
rect 8852 9590 8904 9596
rect 8766 9276 9074 9296
rect 8766 9274 8772 9276
rect 8828 9274 8852 9276
rect 8908 9274 8932 9276
rect 8988 9274 9012 9276
rect 9068 9274 9074 9276
rect 8828 9222 8830 9274
rect 9010 9222 9012 9274
rect 8766 9220 8772 9222
rect 8828 9220 8852 9222
rect 8908 9220 8932 9222
rect 8988 9220 9012 9222
rect 9068 9220 9074 9222
rect 8766 9200 9074 9220
rect 8760 9104 8812 9110
rect 8760 9046 8812 9052
rect 8772 8906 8800 9046
rect 8760 8900 8812 8906
rect 8760 8842 8812 8848
rect 9140 8498 9168 11630
rect 9232 11150 9260 11766
rect 9312 11620 9364 11626
rect 9312 11562 9364 11568
rect 9220 11144 9272 11150
rect 9220 11086 9272 11092
rect 9218 9616 9274 9625
rect 9218 9551 9274 9560
rect 9232 9217 9260 9551
rect 9218 9208 9274 9217
rect 9324 9178 9352 11562
rect 13726 11520 13782 11529
rect 13726 11455 13782 11464
rect 13740 11218 13768 11455
rect 13820 11280 13872 11286
rect 13820 11222 13872 11228
rect 13728 11212 13780 11218
rect 13728 11154 13780 11160
rect 13832 11121 13860 11222
rect 13818 11112 13874 11121
rect 13818 11047 13874 11056
rect 9404 11008 9456 11014
rect 9404 10950 9456 10956
rect 9416 10305 9444 10950
rect 16580 10464 16632 10470
rect 16580 10406 16632 10412
rect 9402 10296 9458 10305
rect 9402 10231 9458 10240
rect 9496 10056 9548 10062
rect 9496 9998 9548 10004
rect 9404 9648 9456 9654
rect 9404 9590 9456 9596
rect 9218 9143 9274 9152
rect 9312 9172 9364 9178
rect 9312 9114 9364 9120
rect 9416 9110 9444 9590
rect 9404 9104 9456 9110
rect 9404 9046 9456 9052
rect 9220 8968 9272 8974
rect 9220 8910 9272 8916
rect 9128 8492 9180 8498
rect 9128 8434 9180 8440
rect 9128 8288 9180 8294
rect 9128 8230 9180 8236
rect 8766 8188 9074 8208
rect 8766 8186 8772 8188
rect 8828 8186 8852 8188
rect 8908 8186 8932 8188
rect 8988 8186 9012 8188
rect 9068 8186 9074 8188
rect 8828 8134 8830 8186
rect 9010 8134 9012 8186
rect 8766 8132 8772 8134
rect 8828 8132 8852 8134
rect 8908 8132 8932 8134
rect 8988 8132 9012 8134
rect 9068 8132 9074 8134
rect 8766 8112 9074 8132
rect 9034 7984 9090 7993
rect 9034 7919 9090 7928
rect 9048 7886 9076 7919
rect 9036 7880 9088 7886
rect 9036 7822 9088 7828
rect 8668 7336 8720 7342
rect 8668 7278 8720 7284
rect 8576 6996 8628 7002
rect 8576 6938 8628 6944
rect 8680 6866 8708 7278
rect 9048 7188 9076 7822
rect 9140 7546 9168 8230
rect 9232 7546 9260 8910
rect 9312 8900 9364 8906
rect 9312 8842 9364 8848
rect 9324 8265 9352 8842
rect 9404 8832 9456 8838
rect 9404 8774 9456 8780
rect 9310 8256 9366 8265
rect 9310 8191 9366 8200
rect 9128 7540 9180 7546
rect 9128 7482 9180 7488
rect 9220 7540 9272 7546
rect 9220 7482 9272 7488
rect 9048 7160 9168 7188
rect 8766 7100 9074 7120
rect 8766 7098 8772 7100
rect 8828 7098 8852 7100
rect 8908 7098 8932 7100
rect 8988 7098 9012 7100
rect 9068 7098 9074 7100
rect 8828 7046 8830 7098
rect 9010 7046 9012 7098
rect 8766 7044 8772 7046
rect 8828 7044 8852 7046
rect 8908 7044 8932 7046
rect 8988 7044 9012 7046
rect 9068 7044 9074 7046
rect 8766 7024 9074 7044
rect 8668 6860 8720 6866
rect 8668 6802 8720 6808
rect 9140 6798 9168 7160
rect 9416 7041 9444 8774
rect 9508 8634 9536 9998
rect 10876 9920 10928 9926
rect 10876 9862 10928 9868
rect 9496 8628 9548 8634
rect 9496 8570 9548 8576
rect 9588 8016 9640 8022
rect 9588 7958 9640 7964
rect 9496 7404 9548 7410
rect 9496 7346 9548 7352
rect 9402 7032 9458 7041
rect 9402 6967 9458 6976
rect 9128 6792 9180 6798
rect 9128 6734 9180 6740
rect 8668 6724 8720 6730
rect 8668 6666 8720 6672
rect 8404 6446 8524 6474
rect 8300 4752 8352 4758
rect 8300 4694 8352 4700
rect 8404 4690 8432 6446
rect 8484 6316 8536 6322
rect 8484 6258 8536 6264
rect 8496 4826 8524 6258
rect 8680 5710 8708 6666
rect 9128 6656 9180 6662
rect 9128 6598 9180 6604
rect 9220 6656 9272 6662
rect 9220 6598 9272 6604
rect 9140 6458 9168 6598
rect 9128 6452 9180 6458
rect 9128 6394 9180 6400
rect 9128 6112 9180 6118
rect 9128 6054 9180 6060
rect 8766 6012 9074 6032
rect 8766 6010 8772 6012
rect 8828 6010 8852 6012
rect 8908 6010 8932 6012
rect 8988 6010 9012 6012
rect 9068 6010 9074 6012
rect 8828 5958 8830 6010
rect 9010 5958 9012 6010
rect 8766 5956 8772 5958
rect 8828 5956 8852 5958
rect 8908 5956 8932 5958
rect 8988 5956 9012 5958
rect 9068 5956 9074 5958
rect 8766 5936 9074 5956
rect 8668 5704 8720 5710
rect 9140 5658 9168 6054
rect 8668 5646 8720 5652
rect 9048 5642 9168 5658
rect 9036 5636 9168 5642
rect 9088 5630 9168 5636
rect 9036 5578 9088 5584
rect 9128 5568 9180 5574
rect 9128 5510 9180 5516
rect 8576 5160 8628 5166
rect 8760 5160 8812 5166
rect 8576 5102 8628 5108
rect 8680 5108 8760 5114
rect 8680 5102 8812 5108
rect 8484 4820 8536 4826
rect 8484 4762 8536 4768
rect 8208 4684 8260 4690
rect 8208 4626 8260 4632
rect 8392 4684 8444 4690
rect 8392 4626 8444 4632
rect 8116 3052 8168 3058
rect 6368 2984 6420 2990
rect 6368 2926 6420 2932
rect 5666 2748 5974 2768
rect 5666 2746 5672 2748
rect 5728 2746 5752 2748
rect 5808 2746 5832 2748
rect 5888 2746 5912 2748
rect 5968 2746 5974 2748
rect 5728 2694 5730 2746
rect 5910 2694 5912 2746
rect 5666 2692 5672 2694
rect 5728 2692 5752 2694
rect 5808 2692 5832 2694
rect 5888 2692 5912 2694
rect 5968 2692 5974 2694
rect 5666 2672 5974 2692
rect 4116 2204 4424 2224
rect 4116 2202 4122 2204
rect 4178 2202 4202 2204
rect 4258 2202 4282 2204
rect 4338 2202 4362 2204
rect 4418 2202 4424 2204
rect 4178 2150 4180 2202
rect 4360 2150 4362 2202
rect 4116 2148 4122 2150
rect 4178 2148 4202 2150
rect 4258 2148 4282 2150
rect 4338 2148 4362 2150
rect 4418 2148 4424 2150
rect 4116 2128 4424 2148
rect 7216 2204 7524 2224
rect 7216 2202 7222 2204
rect 7278 2202 7302 2204
rect 7358 2202 7382 2204
rect 7438 2202 7462 2204
rect 7518 2202 7524 2204
rect 7278 2150 7280 2202
rect 7460 2150 7462 2202
rect 7216 2148 7222 2150
rect 7278 2148 7302 2150
rect 7358 2148 7382 2150
rect 7438 2148 7462 2150
rect 7518 2148 7524 2150
rect 7216 2128 7524 2148
rect 7852 1902 7880 3046
rect 8116 2994 8168 3000
rect 8128 2774 8156 2994
rect 7944 2746 8156 2774
rect 7944 2650 7972 2746
rect 7932 2644 7984 2650
rect 7932 2586 7984 2592
rect 8220 2106 8248 4626
rect 8392 4548 8444 4554
rect 8392 4490 8444 4496
rect 8300 4276 8352 4282
rect 8300 4218 8352 4224
rect 8312 3058 8340 4218
rect 8404 3194 8432 4490
rect 8588 4282 8616 5102
rect 8680 5086 8800 5102
rect 8576 4276 8628 4282
rect 8576 4218 8628 4224
rect 8484 4208 8536 4214
rect 8484 4150 8536 4156
rect 8496 3398 8524 4150
rect 8576 4140 8628 4146
rect 8576 4082 8628 4088
rect 8588 3738 8616 4082
rect 8576 3732 8628 3738
rect 8576 3674 8628 3680
rect 8484 3392 8536 3398
rect 8484 3334 8536 3340
rect 8680 3194 8708 5086
rect 8766 4924 9074 4944
rect 8766 4922 8772 4924
rect 8828 4922 8852 4924
rect 8908 4922 8932 4924
rect 8988 4922 9012 4924
rect 9068 4922 9074 4924
rect 8828 4870 8830 4922
rect 9010 4870 9012 4922
rect 8766 4868 8772 4870
rect 8828 4868 8852 4870
rect 8908 4868 8932 4870
rect 8988 4868 9012 4870
rect 9068 4868 9074 4870
rect 8766 4848 9074 4868
rect 8944 4480 8996 4486
rect 8944 4422 8996 4428
rect 8956 4282 8984 4422
rect 8944 4276 8996 4282
rect 8944 4218 8996 4224
rect 8766 3836 9074 3856
rect 8766 3834 8772 3836
rect 8828 3834 8852 3836
rect 8908 3834 8932 3836
rect 8988 3834 9012 3836
rect 9068 3834 9074 3836
rect 8828 3782 8830 3834
rect 9010 3782 9012 3834
rect 8766 3780 8772 3782
rect 8828 3780 8852 3782
rect 8908 3780 8932 3782
rect 8988 3780 9012 3782
rect 9068 3780 9074 3782
rect 8766 3760 9074 3780
rect 9140 3482 9168 5510
rect 9232 4826 9260 6598
rect 9312 6384 9364 6390
rect 9312 6326 9364 6332
rect 9324 5914 9352 6326
rect 9404 6112 9456 6118
rect 9404 6054 9456 6060
rect 9312 5908 9364 5914
rect 9312 5850 9364 5856
rect 9312 5636 9364 5642
rect 9312 5578 9364 5584
rect 9220 4820 9272 4826
rect 9220 4762 9272 4768
rect 9324 4570 9352 5578
rect 9416 5001 9444 6054
rect 9508 5846 9536 7346
rect 9496 5840 9548 5846
rect 9496 5782 9548 5788
rect 9496 5228 9548 5234
rect 9496 5170 9548 5176
rect 9402 4992 9458 5001
rect 9402 4927 9458 4936
rect 9324 4542 9444 4570
rect 9312 4480 9364 4486
rect 9312 4422 9364 4428
rect 9324 4146 9352 4422
rect 9312 4140 9364 4146
rect 9312 4082 9364 4088
rect 9220 4072 9272 4078
rect 9220 4014 9272 4020
rect 9048 3454 9168 3482
rect 8392 3188 8444 3194
rect 8392 3130 8444 3136
rect 8668 3188 8720 3194
rect 8668 3130 8720 3136
rect 9048 3126 9076 3454
rect 9128 3392 9180 3398
rect 9128 3334 9180 3340
rect 9036 3120 9088 3126
rect 9036 3062 9088 3068
rect 8300 3052 8352 3058
rect 8300 2994 8352 3000
rect 8300 2916 8352 2922
rect 8300 2858 8352 2864
rect 8312 2514 8340 2858
rect 8766 2748 9074 2768
rect 8766 2746 8772 2748
rect 8828 2746 8852 2748
rect 8908 2746 8932 2748
rect 8988 2746 9012 2748
rect 9068 2746 9074 2748
rect 8828 2694 8830 2746
rect 9010 2694 9012 2746
rect 8766 2692 8772 2694
rect 8828 2692 8852 2694
rect 8908 2692 8932 2694
rect 8988 2692 9012 2694
rect 9068 2692 9074 2694
rect 8766 2672 9074 2692
rect 8300 2508 8352 2514
rect 8300 2450 8352 2456
rect 9140 2446 9168 3334
rect 9232 2650 9260 4014
rect 9220 2644 9272 2650
rect 9220 2586 9272 2592
rect 9324 2582 9352 4082
rect 9416 4010 9444 4542
rect 9404 4004 9456 4010
rect 9404 3946 9456 3952
rect 9416 3738 9444 3946
rect 9404 3732 9456 3738
rect 9404 3674 9456 3680
rect 9508 3534 9536 5170
rect 9600 5114 9628 7958
rect 10888 7857 10916 9862
rect 13818 9208 13874 9217
rect 13818 9143 13820 9152
rect 13872 9143 13874 9152
rect 13820 9114 13872 9120
rect 16592 8673 16620 10406
rect 16684 9178 16712 11863
rect 16672 9172 16724 9178
rect 16672 9114 16724 9120
rect 16578 8664 16634 8673
rect 16578 8599 16634 8608
rect 10874 7848 10930 7857
rect 10874 7783 10930 7792
rect 12256 7744 12308 7750
rect 12256 7686 12308 7692
rect 11060 7200 11112 7206
rect 11060 7142 11112 7148
rect 11072 6225 11100 7142
rect 11058 6216 11114 6225
rect 11058 6151 11114 6160
rect 12268 5409 12296 7686
rect 12254 5400 12310 5409
rect 12254 5335 12310 5344
rect 9600 5086 9720 5114
rect 9588 5024 9640 5030
rect 9588 4966 9640 4972
rect 9496 3528 9548 3534
rect 9496 3470 9548 3476
rect 9494 3360 9550 3369
rect 9494 3295 9550 3304
rect 9404 2848 9456 2854
rect 9404 2790 9456 2796
rect 9312 2576 9364 2582
rect 9416 2553 9444 2790
rect 9508 2650 9536 3295
rect 9496 2644 9548 2650
rect 9496 2586 9548 2592
rect 9312 2518 9364 2524
rect 9402 2544 9458 2553
rect 9402 2479 9458 2488
rect 9128 2440 9180 2446
rect 9128 2382 9180 2388
rect 8208 2100 8260 2106
rect 8208 2042 8260 2048
rect 7840 1896 7892 1902
rect 7840 1838 7892 1844
rect 9220 1896 9272 1902
rect 9220 1838 9272 1844
rect 9128 1760 9180 1766
rect 9128 1702 9180 1708
rect 5666 1660 5974 1680
rect 5666 1658 5672 1660
rect 5728 1658 5752 1660
rect 5808 1658 5832 1660
rect 5888 1658 5912 1660
rect 5968 1658 5974 1660
rect 5728 1606 5730 1658
rect 5910 1606 5912 1658
rect 5666 1604 5672 1606
rect 5728 1604 5752 1606
rect 5808 1604 5832 1606
rect 5888 1604 5912 1606
rect 5968 1604 5974 1606
rect 5666 1584 5974 1604
rect 8766 1660 9074 1680
rect 8766 1658 8772 1660
rect 8828 1658 8852 1660
rect 8908 1658 8932 1660
rect 8988 1658 9012 1660
rect 9068 1658 9074 1660
rect 8828 1606 8830 1658
rect 9010 1606 9012 1658
rect 8766 1604 8772 1606
rect 8828 1604 8852 1606
rect 8908 1604 8932 1606
rect 8988 1604 9012 1606
rect 9068 1604 9074 1606
rect 8766 1584 9074 1604
rect 4116 1116 4424 1136
rect 4116 1114 4122 1116
rect 4178 1114 4202 1116
rect 4258 1114 4282 1116
rect 4338 1114 4362 1116
rect 4418 1114 4424 1116
rect 4178 1062 4180 1114
rect 4360 1062 4362 1114
rect 4116 1060 4122 1062
rect 4178 1060 4202 1062
rect 4258 1060 4282 1062
rect 4338 1060 4362 1062
rect 4418 1060 4424 1062
rect 4116 1040 4424 1060
rect 7216 1116 7524 1136
rect 7216 1114 7222 1116
rect 7278 1114 7302 1116
rect 7358 1114 7382 1116
rect 7438 1114 7462 1116
rect 7518 1114 7524 1116
rect 7278 1062 7280 1114
rect 7460 1062 7462 1114
rect 7216 1060 7222 1062
rect 7278 1060 7302 1062
rect 7358 1060 7382 1062
rect 7438 1060 7462 1062
rect 7518 1060 7524 1062
rect 7216 1040 7524 1060
rect 9140 513 9168 1702
rect 9232 921 9260 1838
rect 9600 1329 9628 4966
rect 9692 3126 9720 5086
rect 16580 5092 16632 5098
rect 16580 5034 16632 5040
rect 16592 4185 16620 5034
rect 16578 4176 16634 4185
rect 16578 4111 16634 4120
rect 16580 3936 16632 3942
rect 16580 3878 16632 3884
rect 16592 3777 16620 3878
rect 16578 3768 16634 3777
rect 16578 3703 16634 3712
rect 9680 3120 9732 3126
rect 9680 3062 9732 3068
rect 16580 2984 16632 2990
rect 16578 2952 16580 2961
rect 16632 2952 16634 2961
rect 16578 2887 16634 2896
rect 16580 2372 16632 2378
rect 16580 2314 16632 2320
rect 16592 2145 16620 2314
rect 16578 2136 16634 2145
rect 16578 2071 16634 2080
rect 16580 1828 16632 1834
rect 16580 1770 16632 1776
rect 16592 1737 16620 1770
rect 16578 1728 16634 1737
rect 16578 1663 16634 1672
rect 9586 1320 9642 1329
rect 9586 1255 9642 1264
rect 9218 912 9274 921
rect 9218 847 9274 856
rect 9126 504 9182 513
rect 9126 439 9182 448
<< via2 >>
rect 1674 11600 1730 11656
rect 1398 10920 1454 10976
rect 1214 10104 1270 10160
rect 1398 10004 1400 10024
rect 1400 10004 1452 10024
rect 1452 10004 1454 10024
rect 1398 9968 1454 10004
rect 1398 9832 1454 9888
rect 1306 9424 1362 9480
rect 1214 9016 1270 9072
rect 1766 9560 1822 9616
rect 2410 12144 2466 12200
rect 2042 11056 2098 11112
rect 1950 9968 2006 10024
rect 1582 9016 1638 9072
rect 1674 7520 1730 7576
rect 2134 10668 2190 10704
rect 2134 10648 2136 10668
rect 2136 10648 2188 10668
rect 2188 10648 2190 10668
rect 2134 10532 2190 10568
rect 2134 10512 2136 10532
rect 2136 10512 2188 10532
rect 2188 10512 2190 10532
rect 2870 11736 2926 11792
rect 2572 11450 2628 11452
rect 2652 11450 2708 11452
rect 2732 11450 2788 11452
rect 2812 11450 2868 11452
rect 2572 11398 2618 11450
rect 2618 11398 2628 11450
rect 2652 11398 2682 11450
rect 2682 11398 2694 11450
rect 2694 11398 2708 11450
rect 2732 11398 2746 11450
rect 2746 11398 2758 11450
rect 2758 11398 2788 11450
rect 2812 11398 2822 11450
rect 2822 11398 2868 11450
rect 2572 11396 2628 11398
rect 2652 11396 2708 11398
rect 2732 11396 2788 11398
rect 2812 11396 2868 11398
rect 2594 11192 2650 11248
rect 2410 11056 2466 11112
rect 2778 10784 2834 10840
rect 3054 10376 3110 10432
rect 2572 10362 2628 10364
rect 2652 10362 2708 10364
rect 2732 10362 2788 10364
rect 2812 10362 2868 10364
rect 2572 10310 2618 10362
rect 2618 10310 2628 10362
rect 2652 10310 2682 10362
rect 2682 10310 2694 10362
rect 2694 10310 2708 10362
rect 2732 10310 2746 10362
rect 2746 10310 2758 10362
rect 2758 10310 2788 10362
rect 2812 10310 2822 10362
rect 2822 10310 2868 10362
rect 2572 10308 2628 10310
rect 2652 10308 2708 10310
rect 2732 10308 2788 10310
rect 2812 10308 2868 10310
rect 2962 10240 3018 10296
rect 2042 9424 2098 9480
rect 2134 9016 2190 9072
rect 2042 8880 2098 8936
rect 1950 8356 2006 8392
rect 1950 8336 1952 8356
rect 1952 8336 2004 8356
rect 2004 8336 2006 8356
rect 2318 9832 2374 9888
rect 2318 9424 2374 9480
rect 2594 9580 2650 9616
rect 2594 9560 2596 9580
rect 2596 9560 2648 9580
rect 2648 9560 2650 9580
rect 2962 9424 3018 9480
rect 2572 9274 2628 9276
rect 2652 9274 2708 9276
rect 2732 9274 2788 9276
rect 2812 9274 2868 9276
rect 2572 9222 2618 9274
rect 2618 9222 2628 9274
rect 2652 9222 2682 9274
rect 2682 9222 2694 9274
rect 2694 9222 2708 9274
rect 2732 9222 2746 9274
rect 2746 9222 2758 9274
rect 2758 9222 2788 9274
rect 2812 9222 2822 9274
rect 2822 9222 2868 9274
rect 2572 9220 2628 9222
rect 2652 9220 2708 9222
rect 2732 9220 2788 9222
rect 2812 9220 2868 9222
rect 2572 8186 2628 8188
rect 2652 8186 2708 8188
rect 2732 8186 2788 8188
rect 2812 8186 2868 8188
rect 2572 8134 2618 8186
rect 2618 8134 2628 8186
rect 2652 8134 2682 8186
rect 2682 8134 2694 8186
rect 2694 8134 2708 8186
rect 2732 8134 2746 8186
rect 2746 8134 2758 8186
rect 2758 8134 2788 8186
rect 2812 8134 2822 8186
rect 2822 8134 2868 8186
rect 2572 8132 2628 8134
rect 2652 8132 2708 8134
rect 2732 8132 2788 8134
rect 2812 8132 2868 8134
rect 2686 7928 2742 7984
rect 2778 7520 2834 7576
rect 3054 8064 3110 8120
rect 3054 7928 3110 7984
rect 2410 7248 2466 7304
rect 2962 7248 3018 7304
rect 2572 7098 2628 7100
rect 2652 7098 2708 7100
rect 2732 7098 2788 7100
rect 2812 7098 2868 7100
rect 2572 7046 2618 7098
rect 2618 7046 2628 7098
rect 2652 7046 2682 7098
rect 2682 7046 2694 7098
rect 2694 7046 2708 7098
rect 2732 7046 2746 7098
rect 2746 7046 2758 7098
rect 2758 7046 2788 7098
rect 2812 7046 2822 7098
rect 2822 7046 2868 7098
rect 2572 7044 2628 7046
rect 2652 7044 2708 7046
rect 2732 7044 2788 7046
rect 2812 7044 2868 7046
rect 2572 6010 2628 6012
rect 2652 6010 2708 6012
rect 2732 6010 2788 6012
rect 2812 6010 2868 6012
rect 2572 5958 2618 6010
rect 2618 5958 2628 6010
rect 2652 5958 2682 6010
rect 2682 5958 2694 6010
rect 2694 5958 2708 6010
rect 2732 5958 2746 6010
rect 2746 5958 2758 6010
rect 2758 5958 2788 6010
rect 2812 5958 2822 6010
rect 2822 5958 2868 6010
rect 2572 5956 2628 5958
rect 2652 5956 2708 5958
rect 2732 5956 2788 5958
rect 2812 5956 2868 5958
rect 3514 11328 3570 11384
rect 3514 10784 3570 10840
rect 3330 9424 3386 9480
rect 3422 8916 3424 8936
rect 3424 8916 3476 8936
rect 3476 8916 3478 8936
rect 3422 8880 3478 8916
rect 4122 10906 4178 10908
rect 4202 10906 4258 10908
rect 4282 10906 4338 10908
rect 4362 10906 4418 10908
rect 4122 10854 4168 10906
rect 4168 10854 4178 10906
rect 4202 10854 4232 10906
rect 4232 10854 4244 10906
rect 4244 10854 4258 10906
rect 4282 10854 4296 10906
rect 4296 10854 4308 10906
rect 4308 10854 4338 10906
rect 4362 10854 4372 10906
rect 4372 10854 4418 10906
rect 4122 10852 4178 10854
rect 4202 10852 4258 10854
rect 4282 10852 4338 10854
rect 4362 10852 4418 10854
rect 5170 11600 5226 11656
rect 4526 10648 4582 10704
rect 3514 8472 3570 8528
rect 3422 8084 3478 8120
rect 3422 8064 3424 8084
rect 3424 8064 3476 8084
rect 3476 8064 3478 8084
rect 4158 10376 4214 10432
rect 3882 10240 3938 10296
rect 3790 8744 3846 8800
rect 3790 8064 3846 8120
rect 4122 9818 4178 9820
rect 4202 9818 4258 9820
rect 4282 9818 4338 9820
rect 4362 9818 4418 9820
rect 4122 9766 4168 9818
rect 4168 9766 4178 9818
rect 4202 9766 4232 9818
rect 4232 9766 4244 9818
rect 4244 9766 4258 9818
rect 4282 9766 4296 9818
rect 4296 9766 4308 9818
rect 4308 9766 4338 9818
rect 4362 9766 4372 9818
rect 4372 9766 4418 9818
rect 4122 9764 4178 9766
rect 4202 9764 4258 9766
rect 4282 9764 4338 9766
rect 4362 9764 4418 9766
rect 4342 8900 4398 8936
rect 4342 8880 4344 8900
rect 4344 8880 4396 8900
rect 4396 8880 4398 8900
rect 4122 8730 4178 8732
rect 4202 8730 4258 8732
rect 4282 8730 4338 8732
rect 4362 8730 4418 8732
rect 4122 8678 4168 8730
rect 4168 8678 4178 8730
rect 4202 8678 4232 8730
rect 4232 8678 4244 8730
rect 4244 8678 4258 8730
rect 4282 8678 4296 8730
rect 4296 8678 4308 8730
rect 4308 8678 4338 8730
rect 4362 8678 4372 8730
rect 4372 8678 4418 8730
rect 4122 8676 4178 8678
rect 4202 8676 4258 8678
rect 4282 8676 4338 8678
rect 4362 8676 4418 8678
rect 5078 11056 5134 11112
rect 5672 11450 5728 11452
rect 5752 11450 5808 11452
rect 5832 11450 5888 11452
rect 5912 11450 5968 11452
rect 5672 11398 5718 11450
rect 5718 11398 5728 11450
rect 5752 11398 5782 11450
rect 5782 11398 5794 11450
rect 5794 11398 5808 11450
rect 5832 11398 5846 11450
rect 5846 11398 5858 11450
rect 5858 11398 5888 11450
rect 5912 11398 5922 11450
rect 5922 11398 5968 11450
rect 5672 11396 5728 11398
rect 5752 11396 5808 11398
rect 5832 11396 5888 11398
rect 5912 11396 5968 11398
rect 5538 11328 5594 11384
rect 5446 11192 5502 11248
rect 5262 11092 5264 11112
rect 5264 11092 5316 11112
rect 5316 11092 5318 11112
rect 5262 11056 5318 11092
rect 5998 11056 6054 11112
rect 5672 10362 5728 10364
rect 5752 10362 5808 10364
rect 5832 10362 5888 10364
rect 5912 10362 5968 10364
rect 5672 10310 5718 10362
rect 5718 10310 5728 10362
rect 5752 10310 5782 10362
rect 5782 10310 5794 10362
rect 5794 10310 5808 10362
rect 5832 10310 5846 10362
rect 5846 10310 5858 10362
rect 5858 10310 5888 10362
rect 5912 10310 5922 10362
rect 5922 10310 5968 10362
rect 5672 10308 5728 10310
rect 5752 10308 5808 10310
rect 5832 10308 5888 10310
rect 5912 10308 5968 10310
rect 5998 9580 6054 9616
rect 5998 9560 6000 9580
rect 6000 9560 6052 9580
rect 6052 9560 6054 9580
rect 4066 8084 4122 8120
rect 4066 8064 4068 8084
rect 4068 8064 4120 8084
rect 4120 8064 4122 8084
rect 4122 7642 4178 7644
rect 4202 7642 4258 7644
rect 4282 7642 4338 7644
rect 4362 7642 4418 7644
rect 4122 7590 4168 7642
rect 4168 7590 4178 7642
rect 4202 7590 4232 7642
rect 4232 7590 4244 7642
rect 4244 7590 4258 7642
rect 4282 7590 4296 7642
rect 4296 7590 4308 7642
rect 4308 7590 4338 7642
rect 4362 7590 4372 7642
rect 4372 7590 4418 7642
rect 4122 7588 4178 7590
rect 4202 7588 4258 7590
rect 4282 7588 4338 7590
rect 4362 7588 4418 7590
rect 4122 6554 4178 6556
rect 4202 6554 4258 6556
rect 4282 6554 4338 6556
rect 4362 6554 4418 6556
rect 4122 6502 4168 6554
rect 4168 6502 4178 6554
rect 4202 6502 4232 6554
rect 4232 6502 4244 6554
rect 4244 6502 4258 6554
rect 4282 6502 4296 6554
rect 4296 6502 4308 6554
rect 4308 6502 4338 6554
rect 4362 6502 4372 6554
rect 4372 6502 4418 6554
rect 4122 6500 4178 6502
rect 4202 6500 4258 6502
rect 4282 6500 4338 6502
rect 4362 6500 4418 6502
rect 4122 5466 4178 5468
rect 4202 5466 4258 5468
rect 4282 5466 4338 5468
rect 4362 5466 4418 5468
rect 4122 5414 4168 5466
rect 4168 5414 4178 5466
rect 4202 5414 4232 5466
rect 4232 5414 4244 5466
rect 4244 5414 4258 5466
rect 4282 5414 4296 5466
rect 4296 5414 4308 5466
rect 4308 5414 4338 5466
rect 4362 5414 4372 5466
rect 4372 5414 4418 5466
rect 4122 5412 4178 5414
rect 4202 5412 4258 5414
rect 4282 5412 4338 5414
rect 4362 5412 4418 5414
rect 5078 7384 5134 7440
rect 5672 9274 5728 9276
rect 5752 9274 5808 9276
rect 5832 9274 5888 9276
rect 5912 9274 5968 9276
rect 5672 9222 5718 9274
rect 5718 9222 5728 9274
rect 5752 9222 5782 9274
rect 5782 9222 5794 9274
rect 5794 9222 5808 9274
rect 5832 9222 5846 9274
rect 5846 9222 5858 9274
rect 5858 9222 5888 9274
rect 5912 9222 5922 9274
rect 5922 9222 5968 9274
rect 5672 9220 5728 9222
rect 5752 9220 5808 9222
rect 5832 9220 5888 9222
rect 5912 9220 5968 9222
rect 5538 8880 5594 8936
rect 5722 8508 5724 8528
rect 5724 8508 5776 8528
rect 5776 8508 5778 8528
rect 5722 8472 5778 8508
rect 5672 8186 5728 8188
rect 5752 8186 5808 8188
rect 5832 8186 5888 8188
rect 5912 8186 5968 8188
rect 5672 8134 5718 8186
rect 5718 8134 5728 8186
rect 5752 8134 5782 8186
rect 5782 8134 5794 8186
rect 5794 8134 5808 8186
rect 5832 8134 5846 8186
rect 5846 8134 5858 8186
rect 5858 8134 5888 8186
rect 5912 8134 5922 8186
rect 5922 8134 5968 8186
rect 5672 8132 5728 8134
rect 5752 8132 5808 8134
rect 5832 8132 5888 8134
rect 5912 8132 5968 8134
rect 6366 7928 6422 7984
rect 5672 7098 5728 7100
rect 5752 7098 5808 7100
rect 5832 7098 5888 7100
rect 5912 7098 5968 7100
rect 5672 7046 5718 7098
rect 5718 7046 5728 7098
rect 5752 7046 5782 7098
rect 5782 7046 5794 7098
rect 5794 7046 5808 7098
rect 5832 7046 5846 7098
rect 5846 7046 5858 7098
rect 5858 7046 5888 7098
rect 5912 7046 5922 7098
rect 5922 7046 5968 7098
rect 5672 7044 5728 7046
rect 5752 7044 5808 7046
rect 5832 7044 5888 7046
rect 5912 7044 5968 7046
rect 6642 11348 6698 11384
rect 6642 11328 6644 11348
rect 6644 11328 6696 11348
rect 6696 11328 6698 11348
rect 6734 9016 6790 9072
rect 5672 6010 5728 6012
rect 5752 6010 5808 6012
rect 5832 6010 5888 6012
rect 5912 6010 5968 6012
rect 5672 5958 5718 6010
rect 5718 5958 5728 6010
rect 5752 5958 5782 6010
rect 5782 5958 5794 6010
rect 5794 5958 5808 6010
rect 5832 5958 5846 6010
rect 5846 5958 5858 6010
rect 5858 5958 5888 6010
rect 5912 5958 5922 6010
rect 5922 5958 5968 6010
rect 5672 5956 5728 5958
rect 5752 5956 5808 5958
rect 5832 5956 5888 5958
rect 5912 5956 5968 5958
rect 3698 4564 3700 4584
rect 3700 4564 3752 4584
rect 3752 4564 3754 4584
rect 3698 4528 3754 4564
rect 4122 4378 4178 4380
rect 4202 4378 4258 4380
rect 4282 4378 4338 4380
rect 4362 4378 4418 4380
rect 4122 4326 4168 4378
rect 4168 4326 4178 4378
rect 4202 4326 4232 4378
rect 4232 4326 4244 4378
rect 4244 4326 4258 4378
rect 4282 4326 4296 4378
rect 4296 4326 4308 4378
rect 4308 4326 4338 4378
rect 4362 4326 4372 4378
rect 4372 4326 4418 4378
rect 4122 4324 4178 4326
rect 4202 4324 4258 4326
rect 4282 4324 4338 4326
rect 4362 4324 4418 4326
rect 2686 3304 2742 3360
rect 4122 3290 4178 3292
rect 4202 3290 4258 3292
rect 4282 3290 4338 3292
rect 4362 3290 4418 3292
rect 4122 3238 4168 3290
rect 4168 3238 4178 3290
rect 4202 3238 4232 3290
rect 4232 3238 4244 3290
rect 4244 3238 4258 3290
rect 4282 3238 4296 3290
rect 4296 3238 4308 3290
rect 4308 3238 4338 3290
rect 4362 3238 4372 3290
rect 4372 3238 4418 3290
rect 4122 3236 4178 3238
rect 4202 3236 4258 3238
rect 4282 3236 4338 3238
rect 4362 3236 4418 3238
rect 5672 4922 5728 4924
rect 5752 4922 5808 4924
rect 5832 4922 5888 4924
rect 5912 4922 5968 4924
rect 5672 4870 5718 4922
rect 5718 4870 5728 4922
rect 5752 4870 5782 4922
rect 5782 4870 5794 4922
rect 5794 4870 5808 4922
rect 5832 4870 5846 4922
rect 5846 4870 5858 4922
rect 5858 4870 5888 4922
rect 5912 4870 5922 4922
rect 5922 4870 5968 4922
rect 5672 4868 5728 4870
rect 5752 4868 5808 4870
rect 5832 4868 5888 4870
rect 5912 4868 5968 4870
rect 5722 4564 5724 4584
rect 5724 4564 5776 4584
rect 5776 4564 5778 4584
rect 5722 4528 5778 4564
rect 5672 3834 5728 3836
rect 5752 3834 5808 3836
rect 5832 3834 5888 3836
rect 5912 3834 5968 3836
rect 5672 3782 5718 3834
rect 5718 3782 5728 3834
rect 5752 3782 5782 3834
rect 5782 3782 5794 3834
rect 5794 3782 5808 3834
rect 5832 3782 5846 3834
rect 5846 3782 5858 3834
rect 5858 3782 5888 3834
rect 5912 3782 5922 3834
rect 5922 3782 5968 3834
rect 5672 3780 5728 3782
rect 5752 3780 5808 3782
rect 5832 3780 5888 3782
rect 5912 3780 5968 3782
rect 7222 10906 7278 10908
rect 7302 10906 7358 10908
rect 7382 10906 7438 10908
rect 7462 10906 7518 10908
rect 7222 10854 7268 10906
rect 7268 10854 7278 10906
rect 7302 10854 7332 10906
rect 7332 10854 7344 10906
rect 7344 10854 7358 10906
rect 7382 10854 7396 10906
rect 7396 10854 7408 10906
rect 7408 10854 7438 10906
rect 7462 10854 7472 10906
rect 7472 10854 7518 10906
rect 7222 10852 7278 10854
rect 7302 10852 7358 10854
rect 7382 10852 7438 10854
rect 7462 10852 7518 10854
rect 7470 10512 7526 10568
rect 7222 9818 7278 9820
rect 7302 9818 7358 9820
rect 7382 9818 7438 9820
rect 7462 9818 7518 9820
rect 7222 9766 7268 9818
rect 7268 9766 7278 9818
rect 7302 9766 7332 9818
rect 7332 9766 7344 9818
rect 7344 9766 7358 9818
rect 7382 9766 7396 9818
rect 7396 9766 7408 9818
rect 7408 9766 7438 9818
rect 7462 9766 7472 9818
rect 7472 9766 7518 9818
rect 7222 9764 7278 9766
rect 7302 9764 7358 9766
rect 7382 9764 7438 9766
rect 7462 9764 7518 9766
rect 8022 11736 8078 11792
rect 8206 11348 8262 11384
rect 8206 11328 8208 11348
rect 8208 11328 8260 11348
rect 8260 11328 8262 11348
rect 16670 11872 16726 11928
rect 7222 8730 7278 8732
rect 7302 8730 7358 8732
rect 7382 8730 7438 8732
rect 7462 8730 7518 8732
rect 7222 8678 7268 8730
rect 7268 8678 7278 8730
rect 7302 8678 7332 8730
rect 7332 8678 7344 8730
rect 7344 8678 7358 8730
rect 7382 8678 7396 8730
rect 7396 8678 7408 8730
rect 7408 8678 7438 8730
rect 7462 8678 7472 8730
rect 7472 8678 7518 8730
rect 7222 8676 7278 8678
rect 7302 8676 7358 8678
rect 7382 8676 7438 8678
rect 7462 8676 7518 8678
rect 7222 7642 7278 7644
rect 7302 7642 7358 7644
rect 7382 7642 7438 7644
rect 7462 7642 7518 7644
rect 7222 7590 7268 7642
rect 7268 7590 7278 7642
rect 7302 7590 7332 7642
rect 7332 7590 7344 7642
rect 7344 7590 7358 7642
rect 7382 7590 7396 7642
rect 7396 7590 7408 7642
rect 7408 7590 7438 7642
rect 7462 7590 7472 7642
rect 7472 7590 7518 7642
rect 7222 7588 7278 7590
rect 7302 7588 7358 7590
rect 7382 7588 7438 7590
rect 7462 7588 7518 7590
rect 8206 9424 8262 9480
rect 8206 8336 8262 8392
rect 7222 6554 7278 6556
rect 7302 6554 7358 6556
rect 7382 6554 7438 6556
rect 7462 6554 7518 6556
rect 7222 6502 7268 6554
rect 7268 6502 7278 6554
rect 7302 6502 7332 6554
rect 7332 6502 7344 6554
rect 7344 6502 7358 6554
rect 7382 6502 7396 6554
rect 7396 6502 7408 6554
rect 7408 6502 7438 6554
rect 7462 6502 7472 6554
rect 7472 6502 7518 6554
rect 7222 6500 7278 6502
rect 7302 6500 7358 6502
rect 7382 6500 7438 6502
rect 7462 6500 7518 6502
rect 7222 5466 7278 5468
rect 7302 5466 7358 5468
rect 7382 5466 7438 5468
rect 7462 5466 7518 5468
rect 7222 5414 7268 5466
rect 7268 5414 7278 5466
rect 7302 5414 7332 5466
rect 7332 5414 7344 5466
rect 7344 5414 7358 5466
rect 7382 5414 7396 5466
rect 7396 5414 7408 5466
rect 7408 5414 7438 5466
rect 7462 5414 7472 5466
rect 7472 5414 7518 5466
rect 7222 5412 7278 5414
rect 7302 5412 7358 5414
rect 7382 5412 7438 5414
rect 7462 5412 7518 5414
rect 8114 5752 8170 5808
rect 7222 4378 7278 4380
rect 7302 4378 7358 4380
rect 7382 4378 7438 4380
rect 7462 4378 7518 4380
rect 7222 4326 7268 4378
rect 7268 4326 7278 4378
rect 7302 4326 7332 4378
rect 7332 4326 7344 4378
rect 7344 4326 7358 4378
rect 7382 4326 7396 4378
rect 7396 4326 7408 4378
rect 7408 4326 7438 4378
rect 7462 4326 7472 4378
rect 7472 4326 7518 4378
rect 7222 4324 7278 4326
rect 7302 4324 7358 4326
rect 7382 4324 7438 4326
rect 7462 4324 7518 4326
rect 7930 4528 7986 4584
rect 7222 3290 7278 3292
rect 7302 3290 7358 3292
rect 7382 3290 7438 3292
rect 7462 3290 7518 3292
rect 7222 3238 7268 3290
rect 7268 3238 7278 3290
rect 7302 3238 7332 3290
rect 7332 3238 7344 3290
rect 7344 3238 7358 3290
rect 7382 3238 7396 3290
rect 7396 3238 7408 3290
rect 7408 3238 7438 3290
rect 7462 3238 7472 3290
rect 7472 3238 7518 3290
rect 7222 3236 7278 3238
rect 7302 3236 7358 3238
rect 7382 3236 7438 3238
rect 7462 3236 7518 3238
rect 8772 11450 8828 11452
rect 8852 11450 8908 11452
rect 8932 11450 8988 11452
rect 9012 11450 9068 11452
rect 8772 11398 8818 11450
rect 8818 11398 8828 11450
rect 8852 11398 8882 11450
rect 8882 11398 8894 11450
rect 8894 11398 8908 11450
rect 8932 11398 8946 11450
rect 8946 11398 8958 11450
rect 8958 11398 8988 11450
rect 9012 11398 9022 11450
rect 9022 11398 9068 11450
rect 8772 11396 8828 11398
rect 8852 11396 8908 11398
rect 8932 11396 8988 11398
rect 9012 11396 9068 11398
rect 8390 6568 8446 6624
rect 8772 10362 8828 10364
rect 8852 10362 8908 10364
rect 8932 10362 8988 10364
rect 9012 10362 9068 10364
rect 8772 10310 8818 10362
rect 8818 10310 8828 10362
rect 8852 10310 8882 10362
rect 8882 10310 8894 10362
rect 8894 10310 8908 10362
rect 8932 10310 8946 10362
rect 8946 10310 8958 10362
rect 8958 10310 8988 10362
rect 9012 10310 9022 10362
rect 9022 10310 9068 10362
rect 8772 10308 8828 10310
rect 8852 10308 8908 10310
rect 8932 10308 8988 10310
rect 9012 10308 9068 10310
rect 8772 9274 8828 9276
rect 8852 9274 8908 9276
rect 8932 9274 8988 9276
rect 9012 9274 9068 9276
rect 8772 9222 8818 9274
rect 8818 9222 8828 9274
rect 8852 9222 8882 9274
rect 8882 9222 8894 9274
rect 8894 9222 8908 9274
rect 8932 9222 8946 9274
rect 8946 9222 8958 9274
rect 8958 9222 8988 9274
rect 9012 9222 9022 9274
rect 9022 9222 9068 9274
rect 8772 9220 8828 9222
rect 8852 9220 8908 9222
rect 8932 9220 8988 9222
rect 9012 9220 9068 9222
rect 9218 9560 9274 9616
rect 9218 9152 9274 9208
rect 13726 11464 13782 11520
rect 13818 11056 13874 11112
rect 9402 10240 9458 10296
rect 8772 8186 8828 8188
rect 8852 8186 8908 8188
rect 8932 8186 8988 8188
rect 9012 8186 9068 8188
rect 8772 8134 8818 8186
rect 8818 8134 8828 8186
rect 8852 8134 8882 8186
rect 8882 8134 8894 8186
rect 8894 8134 8908 8186
rect 8932 8134 8946 8186
rect 8946 8134 8958 8186
rect 8958 8134 8988 8186
rect 9012 8134 9022 8186
rect 9022 8134 9068 8186
rect 8772 8132 8828 8134
rect 8852 8132 8908 8134
rect 8932 8132 8988 8134
rect 9012 8132 9068 8134
rect 9034 7928 9090 7984
rect 9310 8200 9366 8256
rect 8772 7098 8828 7100
rect 8852 7098 8908 7100
rect 8932 7098 8988 7100
rect 9012 7098 9068 7100
rect 8772 7046 8818 7098
rect 8818 7046 8828 7098
rect 8852 7046 8882 7098
rect 8882 7046 8894 7098
rect 8894 7046 8908 7098
rect 8932 7046 8946 7098
rect 8946 7046 8958 7098
rect 8958 7046 8988 7098
rect 9012 7046 9022 7098
rect 9022 7046 9068 7098
rect 8772 7044 8828 7046
rect 8852 7044 8908 7046
rect 8932 7044 8988 7046
rect 9012 7044 9068 7046
rect 9402 6976 9458 7032
rect 8772 6010 8828 6012
rect 8852 6010 8908 6012
rect 8932 6010 8988 6012
rect 9012 6010 9068 6012
rect 8772 5958 8818 6010
rect 8818 5958 8828 6010
rect 8852 5958 8882 6010
rect 8882 5958 8894 6010
rect 8894 5958 8908 6010
rect 8932 5958 8946 6010
rect 8946 5958 8958 6010
rect 8958 5958 8988 6010
rect 9012 5958 9022 6010
rect 9022 5958 9068 6010
rect 8772 5956 8828 5958
rect 8852 5956 8908 5958
rect 8932 5956 8988 5958
rect 9012 5956 9068 5958
rect 5672 2746 5728 2748
rect 5752 2746 5808 2748
rect 5832 2746 5888 2748
rect 5912 2746 5968 2748
rect 5672 2694 5718 2746
rect 5718 2694 5728 2746
rect 5752 2694 5782 2746
rect 5782 2694 5794 2746
rect 5794 2694 5808 2746
rect 5832 2694 5846 2746
rect 5846 2694 5858 2746
rect 5858 2694 5888 2746
rect 5912 2694 5922 2746
rect 5922 2694 5968 2746
rect 5672 2692 5728 2694
rect 5752 2692 5808 2694
rect 5832 2692 5888 2694
rect 5912 2692 5968 2694
rect 4122 2202 4178 2204
rect 4202 2202 4258 2204
rect 4282 2202 4338 2204
rect 4362 2202 4418 2204
rect 4122 2150 4168 2202
rect 4168 2150 4178 2202
rect 4202 2150 4232 2202
rect 4232 2150 4244 2202
rect 4244 2150 4258 2202
rect 4282 2150 4296 2202
rect 4296 2150 4308 2202
rect 4308 2150 4338 2202
rect 4362 2150 4372 2202
rect 4372 2150 4418 2202
rect 4122 2148 4178 2150
rect 4202 2148 4258 2150
rect 4282 2148 4338 2150
rect 4362 2148 4418 2150
rect 7222 2202 7278 2204
rect 7302 2202 7358 2204
rect 7382 2202 7438 2204
rect 7462 2202 7518 2204
rect 7222 2150 7268 2202
rect 7268 2150 7278 2202
rect 7302 2150 7332 2202
rect 7332 2150 7344 2202
rect 7344 2150 7358 2202
rect 7382 2150 7396 2202
rect 7396 2150 7408 2202
rect 7408 2150 7438 2202
rect 7462 2150 7472 2202
rect 7472 2150 7518 2202
rect 7222 2148 7278 2150
rect 7302 2148 7358 2150
rect 7382 2148 7438 2150
rect 7462 2148 7518 2150
rect 8772 4922 8828 4924
rect 8852 4922 8908 4924
rect 8932 4922 8988 4924
rect 9012 4922 9068 4924
rect 8772 4870 8818 4922
rect 8818 4870 8828 4922
rect 8852 4870 8882 4922
rect 8882 4870 8894 4922
rect 8894 4870 8908 4922
rect 8932 4870 8946 4922
rect 8946 4870 8958 4922
rect 8958 4870 8988 4922
rect 9012 4870 9022 4922
rect 9022 4870 9068 4922
rect 8772 4868 8828 4870
rect 8852 4868 8908 4870
rect 8932 4868 8988 4870
rect 9012 4868 9068 4870
rect 8772 3834 8828 3836
rect 8852 3834 8908 3836
rect 8932 3834 8988 3836
rect 9012 3834 9068 3836
rect 8772 3782 8818 3834
rect 8818 3782 8828 3834
rect 8852 3782 8882 3834
rect 8882 3782 8894 3834
rect 8894 3782 8908 3834
rect 8932 3782 8946 3834
rect 8946 3782 8958 3834
rect 8958 3782 8988 3834
rect 9012 3782 9022 3834
rect 9022 3782 9068 3834
rect 8772 3780 8828 3782
rect 8852 3780 8908 3782
rect 8932 3780 8988 3782
rect 9012 3780 9068 3782
rect 9402 4936 9458 4992
rect 8772 2746 8828 2748
rect 8852 2746 8908 2748
rect 8932 2746 8988 2748
rect 9012 2746 9068 2748
rect 8772 2694 8818 2746
rect 8818 2694 8828 2746
rect 8852 2694 8882 2746
rect 8882 2694 8894 2746
rect 8894 2694 8908 2746
rect 8932 2694 8946 2746
rect 8946 2694 8958 2746
rect 8958 2694 8988 2746
rect 9012 2694 9022 2746
rect 9022 2694 9068 2746
rect 8772 2692 8828 2694
rect 8852 2692 8908 2694
rect 8932 2692 8988 2694
rect 9012 2692 9068 2694
rect 13818 9172 13874 9208
rect 13818 9152 13820 9172
rect 13820 9152 13872 9172
rect 13872 9152 13874 9172
rect 16578 8608 16634 8664
rect 10874 7792 10930 7848
rect 11058 6160 11114 6216
rect 12254 5344 12310 5400
rect 9494 3304 9550 3360
rect 9402 2488 9458 2544
rect 5672 1658 5728 1660
rect 5752 1658 5808 1660
rect 5832 1658 5888 1660
rect 5912 1658 5968 1660
rect 5672 1606 5718 1658
rect 5718 1606 5728 1658
rect 5752 1606 5782 1658
rect 5782 1606 5794 1658
rect 5794 1606 5808 1658
rect 5832 1606 5846 1658
rect 5846 1606 5858 1658
rect 5858 1606 5888 1658
rect 5912 1606 5922 1658
rect 5922 1606 5968 1658
rect 5672 1604 5728 1606
rect 5752 1604 5808 1606
rect 5832 1604 5888 1606
rect 5912 1604 5968 1606
rect 8772 1658 8828 1660
rect 8852 1658 8908 1660
rect 8932 1658 8988 1660
rect 9012 1658 9068 1660
rect 8772 1606 8818 1658
rect 8818 1606 8828 1658
rect 8852 1606 8882 1658
rect 8882 1606 8894 1658
rect 8894 1606 8908 1658
rect 8932 1606 8946 1658
rect 8946 1606 8958 1658
rect 8958 1606 8988 1658
rect 9012 1606 9022 1658
rect 9022 1606 9068 1658
rect 8772 1604 8828 1606
rect 8852 1604 8908 1606
rect 8932 1604 8988 1606
rect 9012 1604 9068 1606
rect 4122 1114 4178 1116
rect 4202 1114 4258 1116
rect 4282 1114 4338 1116
rect 4362 1114 4418 1116
rect 4122 1062 4168 1114
rect 4168 1062 4178 1114
rect 4202 1062 4232 1114
rect 4232 1062 4244 1114
rect 4244 1062 4258 1114
rect 4282 1062 4296 1114
rect 4296 1062 4308 1114
rect 4308 1062 4338 1114
rect 4362 1062 4372 1114
rect 4372 1062 4418 1114
rect 4122 1060 4178 1062
rect 4202 1060 4258 1062
rect 4282 1060 4338 1062
rect 4362 1060 4418 1062
rect 7222 1114 7278 1116
rect 7302 1114 7358 1116
rect 7382 1114 7438 1116
rect 7462 1114 7518 1116
rect 7222 1062 7268 1114
rect 7268 1062 7278 1114
rect 7302 1062 7332 1114
rect 7332 1062 7344 1114
rect 7344 1062 7358 1114
rect 7382 1062 7396 1114
rect 7396 1062 7408 1114
rect 7408 1062 7438 1114
rect 7462 1062 7472 1114
rect 7472 1062 7518 1114
rect 7222 1060 7278 1062
rect 7302 1060 7358 1062
rect 7382 1060 7438 1062
rect 7462 1060 7518 1062
rect 16578 4120 16634 4176
rect 16578 3712 16634 3768
rect 16578 2932 16580 2952
rect 16580 2932 16632 2952
rect 16632 2932 16634 2952
rect 16578 2896 16634 2932
rect 16578 2080 16634 2136
rect 16578 1672 16634 1728
rect 9586 1264 9642 1320
rect 9218 856 9274 912
rect 9126 448 9182 504
<< metal3 >>
rect 14000 12338 34000 12368
rect 2730 12278 34000 12338
rect 2405 12202 2471 12205
rect 2730 12202 2790 12278
rect 14000 12248 34000 12278
rect 2405 12200 2790 12202
rect 2405 12144 2410 12200
rect 2466 12144 2790 12200
rect 2405 12142 2790 12144
rect 2405 12139 2471 12142
rect 14000 11928 34000 11960
rect 14000 11872 16670 11928
rect 16726 11872 34000 11928
rect 14000 11840 34000 11872
rect 2865 11794 2931 11797
rect 8017 11794 8083 11797
rect 2865 11792 8083 11794
rect 2865 11736 2870 11792
rect 2926 11736 8022 11792
rect 8078 11736 8083 11792
rect 2865 11734 8083 11736
rect 2865 11731 2931 11734
rect 8017 11731 8083 11734
rect 1669 11658 1735 11661
rect 5165 11658 5231 11661
rect 1669 11656 5231 11658
rect 1669 11600 1674 11656
rect 1730 11600 5170 11656
rect 5226 11600 5231 11656
rect 1669 11598 5231 11600
rect 1669 11595 1735 11598
rect 5165 11595 5231 11598
rect 13721 11522 13787 11525
rect 14000 11522 34000 11552
rect 13721 11520 34000 11522
rect 13721 11464 13726 11520
rect 13782 11464 34000 11520
rect 13721 11462 34000 11464
rect 13721 11459 13787 11462
rect 2560 11456 2880 11457
rect 2560 11392 2568 11456
rect 2632 11392 2648 11456
rect 2712 11392 2728 11456
rect 2792 11392 2808 11456
rect 2872 11392 2880 11456
rect 2560 11391 2880 11392
rect 5660 11456 5980 11457
rect 5660 11392 5668 11456
rect 5732 11392 5748 11456
rect 5812 11392 5828 11456
rect 5892 11392 5908 11456
rect 5972 11392 5980 11456
rect 5660 11391 5980 11392
rect 8760 11456 9080 11457
rect 8760 11392 8768 11456
rect 8832 11392 8848 11456
rect 8912 11392 8928 11456
rect 8992 11392 9008 11456
rect 9072 11392 9080 11456
rect 14000 11432 34000 11462
rect 8760 11391 9080 11392
rect 3509 11386 3575 11389
rect 5533 11386 5599 11389
rect 3509 11384 5599 11386
rect 3509 11328 3514 11384
rect 3570 11328 5538 11384
rect 5594 11328 5599 11384
rect 3509 11326 5599 11328
rect 3509 11323 3575 11326
rect 5533 11323 5599 11326
rect 6637 11386 6703 11389
rect 8201 11386 8267 11389
rect 6637 11384 8267 11386
rect 6637 11328 6642 11384
rect 6698 11328 8206 11384
rect 8262 11328 8267 11384
rect 6637 11326 8267 11328
rect 6637 11323 6703 11326
rect 8201 11323 8267 11326
rect 2589 11250 2655 11253
rect 5441 11250 5507 11253
rect 2589 11248 5507 11250
rect 2589 11192 2594 11248
rect 2650 11192 5446 11248
rect 5502 11192 5507 11248
rect 2589 11190 5507 11192
rect 2589 11187 2655 11190
rect 5441 11187 5507 11190
rect 2037 11114 2103 11117
rect 2405 11114 2471 11117
rect 5073 11114 5139 11117
rect 2037 11112 2471 11114
rect 2037 11056 2042 11112
rect 2098 11056 2410 11112
rect 2466 11056 2471 11112
rect 2037 11054 2471 11056
rect 2037 11051 2103 11054
rect 2405 11051 2471 11054
rect 2730 11112 5139 11114
rect 2730 11056 5078 11112
rect 5134 11056 5139 11112
rect 2730 11054 5139 11056
rect 1393 10978 1459 10981
rect 2730 10978 2790 11054
rect 5073 11051 5139 11054
rect 5257 11114 5323 11117
rect 5993 11114 6059 11117
rect 5257 11112 6059 11114
rect 5257 11056 5262 11112
rect 5318 11056 5998 11112
rect 6054 11056 6059 11112
rect 5257 11054 6059 11056
rect 5257 11051 5323 11054
rect 5993 11051 6059 11054
rect 13813 11114 13879 11117
rect 14000 11114 34000 11144
rect 13813 11112 34000 11114
rect 13813 11056 13818 11112
rect 13874 11056 34000 11112
rect 13813 11054 34000 11056
rect 13813 11051 13879 11054
rect 14000 11024 34000 11054
rect 1393 10976 2790 10978
rect 1393 10920 1398 10976
rect 1454 10920 2790 10976
rect 1393 10918 2790 10920
rect 1393 10915 1459 10918
rect 4110 10912 4430 10913
rect 4110 10848 4118 10912
rect 4182 10848 4198 10912
rect 4262 10848 4278 10912
rect 4342 10848 4358 10912
rect 4422 10848 4430 10912
rect 4110 10847 4430 10848
rect 7210 10912 7530 10913
rect 7210 10848 7218 10912
rect 7282 10848 7298 10912
rect 7362 10848 7378 10912
rect 7442 10848 7458 10912
rect 7522 10848 7530 10912
rect 7210 10847 7530 10848
rect 2773 10842 2839 10845
rect 3509 10842 3575 10845
rect 2773 10840 3575 10842
rect 2773 10784 2778 10840
rect 2834 10784 3514 10840
rect 3570 10784 3575 10840
rect 2773 10782 3575 10784
rect 2773 10779 2839 10782
rect 3509 10779 3575 10782
rect 2129 10706 2195 10709
rect 4521 10706 4587 10709
rect 14000 10706 34000 10736
rect 2129 10704 4587 10706
rect 2129 10648 2134 10704
rect 2190 10648 4526 10704
rect 4582 10648 4587 10704
rect 2129 10646 4587 10648
rect 2129 10643 2195 10646
rect 4521 10643 4587 10646
rect 12390 10646 34000 10706
rect 2129 10570 2195 10573
rect 7465 10570 7531 10573
rect 12390 10570 12450 10646
rect 14000 10616 34000 10646
rect 2129 10568 7531 10570
rect 2129 10512 2134 10568
rect 2190 10512 7470 10568
rect 7526 10512 7531 10568
rect 2129 10510 7531 10512
rect 2129 10507 2195 10510
rect 7465 10507 7531 10510
rect 7606 10510 12450 10570
rect 3049 10434 3115 10437
rect 4153 10434 4219 10437
rect 3049 10432 4219 10434
rect 3049 10376 3054 10432
rect 3110 10376 4158 10432
rect 4214 10376 4219 10432
rect 3049 10374 4219 10376
rect 3049 10371 3115 10374
rect 4153 10371 4219 10374
rect 2560 10368 2880 10369
rect 2560 10304 2568 10368
rect 2632 10304 2648 10368
rect 2712 10304 2728 10368
rect 2792 10304 2808 10368
rect 2872 10304 2880 10368
rect 2560 10303 2880 10304
rect 5660 10368 5980 10369
rect 5660 10304 5668 10368
rect 5732 10304 5748 10368
rect 5812 10304 5828 10368
rect 5892 10304 5908 10368
rect 5972 10304 5980 10368
rect 5660 10303 5980 10304
rect 2957 10298 3023 10301
rect 3877 10298 3943 10301
rect 2957 10296 3943 10298
rect 2957 10240 2962 10296
rect 3018 10240 3882 10296
rect 3938 10240 3943 10296
rect 2957 10238 3943 10240
rect 2957 10235 3023 10238
rect 3877 10235 3943 10238
rect 1209 10162 1275 10165
rect 7606 10162 7666 10510
rect 8760 10368 9080 10369
rect 8760 10304 8768 10368
rect 8832 10304 8848 10368
rect 8912 10304 8928 10368
rect 8992 10304 9008 10368
rect 9072 10304 9080 10368
rect 8760 10303 9080 10304
rect 9397 10298 9463 10301
rect 14000 10298 34000 10328
rect 9397 10296 34000 10298
rect 9397 10240 9402 10296
rect 9458 10240 34000 10296
rect 9397 10238 34000 10240
rect 9397 10235 9463 10238
rect 14000 10208 34000 10238
rect 1209 10160 7666 10162
rect 1209 10104 1214 10160
rect 1270 10104 7666 10160
rect 1209 10102 7666 10104
rect 1209 10099 1275 10102
rect 1393 10026 1459 10029
rect 1945 10026 2011 10029
rect 1393 10024 12450 10026
rect 1393 9968 1398 10024
rect 1454 9968 1950 10024
rect 2006 9968 12450 10024
rect 1393 9966 12450 9968
rect 1393 9963 1459 9966
rect 1945 9963 2011 9966
rect 1393 9890 1459 9893
rect 2313 9890 2379 9893
rect 1393 9888 2379 9890
rect 1393 9832 1398 9888
rect 1454 9832 2318 9888
rect 2374 9832 2379 9888
rect 1393 9830 2379 9832
rect 12390 9890 12450 9966
rect 14000 9890 34000 9920
rect 12390 9830 34000 9890
rect 1393 9827 1459 9830
rect 2313 9827 2379 9830
rect 4110 9824 4430 9825
rect 4110 9760 4118 9824
rect 4182 9760 4198 9824
rect 4262 9760 4278 9824
rect 4342 9760 4358 9824
rect 4422 9760 4430 9824
rect 4110 9759 4430 9760
rect 7210 9824 7530 9825
rect 7210 9760 7218 9824
rect 7282 9760 7298 9824
rect 7362 9760 7378 9824
rect 7442 9760 7458 9824
rect 7522 9760 7530 9824
rect 14000 9800 34000 9830
rect 7210 9759 7530 9760
rect 1761 9618 1827 9621
rect 2589 9618 2655 9621
rect 5993 9618 6059 9621
rect 9213 9618 9279 9621
rect 1761 9616 6059 9618
rect 1761 9560 1766 9616
rect 1822 9560 2594 9616
rect 2650 9560 5998 9616
rect 6054 9560 6059 9616
rect 1761 9558 6059 9560
rect 1761 9555 1827 9558
rect 2589 9555 2655 9558
rect 5993 9555 6059 9558
rect 6502 9616 9279 9618
rect 6502 9560 9218 9616
rect 9274 9560 9279 9616
rect 6502 9558 9279 9560
rect 1301 9482 1367 9485
rect 2037 9482 2103 9485
rect 1301 9480 2103 9482
rect 1301 9424 1306 9480
rect 1362 9424 2042 9480
rect 2098 9424 2103 9480
rect 1301 9422 2103 9424
rect 1301 9419 1367 9422
rect 2037 9419 2103 9422
rect 2313 9482 2379 9485
rect 2957 9482 3023 9485
rect 3325 9482 3391 9485
rect 2313 9480 3391 9482
rect 2313 9424 2318 9480
rect 2374 9424 2962 9480
rect 3018 9424 3330 9480
rect 3386 9424 3391 9480
rect 2313 9422 3391 9424
rect 2313 9419 2379 9422
rect 2957 9419 3023 9422
rect 3325 9419 3391 9422
rect 2560 9280 2880 9281
rect 2560 9216 2568 9280
rect 2632 9216 2648 9280
rect 2712 9216 2728 9280
rect 2792 9216 2808 9280
rect 2872 9216 2880 9280
rect 2560 9215 2880 9216
rect 5660 9280 5980 9281
rect 5660 9216 5668 9280
rect 5732 9216 5748 9280
rect 5812 9216 5828 9280
rect 5892 9216 5908 9280
rect 5972 9216 5980 9280
rect 5660 9215 5980 9216
rect 1209 9074 1275 9077
rect 1577 9074 1643 9077
rect 1209 9072 1643 9074
rect 1209 9016 1214 9072
rect 1270 9016 1582 9072
rect 1638 9016 1643 9072
rect 1209 9014 1643 9016
rect 1209 9011 1275 9014
rect 1577 9011 1643 9014
rect 2129 9074 2195 9077
rect 6502 9074 6562 9558
rect 9213 9555 9279 9558
rect 8201 9482 8267 9485
rect 14000 9482 34000 9512
rect 8201 9480 34000 9482
rect 8201 9424 8206 9480
rect 8262 9424 34000 9480
rect 8201 9422 34000 9424
rect 8201 9419 8267 9422
rect 14000 9392 34000 9422
rect 8760 9280 9080 9281
rect 8760 9216 8768 9280
rect 8832 9216 8848 9280
rect 8912 9216 8928 9280
rect 8992 9216 9008 9280
rect 9072 9216 9080 9280
rect 8760 9215 9080 9216
rect 9213 9210 9279 9213
rect 13813 9210 13879 9213
rect 9213 9208 13879 9210
rect 9213 9152 9218 9208
rect 9274 9152 13818 9208
rect 13874 9152 13879 9208
rect 9213 9150 13879 9152
rect 9213 9147 9279 9150
rect 13813 9147 13879 9150
rect 2129 9072 6562 9074
rect 2129 9016 2134 9072
rect 2190 9016 6562 9072
rect 2129 9014 6562 9016
rect 6729 9074 6795 9077
rect 14000 9074 34000 9104
rect 6729 9072 34000 9074
rect 6729 9016 6734 9072
rect 6790 9016 34000 9072
rect 6729 9014 34000 9016
rect 2129 9011 2195 9014
rect 6729 9011 6795 9014
rect 14000 8984 34000 9014
rect 2037 8938 2103 8941
rect 3417 8938 3483 8941
rect 4337 8938 4403 8941
rect 5533 8938 5599 8941
rect 2037 8936 3483 8938
rect 2037 8880 2042 8936
rect 2098 8880 3422 8936
rect 3478 8880 3483 8936
rect 2037 8878 3483 8880
rect 2037 8875 2103 8878
rect 3417 8875 3483 8878
rect 3788 8936 5599 8938
rect 3788 8880 4342 8936
rect 4398 8880 5538 8936
rect 5594 8880 5599 8936
rect 3788 8878 5599 8880
rect 3788 8805 3848 8878
rect 4337 8875 4403 8878
rect 5533 8875 5599 8878
rect 3785 8800 3851 8805
rect 3785 8744 3790 8800
rect 3846 8744 3851 8800
rect 3785 8739 3851 8744
rect 4110 8736 4430 8737
rect 4110 8672 4118 8736
rect 4182 8672 4198 8736
rect 4262 8672 4278 8736
rect 4342 8672 4358 8736
rect 4422 8672 4430 8736
rect 4110 8671 4430 8672
rect 7210 8736 7530 8737
rect 7210 8672 7218 8736
rect 7282 8672 7298 8736
rect 7362 8672 7378 8736
rect 7442 8672 7458 8736
rect 7522 8672 7530 8736
rect 7210 8671 7530 8672
rect 14000 8664 34000 8696
rect 14000 8608 16578 8664
rect 16634 8608 34000 8664
rect 14000 8576 34000 8608
rect 3509 8530 3575 8533
rect 5717 8530 5783 8533
rect 3509 8528 5783 8530
rect 3509 8472 3514 8528
rect 3570 8472 5722 8528
rect 5778 8472 5783 8528
rect 3509 8470 5783 8472
rect 3509 8467 3575 8470
rect 5717 8467 5783 8470
rect 1945 8394 2011 8397
rect 8201 8394 8267 8397
rect 1945 8392 8267 8394
rect 1945 8336 1950 8392
rect 2006 8336 8206 8392
rect 8262 8336 8267 8392
rect 1945 8334 8267 8336
rect 1945 8331 2011 8334
rect 8201 8331 8267 8334
rect 9305 8258 9371 8261
rect 14000 8258 34000 8288
rect 9305 8256 34000 8258
rect 9305 8200 9310 8256
rect 9366 8200 34000 8256
rect 9305 8198 34000 8200
rect 9305 8195 9371 8198
rect 2560 8192 2880 8193
rect 2560 8128 2568 8192
rect 2632 8128 2648 8192
rect 2712 8128 2728 8192
rect 2792 8128 2808 8192
rect 2872 8128 2880 8192
rect 2560 8127 2880 8128
rect 5660 8192 5980 8193
rect 5660 8128 5668 8192
rect 5732 8128 5748 8192
rect 5812 8128 5828 8192
rect 5892 8128 5908 8192
rect 5972 8128 5980 8192
rect 5660 8127 5980 8128
rect 8760 8192 9080 8193
rect 8760 8128 8768 8192
rect 8832 8128 8848 8192
rect 8912 8128 8928 8192
rect 8992 8128 9008 8192
rect 9072 8128 9080 8192
rect 14000 8168 34000 8198
rect 8760 8127 9080 8128
rect 3049 8122 3115 8125
rect 3417 8122 3483 8125
rect 3785 8122 3851 8125
rect 4061 8122 4127 8125
rect 3049 8120 3483 8122
rect 3049 8064 3054 8120
rect 3110 8064 3422 8120
rect 3478 8064 3483 8120
rect 3049 8062 3483 8064
rect 3049 8059 3115 8062
rect 3417 8059 3483 8062
rect 3558 8120 4127 8122
rect 3558 8064 3790 8120
rect 3846 8064 4066 8120
rect 4122 8064 4127 8120
rect 3558 8062 4127 8064
rect 2681 7986 2747 7989
rect 3049 7986 3115 7989
rect 3558 7986 3618 8062
rect 3785 8059 3851 8062
rect 4061 8059 4127 8062
rect 2681 7984 3618 7986
rect 2681 7928 2686 7984
rect 2742 7928 3054 7984
rect 3110 7928 3618 7984
rect 2681 7926 3618 7928
rect 6361 7986 6427 7989
rect 9029 7986 9095 7989
rect 6361 7984 9095 7986
rect 6361 7928 6366 7984
rect 6422 7928 9034 7984
rect 9090 7928 9095 7984
rect 6361 7926 9095 7928
rect 2681 7923 2747 7926
rect 3049 7923 3115 7926
rect 6361 7923 6427 7926
rect 9029 7923 9095 7926
rect 10869 7850 10935 7853
rect 14000 7850 34000 7880
rect 10869 7848 34000 7850
rect 10869 7792 10874 7848
rect 10930 7792 34000 7848
rect 10869 7790 34000 7792
rect 10869 7787 10935 7790
rect 14000 7760 34000 7790
rect 4110 7648 4430 7649
rect 4110 7584 4118 7648
rect 4182 7584 4198 7648
rect 4262 7584 4278 7648
rect 4342 7584 4358 7648
rect 4422 7584 4430 7648
rect 4110 7583 4430 7584
rect 7210 7648 7530 7649
rect 7210 7584 7218 7648
rect 7282 7584 7298 7648
rect 7362 7584 7378 7648
rect 7442 7584 7458 7648
rect 7522 7584 7530 7648
rect 7210 7583 7530 7584
rect 1669 7578 1735 7581
rect 2773 7578 2839 7581
rect 1669 7576 2839 7578
rect 1669 7520 1674 7576
rect 1730 7520 2778 7576
rect 2834 7520 2839 7576
rect 1669 7518 2839 7520
rect 1669 7515 1735 7518
rect 2773 7515 2839 7518
rect 5073 7442 5139 7445
rect 14000 7442 34000 7472
rect 5073 7440 34000 7442
rect 5073 7384 5078 7440
rect 5134 7384 34000 7440
rect 5073 7382 34000 7384
rect 5073 7379 5139 7382
rect 14000 7352 34000 7382
rect 2405 7306 2471 7309
rect 2957 7306 3023 7309
rect 2405 7304 3023 7306
rect 2405 7248 2410 7304
rect 2466 7248 2962 7304
rect 3018 7248 3023 7304
rect 2405 7246 3023 7248
rect 2405 7243 2471 7246
rect 2957 7243 3023 7246
rect 2560 7104 2880 7105
rect 2560 7040 2568 7104
rect 2632 7040 2648 7104
rect 2712 7040 2728 7104
rect 2792 7040 2808 7104
rect 2872 7040 2880 7104
rect 2560 7039 2880 7040
rect 5660 7104 5980 7105
rect 5660 7040 5668 7104
rect 5732 7040 5748 7104
rect 5812 7040 5828 7104
rect 5892 7040 5908 7104
rect 5972 7040 5980 7104
rect 5660 7039 5980 7040
rect 8760 7104 9080 7105
rect 8760 7040 8768 7104
rect 8832 7040 8848 7104
rect 8912 7040 8928 7104
rect 8992 7040 9008 7104
rect 9072 7040 9080 7104
rect 8760 7039 9080 7040
rect 9397 7034 9463 7037
rect 14000 7034 34000 7064
rect 9397 7032 34000 7034
rect 9397 6976 9402 7032
rect 9458 6976 34000 7032
rect 9397 6974 34000 6976
rect 9397 6971 9463 6974
rect 14000 6944 34000 6974
rect 8385 6626 8451 6629
rect 14000 6626 34000 6656
rect 8385 6624 34000 6626
rect 8385 6568 8390 6624
rect 8446 6568 34000 6624
rect 8385 6566 34000 6568
rect 8385 6563 8451 6566
rect 4110 6560 4430 6561
rect 4110 6496 4118 6560
rect 4182 6496 4198 6560
rect 4262 6496 4278 6560
rect 4342 6496 4358 6560
rect 4422 6496 4430 6560
rect 4110 6495 4430 6496
rect 7210 6560 7530 6561
rect 7210 6496 7218 6560
rect 7282 6496 7298 6560
rect 7362 6496 7378 6560
rect 7442 6496 7458 6560
rect 7522 6496 7530 6560
rect 14000 6536 34000 6566
rect 7210 6495 7530 6496
rect 11053 6218 11119 6221
rect 14000 6218 34000 6248
rect 11053 6216 34000 6218
rect 11053 6160 11058 6216
rect 11114 6160 34000 6216
rect 11053 6158 34000 6160
rect 11053 6155 11119 6158
rect 14000 6128 34000 6158
rect 2560 6016 2880 6017
rect 2560 5952 2568 6016
rect 2632 5952 2648 6016
rect 2712 5952 2728 6016
rect 2792 5952 2808 6016
rect 2872 5952 2880 6016
rect 2560 5951 2880 5952
rect 5660 6016 5980 6017
rect 5660 5952 5668 6016
rect 5732 5952 5748 6016
rect 5812 5952 5828 6016
rect 5892 5952 5908 6016
rect 5972 5952 5980 6016
rect 5660 5951 5980 5952
rect 8760 6016 9080 6017
rect 8760 5952 8768 6016
rect 8832 5952 8848 6016
rect 8912 5952 8928 6016
rect 8992 5952 9008 6016
rect 9072 5952 9080 6016
rect 8760 5951 9080 5952
rect 8109 5810 8175 5813
rect 14000 5810 34000 5840
rect 8109 5808 34000 5810
rect 8109 5752 8114 5808
rect 8170 5752 34000 5808
rect 8109 5750 34000 5752
rect 8109 5747 8175 5750
rect 14000 5720 34000 5750
rect 4110 5472 4430 5473
rect 4110 5408 4118 5472
rect 4182 5408 4198 5472
rect 4262 5408 4278 5472
rect 4342 5408 4358 5472
rect 4422 5408 4430 5472
rect 4110 5407 4430 5408
rect 7210 5472 7530 5473
rect 7210 5408 7218 5472
rect 7282 5408 7298 5472
rect 7362 5408 7378 5472
rect 7442 5408 7458 5472
rect 7522 5408 7530 5472
rect 7210 5407 7530 5408
rect 12249 5402 12315 5405
rect 14000 5402 34000 5432
rect 12249 5400 34000 5402
rect 12249 5344 12254 5400
rect 12310 5344 34000 5400
rect 12249 5342 34000 5344
rect 12249 5339 12315 5342
rect 14000 5312 34000 5342
rect 9397 4994 9463 4997
rect 14000 4994 34000 5024
rect 9397 4992 34000 4994
rect 9397 4936 9402 4992
rect 9458 4936 34000 4992
rect 9397 4934 34000 4936
rect 9397 4931 9463 4934
rect 5660 4928 5980 4929
rect 5660 4864 5668 4928
rect 5732 4864 5748 4928
rect 5812 4864 5828 4928
rect 5892 4864 5908 4928
rect 5972 4864 5980 4928
rect 5660 4863 5980 4864
rect 8760 4928 9080 4929
rect 8760 4864 8768 4928
rect 8832 4864 8848 4928
rect 8912 4864 8928 4928
rect 8992 4864 9008 4928
rect 9072 4864 9080 4928
rect 14000 4904 34000 4934
rect 8760 4863 9080 4864
rect 3693 4586 3759 4589
rect 5717 4586 5783 4589
rect 3693 4584 5783 4586
rect 3693 4528 3698 4584
rect 3754 4528 5722 4584
rect 5778 4528 5783 4584
rect 3693 4526 5783 4528
rect 3693 4523 3759 4526
rect 5717 4523 5783 4526
rect 7925 4586 7991 4589
rect 14000 4586 34000 4616
rect 7925 4584 34000 4586
rect 7925 4528 7930 4584
rect 7986 4528 34000 4584
rect 7925 4526 34000 4528
rect 7925 4523 7991 4526
rect 14000 4496 34000 4526
rect 4110 4384 4430 4385
rect 4110 4320 4118 4384
rect 4182 4320 4198 4384
rect 4262 4320 4278 4384
rect 4342 4320 4358 4384
rect 4422 4320 4430 4384
rect 4110 4319 4430 4320
rect 7210 4384 7530 4385
rect 7210 4320 7218 4384
rect 7282 4320 7298 4384
rect 7362 4320 7378 4384
rect 7442 4320 7458 4384
rect 7522 4320 7530 4384
rect 7210 4319 7530 4320
rect 14000 4176 34000 4208
rect 14000 4120 16578 4176
rect 16634 4120 34000 4176
rect 14000 4088 34000 4120
rect 5660 3840 5980 3841
rect 5660 3776 5668 3840
rect 5732 3776 5748 3840
rect 5812 3776 5828 3840
rect 5892 3776 5908 3840
rect 5972 3776 5980 3840
rect 5660 3775 5980 3776
rect 8760 3840 9080 3841
rect 8760 3776 8768 3840
rect 8832 3776 8848 3840
rect 8912 3776 8928 3840
rect 8992 3776 9008 3840
rect 9072 3776 9080 3840
rect 8760 3775 9080 3776
rect 14000 3768 34000 3800
rect 14000 3712 16578 3768
rect 16634 3712 34000 3768
rect 14000 3680 34000 3712
rect 2681 3362 2747 3365
rect 2484 3360 2747 3362
rect 2484 3304 2686 3360
rect 2742 3304 2747 3360
rect 2484 3302 2747 3304
rect 2681 3299 2747 3302
rect 9489 3362 9555 3365
rect 14000 3362 34000 3392
rect 9489 3360 34000 3362
rect 9489 3304 9494 3360
rect 9550 3304 34000 3360
rect 9489 3302 34000 3304
rect 9489 3299 9555 3302
rect 4110 3296 4430 3297
rect 4110 3232 4118 3296
rect 4182 3232 4198 3296
rect 4262 3232 4278 3296
rect 4342 3232 4358 3296
rect 4422 3232 4430 3296
rect 4110 3231 4430 3232
rect 7210 3296 7530 3297
rect 7210 3232 7218 3296
rect 7282 3232 7298 3296
rect 7362 3232 7378 3296
rect 7442 3232 7458 3296
rect 7522 3232 7530 3296
rect 14000 3272 34000 3302
rect 7210 3231 7530 3232
rect 14000 2952 34000 2984
rect 14000 2896 16578 2952
rect 16634 2896 34000 2952
rect 14000 2864 34000 2896
rect 5660 2752 5980 2753
rect 5660 2688 5668 2752
rect 5732 2688 5748 2752
rect 5812 2688 5828 2752
rect 5892 2688 5908 2752
rect 5972 2688 5980 2752
rect 5660 2687 5980 2688
rect 8760 2752 9080 2753
rect 8760 2688 8768 2752
rect 8832 2688 8848 2752
rect 8912 2688 8928 2752
rect 8992 2688 9008 2752
rect 9072 2688 9080 2752
rect 8760 2687 9080 2688
rect 9397 2546 9463 2549
rect 14000 2546 34000 2576
rect 9397 2544 34000 2546
rect 9397 2488 9402 2544
rect 9458 2488 34000 2544
rect 9397 2486 34000 2488
rect 9397 2483 9463 2486
rect 14000 2456 34000 2486
rect 4110 2208 4430 2209
rect 4110 2144 4118 2208
rect 4182 2144 4198 2208
rect 4262 2144 4278 2208
rect 4342 2144 4358 2208
rect 4422 2144 4430 2208
rect 4110 2143 4430 2144
rect 7210 2208 7530 2209
rect 7210 2144 7218 2208
rect 7282 2144 7298 2208
rect 7362 2144 7378 2208
rect 7442 2144 7458 2208
rect 7522 2144 7530 2208
rect 7210 2143 7530 2144
rect 14000 2136 34000 2168
rect 14000 2080 16578 2136
rect 16634 2080 34000 2136
rect 14000 2048 34000 2080
rect 14000 1728 34000 1760
rect 14000 1672 16578 1728
rect 16634 1672 34000 1728
rect 5660 1664 5980 1665
rect 5660 1600 5668 1664
rect 5732 1600 5748 1664
rect 5812 1600 5828 1664
rect 5892 1600 5908 1664
rect 5972 1600 5980 1664
rect 5660 1599 5980 1600
rect 8760 1664 9080 1665
rect 8760 1600 8768 1664
rect 8832 1600 8848 1664
rect 8912 1600 8928 1664
rect 8992 1600 9008 1664
rect 9072 1600 9080 1664
rect 14000 1640 34000 1672
rect 8760 1599 9080 1600
rect 9581 1322 9647 1325
rect 14000 1322 34000 1352
rect 9581 1320 34000 1322
rect 9581 1264 9586 1320
rect 9642 1264 34000 1320
rect 9581 1262 34000 1264
rect 9581 1259 9647 1262
rect 14000 1232 34000 1262
rect 4110 1120 4430 1121
rect 4110 1056 4118 1120
rect 4182 1056 4198 1120
rect 4262 1056 4278 1120
rect 4342 1056 4358 1120
rect 4422 1056 4430 1120
rect 4110 1055 4430 1056
rect 7210 1120 7530 1121
rect 7210 1056 7218 1120
rect 7282 1056 7298 1120
rect 7362 1056 7378 1120
rect 7442 1056 7458 1120
rect 7522 1056 7530 1120
rect 7210 1055 7530 1056
rect 9213 914 9279 917
rect 14000 914 34000 944
rect 9213 912 34000 914
rect 9213 856 9218 912
rect 9274 856 34000 912
rect 9213 854 34000 856
rect 9213 851 9279 854
rect 14000 824 34000 854
rect 9121 506 9187 509
rect 14000 506 34000 536
rect 9121 504 34000 506
rect 9121 448 9126 504
rect 9182 448 34000 504
rect 9121 446 34000 448
rect 9121 443 9187 446
rect 14000 416 34000 446
<< via3 >>
rect 2568 11452 2632 11456
rect 2568 11396 2572 11452
rect 2572 11396 2628 11452
rect 2628 11396 2632 11452
rect 2568 11392 2632 11396
rect 2648 11452 2712 11456
rect 2648 11396 2652 11452
rect 2652 11396 2708 11452
rect 2708 11396 2712 11452
rect 2648 11392 2712 11396
rect 2728 11452 2792 11456
rect 2728 11396 2732 11452
rect 2732 11396 2788 11452
rect 2788 11396 2792 11452
rect 2728 11392 2792 11396
rect 2808 11452 2872 11456
rect 2808 11396 2812 11452
rect 2812 11396 2868 11452
rect 2868 11396 2872 11452
rect 2808 11392 2872 11396
rect 5668 11452 5732 11456
rect 5668 11396 5672 11452
rect 5672 11396 5728 11452
rect 5728 11396 5732 11452
rect 5668 11392 5732 11396
rect 5748 11452 5812 11456
rect 5748 11396 5752 11452
rect 5752 11396 5808 11452
rect 5808 11396 5812 11452
rect 5748 11392 5812 11396
rect 5828 11452 5892 11456
rect 5828 11396 5832 11452
rect 5832 11396 5888 11452
rect 5888 11396 5892 11452
rect 5828 11392 5892 11396
rect 5908 11452 5972 11456
rect 5908 11396 5912 11452
rect 5912 11396 5968 11452
rect 5968 11396 5972 11452
rect 5908 11392 5972 11396
rect 8768 11452 8832 11456
rect 8768 11396 8772 11452
rect 8772 11396 8828 11452
rect 8828 11396 8832 11452
rect 8768 11392 8832 11396
rect 8848 11452 8912 11456
rect 8848 11396 8852 11452
rect 8852 11396 8908 11452
rect 8908 11396 8912 11452
rect 8848 11392 8912 11396
rect 8928 11452 8992 11456
rect 8928 11396 8932 11452
rect 8932 11396 8988 11452
rect 8988 11396 8992 11452
rect 8928 11392 8992 11396
rect 9008 11452 9072 11456
rect 9008 11396 9012 11452
rect 9012 11396 9068 11452
rect 9068 11396 9072 11452
rect 9008 11392 9072 11396
rect 4118 10908 4182 10912
rect 4118 10852 4122 10908
rect 4122 10852 4178 10908
rect 4178 10852 4182 10908
rect 4118 10848 4182 10852
rect 4198 10908 4262 10912
rect 4198 10852 4202 10908
rect 4202 10852 4258 10908
rect 4258 10852 4262 10908
rect 4198 10848 4262 10852
rect 4278 10908 4342 10912
rect 4278 10852 4282 10908
rect 4282 10852 4338 10908
rect 4338 10852 4342 10908
rect 4278 10848 4342 10852
rect 4358 10908 4422 10912
rect 4358 10852 4362 10908
rect 4362 10852 4418 10908
rect 4418 10852 4422 10908
rect 4358 10848 4422 10852
rect 7218 10908 7282 10912
rect 7218 10852 7222 10908
rect 7222 10852 7278 10908
rect 7278 10852 7282 10908
rect 7218 10848 7282 10852
rect 7298 10908 7362 10912
rect 7298 10852 7302 10908
rect 7302 10852 7358 10908
rect 7358 10852 7362 10908
rect 7298 10848 7362 10852
rect 7378 10908 7442 10912
rect 7378 10852 7382 10908
rect 7382 10852 7438 10908
rect 7438 10852 7442 10908
rect 7378 10848 7442 10852
rect 7458 10908 7522 10912
rect 7458 10852 7462 10908
rect 7462 10852 7518 10908
rect 7518 10852 7522 10908
rect 7458 10848 7522 10852
rect 2568 10364 2632 10368
rect 2568 10308 2572 10364
rect 2572 10308 2628 10364
rect 2628 10308 2632 10364
rect 2568 10304 2632 10308
rect 2648 10364 2712 10368
rect 2648 10308 2652 10364
rect 2652 10308 2708 10364
rect 2708 10308 2712 10364
rect 2648 10304 2712 10308
rect 2728 10364 2792 10368
rect 2728 10308 2732 10364
rect 2732 10308 2788 10364
rect 2788 10308 2792 10364
rect 2728 10304 2792 10308
rect 2808 10364 2872 10368
rect 2808 10308 2812 10364
rect 2812 10308 2868 10364
rect 2868 10308 2872 10364
rect 2808 10304 2872 10308
rect 5668 10364 5732 10368
rect 5668 10308 5672 10364
rect 5672 10308 5728 10364
rect 5728 10308 5732 10364
rect 5668 10304 5732 10308
rect 5748 10364 5812 10368
rect 5748 10308 5752 10364
rect 5752 10308 5808 10364
rect 5808 10308 5812 10364
rect 5748 10304 5812 10308
rect 5828 10364 5892 10368
rect 5828 10308 5832 10364
rect 5832 10308 5888 10364
rect 5888 10308 5892 10364
rect 5828 10304 5892 10308
rect 5908 10364 5972 10368
rect 5908 10308 5912 10364
rect 5912 10308 5968 10364
rect 5968 10308 5972 10364
rect 5908 10304 5972 10308
rect 8768 10364 8832 10368
rect 8768 10308 8772 10364
rect 8772 10308 8828 10364
rect 8828 10308 8832 10364
rect 8768 10304 8832 10308
rect 8848 10364 8912 10368
rect 8848 10308 8852 10364
rect 8852 10308 8908 10364
rect 8908 10308 8912 10364
rect 8848 10304 8912 10308
rect 8928 10364 8992 10368
rect 8928 10308 8932 10364
rect 8932 10308 8988 10364
rect 8988 10308 8992 10364
rect 8928 10304 8992 10308
rect 9008 10364 9072 10368
rect 9008 10308 9012 10364
rect 9012 10308 9068 10364
rect 9068 10308 9072 10364
rect 9008 10304 9072 10308
rect 4118 9820 4182 9824
rect 4118 9764 4122 9820
rect 4122 9764 4178 9820
rect 4178 9764 4182 9820
rect 4118 9760 4182 9764
rect 4198 9820 4262 9824
rect 4198 9764 4202 9820
rect 4202 9764 4258 9820
rect 4258 9764 4262 9820
rect 4198 9760 4262 9764
rect 4278 9820 4342 9824
rect 4278 9764 4282 9820
rect 4282 9764 4338 9820
rect 4338 9764 4342 9820
rect 4278 9760 4342 9764
rect 4358 9820 4422 9824
rect 4358 9764 4362 9820
rect 4362 9764 4418 9820
rect 4418 9764 4422 9820
rect 4358 9760 4422 9764
rect 7218 9820 7282 9824
rect 7218 9764 7222 9820
rect 7222 9764 7278 9820
rect 7278 9764 7282 9820
rect 7218 9760 7282 9764
rect 7298 9820 7362 9824
rect 7298 9764 7302 9820
rect 7302 9764 7358 9820
rect 7358 9764 7362 9820
rect 7298 9760 7362 9764
rect 7378 9820 7442 9824
rect 7378 9764 7382 9820
rect 7382 9764 7438 9820
rect 7438 9764 7442 9820
rect 7378 9760 7442 9764
rect 7458 9820 7522 9824
rect 7458 9764 7462 9820
rect 7462 9764 7518 9820
rect 7518 9764 7522 9820
rect 7458 9760 7522 9764
rect 2568 9276 2632 9280
rect 2568 9220 2572 9276
rect 2572 9220 2628 9276
rect 2628 9220 2632 9276
rect 2568 9216 2632 9220
rect 2648 9276 2712 9280
rect 2648 9220 2652 9276
rect 2652 9220 2708 9276
rect 2708 9220 2712 9276
rect 2648 9216 2712 9220
rect 2728 9276 2792 9280
rect 2728 9220 2732 9276
rect 2732 9220 2788 9276
rect 2788 9220 2792 9276
rect 2728 9216 2792 9220
rect 2808 9276 2872 9280
rect 2808 9220 2812 9276
rect 2812 9220 2868 9276
rect 2868 9220 2872 9276
rect 2808 9216 2872 9220
rect 5668 9276 5732 9280
rect 5668 9220 5672 9276
rect 5672 9220 5728 9276
rect 5728 9220 5732 9276
rect 5668 9216 5732 9220
rect 5748 9276 5812 9280
rect 5748 9220 5752 9276
rect 5752 9220 5808 9276
rect 5808 9220 5812 9276
rect 5748 9216 5812 9220
rect 5828 9276 5892 9280
rect 5828 9220 5832 9276
rect 5832 9220 5888 9276
rect 5888 9220 5892 9276
rect 5828 9216 5892 9220
rect 5908 9276 5972 9280
rect 5908 9220 5912 9276
rect 5912 9220 5968 9276
rect 5968 9220 5972 9276
rect 5908 9216 5972 9220
rect 8768 9276 8832 9280
rect 8768 9220 8772 9276
rect 8772 9220 8828 9276
rect 8828 9220 8832 9276
rect 8768 9216 8832 9220
rect 8848 9276 8912 9280
rect 8848 9220 8852 9276
rect 8852 9220 8908 9276
rect 8908 9220 8912 9276
rect 8848 9216 8912 9220
rect 8928 9276 8992 9280
rect 8928 9220 8932 9276
rect 8932 9220 8988 9276
rect 8988 9220 8992 9276
rect 8928 9216 8992 9220
rect 9008 9276 9072 9280
rect 9008 9220 9012 9276
rect 9012 9220 9068 9276
rect 9068 9220 9072 9276
rect 9008 9216 9072 9220
rect 4118 8732 4182 8736
rect 4118 8676 4122 8732
rect 4122 8676 4178 8732
rect 4178 8676 4182 8732
rect 4118 8672 4182 8676
rect 4198 8732 4262 8736
rect 4198 8676 4202 8732
rect 4202 8676 4258 8732
rect 4258 8676 4262 8732
rect 4198 8672 4262 8676
rect 4278 8732 4342 8736
rect 4278 8676 4282 8732
rect 4282 8676 4338 8732
rect 4338 8676 4342 8732
rect 4278 8672 4342 8676
rect 4358 8732 4422 8736
rect 4358 8676 4362 8732
rect 4362 8676 4418 8732
rect 4418 8676 4422 8732
rect 4358 8672 4422 8676
rect 7218 8732 7282 8736
rect 7218 8676 7222 8732
rect 7222 8676 7278 8732
rect 7278 8676 7282 8732
rect 7218 8672 7282 8676
rect 7298 8732 7362 8736
rect 7298 8676 7302 8732
rect 7302 8676 7358 8732
rect 7358 8676 7362 8732
rect 7298 8672 7362 8676
rect 7378 8732 7442 8736
rect 7378 8676 7382 8732
rect 7382 8676 7438 8732
rect 7438 8676 7442 8732
rect 7378 8672 7442 8676
rect 7458 8732 7522 8736
rect 7458 8676 7462 8732
rect 7462 8676 7518 8732
rect 7518 8676 7522 8732
rect 7458 8672 7522 8676
rect 2568 8188 2632 8192
rect 2568 8132 2572 8188
rect 2572 8132 2628 8188
rect 2628 8132 2632 8188
rect 2568 8128 2632 8132
rect 2648 8188 2712 8192
rect 2648 8132 2652 8188
rect 2652 8132 2708 8188
rect 2708 8132 2712 8188
rect 2648 8128 2712 8132
rect 2728 8188 2792 8192
rect 2728 8132 2732 8188
rect 2732 8132 2788 8188
rect 2788 8132 2792 8188
rect 2728 8128 2792 8132
rect 2808 8188 2872 8192
rect 2808 8132 2812 8188
rect 2812 8132 2868 8188
rect 2868 8132 2872 8188
rect 2808 8128 2872 8132
rect 5668 8188 5732 8192
rect 5668 8132 5672 8188
rect 5672 8132 5728 8188
rect 5728 8132 5732 8188
rect 5668 8128 5732 8132
rect 5748 8188 5812 8192
rect 5748 8132 5752 8188
rect 5752 8132 5808 8188
rect 5808 8132 5812 8188
rect 5748 8128 5812 8132
rect 5828 8188 5892 8192
rect 5828 8132 5832 8188
rect 5832 8132 5888 8188
rect 5888 8132 5892 8188
rect 5828 8128 5892 8132
rect 5908 8188 5972 8192
rect 5908 8132 5912 8188
rect 5912 8132 5968 8188
rect 5968 8132 5972 8188
rect 5908 8128 5972 8132
rect 8768 8188 8832 8192
rect 8768 8132 8772 8188
rect 8772 8132 8828 8188
rect 8828 8132 8832 8188
rect 8768 8128 8832 8132
rect 8848 8188 8912 8192
rect 8848 8132 8852 8188
rect 8852 8132 8908 8188
rect 8908 8132 8912 8188
rect 8848 8128 8912 8132
rect 8928 8188 8992 8192
rect 8928 8132 8932 8188
rect 8932 8132 8988 8188
rect 8988 8132 8992 8188
rect 8928 8128 8992 8132
rect 9008 8188 9072 8192
rect 9008 8132 9012 8188
rect 9012 8132 9068 8188
rect 9068 8132 9072 8188
rect 9008 8128 9072 8132
rect 4118 7644 4182 7648
rect 4118 7588 4122 7644
rect 4122 7588 4178 7644
rect 4178 7588 4182 7644
rect 4118 7584 4182 7588
rect 4198 7644 4262 7648
rect 4198 7588 4202 7644
rect 4202 7588 4258 7644
rect 4258 7588 4262 7644
rect 4198 7584 4262 7588
rect 4278 7644 4342 7648
rect 4278 7588 4282 7644
rect 4282 7588 4338 7644
rect 4338 7588 4342 7644
rect 4278 7584 4342 7588
rect 4358 7644 4422 7648
rect 4358 7588 4362 7644
rect 4362 7588 4418 7644
rect 4418 7588 4422 7644
rect 4358 7584 4422 7588
rect 7218 7644 7282 7648
rect 7218 7588 7222 7644
rect 7222 7588 7278 7644
rect 7278 7588 7282 7644
rect 7218 7584 7282 7588
rect 7298 7644 7362 7648
rect 7298 7588 7302 7644
rect 7302 7588 7358 7644
rect 7358 7588 7362 7644
rect 7298 7584 7362 7588
rect 7378 7644 7442 7648
rect 7378 7588 7382 7644
rect 7382 7588 7438 7644
rect 7438 7588 7442 7644
rect 7378 7584 7442 7588
rect 7458 7644 7522 7648
rect 7458 7588 7462 7644
rect 7462 7588 7518 7644
rect 7518 7588 7522 7644
rect 7458 7584 7522 7588
rect 2568 7100 2632 7104
rect 2568 7044 2572 7100
rect 2572 7044 2628 7100
rect 2628 7044 2632 7100
rect 2568 7040 2632 7044
rect 2648 7100 2712 7104
rect 2648 7044 2652 7100
rect 2652 7044 2708 7100
rect 2708 7044 2712 7100
rect 2648 7040 2712 7044
rect 2728 7100 2792 7104
rect 2728 7044 2732 7100
rect 2732 7044 2788 7100
rect 2788 7044 2792 7100
rect 2728 7040 2792 7044
rect 2808 7100 2872 7104
rect 2808 7044 2812 7100
rect 2812 7044 2868 7100
rect 2868 7044 2872 7100
rect 2808 7040 2872 7044
rect 5668 7100 5732 7104
rect 5668 7044 5672 7100
rect 5672 7044 5728 7100
rect 5728 7044 5732 7100
rect 5668 7040 5732 7044
rect 5748 7100 5812 7104
rect 5748 7044 5752 7100
rect 5752 7044 5808 7100
rect 5808 7044 5812 7100
rect 5748 7040 5812 7044
rect 5828 7100 5892 7104
rect 5828 7044 5832 7100
rect 5832 7044 5888 7100
rect 5888 7044 5892 7100
rect 5828 7040 5892 7044
rect 5908 7100 5972 7104
rect 5908 7044 5912 7100
rect 5912 7044 5968 7100
rect 5968 7044 5972 7100
rect 5908 7040 5972 7044
rect 8768 7100 8832 7104
rect 8768 7044 8772 7100
rect 8772 7044 8828 7100
rect 8828 7044 8832 7100
rect 8768 7040 8832 7044
rect 8848 7100 8912 7104
rect 8848 7044 8852 7100
rect 8852 7044 8908 7100
rect 8908 7044 8912 7100
rect 8848 7040 8912 7044
rect 8928 7100 8992 7104
rect 8928 7044 8932 7100
rect 8932 7044 8988 7100
rect 8988 7044 8992 7100
rect 8928 7040 8992 7044
rect 9008 7100 9072 7104
rect 9008 7044 9012 7100
rect 9012 7044 9068 7100
rect 9068 7044 9072 7100
rect 9008 7040 9072 7044
rect 4118 6556 4182 6560
rect 4118 6500 4122 6556
rect 4122 6500 4178 6556
rect 4178 6500 4182 6556
rect 4118 6496 4182 6500
rect 4198 6556 4262 6560
rect 4198 6500 4202 6556
rect 4202 6500 4258 6556
rect 4258 6500 4262 6556
rect 4198 6496 4262 6500
rect 4278 6556 4342 6560
rect 4278 6500 4282 6556
rect 4282 6500 4338 6556
rect 4338 6500 4342 6556
rect 4278 6496 4342 6500
rect 4358 6556 4422 6560
rect 4358 6500 4362 6556
rect 4362 6500 4418 6556
rect 4418 6500 4422 6556
rect 4358 6496 4422 6500
rect 7218 6556 7282 6560
rect 7218 6500 7222 6556
rect 7222 6500 7278 6556
rect 7278 6500 7282 6556
rect 7218 6496 7282 6500
rect 7298 6556 7362 6560
rect 7298 6500 7302 6556
rect 7302 6500 7358 6556
rect 7358 6500 7362 6556
rect 7298 6496 7362 6500
rect 7378 6556 7442 6560
rect 7378 6500 7382 6556
rect 7382 6500 7438 6556
rect 7438 6500 7442 6556
rect 7378 6496 7442 6500
rect 7458 6556 7522 6560
rect 7458 6500 7462 6556
rect 7462 6500 7518 6556
rect 7518 6500 7522 6556
rect 7458 6496 7522 6500
rect 2568 6012 2632 6016
rect 2568 5956 2572 6012
rect 2572 5956 2628 6012
rect 2628 5956 2632 6012
rect 2568 5952 2632 5956
rect 2648 6012 2712 6016
rect 2648 5956 2652 6012
rect 2652 5956 2708 6012
rect 2708 5956 2712 6012
rect 2648 5952 2712 5956
rect 2728 6012 2792 6016
rect 2728 5956 2732 6012
rect 2732 5956 2788 6012
rect 2788 5956 2792 6012
rect 2728 5952 2792 5956
rect 2808 6012 2872 6016
rect 2808 5956 2812 6012
rect 2812 5956 2868 6012
rect 2868 5956 2872 6012
rect 2808 5952 2872 5956
rect 5668 6012 5732 6016
rect 5668 5956 5672 6012
rect 5672 5956 5728 6012
rect 5728 5956 5732 6012
rect 5668 5952 5732 5956
rect 5748 6012 5812 6016
rect 5748 5956 5752 6012
rect 5752 5956 5808 6012
rect 5808 5956 5812 6012
rect 5748 5952 5812 5956
rect 5828 6012 5892 6016
rect 5828 5956 5832 6012
rect 5832 5956 5888 6012
rect 5888 5956 5892 6012
rect 5828 5952 5892 5956
rect 5908 6012 5972 6016
rect 5908 5956 5912 6012
rect 5912 5956 5968 6012
rect 5968 5956 5972 6012
rect 5908 5952 5972 5956
rect 8768 6012 8832 6016
rect 8768 5956 8772 6012
rect 8772 5956 8828 6012
rect 8828 5956 8832 6012
rect 8768 5952 8832 5956
rect 8848 6012 8912 6016
rect 8848 5956 8852 6012
rect 8852 5956 8908 6012
rect 8908 5956 8912 6012
rect 8848 5952 8912 5956
rect 8928 6012 8992 6016
rect 8928 5956 8932 6012
rect 8932 5956 8988 6012
rect 8988 5956 8992 6012
rect 8928 5952 8992 5956
rect 9008 6012 9072 6016
rect 9008 5956 9012 6012
rect 9012 5956 9068 6012
rect 9068 5956 9072 6012
rect 9008 5952 9072 5956
rect 4118 5468 4182 5472
rect 4118 5412 4122 5468
rect 4122 5412 4178 5468
rect 4178 5412 4182 5468
rect 4118 5408 4182 5412
rect 4198 5468 4262 5472
rect 4198 5412 4202 5468
rect 4202 5412 4258 5468
rect 4258 5412 4262 5468
rect 4198 5408 4262 5412
rect 4278 5468 4342 5472
rect 4278 5412 4282 5468
rect 4282 5412 4338 5468
rect 4338 5412 4342 5468
rect 4278 5408 4342 5412
rect 4358 5468 4422 5472
rect 4358 5412 4362 5468
rect 4362 5412 4418 5468
rect 4418 5412 4422 5468
rect 4358 5408 4422 5412
rect 7218 5468 7282 5472
rect 7218 5412 7222 5468
rect 7222 5412 7278 5468
rect 7278 5412 7282 5468
rect 7218 5408 7282 5412
rect 7298 5468 7362 5472
rect 7298 5412 7302 5468
rect 7302 5412 7358 5468
rect 7358 5412 7362 5468
rect 7298 5408 7362 5412
rect 7378 5468 7442 5472
rect 7378 5412 7382 5468
rect 7382 5412 7438 5468
rect 7438 5412 7442 5468
rect 7378 5408 7442 5412
rect 7458 5468 7522 5472
rect 7458 5412 7462 5468
rect 7462 5412 7518 5468
rect 7518 5412 7522 5468
rect 7458 5408 7522 5412
rect 5668 4924 5732 4928
rect 5668 4868 5672 4924
rect 5672 4868 5728 4924
rect 5728 4868 5732 4924
rect 5668 4864 5732 4868
rect 5748 4924 5812 4928
rect 5748 4868 5752 4924
rect 5752 4868 5808 4924
rect 5808 4868 5812 4924
rect 5748 4864 5812 4868
rect 5828 4924 5892 4928
rect 5828 4868 5832 4924
rect 5832 4868 5888 4924
rect 5888 4868 5892 4924
rect 5828 4864 5892 4868
rect 5908 4924 5972 4928
rect 5908 4868 5912 4924
rect 5912 4868 5968 4924
rect 5968 4868 5972 4924
rect 5908 4864 5972 4868
rect 8768 4924 8832 4928
rect 8768 4868 8772 4924
rect 8772 4868 8828 4924
rect 8828 4868 8832 4924
rect 8768 4864 8832 4868
rect 8848 4924 8912 4928
rect 8848 4868 8852 4924
rect 8852 4868 8908 4924
rect 8908 4868 8912 4924
rect 8848 4864 8912 4868
rect 8928 4924 8992 4928
rect 8928 4868 8932 4924
rect 8932 4868 8988 4924
rect 8988 4868 8992 4924
rect 8928 4864 8992 4868
rect 9008 4924 9072 4928
rect 9008 4868 9012 4924
rect 9012 4868 9068 4924
rect 9068 4868 9072 4924
rect 9008 4864 9072 4868
rect 4118 4380 4182 4384
rect 4118 4324 4122 4380
rect 4122 4324 4178 4380
rect 4178 4324 4182 4380
rect 4118 4320 4182 4324
rect 4198 4380 4262 4384
rect 4198 4324 4202 4380
rect 4202 4324 4258 4380
rect 4258 4324 4262 4380
rect 4198 4320 4262 4324
rect 4278 4380 4342 4384
rect 4278 4324 4282 4380
rect 4282 4324 4338 4380
rect 4338 4324 4342 4380
rect 4278 4320 4342 4324
rect 4358 4380 4422 4384
rect 4358 4324 4362 4380
rect 4362 4324 4418 4380
rect 4418 4324 4422 4380
rect 4358 4320 4422 4324
rect 7218 4380 7282 4384
rect 7218 4324 7222 4380
rect 7222 4324 7278 4380
rect 7278 4324 7282 4380
rect 7218 4320 7282 4324
rect 7298 4380 7362 4384
rect 7298 4324 7302 4380
rect 7302 4324 7358 4380
rect 7358 4324 7362 4380
rect 7298 4320 7362 4324
rect 7378 4380 7442 4384
rect 7378 4324 7382 4380
rect 7382 4324 7438 4380
rect 7438 4324 7442 4380
rect 7378 4320 7442 4324
rect 7458 4380 7522 4384
rect 7458 4324 7462 4380
rect 7462 4324 7518 4380
rect 7518 4324 7522 4380
rect 7458 4320 7522 4324
rect 5668 3836 5732 3840
rect 5668 3780 5672 3836
rect 5672 3780 5728 3836
rect 5728 3780 5732 3836
rect 5668 3776 5732 3780
rect 5748 3836 5812 3840
rect 5748 3780 5752 3836
rect 5752 3780 5808 3836
rect 5808 3780 5812 3836
rect 5748 3776 5812 3780
rect 5828 3836 5892 3840
rect 5828 3780 5832 3836
rect 5832 3780 5888 3836
rect 5888 3780 5892 3836
rect 5828 3776 5892 3780
rect 5908 3836 5972 3840
rect 5908 3780 5912 3836
rect 5912 3780 5968 3836
rect 5968 3780 5972 3836
rect 5908 3776 5972 3780
rect 8768 3836 8832 3840
rect 8768 3780 8772 3836
rect 8772 3780 8828 3836
rect 8828 3780 8832 3836
rect 8768 3776 8832 3780
rect 8848 3836 8912 3840
rect 8848 3780 8852 3836
rect 8852 3780 8908 3836
rect 8908 3780 8912 3836
rect 8848 3776 8912 3780
rect 8928 3836 8992 3840
rect 8928 3780 8932 3836
rect 8932 3780 8988 3836
rect 8988 3780 8992 3836
rect 8928 3776 8992 3780
rect 9008 3836 9072 3840
rect 9008 3780 9012 3836
rect 9012 3780 9068 3836
rect 9068 3780 9072 3836
rect 9008 3776 9072 3780
rect 4118 3292 4182 3296
rect 4118 3236 4122 3292
rect 4122 3236 4178 3292
rect 4178 3236 4182 3292
rect 4118 3232 4182 3236
rect 4198 3292 4262 3296
rect 4198 3236 4202 3292
rect 4202 3236 4258 3292
rect 4258 3236 4262 3292
rect 4198 3232 4262 3236
rect 4278 3292 4342 3296
rect 4278 3236 4282 3292
rect 4282 3236 4338 3292
rect 4338 3236 4342 3292
rect 4278 3232 4342 3236
rect 4358 3292 4422 3296
rect 4358 3236 4362 3292
rect 4362 3236 4418 3292
rect 4418 3236 4422 3292
rect 4358 3232 4422 3236
rect 7218 3292 7282 3296
rect 7218 3236 7222 3292
rect 7222 3236 7278 3292
rect 7278 3236 7282 3292
rect 7218 3232 7282 3236
rect 7298 3292 7362 3296
rect 7298 3236 7302 3292
rect 7302 3236 7358 3292
rect 7358 3236 7362 3292
rect 7298 3232 7362 3236
rect 7378 3292 7442 3296
rect 7378 3236 7382 3292
rect 7382 3236 7438 3292
rect 7438 3236 7442 3292
rect 7378 3232 7442 3236
rect 7458 3292 7522 3296
rect 7458 3236 7462 3292
rect 7462 3236 7518 3292
rect 7518 3236 7522 3292
rect 7458 3232 7522 3236
rect 5668 2748 5732 2752
rect 5668 2692 5672 2748
rect 5672 2692 5728 2748
rect 5728 2692 5732 2748
rect 5668 2688 5732 2692
rect 5748 2748 5812 2752
rect 5748 2692 5752 2748
rect 5752 2692 5808 2748
rect 5808 2692 5812 2748
rect 5748 2688 5812 2692
rect 5828 2748 5892 2752
rect 5828 2692 5832 2748
rect 5832 2692 5888 2748
rect 5888 2692 5892 2748
rect 5828 2688 5892 2692
rect 5908 2748 5972 2752
rect 5908 2692 5912 2748
rect 5912 2692 5968 2748
rect 5968 2692 5972 2748
rect 5908 2688 5972 2692
rect 8768 2748 8832 2752
rect 8768 2692 8772 2748
rect 8772 2692 8828 2748
rect 8828 2692 8832 2748
rect 8768 2688 8832 2692
rect 8848 2748 8912 2752
rect 8848 2692 8852 2748
rect 8852 2692 8908 2748
rect 8908 2692 8912 2748
rect 8848 2688 8912 2692
rect 8928 2748 8992 2752
rect 8928 2692 8932 2748
rect 8932 2692 8988 2748
rect 8988 2692 8992 2748
rect 8928 2688 8992 2692
rect 9008 2748 9072 2752
rect 9008 2692 9012 2748
rect 9012 2692 9068 2748
rect 9068 2692 9072 2748
rect 9008 2688 9072 2692
rect 4118 2204 4182 2208
rect 4118 2148 4122 2204
rect 4122 2148 4178 2204
rect 4178 2148 4182 2204
rect 4118 2144 4182 2148
rect 4198 2204 4262 2208
rect 4198 2148 4202 2204
rect 4202 2148 4258 2204
rect 4258 2148 4262 2204
rect 4198 2144 4262 2148
rect 4278 2204 4342 2208
rect 4278 2148 4282 2204
rect 4282 2148 4338 2204
rect 4338 2148 4342 2204
rect 4278 2144 4342 2148
rect 4358 2204 4422 2208
rect 4358 2148 4362 2204
rect 4362 2148 4418 2204
rect 4418 2148 4422 2204
rect 4358 2144 4422 2148
rect 7218 2204 7282 2208
rect 7218 2148 7222 2204
rect 7222 2148 7278 2204
rect 7278 2148 7282 2204
rect 7218 2144 7282 2148
rect 7298 2204 7362 2208
rect 7298 2148 7302 2204
rect 7302 2148 7358 2204
rect 7358 2148 7362 2204
rect 7298 2144 7362 2148
rect 7378 2204 7442 2208
rect 7378 2148 7382 2204
rect 7382 2148 7438 2204
rect 7438 2148 7442 2204
rect 7378 2144 7442 2148
rect 7458 2204 7522 2208
rect 7458 2148 7462 2204
rect 7462 2148 7518 2204
rect 7518 2148 7522 2204
rect 7458 2144 7522 2148
rect 5668 1660 5732 1664
rect 5668 1604 5672 1660
rect 5672 1604 5728 1660
rect 5728 1604 5732 1660
rect 5668 1600 5732 1604
rect 5748 1660 5812 1664
rect 5748 1604 5752 1660
rect 5752 1604 5808 1660
rect 5808 1604 5812 1660
rect 5748 1600 5812 1604
rect 5828 1660 5892 1664
rect 5828 1604 5832 1660
rect 5832 1604 5888 1660
rect 5888 1604 5892 1660
rect 5828 1600 5892 1604
rect 5908 1660 5972 1664
rect 5908 1604 5912 1660
rect 5912 1604 5968 1660
rect 5968 1604 5972 1660
rect 5908 1600 5972 1604
rect 8768 1660 8832 1664
rect 8768 1604 8772 1660
rect 8772 1604 8828 1660
rect 8828 1604 8832 1660
rect 8768 1600 8832 1604
rect 8848 1660 8912 1664
rect 8848 1604 8852 1660
rect 8852 1604 8908 1660
rect 8908 1604 8912 1660
rect 8848 1600 8912 1604
rect 8928 1660 8992 1664
rect 8928 1604 8932 1660
rect 8932 1604 8988 1660
rect 8988 1604 8992 1660
rect 8928 1600 8992 1604
rect 9008 1660 9072 1664
rect 9008 1604 9012 1660
rect 9012 1604 9068 1660
rect 9068 1604 9072 1660
rect 9008 1600 9072 1604
rect 4118 1116 4182 1120
rect 4118 1060 4122 1116
rect 4122 1060 4178 1116
rect 4178 1060 4182 1116
rect 4118 1056 4182 1060
rect 4198 1116 4262 1120
rect 4198 1060 4202 1116
rect 4202 1060 4258 1116
rect 4258 1060 4262 1116
rect 4198 1056 4262 1060
rect 4278 1116 4342 1120
rect 4278 1060 4282 1116
rect 4282 1060 4338 1116
rect 4338 1060 4342 1116
rect 4278 1056 4342 1060
rect 4358 1116 4422 1120
rect 4358 1060 4362 1116
rect 4362 1060 4418 1116
rect 4418 1060 4422 1116
rect 4358 1056 4422 1060
rect 7218 1116 7282 1120
rect 7218 1060 7222 1116
rect 7222 1060 7278 1116
rect 7278 1060 7282 1116
rect 7218 1056 7282 1060
rect 7298 1116 7362 1120
rect 7298 1060 7302 1116
rect 7302 1060 7358 1116
rect 7358 1060 7362 1116
rect 7298 1056 7362 1060
rect 7378 1116 7442 1120
rect 7378 1060 7382 1116
rect 7382 1060 7438 1116
rect 7438 1060 7442 1116
rect 7378 1056 7442 1060
rect 7458 1116 7522 1120
rect 7458 1060 7462 1116
rect 7462 1060 7518 1116
rect 7518 1060 7522 1116
rect 7458 1056 7522 1060
<< metal4 >>
rect 2560 11456 2880 11472
rect 2560 11392 2568 11456
rect 2632 11392 2648 11456
rect 2712 11392 2728 11456
rect 2792 11392 2808 11456
rect 2872 11392 2880 11456
rect 2560 10368 2880 11392
rect 2560 10304 2568 10368
rect 2632 10304 2648 10368
rect 2712 10304 2728 10368
rect 2792 10304 2808 10368
rect 2872 10304 2880 10368
rect 2560 9280 2880 10304
rect 2560 9216 2568 9280
rect 2632 9216 2648 9280
rect 2712 9216 2728 9280
rect 2792 9216 2808 9280
rect 2872 9216 2880 9280
rect 2560 8218 2880 9216
rect 2560 8192 2602 8218
rect 2838 8192 2880 8218
rect 2560 8128 2568 8192
rect 2872 8128 2880 8192
rect 2560 7982 2602 8128
rect 2838 7982 2880 8128
rect 2560 7104 2880 7982
rect 2560 7040 2568 7104
rect 2632 7040 2648 7104
rect 2712 7040 2728 7104
rect 2792 7040 2808 7104
rect 2872 7040 2880 7104
rect 2560 6016 2880 7040
rect 2560 5952 2568 6016
rect 2632 5952 2648 6016
rect 2712 5952 2728 6016
rect 2792 5952 2808 6016
rect 2872 5952 2880 6016
rect 2560 4838 2880 5952
rect 2560 4602 2602 4838
rect 2838 4602 2880 4838
rect 1996 4196 2276 4238
rect 1996 3960 2018 4196
rect 2254 3960 2276 4196
rect 1996 3918 2276 3960
rect 1256 2506 1536 2548
rect 1256 2270 1278 2506
rect 1514 2270 1536 2506
rect 1256 2228 1536 2270
rect 2560 1458 2880 4602
rect 2560 1222 2602 1458
rect 2838 1222 2880 1458
rect 2560 1088 2880 1222
rect 3560 9266 3880 11424
rect 3560 9030 3602 9266
rect 3838 9030 3880 9266
rect 3560 5886 3880 9030
rect 3560 5650 3602 5886
rect 3838 5650 3880 5886
rect 3560 2506 3880 5650
rect 3560 2270 3602 2506
rect 3838 2270 3880 2506
rect 3560 1088 3880 2270
rect 4110 10912 4430 11472
rect 5660 11456 5980 11472
rect 4110 10848 4118 10912
rect 4182 10848 4198 10912
rect 4262 10848 4278 10912
rect 4342 10848 4358 10912
rect 4422 10848 4430 10912
rect 4110 9908 4430 10848
rect 4110 9824 4152 9908
rect 4388 9824 4430 9908
rect 4110 9760 4118 9824
rect 4422 9760 4430 9824
rect 4110 9672 4152 9760
rect 4388 9672 4430 9760
rect 4110 8736 4430 9672
rect 4110 8672 4118 8736
rect 4182 8672 4198 8736
rect 4262 8672 4278 8736
rect 4342 8672 4358 8736
rect 4422 8672 4430 8736
rect 4110 7648 4430 8672
rect 4110 7584 4118 7648
rect 4182 7584 4198 7648
rect 4262 7584 4278 7648
rect 4342 7584 4358 7648
rect 4422 7584 4430 7648
rect 4110 6560 4430 7584
rect 4110 6496 4118 6560
rect 4182 6528 4198 6560
rect 4262 6528 4278 6560
rect 4342 6528 4358 6560
rect 4422 6496 4430 6560
rect 4110 6292 4152 6496
rect 4388 6292 4430 6496
rect 4110 5472 4430 6292
rect 4110 5408 4118 5472
rect 4182 5408 4198 5472
rect 4262 5408 4278 5472
rect 4342 5408 4358 5472
rect 4422 5408 4430 5472
rect 4110 4384 4430 5408
rect 4110 4320 4118 4384
rect 4182 4320 4198 4384
rect 4262 4320 4278 4384
rect 4342 4320 4358 4384
rect 4422 4320 4430 4384
rect 4110 3296 4430 4320
rect 4110 3232 4118 3296
rect 4182 3232 4198 3296
rect 4262 3232 4278 3296
rect 4342 3232 4358 3296
rect 4422 3232 4430 3296
rect 4110 3148 4430 3232
rect 4110 2912 4152 3148
rect 4388 2912 4430 3148
rect 4110 2208 4430 2912
rect 4110 2144 4118 2208
rect 4182 2144 4198 2208
rect 4262 2144 4278 2208
rect 4342 2144 4358 2208
rect 4422 2144 4430 2208
rect 4110 1120 4430 2144
rect 4110 1056 4118 1120
rect 4182 1056 4198 1120
rect 4262 1056 4278 1120
rect 4342 1056 4358 1120
rect 4422 1056 4430 1120
rect 5110 10956 5430 11424
rect 5110 10720 5152 10956
rect 5388 10720 5430 10956
rect 5110 7576 5430 10720
rect 5110 7340 5152 7576
rect 5388 7340 5430 7576
rect 5110 4196 5430 7340
rect 5110 3960 5152 4196
rect 5388 3960 5430 4196
rect 5110 1088 5430 3960
rect 5660 11392 5668 11456
rect 5732 11392 5748 11456
rect 5812 11392 5828 11456
rect 5892 11392 5908 11456
rect 5972 11392 5980 11456
rect 5660 10368 5980 11392
rect 5660 10304 5668 10368
rect 5732 10304 5748 10368
rect 5812 10304 5828 10368
rect 5892 10304 5908 10368
rect 5972 10304 5980 10368
rect 5660 9280 5980 10304
rect 5660 9216 5668 9280
rect 5732 9216 5748 9280
rect 5812 9216 5828 9280
rect 5892 9216 5908 9280
rect 5972 9216 5980 9280
rect 5660 8218 5980 9216
rect 5660 8192 5702 8218
rect 5938 8192 5980 8218
rect 5660 8128 5668 8192
rect 5972 8128 5980 8192
rect 5660 7982 5702 8128
rect 5938 7982 5980 8128
rect 5660 7104 5980 7982
rect 5660 7040 5668 7104
rect 5732 7040 5748 7104
rect 5812 7040 5828 7104
rect 5892 7040 5908 7104
rect 5972 7040 5980 7104
rect 5660 6016 5980 7040
rect 5660 5952 5668 6016
rect 5732 5952 5748 6016
rect 5812 5952 5828 6016
rect 5892 5952 5908 6016
rect 5972 5952 5980 6016
rect 5660 4928 5980 5952
rect 5660 4864 5668 4928
rect 5732 4864 5748 4928
rect 5812 4864 5828 4928
rect 5892 4864 5908 4928
rect 5972 4864 5980 4928
rect 5660 4838 5980 4864
rect 5660 4602 5702 4838
rect 5938 4602 5980 4838
rect 5660 3840 5980 4602
rect 5660 3776 5668 3840
rect 5732 3776 5748 3840
rect 5812 3776 5828 3840
rect 5892 3776 5908 3840
rect 5972 3776 5980 3840
rect 5660 2752 5980 3776
rect 5660 2688 5668 2752
rect 5732 2688 5748 2752
rect 5812 2688 5828 2752
rect 5892 2688 5908 2752
rect 5972 2688 5980 2752
rect 5660 1664 5980 2688
rect 5660 1600 5668 1664
rect 5732 1600 5748 1664
rect 5812 1600 5828 1664
rect 5892 1600 5908 1664
rect 5972 1600 5980 1664
rect 5660 1458 5980 1600
rect 5660 1222 5702 1458
rect 5938 1222 5980 1458
rect 4110 1040 4430 1056
rect 5660 1040 5980 1222
rect 6660 9266 6980 11424
rect 6660 9030 6702 9266
rect 6938 9030 6980 9266
rect 6660 5886 6980 9030
rect 6660 5650 6702 5886
rect 6938 5650 6980 5886
rect 6660 2506 6980 5650
rect 6660 2270 6702 2506
rect 6938 2270 6980 2506
rect 6660 1088 6980 2270
rect 7210 10912 7530 11472
rect 8760 11456 9080 11472
rect 7210 10848 7218 10912
rect 7282 10848 7298 10912
rect 7362 10848 7378 10912
rect 7442 10848 7458 10912
rect 7522 10848 7530 10912
rect 7210 9908 7530 10848
rect 7210 9824 7252 9908
rect 7488 9824 7530 9908
rect 7210 9760 7218 9824
rect 7522 9760 7530 9824
rect 7210 9672 7252 9760
rect 7488 9672 7530 9760
rect 7210 8736 7530 9672
rect 7210 8672 7218 8736
rect 7282 8672 7298 8736
rect 7362 8672 7378 8736
rect 7442 8672 7458 8736
rect 7522 8672 7530 8736
rect 7210 7648 7530 8672
rect 7210 7584 7218 7648
rect 7282 7584 7298 7648
rect 7362 7584 7378 7648
rect 7442 7584 7458 7648
rect 7522 7584 7530 7648
rect 7210 6560 7530 7584
rect 7210 6496 7218 6560
rect 7282 6528 7298 6560
rect 7362 6528 7378 6560
rect 7442 6528 7458 6560
rect 7522 6496 7530 6560
rect 7210 6292 7252 6496
rect 7488 6292 7530 6496
rect 7210 5472 7530 6292
rect 7210 5408 7218 5472
rect 7282 5408 7298 5472
rect 7362 5408 7378 5472
rect 7442 5408 7458 5472
rect 7522 5408 7530 5472
rect 7210 4384 7530 5408
rect 7210 4320 7218 4384
rect 7282 4320 7298 4384
rect 7362 4320 7378 4384
rect 7442 4320 7458 4384
rect 7522 4320 7530 4384
rect 7210 3296 7530 4320
rect 7210 3232 7218 3296
rect 7282 3232 7298 3296
rect 7362 3232 7378 3296
rect 7442 3232 7458 3296
rect 7522 3232 7530 3296
rect 7210 3148 7530 3232
rect 7210 2912 7252 3148
rect 7488 2912 7530 3148
rect 7210 2208 7530 2912
rect 7210 2144 7218 2208
rect 7282 2144 7298 2208
rect 7362 2144 7378 2208
rect 7442 2144 7458 2208
rect 7522 2144 7530 2208
rect 7210 1120 7530 2144
rect 7210 1056 7218 1120
rect 7282 1056 7298 1120
rect 7362 1056 7378 1120
rect 7442 1056 7458 1120
rect 7522 1056 7530 1120
rect 8210 10956 8530 11424
rect 8210 10720 8252 10956
rect 8488 10720 8530 10956
rect 8210 7576 8530 10720
rect 8210 7340 8252 7576
rect 8488 7340 8530 7576
rect 8210 4196 8530 7340
rect 8210 3960 8252 4196
rect 8488 3960 8530 4196
rect 8210 1088 8530 3960
rect 8760 11392 8768 11456
rect 8832 11392 8848 11456
rect 8912 11392 8928 11456
rect 8992 11392 9008 11456
rect 9072 11392 9080 11456
rect 8760 10368 9080 11392
rect 8760 10304 8768 10368
rect 8832 10304 8848 10368
rect 8912 10304 8928 10368
rect 8992 10304 9008 10368
rect 9072 10304 9080 10368
rect 8760 9280 9080 10304
rect 8760 9216 8768 9280
rect 8832 9216 8848 9280
rect 8912 9216 8928 9280
rect 8992 9216 9008 9280
rect 9072 9216 9080 9280
rect 8760 8218 9080 9216
rect 8760 8192 8802 8218
rect 9038 8192 9080 8218
rect 8760 8128 8768 8192
rect 9072 8128 9080 8192
rect 8760 7982 8802 8128
rect 9038 7982 9080 8128
rect 8760 7104 9080 7982
rect 8760 7040 8768 7104
rect 8832 7040 8848 7104
rect 8912 7040 8928 7104
rect 8992 7040 9008 7104
rect 9072 7040 9080 7104
rect 8760 6016 9080 7040
rect 8760 5952 8768 6016
rect 8832 5952 8848 6016
rect 8912 5952 8928 6016
rect 8992 5952 9008 6016
rect 9072 5952 9080 6016
rect 8760 4928 9080 5952
rect 8760 4864 8768 4928
rect 8832 4864 8848 4928
rect 8912 4864 8928 4928
rect 8992 4864 9008 4928
rect 9072 4864 9080 4928
rect 8760 4838 9080 4864
rect 8760 4602 8802 4838
rect 9038 4602 9080 4838
rect 8760 3840 9080 4602
rect 8760 3776 8768 3840
rect 8832 3776 8848 3840
rect 8912 3776 8928 3840
rect 8992 3776 9008 3840
rect 9072 3776 9080 3840
rect 8760 2752 9080 3776
rect 8760 2688 8768 2752
rect 8832 2688 8848 2752
rect 8912 2688 8928 2752
rect 8992 2688 9008 2752
rect 9072 2688 9080 2752
rect 8760 1664 9080 2688
rect 8760 1600 8768 1664
rect 8832 1600 8848 1664
rect 8912 1600 8928 1664
rect 8992 1600 9008 1664
rect 9072 1600 9080 1664
rect 8760 1458 9080 1600
rect 8760 1222 8802 1458
rect 9038 1222 9080 1458
rect 7210 1040 7530 1056
rect 8760 1040 9080 1222
<< via4 >>
rect 2602 8192 2838 8218
rect 2602 8128 2632 8192
rect 2632 8128 2648 8192
rect 2648 8128 2712 8192
rect 2712 8128 2728 8192
rect 2728 8128 2792 8192
rect 2792 8128 2808 8192
rect 2808 8128 2838 8192
rect 2602 7982 2838 8128
rect 2602 4602 2838 4838
rect 2018 3960 2254 4196
rect 1278 2270 1514 2506
rect 2602 1222 2838 1458
rect 3602 9030 3838 9266
rect 3602 5650 3838 5886
rect 3602 2270 3838 2506
rect 4152 9824 4388 9908
rect 4152 9760 4182 9824
rect 4182 9760 4198 9824
rect 4198 9760 4262 9824
rect 4262 9760 4278 9824
rect 4278 9760 4342 9824
rect 4342 9760 4358 9824
rect 4358 9760 4388 9824
rect 4152 9672 4388 9760
rect 4152 6496 4182 6528
rect 4182 6496 4198 6528
rect 4198 6496 4262 6528
rect 4262 6496 4278 6528
rect 4278 6496 4342 6528
rect 4342 6496 4358 6528
rect 4358 6496 4388 6528
rect 4152 6292 4388 6496
rect 4152 2912 4388 3148
rect 5152 10720 5388 10956
rect 5152 7340 5388 7576
rect 5152 3960 5388 4196
rect 5702 8192 5938 8218
rect 5702 8128 5732 8192
rect 5732 8128 5748 8192
rect 5748 8128 5812 8192
rect 5812 8128 5828 8192
rect 5828 8128 5892 8192
rect 5892 8128 5908 8192
rect 5908 8128 5938 8192
rect 5702 7982 5938 8128
rect 5702 4602 5938 4838
rect 5702 1222 5938 1458
rect 6702 9030 6938 9266
rect 6702 5650 6938 5886
rect 6702 2270 6938 2506
rect 7252 9824 7488 9908
rect 7252 9760 7282 9824
rect 7282 9760 7298 9824
rect 7298 9760 7362 9824
rect 7362 9760 7378 9824
rect 7378 9760 7442 9824
rect 7442 9760 7458 9824
rect 7458 9760 7488 9824
rect 7252 9672 7488 9760
rect 7252 6496 7282 6528
rect 7282 6496 7298 6528
rect 7298 6496 7362 6528
rect 7362 6496 7378 6528
rect 7378 6496 7442 6528
rect 7442 6496 7458 6528
rect 7458 6496 7488 6528
rect 7252 6292 7488 6496
rect 7252 2912 7488 3148
rect 8252 10720 8488 10956
rect 8252 7340 8488 7576
rect 8252 3960 8488 4196
rect 8802 8192 9038 8218
rect 8802 8128 8832 8192
rect 8832 8128 8848 8192
rect 8848 8128 8912 8192
rect 8912 8128 8928 8192
rect 8928 8128 8992 8192
rect 8992 8128 9008 8192
rect 9008 8128 9038 8192
rect 8802 7982 9038 8128
rect 8802 4602 9038 4838
rect 8802 1222 9038 1458
<< metal5 >>
rect 920 10956 9844 10998
rect 920 10720 5152 10956
rect 5388 10720 8252 10956
rect 8488 10720 9844 10956
rect 920 10678 9844 10720
rect 920 9908 9844 9950
rect 920 9672 4152 9908
rect 4388 9672 7252 9908
rect 7488 9672 9844 9908
rect 920 9630 9844 9672
rect 920 9266 9844 9308
rect 920 9030 3602 9266
rect 3838 9030 6702 9266
rect 6938 9030 9844 9266
rect 920 8988 9844 9030
rect 920 8218 9844 8260
rect 920 7982 2602 8218
rect 2838 7982 5702 8218
rect 5938 7982 8802 8218
rect 9038 7982 9844 8218
rect 920 7940 9844 7982
rect 920 7576 9844 7618
rect 920 7340 5152 7576
rect 5388 7340 8252 7576
rect 8488 7340 9844 7576
rect 920 7298 9844 7340
rect 920 6528 9844 6570
rect 920 6292 4152 6528
rect 4388 6292 7252 6528
rect 7488 6292 9844 6528
rect 920 6250 9844 6292
rect 920 5886 9844 5928
rect 920 5650 3602 5886
rect 3838 5650 6702 5886
rect 6938 5650 9844 5886
rect 920 5608 9844 5650
rect 920 4838 9844 4880
rect 920 4602 2602 4838
rect 2838 4602 5702 4838
rect 5938 4602 8802 4838
rect 9038 4602 9844 4838
rect 920 4560 9844 4602
rect 920 4196 9844 4238
rect 920 3960 2018 4196
rect 2254 3960 5152 4196
rect 5388 3960 8252 4196
rect 8488 3960 9844 4196
rect 920 3918 9844 3960
rect 920 3148 9844 3190
rect 920 2912 4152 3148
rect 4388 2912 7252 3148
rect 7488 2912 9844 3148
rect 920 2870 9844 2912
rect 920 2506 9844 2548
rect 920 2270 1278 2506
rect 1514 2270 3602 2506
rect 3838 2270 6702 2506
rect 6938 2270 9844 2506
rect 920 2228 9844 2270
rect 920 1458 9844 1500
rect 920 1222 2602 1458
rect 2838 1222 5702 1458
rect 5938 1222 8802 1458
rect 9038 1222 9844 1458
rect 920 1180 9844 1222
use sky130_fd_sc_hd__decap_3  PHY_4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 3036 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1635271187
transform 1 0 3036 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1635271187
transform 1 0 3036 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_26 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 3312 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_26
timestamp 1635271187
transform 1 0 3312 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_26
timestamp 1635271187
transform 1 0 3312 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _113_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform -1 0 3588 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1635271187
transform 1 0 3036 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1635271187
transform 1 0 3036 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1635271187
transform 1 0 3036 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_26 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 3312 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_26
timestamp 1635271187
transform 1 0 3312 0 -1 3264
box -38 -48 774 592
use gpio_logic_high  gpio_logic_high
timestamp 1636122974
transform 1 0 1196 0 1 1680
box -38 -48 1418 2768
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 5612 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_50
timestamp 1635271187
transform 1 0 5520 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_38
timestamp 1635271187
transform 1 0 4416 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_52
timestamp 1635271187
transform 1 0 5704 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 5520 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_38
timestamp 1635271187
transform 1 0 4416 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1635271187
transform 1 0 5612 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_52
timestamp 1635271187
transform 1 0 5704 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_50
timestamp 1635271187
transform 1 0 5520 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_38
timestamp 1635271187
transform 1 0 4416 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__dfbbn_1  _209_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 4232 0 -1 3264
box -38 -48 2430 592
use sky130_fd_sc_hd__fill_2  FILLER_3_34 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 4048 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _117_
timestamp 1635271187
transform -1 0 4968 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _115_
timestamp 1635271187
transform -1 0 4600 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _109_
timestamp 1635271187
transform -1 0 5244 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1635271187
transform 1 0 5612 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_52
timestamp 1635271187
transform 1 0 5704 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_47 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 5244 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_40
timestamp 1635271187
transform 1 0 4600 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_34
timestamp 1635271187
transform 1 0 4048 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dfbbn_1  _208_
timestamp 1635271187
transform 1 0 3588 0 -1 4352
box -38 -48 2430 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1635271187
transform 1 0 8188 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1635271187
transform 1 0 8188 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_80
timestamp 1635271187
transform 1 0 8280 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_78
timestamp 1635271187
transform 1 0 8096 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_74
timestamp 1635271187
transform 1 0 7728 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1635271187
transform 1 0 6624 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_80
timestamp 1635271187
transform 1 0 8280 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_76
timestamp 1635271187
transform 1 0 7912 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_64
timestamp 1635271187
transform 1 0 6808 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_76
timestamp 1635271187
transform 1 0 7912 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_64
timestamp 1635271187
transform 1 0 6808 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform -1 0 8372 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1635271187
transform -1 0 8188 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _185_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 8280 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _135_
timestamp 1635271187
transform -1 0 7912 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1635271187
transform 1 0 8188 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_70
timestamp 1635271187
transform 1 0 7360 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_62
timestamp 1635271187
transform 1 0 6624 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dfbbn_1  _205_
timestamp 1635271187
transform 1 0 6532 0 1 3264
box -38 -48 2430 592
use sky130_fd_sc_hd__fill_1  FILLER_4_60
timestamp 1635271187
transform 1 0 6440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output28 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform -1 0 8188 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp 1635271187
transform -1 0 8648 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _134_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 7084 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _133_
timestamp 1635271187
transform -1 0 7820 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _132_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 6532 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _131_
timestamp 1635271187
transform -1 0 6532 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _130_
timestamp 1635271187
transform -1 0 6256 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1635271187
transform 1 0 8188 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  const_source $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 8924 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_90
timestamp 1635271187
transform 1 0 9200 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_84
timestamp 1635271187
transform 1 0 8648 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1635271187
transform -1 0 8924 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1635271187
transform 1 0 9292 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1635271187
transform -1 0 9844 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1635271187
transform -1 0 9844 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_92
timestamp 1635271187
transform 1 0 9384 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  output25
timestamp 1635271187
transform 1 0 9200 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1635271187
transform -1 0 8924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _184_
timestamp 1635271187
transform 1 0 8924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_81
timestamp 1635271187
transform 1 0 8372 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1635271187
transform -1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1635271187
transform -1 0 9844 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output24
timestamp 1635271187
transform 1 0 8832 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 1635271187
transform 1 0 9200 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _180_
timestamp 1635271187
transform -1 0 8832 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1635271187
transform -1 0 9844 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _183_
timestamp 1635271187
transform 1 0 8924 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1635271187
transform -1 0 9844 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_93
timestamp 1635271187
transform 1 0 9476 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _194_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 8648 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1635271187
transform -1 0 9844 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_93
timestamp 1635271187
transform 1 0 9476 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1635271187
transform 1 0 3036 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_26
timestamp 1635271187
transform 1 0 3312 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _217_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 3312 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1635271187
transform 1 0 3036 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _147_
timestamp 1635271187
transform -1 0 3496 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _146_
timestamp 1635271187
transform -1 0 2760 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _144_
timestamp 1635271187
transform -1 0 3036 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1635271187
transform 1 0 920 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1635271187
transform 1 0 1196 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_15
timestamp 1635271187
transform 1 0 2300 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_1  _216_
timestamp 1635271187
transform 1 0 2392 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1635271187
transform 1 0 920 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_7
timestamp 1635271187
transform 1 0 1564 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_3
timestamp 1635271187
transform 1 0 1196 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_9_13
timestamp 1635271187
transform 1 0 2116 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_10
timestamp 1635271187
transform 1 0 1840 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1635271187
transform -1 0 1840 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1635271187
transform -1 0 2116 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_1  _215_
timestamp 1635271187
transform 1 0 1656 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  _148_
timestamp 1635271187
transform -1 0 1656 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1635271187
transform 1 0 920 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1635271187
transform -1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _125_
timestamp 1635271187
transform -1 0 5612 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _116_
timestamp 1635271187
transform 1 0 5704 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _114_
timestamp 1635271187
transform 1 0 3680 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _112_
timestamp 1635271187
transform 1 0 3404 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _110_
timestamp 1635271187
transform 1 0 4876 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _108_
timestamp 1635271187
transform 1 0 4324 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1635271187
transform 1 0 5612 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_36
timestamp 1635271187
transform 1 0 4232 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__dfbbn_1  _206_
timestamp 1635271187
transform 1 0 5796 0 -1 5440
box -38 -48 2430 592
use sky130_fd_sc_hd__clkbuf_1  _124_
timestamp 1635271187
transform 1 0 5428 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _119_
timestamp 1635271187
transform -1 0 5428 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_52
timestamp 1635271187
transform 1 0 5704 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _222_
timestamp 1635271187
transform 1 0 4232 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__or2b_1  _145_
timestamp 1635271187
transform -1 0 4140 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1635271187
transform 1 0 3496 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_35
timestamp 1635271187
transform 1 0 4140 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_serial_clock $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform -1 0 6072 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfbbn_1  _203_
timestamp 1635271187
transform 1 0 3588 0 1 6528
box -38 -48 2430 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1635271187
transform 1 0 3496 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_2  gpio_in_buf $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 7820 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _186_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform -1 0 7820 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _129_
timestamp 1635271187
transform -1 0 6808 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _127_
timestamp 1635271187
transform -1 0 7084 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _123_
timestamp 1635271187
transform -1 0 7360 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _111_
timestamp 1635271187
transform 1 0 6164 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_60
timestamp 1635271187
transform 1 0 6440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 1635271187
transform 1 0 8280 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1635271187
transform 1 0 8188 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _223_
timestamp 1635271187
transform 1 0 6256 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__or2_1  _128_
timestamp 1635271187
transform 1 0 8096 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1635271187
transform 1 0 6072 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_57
timestamp 1635271187
transform 1 0 6164 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__dfbbn_1  _207_
timestamp 1635271187
transform 1 0 6808 0 -1 6528
box -38 -48 2430 592
use sky130_fd_sc_hd__or2b_1  _126_
timestamp 1635271187
transform 1 0 6256 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1635271187
transform 1 0 6072 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_57
timestamp 1635271187
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _221_
timestamp 1635271187
transform -1 0 8648 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__or2b_1  _120_
timestamp 1635271187
transform 1 0 6256 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _118_
timestamp 1635271187
transform 1 0 5980 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _195_
timestamp 1635271187
transform -1 0 9476 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__186__A
timestamp 1635271187
transform -1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1635271187
transform -1 0 9844 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_93
timestamp 1635271187
transform 1 0 9476 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__ebufn_1  _197_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 8648 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1635271187
transform -1 0 9844 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_92
timestamp 1635271187
transform 1 0 9384 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__or2b_1  _179_
timestamp 1635271187
transform -1 0 9292 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1635271187
transform 1 0 8648 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1635271187
transform 1 0 8556 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _121_
timestamp 1635271187
transform 1 0 9292 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1635271187
transform -1 0 9844 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output29
timestamp 1635271187
transform 1 0 9200 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1635271187
transform -1 0 9844 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _196_
timestamp 1635271187
transform 1 0 8740 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1635271187
transform 1 0 8648 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1635271187
transform -1 0 9844 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_serial_clock $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform -1 0 2576 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dfbbn_1  _202_
timestamp 1635271187
transform 1 0 2576 0 -1 7616
box -38 -48 2430 592
use sky130_fd_sc_hd__clkbuf_1  _182_
timestamp 1635271187
transform -1 0 1656 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _149_
timestamp 1635271187
transform -1 0 1932 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _143_
timestamp 1635271187
transform -1 0 2208 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1635271187
transform 1 0 920 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1635271187
transform -1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_1  _214_
timestamp 1635271187
transform -1 0 3496 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  _188_
timestamp 1635271187
transform -1 0 1656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1635271187
transform 1 0 920 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1635271187
transform -1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  output37
timestamp 1635271187
transform -1 0 2024 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _213_
timestamp 1635271187
transform 1 0 2300 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  _150_
timestamp 1635271187
transform -1 0 2300 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1635271187
transform 1 0 920 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1635271187
transform -1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1635271187
transform -1 0 1564 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1635271187
transform -1 0 1748 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1635271187
transform 1 0 920 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1635271187
transform 1 0 920 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1635271187
transform -1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1635271187
transform -1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1635271187
transform -1 0 1656 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1635271187
transform -1 0 1656 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1635271187
transform -1 0 1932 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1635271187
transform -1 0 1932 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1635271187
transform -1 0 2208 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1635271187
transform -1 0 2116 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1635271187
transform -1 0 2392 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _137_
timestamp 1635271187
transform 1 0 2484 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _138_
timestamp 1635271187
transform -1 0 2484 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _140_
timestamp 1635271187
transform -1 0 3496 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _172_
timestamp 1635271187
transform -1 0 3220 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _189_
timestamp 1635271187
transform -1 0 2944 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _190_
timestamp 1635271187
transform -1 0 2668 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfbbn_1  _204_
timestamp 1635271187
transform 1 0 2760 0 -1 9792
box -38 -48 2430 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _107_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform -1 0 5980 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__fill_1  FILLER_11_44
timestamp 1635271187
transform 1 0 4968 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__dfbbn_1  _210_
timestamp 1635271187
transform 1 0 5152 0 1 7616
box -38 -48 2430 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _136_
timestamp 1635271187
transform 1 0 4232 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__or2b_1  _102_
timestamp 1635271187
transform 1 0 3680 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1635271187
transform 1 0 3496 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_29
timestamp 1635271187
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _218_
timestamp 1635271187
transform 1 0 4140 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1635271187
transform 1 0 3496 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _142_
timestamp 1635271187
transform 1 0 4600 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _151_
timestamp 1635271187
transform 1 0 3588 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _153_
timestamp 1635271187
transform 1 0 4140 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_14_43
timestamp 1635271187
transform 1 0 4876 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_52
timestamp 1635271187
transform 1 0 5704 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _152_
timestamp 1635271187
transform 1 0 5152 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _154_
timestamp 1635271187
transform 1 0 5428 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _155_
timestamp 1635271187
transform 1 0 5796 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output34
timestamp 1635271187
transform -1 0 5336 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _219_
timestamp 1635271187
transform 1 0 5336 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_2  output31
timestamp 1635271187
transform 1 0 8280 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _220_
timestamp 1635271187
transform 1 0 6440 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  _103_
timestamp 1635271187
transform -1 0 6440 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1635271187
transform 1 0 6072 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1635271187
transform 1 0 5980 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output32
timestamp 1635271187
transform -1 0 8648 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _122_
timestamp 1635271187
transform 1 0 7544 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _105_
timestamp 1635271187
transform 1 0 8004 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_serial_clock
timestamp 1635271187
transform 1 0 6808 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dfbbn_1  _201_
timestamp 1635271187
transform 1 0 7176 0 -1 8704
box -38 -48 2430 592
use sky130_fd_sc_hd__or2_1  _104_
timestamp 1635271187
transform 1 0 6164 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1635271187
transform 1 0 6072 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1635271187
transform 1 0 5980 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_serial_clock_A
timestamp 1635271187
transform 1 0 6624 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__buf_12  input17 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform -1 0 8648 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform -1 0 6900 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dfbbn_1  _200_
timestamp 1635271187
transform 1 0 7176 0 -1 9792
box -38 -48 2430 592
use sky130_fd_sc_hd__inv_2  _106_
timestamp 1635271187
transform 1 0 6900 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1635271187
transform 1 0 6072 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _193_
timestamp 1635271187
transform -1 0 9476 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1635271187
transform -1 0 9844 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_93
timestamp 1635271187
transform 1 0 9476 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output30
timestamp 1635271187
transform 1 0 9200 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _181_
timestamp 1635271187
transform -1 0 9200 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1635271187
transform 1 0 8648 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1635271187
transform -1 0 9844 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output33
timestamp 1635271187
transform 1 0 9200 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _159_
timestamp 1635271187
transform 1 0 8740 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1635271187
transform 1 0 8648 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1635271187
transform -1 0 9844 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1635271187
transform -1 0 9844 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1635271187
transform -1 0 9844 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1635271187
transform -1 0 1656 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _212_
timestamp 1635271187
transform -1 0 3496 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1635271187
transform 1 0 920 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1635271187
transform -1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1635271187
transform -1 0 2852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1635271187
transform -1 0 1472 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1635271187
transform -1 0 1748 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1635271187
transform -1 0 2024 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1635271187
transform -1 0 2300 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1635271187
transform -1 0 2576 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _139_
timestamp 1635271187
transform 1 0 2852 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1635271187
transform 1 0 920 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1635271187
transform 1 0 920 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1635271187
transform -1 0 1472 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1635271187
transform -1 0 1748 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_9
timestamp 1635271187
transform 1 0 1748 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1635271187
transform -1 0 2116 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1635271187
transform -1 0 2392 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _187_
timestamp 1635271187
transform -1 0 2944 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _192_
timestamp 1635271187
transform -1 0 2668 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _178_
timestamp 1635271187
transform -1 0 3220 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _176_
timestamp 1635271187
transform -1 0 3496 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dfbbn_1  _199_
timestamp 1635271187
transform 1 0 3680 0 1 9792
box -38 -48 2430 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1635271187
transform 1 0 3496 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_29
timestamp 1635271187
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _177_
timestamp 1635271187
transform -1 0 6072 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _171_
timestamp 1635271187
transform 1 0 4416 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _169_
timestamp 1635271187
transform 1 0 3864 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _158_
timestamp 1635271187
transform -1 0 5336 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _156_
timestamp 1635271187
transform -1 0 5612 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _141_
timestamp 1635271187
transform 1 0 3404 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1635271187
transform -1 0 5060 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1635271187
transform 1 0 3588 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1635271187
transform 1 0 3496 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _168_
timestamp 1635271187
transform 1 0 4048 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _174_
timestamp 1635271187
transform -1 0 4048 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1635271187
transform -1 0 4508 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _170_
timestamp 1635271187
transform 1 0 4784 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _173_
timestamp 1635271187
transform 1 0 4508 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _161_
timestamp 1635271187
transform -1 0 5336 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _160_
timestamp 1635271187
transform -1 0 5612 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _167_
timestamp 1635271187
transform 1 0 5612 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _211_
timestamp 1635271187
transform -1 0 7912 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__or2b_1  _157_
timestamp 1635271187
transform -1 0 8464 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__dfbbn_1  _198_
timestamp 1635271187
transform 1 0 6164 0 -1 10880
box -38 -48 2430 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1635271187
transform 1 0 6072 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1635271187
transform -1 0 6072 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_57
timestamp 1635271187
transform 1 0 6164 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1635271187
transform 1 0 6072 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__or2b_1  _175_
timestamp 1635271187
transform -1 0 6808 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _162_
timestamp 1635271187
transform -1 0 7084 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _166_
timestamp 1635271187
transform -1 0 7360 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _163_
timestamp 1635271187
transform -1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _164_
timestamp 1635271187
transform -1 0 7636 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_79
timestamp 1635271187
transform 1 0 8188 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output40
timestamp 1635271187
transform 1 0 8280 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _191_
timestamp 1635271187
transform 1 0 8832 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1635271187
transform 1 0 8648 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_85
timestamp 1635271187
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1635271187
transform -1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  output35
timestamp 1635271187
transform -1 0 9568 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1635271187
transform -1 0 9844 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output39
timestamp 1635271187
transform 1 0 8832 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _165_
timestamp 1635271187
transform 1 0 8556 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1635271187
transform 1 0 8648 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_85
timestamp 1635271187
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output38
timestamp 1635271187
transform 1 0 9200 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output36
timestamp 1635271187
transform 1 0 9200 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1635271187
transform -1 0 9844 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1635271187
transform -1 0 9844 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1635271187
transform -1 0 9200 0 -1 10880
box -38 -48 222 592
<< labels >>
rlabel metal2 s 938 12200 994 13000 6 gpio_defaults[0]
port 0 nsew signal input
rlabel metal2 s 5538 12200 5594 13000 6 gpio_defaults[10]
port 1 nsew signal input
rlabel metal2 s 5998 12200 6054 13000 6 gpio_defaults[11]
port 2 nsew signal input
rlabel metal2 s 6458 12200 6514 13000 6 gpio_defaults[12]
port 3 nsew signal input
rlabel metal2 s 1398 12200 1454 13000 6 gpio_defaults[1]
port 4 nsew signal input
rlabel metal2 s 1858 12200 1914 13000 6 gpio_defaults[2]
port 5 nsew signal input
rlabel metal2 s 2318 12200 2374 13000 6 gpio_defaults[3]
port 6 nsew signal input
rlabel metal2 s 2778 12200 2834 13000 6 gpio_defaults[4]
port 7 nsew signal input
rlabel metal2 s 3238 12200 3294 13000 6 gpio_defaults[5]
port 8 nsew signal input
rlabel metal2 s 3698 12200 3754 13000 6 gpio_defaults[6]
port 9 nsew signal input
rlabel metal2 s 4158 12200 4214 13000 6 gpio_defaults[7]
port 10 nsew signal input
rlabel metal2 s 4618 12200 4674 13000 6 gpio_defaults[8]
port 11 nsew signal input
rlabel metal2 s 5078 12200 5134 13000 6 gpio_defaults[9]
port 12 nsew signal input
rlabel metal3 s 14000 1232 34000 1352 6 mgmt_gpio_in
port 13 nsew signal tristate
rlabel metal3 s 14000 1640 34000 1760 6 mgmt_gpio_oeb
port 14 nsew signal input
rlabel metal3 s 14000 2048 34000 2168 6 mgmt_gpio_out
port 15 nsew signal input
rlabel metal3 s 14000 824 34000 944 6 one
port 16 nsew signal tristate
rlabel metal3 s 14000 2456 34000 2576 6 pad_gpio_ana_en
port 17 nsew signal tristate
rlabel metal3 s 14000 2864 34000 2984 6 pad_gpio_ana_pol
port 18 nsew signal tristate
rlabel metal3 s 14000 3272 34000 3392 6 pad_gpio_ana_sel
port 19 nsew signal tristate
rlabel metal3 s 14000 3680 34000 3800 6 pad_gpio_dm[0]
port 20 nsew signal tristate
rlabel metal3 s 14000 4088 34000 4208 6 pad_gpio_dm[1]
port 21 nsew signal tristate
rlabel metal3 s 14000 4496 34000 4616 6 pad_gpio_dm[2]
port 22 nsew signal tristate
rlabel metal3 s 14000 4904 34000 5024 6 pad_gpio_holdover
port 23 nsew signal tristate
rlabel metal3 s 14000 5312 34000 5432 6 pad_gpio_ib_mode_sel
port 24 nsew signal tristate
rlabel metal3 s 14000 5720 34000 5840 6 pad_gpio_in
port 25 nsew signal input
rlabel metal3 s 14000 6128 34000 6248 6 pad_gpio_inenb
port 26 nsew signal tristate
rlabel metal3 s 14000 6536 34000 6656 6 pad_gpio_out
port 27 nsew signal tristate
rlabel metal3 s 14000 6944 34000 7064 6 pad_gpio_outenb
port 28 nsew signal tristate
rlabel metal3 s 14000 7352 34000 7472 6 pad_gpio_slow_sel
port 29 nsew signal tristate
rlabel metal3 s 14000 7760 34000 7880 6 pad_gpio_vtrip_sel
port 30 nsew signal tristate
rlabel metal3 s 14000 8168 34000 8288 6 resetn
port 31 nsew signal input
rlabel metal3 s 14000 8576 34000 8696 6 resetn_out
port 32 nsew signal tristate
rlabel metal3 s 14000 8984 34000 9104 6 serial_clock
port 33 nsew signal input
rlabel metal3 s 14000 9392 34000 9512 6 serial_clock_out
port 34 nsew signal tristate
rlabel metal3 s 14000 9800 34000 9920 6 serial_data_in
port 35 nsew signal input
rlabel metal3 s 14000 10208 34000 10328 6 serial_data_out
port 36 nsew signal tristate
rlabel metal3 s 14000 10616 34000 10736 6 serial_load
port 37 nsew signal input
rlabel metal3 s 14000 11024 34000 11144 6 serial_load_out
port 38 nsew signal tristate
rlabel metal3 s 14000 11432 34000 11552 6 user_gpio_in
port 39 nsew signal tristate
rlabel metal3 s 14000 11840 34000 11960 6 user_gpio_oeb
port 40 nsew signal input
rlabel metal3 s 14000 12248 34000 12368 6 user_gpio_out
port 41 nsew signal input
rlabel metal5 s 920 1180 9844 1500 6 vccd
port 42 nsew power input
rlabel metal5 s 920 4560 9844 4880 6 vccd
port 42 nsew power input
rlabel metal5 s 920 7940 9844 8260 6 vccd
port 42 nsew power input
rlabel metal4 s 2560 1088 2880 11472 6 vccd
port 42 nsew power input
rlabel metal4 s 5660 1040 5980 11472 6 vccd
port 42 nsew power input
rlabel metal4 s 8760 1040 9080 11472 6 vccd
port 42 nsew power input
rlabel metal5 s 920 2228 9844 2548 6 vccd1
port 43 nsew power input
rlabel metal5 s 920 5608 9844 5928 6 vccd1
port 43 nsew power input
rlabel metal5 s 920 8988 9844 9308 6 vccd1
port 43 nsew power input
rlabel metal4 s 3560 1088 3880 11424 6 vccd1
port 43 nsew power input
rlabel metal4 s 6660 1088 6980 11424 6 vccd1
port 43 nsew power input
rlabel metal5 s 920 2870 9844 3190 6 vssd
port 44 nsew ground input
rlabel metal5 s 920 6250 9844 6570 6 vssd
port 44 nsew ground input
rlabel metal5 s 920 9630 9844 9950 6 vssd
port 44 nsew ground input
rlabel metal4 s 4110 1040 4430 11472 6 vssd
port 44 nsew ground input
rlabel metal4 s 7210 1040 7530 11472 6 vssd
port 44 nsew ground input
rlabel metal5 s 920 3918 9844 4238 6 vssd1
port 45 nsew ground input
rlabel metal5 s 920 7298 9844 7618 6 vssd1
port 45 nsew ground input
rlabel metal5 s 920 10678 9844 10998 6 vssd1
port 45 nsew ground input
rlabel metal4 s 5110 1088 5430 11424 6 vssd1
port 45 nsew ground input
rlabel metal4 s 8210 1088 8530 11424 6 vssd1
port 45 nsew ground input
rlabel metal3 s 14000 416 34000 536 6 zero
port 46 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 34000 13000
<< end >>
