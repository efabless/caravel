magic
tech sky130A
magscale 1 2
timestamp 1675767944
<< nwell >>
rect 1066 26373 382850 26694
rect 1066 25285 382850 25851
rect 1066 24197 382850 24763
rect 1066 23109 382850 23675
rect 1066 22021 382850 22587
rect 1066 20933 382850 21499
rect 1066 19845 382850 20411
rect 1066 18757 382850 19323
rect 1066 17669 382850 18235
rect 1066 16581 382850 17147
rect 1066 15493 382850 16059
rect 1066 14405 382850 14971
rect 1066 13317 250278 13883
rect 1066 12474 250278 12795
rect 1066 12229 133714 12474
rect 1066 11386 133714 11707
rect 1066 11141 64070 11386
rect 1066 10053 64070 10619
rect 1066 8965 64070 9531
rect 1066 7877 64070 8443
rect 1066 6789 64070 7355
rect 1066 5701 64070 6267
rect 1066 4613 133714 5179
rect 1066 3525 133714 4091
rect 1066 2437 382850 3003
rect 1066 1349 382850 1915
<< obsli1 >>
rect 1104 1071 382812 26673
<< obsm1 >>
rect 1104 8 382812 27996
<< metal2 >>
rect 11610 27200 11666 28400
rect 12346 27200 12402 28400
rect 13082 27200 13138 28400
rect 13818 27200 13874 28400
rect 14554 27200 14610 28400
rect 15290 27200 15346 28400
rect 16026 27200 16082 28400
rect 16762 27200 16818 28400
rect 17498 27200 17554 28400
rect 18234 27200 18290 28400
rect 18970 27200 19026 28400
rect 19706 27200 19762 28400
rect 20442 27200 20498 28400
rect 21178 27200 21234 28400
rect 21914 27200 21970 28400
rect 22650 27200 22706 28400
rect 23386 27200 23442 28400
rect 24122 27200 24178 28400
rect 24858 27200 24914 28400
rect 25594 27200 25650 28400
rect 26330 27200 26386 28400
rect 27066 27200 27122 28400
rect 27802 27200 27858 28400
rect 28538 27200 28594 28400
rect 29274 27200 29330 28400
rect 30010 27200 30066 28400
rect 30746 27200 30802 28400
rect 31482 27200 31538 28400
rect 32218 27200 32274 28400
rect 32954 27200 33010 28400
rect 33690 27200 33746 28400
rect 34426 27200 34482 28400
rect 35162 27200 35218 28400
rect 35898 27200 35954 28400
rect 36634 27200 36690 28400
rect 37370 27200 37426 28400
rect 38106 27200 38162 28400
rect 38842 27200 38898 28400
rect 39578 27200 39634 28400
rect 40314 27200 40370 28400
rect 41050 27200 41106 28400
rect 41786 27200 41842 28400
rect 42522 27200 42578 28400
rect 43258 27200 43314 28400
rect 43994 27200 44050 28400
rect 44730 27200 44786 28400
rect 45466 27200 45522 28400
rect 46202 27200 46258 28400
rect 46938 27200 46994 28400
rect 47674 27200 47730 28400
rect 48410 27200 48466 28400
rect 49146 27200 49202 28400
rect 49882 27200 49938 28400
rect 50618 27200 50674 28400
rect 51354 27200 51410 28400
rect 52090 27200 52146 28400
rect 52826 27200 52882 28400
rect 53562 27200 53618 28400
rect 54298 27200 54354 28400
rect 55034 27200 55090 28400
rect 55770 27200 55826 28400
rect 56506 27200 56562 28400
rect 57242 27200 57298 28400
rect 57978 27200 58034 28400
rect 58714 27200 58770 28400
rect 59450 27200 59506 28400
rect 60186 27200 60242 28400
rect 60922 27200 60978 28400
rect 61658 27200 61714 28400
rect 62394 27200 62450 28400
rect 63130 27200 63186 28400
rect 63866 27200 63922 28400
rect 64602 27200 64658 28400
rect 65338 27200 65394 28400
rect 66074 27200 66130 28400
rect 66810 27200 66866 28400
rect 67546 27200 67602 28400
rect 68282 27200 68338 28400
rect 69018 27200 69074 28400
rect 69754 27200 69810 28400
rect 70490 27200 70546 28400
rect 71226 27200 71282 28400
rect 71962 27200 72018 28400
rect 72698 27200 72754 28400
rect 73434 27200 73490 28400
rect 74170 27200 74226 28400
rect 74906 27200 74962 28400
rect 75642 27200 75698 28400
rect 76378 27200 76434 28400
rect 77114 27200 77170 28400
rect 77850 27200 77906 28400
rect 78586 27200 78642 28400
rect 79322 27200 79378 28400
rect 80058 27200 80114 28400
rect 80794 27200 80850 28400
rect 81530 27200 81586 28400
rect 82266 27200 82322 28400
rect 83002 27200 83058 28400
rect 83738 27200 83794 28400
rect 84474 27200 84530 28400
rect 85210 27200 85266 28400
rect 85946 27200 86002 28400
rect 86682 27200 86738 28400
rect 87418 27200 87474 28400
rect 88154 27200 88210 28400
rect 88890 27200 88946 28400
rect 89626 27200 89682 28400
rect 90362 27200 90418 28400
rect 91098 27200 91154 28400
rect 91834 27200 91890 28400
rect 92570 27200 92626 28400
rect 93306 27200 93362 28400
rect 94042 27200 94098 28400
rect 94778 27200 94834 28400
rect 95514 27200 95570 28400
rect 96250 27200 96306 28400
rect 96986 27200 97042 28400
rect 97722 27200 97778 28400
rect 98458 27200 98514 28400
rect 99194 27200 99250 28400
rect 99930 27200 99986 28400
rect 100666 27200 100722 28400
rect 101402 27200 101458 28400
rect 102138 27200 102194 28400
rect 102874 27200 102930 28400
rect 103610 27200 103666 28400
rect 104346 27200 104402 28400
rect 105082 27200 105138 28400
rect 105818 27200 105874 28400
rect 106554 27200 106610 28400
rect 107290 27200 107346 28400
rect 108026 27200 108082 28400
rect 108762 27200 108818 28400
rect 109498 27200 109554 28400
rect 110234 27200 110290 28400
rect 110970 27200 111026 28400
rect 111706 27200 111762 28400
rect 112442 27200 112498 28400
rect 113178 27200 113234 28400
rect 113914 27200 113970 28400
rect 114650 27200 114706 28400
rect 115386 27200 115442 28400
rect 116122 27200 116178 28400
rect 116858 27200 116914 28400
rect 117594 27200 117650 28400
rect 118330 27200 118386 28400
rect 119066 27200 119122 28400
rect 119802 27200 119858 28400
rect 120538 27200 120594 28400
rect 121274 27200 121330 28400
rect 122010 27200 122066 28400
rect 122746 27200 122802 28400
rect 123482 27200 123538 28400
rect 124218 27200 124274 28400
rect 124954 27200 125010 28400
rect 125690 27200 125746 28400
rect 126426 27200 126482 28400
rect 127162 27200 127218 28400
rect 127898 27200 127954 28400
rect 128634 27200 128690 28400
rect 129370 27200 129426 28400
rect 130106 27200 130162 28400
rect 130842 27200 130898 28400
rect 131578 27200 131634 28400
rect 132314 27200 132370 28400
rect 133050 27200 133106 28400
rect 133786 27200 133842 28400
rect 134522 27200 134578 28400
rect 135258 27200 135314 28400
rect 135994 27200 136050 28400
rect 136730 27200 136786 28400
rect 137466 27200 137522 28400
rect 138202 27200 138258 28400
rect 138938 27200 138994 28400
rect 139674 27200 139730 28400
rect 140410 27200 140466 28400
rect 141146 27200 141202 28400
rect 141882 27200 141938 28400
rect 142618 27200 142674 28400
rect 143354 27200 143410 28400
rect 144090 27200 144146 28400
rect 144826 27200 144882 28400
rect 145562 27200 145618 28400
rect 146298 27200 146354 28400
rect 147034 27200 147090 28400
rect 147770 27200 147826 28400
rect 148506 27200 148562 28400
rect 149242 27200 149298 28400
rect 149978 27200 150034 28400
rect 150714 27200 150770 28400
rect 151450 27200 151506 28400
rect 152186 27200 152242 28400
rect 152922 27200 152978 28400
rect 153658 27200 153714 28400
rect 154394 27200 154450 28400
rect 155130 27200 155186 28400
rect 155866 27200 155922 28400
rect 156602 27200 156658 28400
rect 157338 27200 157394 28400
rect 158074 27200 158130 28400
rect 158810 27200 158866 28400
rect 159546 27200 159602 28400
rect 160282 27200 160338 28400
rect 161018 27200 161074 28400
rect 161754 27200 161810 28400
rect 162490 27200 162546 28400
rect 163226 27200 163282 28400
rect 163962 27200 164018 28400
rect 164698 27200 164754 28400
rect 165434 27200 165490 28400
rect 166170 27200 166226 28400
rect 166906 27200 166962 28400
rect 167642 27200 167698 28400
rect 168378 27200 168434 28400
rect 169114 27200 169170 28400
rect 169850 27200 169906 28400
rect 170586 27200 170642 28400
rect 171322 27200 171378 28400
rect 172058 27200 172114 28400
rect 172794 27200 172850 28400
rect 173530 27200 173586 28400
rect 174266 27200 174322 28400
rect 175002 27200 175058 28400
rect 175738 27200 175794 28400
rect 176474 27200 176530 28400
rect 177210 27200 177266 28400
rect 177946 27200 178002 28400
rect 178682 27200 178738 28400
rect 179418 27200 179474 28400
rect 180154 27200 180210 28400
rect 180890 27200 180946 28400
rect 181626 27200 181682 28400
rect 182362 27200 182418 28400
rect 183098 27200 183154 28400
rect 183834 27200 183890 28400
rect 184570 27200 184626 28400
rect 185306 27200 185362 28400
rect 186042 27200 186098 28400
rect 186778 27200 186834 28400
rect 187514 27200 187570 28400
rect 188250 27200 188306 28400
rect 188986 27200 189042 28400
rect 189722 27200 189778 28400
rect 190458 27200 190514 28400
rect 191194 27200 191250 28400
rect 191930 27200 191986 28400
rect 192666 27200 192722 28400
rect 193402 27200 193458 28400
rect 194138 27200 194194 28400
rect 194874 27200 194930 28400
rect 195610 27200 195666 28400
rect 196346 27200 196402 28400
rect 197082 27200 197138 28400
rect 197818 27200 197874 28400
rect 198554 27200 198610 28400
rect 199290 27200 199346 28400
rect 200026 27200 200082 28400
rect 200762 27200 200818 28400
rect 201498 27200 201554 28400
rect 202234 27200 202290 28400
rect 202970 27200 203026 28400
rect 203706 27200 203762 28400
rect 204442 27200 204498 28400
rect 205178 27200 205234 28400
rect 205914 27200 205970 28400
rect 206650 27200 206706 28400
rect 207386 27200 207442 28400
rect 208122 27200 208178 28400
rect 208858 27200 208914 28400
rect 209594 27200 209650 28400
rect 210330 27200 210386 28400
rect 211066 27200 211122 28400
rect 211802 27200 211858 28400
rect 212538 27200 212594 28400
rect 213274 27200 213330 28400
rect 214010 27200 214066 28400
rect 214746 27200 214802 28400
rect 215482 27200 215538 28400
rect 216218 27200 216274 28400
rect 216954 27200 217010 28400
rect 217690 27200 217746 28400
rect 218426 27200 218482 28400
rect 219162 27200 219218 28400
rect 219898 27200 219954 28400
rect 220634 27200 220690 28400
rect 221370 27200 221426 28400
rect 222106 27200 222162 28400
rect 222842 27200 222898 28400
rect 223578 27200 223634 28400
rect 224314 27200 224370 28400
rect 225050 27200 225106 28400
rect 225786 27200 225842 28400
rect 226522 27200 226578 28400
rect 227258 27200 227314 28400
rect 227994 27200 228050 28400
rect 228730 27200 228786 28400
rect 229466 27200 229522 28400
rect 230202 27200 230258 28400
rect 230938 27200 230994 28400
rect 231674 27200 231730 28400
rect 232410 27200 232466 28400
rect 233146 27200 233202 28400
rect 233882 27200 233938 28400
rect 234618 27200 234674 28400
rect 235354 27200 235410 28400
rect 236090 27200 236146 28400
rect 236826 27200 236882 28400
rect 237562 27200 237618 28400
rect 238298 27200 238354 28400
rect 239034 27200 239090 28400
rect 239770 27200 239826 28400
rect 240506 27200 240562 28400
rect 241242 27200 241298 28400
rect 241978 27200 242034 28400
rect 242714 27200 242770 28400
rect 243450 27200 243506 28400
rect 244186 27200 244242 28400
rect 244922 27200 244978 28400
rect 245658 27200 245714 28400
rect 246394 27200 246450 28400
rect 247130 27200 247186 28400
rect 247866 27200 247922 28400
rect 248602 27200 248658 28400
rect 249338 27200 249394 28400
rect 250074 27200 250130 28400
rect 250810 27200 250866 28400
rect 251546 27200 251602 28400
rect 252282 27200 252338 28400
rect 253018 27200 253074 28400
rect 253754 27200 253810 28400
rect 254490 27200 254546 28400
rect 255226 27200 255282 28400
rect 255962 27200 256018 28400
rect 256698 27200 256754 28400
rect 257434 27200 257490 28400
rect 258170 27200 258226 28400
rect 258906 27200 258962 28400
rect 259642 27200 259698 28400
rect 260378 27200 260434 28400
rect 261114 27200 261170 28400
rect 261850 27200 261906 28400
rect 262586 27200 262642 28400
rect 263322 27200 263378 28400
rect 264058 27200 264114 28400
rect 264794 27200 264850 28400
rect 265530 27200 265586 28400
rect 266266 27200 266322 28400
rect 267002 27200 267058 28400
rect 267738 27200 267794 28400
rect 268474 27200 268530 28400
rect 269210 27200 269266 28400
rect 269946 27200 270002 28400
rect 270682 27200 270738 28400
rect 271418 27200 271474 28400
rect 272154 27200 272210 28400
rect 272890 27200 272946 28400
rect 273626 27200 273682 28400
rect 274362 27200 274418 28400
rect 275098 27200 275154 28400
rect 275834 27200 275890 28400
rect 276570 27200 276626 28400
rect 277306 27200 277362 28400
rect 278042 27200 278098 28400
rect 278778 27200 278834 28400
rect 279514 27200 279570 28400
rect 280250 27200 280306 28400
rect 280986 27200 281042 28400
rect 281722 27200 281778 28400
rect 282458 27200 282514 28400
rect 283194 27200 283250 28400
rect 283930 27200 283986 28400
rect 284666 27200 284722 28400
rect 285402 27200 285458 28400
rect 286138 27200 286194 28400
rect 286874 27200 286930 28400
rect 287610 27200 287666 28400
rect 288346 27200 288402 28400
rect 289082 27200 289138 28400
rect 289818 27200 289874 28400
rect 290554 27200 290610 28400
rect 291290 27200 291346 28400
rect 292026 27200 292082 28400
rect 292762 27200 292818 28400
rect 293498 27200 293554 28400
rect 294234 27200 294290 28400
rect 294970 27200 295026 28400
rect 295706 27200 295762 28400
rect 296442 27200 296498 28400
rect 297178 27200 297234 28400
rect 297914 27200 297970 28400
rect 298650 27200 298706 28400
rect 299386 27200 299442 28400
rect 300122 27200 300178 28400
rect 300858 27200 300914 28400
rect 301594 27200 301650 28400
rect 302330 27200 302386 28400
rect 303066 27200 303122 28400
rect 303802 27200 303858 28400
rect 304538 27200 304594 28400
rect 305274 27200 305330 28400
rect 306010 27200 306066 28400
rect 306746 27200 306802 28400
rect 307482 27200 307538 28400
rect 308218 27200 308274 28400
rect 308954 27200 309010 28400
rect 309690 27200 309746 28400
rect 310426 27200 310482 28400
rect 311162 27200 311218 28400
rect 311898 27200 311954 28400
rect 312634 27200 312690 28400
rect 313370 27200 313426 28400
rect 314106 27200 314162 28400
rect 314842 27200 314898 28400
rect 315578 27200 315634 28400
rect 316314 27200 316370 28400
rect 317050 27200 317106 28400
rect 317786 27200 317842 28400
rect 318522 27200 318578 28400
rect 319258 27200 319314 28400
rect 319994 27200 320050 28400
rect 320730 27200 320786 28400
rect 321466 27200 321522 28400
rect 322202 27200 322258 28400
rect 322938 27200 322994 28400
rect 323674 27200 323730 28400
rect 324410 27200 324466 28400
rect 325146 27200 325202 28400
rect 325882 27200 325938 28400
rect 326618 27200 326674 28400
rect 327354 27200 327410 28400
rect 328090 27200 328146 28400
rect 328826 27200 328882 28400
rect 329562 27200 329618 28400
rect 330298 27200 330354 28400
rect 331034 27200 331090 28400
rect 331770 27200 331826 28400
rect 332506 27200 332562 28400
rect 333242 27200 333298 28400
rect 333978 27200 334034 28400
rect 334714 27200 334770 28400
rect 335450 27200 335506 28400
rect 336186 27200 336242 28400
rect 336922 27200 336978 28400
rect 337658 27200 337714 28400
rect 338394 27200 338450 28400
rect 339130 27200 339186 28400
rect 339866 27200 339922 28400
rect 340602 27200 340658 28400
rect 341338 27200 341394 28400
rect 342074 27200 342130 28400
rect 342810 27200 342866 28400
rect 343546 27200 343602 28400
rect 344282 27200 344338 28400
rect 345018 27200 345074 28400
rect 345754 27200 345810 28400
rect 346490 27200 346546 28400
rect 347226 27200 347282 28400
rect 347962 27200 348018 28400
rect 348698 27200 348754 28400
rect 349434 27200 349490 28400
rect 350170 27200 350226 28400
rect 350906 27200 350962 28400
rect 351642 27200 351698 28400
rect 352378 27200 352434 28400
rect 353114 27200 353170 28400
rect 353850 27200 353906 28400
rect 354586 27200 354642 28400
rect 355322 27200 355378 28400
rect 356058 27200 356114 28400
rect 356794 27200 356850 28400
rect 357530 27200 357586 28400
rect 358266 27200 358322 28400
rect 359002 27200 359058 28400
rect 359738 27200 359794 28400
rect 360474 27200 360530 28400
rect 361210 27200 361266 28400
rect 361946 27200 362002 28400
rect 362682 27200 362738 28400
rect 363418 27200 363474 28400
rect 364154 27200 364210 28400
rect 364890 27200 364946 28400
rect 365626 27200 365682 28400
rect 366362 27200 366418 28400
rect 367098 27200 367154 28400
rect 367834 27200 367890 28400
rect 368570 27200 368626 28400
rect 369306 27200 369362 28400
rect 370042 27200 370098 28400
rect 370778 27200 370834 28400
rect 371514 27200 371570 28400
rect 372250 27200 372306 28400
rect 21362 -400 21418 800
rect 21914 -400 21970 800
rect 22466 -400 22522 800
rect 23018 -400 23074 800
rect 23570 -400 23626 800
rect 24122 -400 24178 800
rect 24674 -400 24730 800
rect 25226 -400 25282 800
rect 25778 -400 25834 800
rect 26330 -400 26386 800
rect 26882 -400 26938 800
rect 27434 -400 27490 800
rect 27986 -400 28042 800
rect 28538 -400 28594 800
rect 29090 -400 29146 800
rect 29642 -400 29698 800
rect 30194 -400 30250 800
rect 30746 -400 30802 800
rect 31298 -400 31354 800
rect 31850 -400 31906 800
rect 32402 -400 32458 800
rect 32954 -400 33010 800
rect 33506 -400 33562 800
rect 34058 -400 34114 800
rect 34610 -400 34666 800
rect 35162 -400 35218 800
rect 35714 -400 35770 800
rect 36266 -400 36322 800
rect 36818 -400 36874 800
rect 37370 -400 37426 800
rect 37922 -400 37978 800
rect 38474 -400 38530 800
rect 39026 -400 39082 800
rect 39578 -400 39634 800
rect 40130 -400 40186 800
rect 40682 -400 40738 800
rect 41234 -400 41290 800
rect 41786 -400 41842 800
rect 42338 -400 42394 800
rect 42890 -400 42946 800
rect 43442 -400 43498 800
rect 43994 -400 44050 800
rect 44546 -400 44602 800
rect 45098 -400 45154 800
rect 45650 -400 45706 800
rect 46202 -400 46258 800
rect 46754 -400 46810 800
rect 47306 -400 47362 800
rect 47858 -400 47914 800
rect 48410 -400 48466 800
rect 48962 -400 49018 800
rect 49514 -400 49570 800
rect 50066 -400 50122 800
rect 50618 -400 50674 800
rect 51170 -400 51226 800
rect 51722 -400 51778 800
rect 52274 -400 52330 800
rect 52826 -400 52882 800
rect 53378 -400 53434 800
rect 53930 -400 53986 800
rect 54482 -400 54538 800
rect 55034 -400 55090 800
rect 55586 -400 55642 800
rect 56138 -400 56194 800
rect 56690 -400 56746 800
rect 57242 -400 57298 800
rect 57794 -400 57850 800
rect 58346 -400 58402 800
rect 58898 -400 58954 800
rect 59450 -400 59506 800
rect 60002 -400 60058 800
rect 60554 -400 60610 800
rect 61106 -400 61162 800
rect 61658 -400 61714 800
rect 62210 -400 62266 800
rect 62762 -400 62818 800
rect 63314 -400 63370 800
rect 63866 -400 63922 800
rect 64418 -400 64474 800
rect 64970 -400 65026 800
rect 65522 -400 65578 800
rect 66074 -400 66130 800
rect 66626 -400 66682 800
rect 67178 -400 67234 800
rect 67730 -400 67786 800
rect 68282 -400 68338 800
rect 68834 -400 68890 800
rect 69386 -400 69442 800
rect 69938 -400 69994 800
rect 70490 -400 70546 800
rect 71042 -400 71098 800
rect 71594 -400 71650 800
rect 72146 -400 72202 800
rect 72698 -400 72754 800
rect 73250 -400 73306 800
rect 73802 -400 73858 800
rect 74354 -400 74410 800
rect 74906 -400 74962 800
rect 75458 -400 75514 800
rect 76010 -400 76066 800
rect 76562 -400 76618 800
rect 77114 -400 77170 800
rect 77666 -400 77722 800
rect 78218 -400 78274 800
rect 78770 -400 78826 800
rect 79322 -400 79378 800
rect 79874 -400 79930 800
rect 80426 -400 80482 800
rect 80978 -400 81034 800
rect 81530 -400 81586 800
rect 82082 -400 82138 800
rect 82634 -400 82690 800
rect 83186 -400 83242 800
rect 83738 -400 83794 800
rect 84290 -400 84346 800
rect 84842 -400 84898 800
rect 85394 -400 85450 800
rect 85946 -400 86002 800
rect 86498 -400 86554 800
rect 87050 -400 87106 800
rect 87602 -400 87658 800
rect 88154 -400 88210 800
rect 88706 -400 88762 800
rect 89258 -400 89314 800
rect 89810 -400 89866 800
rect 90362 -400 90418 800
rect 90914 -400 90970 800
rect 91466 -400 91522 800
rect 92018 -400 92074 800
rect 92570 -400 92626 800
rect 93122 -400 93178 800
rect 93674 -400 93730 800
rect 94226 -400 94282 800
rect 94778 -400 94834 800
rect 95330 -400 95386 800
rect 95882 -400 95938 800
rect 96434 -400 96490 800
rect 96986 -400 97042 800
rect 97538 -400 97594 800
rect 98090 -400 98146 800
rect 98642 -400 98698 800
rect 99194 -400 99250 800
rect 99746 -400 99802 800
rect 100298 -400 100354 800
rect 100850 -400 100906 800
rect 101402 -400 101458 800
rect 101954 -400 102010 800
rect 102506 -400 102562 800
rect 103058 -400 103114 800
rect 103610 -400 103666 800
rect 104162 -400 104218 800
rect 104714 -400 104770 800
rect 105266 -400 105322 800
rect 105818 -400 105874 800
rect 106370 -400 106426 800
rect 106922 -400 106978 800
rect 107474 -400 107530 800
rect 108026 -400 108082 800
rect 108578 -400 108634 800
rect 109130 -400 109186 800
rect 109682 -400 109738 800
rect 110234 -400 110290 800
rect 110786 -400 110842 800
rect 111338 -400 111394 800
rect 111890 -400 111946 800
rect 112442 -400 112498 800
rect 112994 -400 113050 800
rect 113546 -400 113602 800
rect 114098 -400 114154 800
rect 114650 -400 114706 800
rect 115202 -400 115258 800
rect 115754 -400 115810 800
rect 116306 -400 116362 800
rect 116858 -400 116914 800
rect 117410 -400 117466 800
rect 117962 -400 118018 800
rect 118514 -400 118570 800
rect 119066 -400 119122 800
rect 119618 -400 119674 800
rect 120170 -400 120226 800
rect 120722 -400 120778 800
rect 121274 -400 121330 800
rect 121826 -400 121882 800
rect 122378 -400 122434 800
rect 122930 -400 122986 800
rect 123482 -400 123538 800
rect 124034 -400 124090 800
rect 124586 -400 124642 800
rect 125138 -400 125194 800
rect 125690 -400 125746 800
rect 126242 -400 126298 800
rect 126794 -400 126850 800
rect 127346 -400 127402 800
rect 127898 -400 127954 800
rect 128450 -400 128506 800
rect 129002 -400 129058 800
rect 129554 -400 129610 800
rect 130106 -400 130162 800
rect 130658 -400 130714 800
rect 131210 -400 131266 800
rect 131762 -400 131818 800
rect 132314 -400 132370 800
rect 132866 -400 132922 800
rect 133418 -400 133474 800
rect 133970 -400 134026 800
rect 134522 -400 134578 800
rect 135074 -400 135130 800
rect 135626 -400 135682 800
rect 136178 -400 136234 800
rect 136730 -400 136786 800
rect 137282 -400 137338 800
rect 137834 -400 137890 800
rect 138386 -400 138442 800
rect 138938 -400 138994 800
rect 139490 -400 139546 800
rect 140042 -400 140098 800
rect 140594 -400 140650 800
rect 141146 -400 141202 800
rect 141698 -400 141754 800
rect 142250 -400 142306 800
rect 142802 -400 142858 800
rect 143354 -400 143410 800
rect 143906 -400 143962 800
rect 144458 -400 144514 800
rect 145010 -400 145066 800
rect 145562 -400 145618 800
rect 146114 -400 146170 800
rect 146666 -400 146722 800
rect 147218 -400 147274 800
rect 147770 -400 147826 800
rect 148322 -400 148378 800
rect 148874 -400 148930 800
rect 149426 -400 149482 800
rect 149978 -400 150034 800
rect 150530 -400 150586 800
rect 151082 -400 151138 800
rect 151634 -400 151690 800
rect 152186 -400 152242 800
rect 152738 -400 152794 800
rect 153290 -400 153346 800
rect 153842 -400 153898 800
rect 154394 -400 154450 800
rect 154946 -400 155002 800
rect 155498 -400 155554 800
rect 156050 -400 156106 800
rect 156602 -400 156658 800
rect 157154 -400 157210 800
rect 157706 -400 157762 800
rect 158258 -400 158314 800
rect 158810 -400 158866 800
rect 159362 -400 159418 800
rect 159914 -400 159970 800
rect 160466 -400 160522 800
rect 161018 -400 161074 800
rect 161570 -400 161626 800
rect 162122 -400 162178 800
rect 162674 -400 162730 800
rect 163226 -400 163282 800
rect 163778 -400 163834 800
rect 164330 -400 164386 800
rect 164882 -400 164938 800
rect 165434 -400 165490 800
rect 165986 -400 166042 800
rect 166538 -400 166594 800
rect 167090 -400 167146 800
rect 167642 -400 167698 800
rect 168194 -400 168250 800
rect 168746 -400 168802 800
rect 169298 -400 169354 800
rect 169850 -400 169906 800
rect 170402 -400 170458 800
rect 170954 -400 171010 800
rect 171506 -400 171562 800
rect 172058 -400 172114 800
rect 172610 -400 172666 800
rect 173162 -400 173218 800
rect 173714 -400 173770 800
rect 174266 -400 174322 800
rect 174818 -400 174874 800
rect 175370 -400 175426 800
rect 175922 -400 175978 800
rect 176474 -400 176530 800
rect 177026 -400 177082 800
rect 177578 -400 177634 800
rect 178130 -400 178186 800
rect 178682 -400 178738 800
rect 179234 -400 179290 800
rect 179786 -400 179842 800
rect 180338 -400 180394 800
rect 180890 -400 180946 800
rect 181442 -400 181498 800
rect 181994 -400 182050 800
rect 182546 -400 182602 800
rect 183098 -400 183154 800
rect 183650 -400 183706 800
rect 184202 -400 184258 800
rect 184754 -400 184810 800
rect 185306 -400 185362 800
rect 185858 -400 185914 800
rect 186410 -400 186466 800
rect 186962 -400 187018 800
rect 187514 -400 187570 800
rect 188066 -400 188122 800
rect 188618 -400 188674 800
rect 189170 -400 189226 800
rect 189722 -400 189778 800
rect 190274 -400 190330 800
rect 190826 -400 190882 800
rect 191378 -400 191434 800
rect 191930 -400 191986 800
rect 192482 -400 192538 800
rect 193034 -400 193090 800
rect 193586 -400 193642 800
rect 194138 -400 194194 800
rect 194690 -400 194746 800
rect 195242 -400 195298 800
rect 195794 -400 195850 800
rect 196346 -400 196402 800
rect 196898 -400 196954 800
rect 197450 -400 197506 800
rect 198002 -400 198058 800
rect 198554 -400 198610 800
rect 199106 -400 199162 800
rect 199658 -400 199714 800
rect 200210 -400 200266 800
rect 200762 -400 200818 800
rect 201314 -400 201370 800
rect 201866 -400 201922 800
rect 202418 -400 202474 800
rect 202970 -400 203026 800
rect 203522 -400 203578 800
rect 204074 -400 204130 800
rect 204626 -400 204682 800
rect 205178 -400 205234 800
rect 205730 -400 205786 800
rect 206282 -400 206338 800
rect 206834 -400 206890 800
rect 207386 -400 207442 800
rect 207938 -400 207994 800
rect 208490 -400 208546 800
rect 209042 -400 209098 800
rect 209594 -400 209650 800
rect 210146 -400 210202 800
rect 210698 -400 210754 800
rect 211250 -400 211306 800
rect 211802 -400 211858 800
rect 212354 -400 212410 800
rect 212906 -400 212962 800
rect 213458 -400 213514 800
rect 214010 -400 214066 800
rect 214562 -400 214618 800
rect 215114 -400 215170 800
rect 215666 -400 215722 800
rect 216218 -400 216274 800
rect 216770 -400 216826 800
rect 217322 -400 217378 800
rect 217874 -400 217930 800
rect 218426 -400 218482 800
rect 218978 -400 219034 800
rect 219530 -400 219586 800
rect 220082 -400 220138 800
rect 220634 -400 220690 800
rect 221186 -400 221242 800
rect 221738 -400 221794 800
rect 222290 -400 222346 800
rect 222842 -400 222898 800
rect 223394 -400 223450 800
rect 223946 -400 224002 800
rect 224498 -400 224554 800
rect 225050 -400 225106 800
rect 225602 -400 225658 800
rect 226154 -400 226210 800
rect 226706 -400 226762 800
rect 227258 -400 227314 800
rect 227810 -400 227866 800
rect 228362 -400 228418 800
rect 228914 -400 228970 800
rect 229466 -400 229522 800
rect 230018 -400 230074 800
rect 230570 -400 230626 800
rect 231122 -400 231178 800
rect 231674 -400 231730 800
rect 232226 -400 232282 800
rect 232778 -400 232834 800
rect 233330 -400 233386 800
rect 233882 -400 233938 800
rect 234434 -400 234490 800
rect 234986 -400 235042 800
rect 235538 -400 235594 800
rect 236090 -400 236146 800
rect 236642 -400 236698 800
rect 237194 -400 237250 800
rect 237746 -400 237802 800
rect 238298 -400 238354 800
rect 238850 -400 238906 800
rect 239402 -400 239458 800
rect 239954 -400 240010 800
rect 240506 -400 240562 800
rect 241058 -400 241114 800
rect 241610 -400 241666 800
rect 242162 -400 242218 800
rect 242714 -400 242770 800
rect 243266 -400 243322 800
rect 243818 -400 243874 800
rect 244370 -400 244426 800
rect 244922 -400 244978 800
rect 245474 -400 245530 800
rect 246026 -400 246082 800
rect 246578 -400 246634 800
rect 247130 -400 247186 800
rect 247682 -400 247738 800
rect 248234 -400 248290 800
rect 248786 -400 248842 800
rect 249338 -400 249394 800
rect 249890 -400 249946 800
rect 250442 -400 250498 800
rect 250994 -400 251050 800
rect 251546 -400 251602 800
rect 252098 -400 252154 800
rect 252650 -400 252706 800
rect 253202 -400 253258 800
rect 253754 -400 253810 800
rect 254306 -400 254362 800
rect 254858 -400 254914 800
rect 255410 -400 255466 800
rect 255962 -400 256018 800
rect 256514 -400 256570 800
rect 257066 -400 257122 800
rect 257618 -400 257674 800
rect 258170 -400 258226 800
rect 258722 -400 258778 800
rect 259274 -400 259330 800
rect 259826 -400 259882 800
rect 260378 -400 260434 800
rect 260930 -400 260986 800
rect 261482 -400 261538 800
rect 262034 -400 262090 800
rect 262586 -400 262642 800
rect 263138 -400 263194 800
rect 263690 -400 263746 800
rect 264242 -400 264298 800
rect 264794 -400 264850 800
rect 265346 -400 265402 800
rect 265898 -400 265954 800
rect 266450 -400 266506 800
rect 267002 -400 267058 800
rect 267554 -400 267610 800
rect 268106 -400 268162 800
rect 268658 -400 268714 800
rect 269210 -400 269266 800
rect 269762 -400 269818 800
rect 270314 -400 270370 800
rect 270866 -400 270922 800
rect 271418 -400 271474 800
rect 271970 -400 272026 800
rect 272522 -400 272578 800
rect 273074 -400 273130 800
rect 273626 -400 273682 800
rect 274178 -400 274234 800
rect 274730 -400 274786 800
rect 275282 -400 275338 800
rect 275834 -400 275890 800
rect 276386 -400 276442 800
rect 276938 -400 276994 800
rect 277490 -400 277546 800
rect 278042 -400 278098 800
rect 278594 -400 278650 800
rect 279146 -400 279202 800
rect 279698 -400 279754 800
rect 280250 -400 280306 800
rect 280802 -400 280858 800
rect 281354 -400 281410 800
rect 281906 -400 281962 800
rect 282458 -400 282514 800
rect 283010 -400 283066 800
rect 283562 -400 283618 800
rect 284114 -400 284170 800
rect 284666 -400 284722 800
rect 285218 -400 285274 800
rect 285770 -400 285826 800
rect 286322 -400 286378 800
rect 286874 -400 286930 800
rect 287426 -400 287482 800
rect 287978 -400 288034 800
rect 288530 -400 288586 800
rect 289082 -400 289138 800
rect 289634 -400 289690 800
rect 290186 -400 290242 800
rect 290738 -400 290794 800
rect 291290 -400 291346 800
rect 291842 -400 291898 800
rect 292394 -400 292450 800
rect 292946 -400 293002 800
rect 293498 -400 293554 800
rect 294050 -400 294106 800
rect 294602 -400 294658 800
rect 295154 -400 295210 800
rect 295706 -400 295762 800
rect 296258 -400 296314 800
rect 296810 -400 296866 800
rect 297362 -400 297418 800
rect 297914 -400 297970 800
rect 298466 -400 298522 800
rect 299018 -400 299074 800
rect 299570 -400 299626 800
rect 300122 -400 300178 800
rect 300674 -400 300730 800
rect 301226 -400 301282 800
rect 301778 -400 301834 800
rect 302330 -400 302386 800
rect 302882 -400 302938 800
rect 303434 -400 303490 800
rect 303986 -400 304042 800
rect 304538 -400 304594 800
rect 305090 -400 305146 800
rect 305642 -400 305698 800
rect 306194 -400 306250 800
rect 306746 -400 306802 800
rect 307298 -400 307354 800
rect 307850 -400 307906 800
rect 308402 -400 308458 800
rect 308954 -400 309010 800
rect 309506 -400 309562 800
rect 310058 -400 310114 800
rect 310610 -400 310666 800
rect 311162 -400 311218 800
rect 311714 -400 311770 800
rect 312266 -400 312322 800
rect 312818 -400 312874 800
rect 313370 -400 313426 800
rect 313922 -400 313978 800
rect 314474 -400 314530 800
rect 315026 -400 315082 800
rect 315578 -400 315634 800
rect 316130 -400 316186 800
rect 316682 -400 316738 800
rect 317234 -400 317290 800
rect 317786 -400 317842 800
rect 318338 -400 318394 800
rect 318890 -400 318946 800
rect 319442 -400 319498 800
rect 319994 -400 320050 800
rect 320546 -400 320602 800
rect 321098 -400 321154 800
rect 321650 -400 321706 800
rect 322202 -400 322258 800
rect 322754 -400 322810 800
rect 323306 -400 323362 800
rect 323858 -400 323914 800
rect 324410 -400 324466 800
rect 324962 -400 325018 800
rect 325514 -400 325570 800
rect 326066 -400 326122 800
rect 326618 -400 326674 800
rect 327170 -400 327226 800
rect 327722 -400 327778 800
rect 328274 -400 328330 800
rect 328826 -400 328882 800
rect 329378 -400 329434 800
rect 329930 -400 329986 800
rect 330482 -400 330538 800
rect 331034 -400 331090 800
rect 331586 -400 331642 800
rect 332138 -400 332194 800
rect 332690 -400 332746 800
rect 333242 -400 333298 800
rect 333794 -400 333850 800
rect 334346 -400 334402 800
rect 334898 -400 334954 800
rect 335450 -400 335506 800
rect 336002 -400 336058 800
rect 336554 -400 336610 800
rect 337106 -400 337162 800
rect 337658 -400 337714 800
rect 338210 -400 338266 800
rect 338762 -400 338818 800
rect 339314 -400 339370 800
rect 339866 -400 339922 800
rect 340418 -400 340474 800
rect 340970 -400 341026 800
rect 341522 -400 341578 800
rect 342074 -400 342130 800
rect 342626 -400 342682 800
rect 343178 -400 343234 800
rect 343730 -400 343786 800
rect 344282 -400 344338 800
rect 344834 -400 344890 800
rect 345386 -400 345442 800
rect 345938 -400 345994 800
rect 346490 -400 346546 800
rect 347042 -400 347098 800
rect 347594 -400 347650 800
rect 348146 -400 348202 800
rect 348698 -400 348754 800
rect 349250 -400 349306 800
rect 349802 -400 349858 800
rect 350354 -400 350410 800
rect 350906 -400 350962 800
rect 351458 -400 351514 800
rect 352010 -400 352066 800
rect 352562 -400 352618 800
rect 353114 -400 353170 800
rect 353666 -400 353722 800
rect 354218 -400 354274 800
rect 354770 -400 354826 800
rect 355322 -400 355378 800
rect 355874 -400 355930 800
rect 356426 -400 356482 800
rect 356978 -400 357034 800
rect 357530 -400 357586 800
rect 358082 -400 358138 800
rect 358634 -400 358690 800
rect 359186 -400 359242 800
rect 359738 -400 359794 800
rect 360290 -400 360346 800
rect 360842 -400 360898 800
rect 361394 -400 361450 800
rect 361946 -400 362002 800
rect 362498 -400 362554 800
<< obsm2 >>
rect 5036 27144 11554 27985
rect 11722 27144 12290 27985
rect 12458 27144 13026 27985
rect 13194 27144 13762 27985
rect 13930 27144 14498 27985
rect 14666 27144 15234 27985
rect 15402 27144 15970 27985
rect 16138 27144 16706 27985
rect 16874 27144 17442 27985
rect 17610 27144 18178 27985
rect 18346 27144 18914 27985
rect 19082 27144 19650 27985
rect 19818 27144 20386 27985
rect 20554 27144 21122 27985
rect 21290 27144 21858 27985
rect 22026 27144 22594 27985
rect 22762 27144 23330 27985
rect 23498 27144 24066 27985
rect 24234 27144 24802 27985
rect 24970 27144 25538 27985
rect 25706 27144 26274 27985
rect 26442 27144 27010 27985
rect 27178 27144 27746 27985
rect 27914 27144 28482 27985
rect 28650 27144 29218 27985
rect 29386 27144 29954 27985
rect 30122 27144 30690 27985
rect 30858 27144 31426 27985
rect 31594 27144 32162 27985
rect 32330 27144 32898 27985
rect 33066 27144 33634 27985
rect 33802 27144 34370 27985
rect 34538 27144 35106 27985
rect 35274 27144 35842 27985
rect 36010 27144 36578 27985
rect 36746 27144 37314 27985
rect 37482 27144 38050 27985
rect 38218 27144 38786 27985
rect 38954 27144 39522 27985
rect 39690 27144 40258 27985
rect 40426 27144 40994 27985
rect 41162 27144 41730 27985
rect 41898 27144 42466 27985
rect 42634 27144 43202 27985
rect 43370 27144 43938 27985
rect 44106 27144 44674 27985
rect 44842 27144 45410 27985
rect 45578 27144 46146 27985
rect 46314 27144 46882 27985
rect 47050 27144 47618 27985
rect 47786 27144 48354 27985
rect 48522 27144 49090 27985
rect 49258 27144 49826 27985
rect 49994 27144 50562 27985
rect 50730 27144 51298 27985
rect 51466 27144 52034 27985
rect 52202 27144 52770 27985
rect 52938 27144 53506 27985
rect 53674 27144 54242 27985
rect 54410 27144 54978 27985
rect 55146 27144 55714 27985
rect 55882 27144 56450 27985
rect 56618 27144 57186 27985
rect 57354 27144 57922 27985
rect 58090 27144 58658 27985
rect 58826 27144 59394 27985
rect 59562 27144 60130 27985
rect 60298 27144 60866 27985
rect 61034 27144 61602 27985
rect 61770 27144 62338 27985
rect 62506 27144 63074 27985
rect 63242 27144 63810 27985
rect 63978 27144 64546 27985
rect 64714 27144 65282 27985
rect 65450 27144 66018 27985
rect 66186 27144 66754 27985
rect 66922 27144 67490 27985
rect 67658 27144 68226 27985
rect 68394 27144 68962 27985
rect 69130 27144 69698 27985
rect 69866 27144 70434 27985
rect 70602 27144 71170 27985
rect 71338 27144 71906 27985
rect 72074 27144 72642 27985
rect 72810 27144 73378 27985
rect 73546 27144 74114 27985
rect 74282 27144 74850 27985
rect 75018 27144 75586 27985
rect 75754 27144 76322 27985
rect 76490 27144 77058 27985
rect 77226 27144 77794 27985
rect 77962 27144 78530 27985
rect 78698 27144 79266 27985
rect 79434 27144 80002 27985
rect 80170 27144 80738 27985
rect 80906 27144 81474 27985
rect 81642 27144 82210 27985
rect 82378 27144 82946 27985
rect 83114 27144 83682 27985
rect 83850 27144 84418 27985
rect 84586 27144 85154 27985
rect 85322 27144 85890 27985
rect 86058 27144 86626 27985
rect 86794 27144 87362 27985
rect 87530 27144 88098 27985
rect 88266 27144 88834 27985
rect 89002 27144 89570 27985
rect 89738 27144 90306 27985
rect 90474 27144 91042 27985
rect 91210 27144 91778 27985
rect 91946 27144 92514 27985
rect 92682 27144 93250 27985
rect 93418 27144 93986 27985
rect 94154 27144 94722 27985
rect 94890 27144 95458 27985
rect 95626 27144 96194 27985
rect 96362 27144 96930 27985
rect 97098 27144 97666 27985
rect 97834 27144 98402 27985
rect 98570 27144 99138 27985
rect 99306 27144 99874 27985
rect 100042 27144 100610 27985
rect 100778 27144 101346 27985
rect 101514 27144 102082 27985
rect 102250 27144 102818 27985
rect 102986 27144 103554 27985
rect 103722 27144 104290 27985
rect 104458 27144 105026 27985
rect 105194 27144 105762 27985
rect 105930 27144 106498 27985
rect 106666 27144 107234 27985
rect 107402 27144 107970 27985
rect 108138 27144 108706 27985
rect 108874 27144 109442 27985
rect 109610 27144 110178 27985
rect 110346 27144 110914 27985
rect 111082 27144 111650 27985
rect 111818 27144 112386 27985
rect 112554 27144 113122 27985
rect 113290 27144 113858 27985
rect 114026 27144 114594 27985
rect 114762 27144 115330 27985
rect 115498 27144 116066 27985
rect 116234 27144 116802 27985
rect 116970 27144 117538 27985
rect 117706 27144 118274 27985
rect 118442 27144 119010 27985
rect 119178 27144 119746 27985
rect 119914 27144 120482 27985
rect 120650 27144 121218 27985
rect 121386 27144 121954 27985
rect 122122 27144 122690 27985
rect 122858 27144 123426 27985
rect 123594 27144 124162 27985
rect 124330 27144 124898 27985
rect 125066 27144 125634 27985
rect 125802 27144 126370 27985
rect 126538 27144 127106 27985
rect 127274 27144 127842 27985
rect 128010 27144 128578 27985
rect 128746 27144 129314 27985
rect 129482 27144 130050 27985
rect 130218 27144 130786 27985
rect 130954 27144 131522 27985
rect 131690 27144 132258 27985
rect 132426 27144 132994 27985
rect 133162 27144 133730 27985
rect 133898 27144 134466 27985
rect 134634 27144 135202 27985
rect 135370 27144 135938 27985
rect 136106 27144 136674 27985
rect 136842 27144 137410 27985
rect 137578 27144 138146 27985
rect 138314 27144 138882 27985
rect 139050 27144 139618 27985
rect 139786 27144 140354 27985
rect 140522 27144 141090 27985
rect 141258 27144 141826 27985
rect 141994 27144 142562 27985
rect 142730 27144 143298 27985
rect 143466 27144 144034 27985
rect 144202 27144 144770 27985
rect 144938 27144 145506 27985
rect 145674 27144 146242 27985
rect 146410 27144 146978 27985
rect 147146 27144 147714 27985
rect 147882 27144 148450 27985
rect 148618 27144 149186 27985
rect 149354 27144 149922 27985
rect 150090 27144 150658 27985
rect 150826 27144 151394 27985
rect 151562 27144 152130 27985
rect 152298 27144 152866 27985
rect 153034 27144 153602 27985
rect 153770 27144 154338 27985
rect 154506 27144 155074 27985
rect 155242 27144 155810 27985
rect 155978 27144 156546 27985
rect 156714 27144 157282 27985
rect 157450 27144 158018 27985
rect 158186 27144 158754 27985
rect 158922 27144 159490 27985
rect 159658 27144 160226 27985
rect 160394 27144 160962 27985
rect 161130 27144 161698 27985
rect 161866 27144 162434 27985
rect 162602 27144 163170 27985
rect 163338 27144 163906 27985
rect 164074 27144 164642 27985
rect 164810 27144 165378 27985
rect 165546 27144 166114 27985
rect 166282 27144 166850 27985
rect 167018 27144 167586 27985
rect 167754 27144 168322 27985
rect 168490 27144 169058 27985
rect 169226 27144 169794 27985
rect 169962 27144 170530 27985
rect 170698 27144 171266 27985
rect 171434 27144 172002 27985
rect 172170 27144 172738 27985
rect 172906 27144 173474 27985
rect 173642 27144 174210 27985
rect 174378 27144 174946 27985
rect 175114 27144 175682 27985
rect 175850 27144 176418 27985
rect 176586 27144 177154 27985
rect 177322 27144 177890 27985
rect 178058 27144 178626 27985
rect 178794 27144 179362 27985
rect 179530 27144 180098 27985
rect 180266 27144 180834 27985
rect 181002 27144 181570 27985
rect 181738 27144 182306 27985
rect 182474 27144 183042 27985
rect 183210 27144 183778 27985
rect 183946 27144 184514 27985
rect 184682 27144 185250 27985
rect 185418 27144 185986 27985
rect 186154 27144 186722 27985
rect 186890 27144 187458 27985
rect 187626 27144 188194 27985
rect 188362 27144 188930 27985
rect 189098 27144 189666 27985
rect 189834 27144 190402 27985
rect 190570 27144 191138 27985
rect 191306 27144 191874 27985
rect 192042 27144 192610 27985
rect 192778 27144 193346 27985
rect 193514 27144 194082 27985
rect 194250 27144 194818 27985
rect 194986 27144 195554 27985
rect 195722 27144 196290 27985
rect 196458 27144 197026 27985
rect 197194 27144 197762 27985
rect 197930 27144 198498 27985
rect 198666 27144 199234 27985
rect 199402 27144 199970 27985
rect 200138 27144 200706 27985
rect 200874 27144 201442 27985
rect 201610 27144 202178 27985
rect 202346 27144 202914 27985
rect 203082 27144 203650 27985
rect 203818 27144 204386 27985
rect 204554 27144 205122 27985
rect 205290 27144 205858 27985
rect 206026 27144 206594 27985
rect 206762 27144 207330 27985
rect 207498 27144 208066 27985
rect 208234 27144 208802 27985
rect 208970 27144 209538 27985
rect 209706 27144 210274 27985
rect 210442 27144 211010 27985
rect 211178 27144 211746 27985
rect 211914 27144 212482 27985
rect 212650 27144 213218 27985
rect 213386 27144 213954 27985
rect 214122 27144 214690 27985
rect 214858 27144 215426 27985
rect 215594 27144 216162 27985
rect 216330 27144 216898 27985
rect 217066 27144 217634 27985
rect 217802 27144 218370 27985
rect 218538 27144 219106 27985
rect 219274 27144 219842 27985
rect 220010 27144 220578 27985
rect 220746 27144 221314 27985
rect 221482 27144 222050 27985
rect 222218 27144 222786 27985
rect 222954 27144 223522 27985
rect 223690 27144 224258 27985
rect 224426 27144 224994 27985
rect 225162 27144 225730 27985
rect 225898 27144 226466 27985
rect 226634 27144 227202 27985
rect 227370 27144 227938 27985
rect 228106 27144 228674 27985
rect 228842 27144 229410 27985
rect 229578 27144 230146 27985
rect 230314 27144 230882 27985
rect 231050 27144 231618 27985
rect 231786 27144 232354 27985
rect 232522 27144 233090 27985
rect 233258 27144 233826 27985
rect 233994 27144 234562 27985
rect 234730 27144 235298 27985
rect 235466 27144 236034 27985
rect 236202 27144 236770 27985
rect 236938 27144 237506 27985
rect 237674 27144 238242 27985
rect 238410 27144 238978 27985
rect 239146 27144 239714 27985
rect 239882 27144 240450 27985
rect 240618 27144 241186 27985
rect 241354 27144 241922 27985
rect 242090 27144 242658 27985
rect 242826 27144 243394 27985
rect 243562 27144 244130 27985
rect 244298 27144 244866 27985
rect 245034 27144 245602 27985
rect 245770 27144 246338 27985
rect 246506 27144 247074 27985
rect 247242 27144 247810 27985
rect 247978 27144 248546 27985
rect 248714 27144 249282 27985
rect 249450 27144 250018 27985
rect 250186 27144 250754 27985
rect 250922 27144 251490 27985
rect 251658 27144 252226 27985
rect 252394 27144 252962 27985
rect 253130 27144 253698 27985
rect 253866 27144 254434 27985
rect 254602 27144 255170 27985
rect 255338 27144 255906 27985
rect 256074 27144 256642 27985
rect 256810 27144 257378 27985
rect 257546 27144 258114 27985
rect 258282 27144 258850 27985
rect 259018 27144 259586 27985
rect 259754 27144 260322 27985
rect 260490 27144 261058 27985
rect 261226 27144 261794 27985
rect 261962 27144 262530 27985
rect 262698 27144 263266 27985
rect 263434 27144 264002 27985
rect 264170 27144 264738 27985
rect 264906 27144 265474 27985
rect 265642 27144 266210 27985
rect 266378 27144 266946 27985
rect 267114 27144 267682 27985
rect 267850 27144 268418 27985
rect 268586 27144 269154 27985
rect 269322 27144 269890 27985
rect 270058 27144 270626 27985
rect 270794 27144 271362 27985
rect 271530 27144 272098 27985
rect 272266 27144 272834 27985
rect 273002 27144 273570 27985
rect 273738 27144 274306 27985
rect 274474 27144 275042 27985
rect 275210 27144 275778 27985
rect 275946 27144 276514 27985
rect 276682 27144 277250 27985
rect 277418 27144 277986 27985
rect 278154 27144 278722 27985
rect 278890 27144 279458 27985
rect 279626 27144 280194 27985
rect 280362 27144 280930 27985
rect 281098 27144 281666 27985
rect 281834 27144 282402 27985
rect 282570 27144 283138 27985
rect 283306 27144 283874 27985
rect 284042 27144 284610 27985
rect 284778 27144 285346 27985
rect 285514 27144 286082 27985
rect 286250 27144 286818 27985
rect 286986 27144 287554 27985
rect 287722 27144 288290 27985
rect 288458 27144 289026 27985
rect 289194 27144 289762 27985
rect 289930 27144 290498 27985
rect 290666 27144 291234 27985
rect 291402 27144 291970 27985
rect 292138 27144 292706 27985
rect 292874 27144 293442 27985
rect 293610 27144 294178 27985
rect 294346 27144 294914 27985
rect 295082 27144 295650 27985
rect 295818 27144 296386 27985
rect 296554 27144 297122 27985
rect 297290 27144 297858 27985
rect 298026 27144 298594 27985
rect 298762 27144 299330 27985
rect 299498 27144 300066 27985
rect 300234 27144 300802 27985
rect 300970 27144 301538 27985
rect 301706 27144 302274 27985
rect 302442 27144 303010 27985
rect 303178 27144 303746 27985
rect 303914 27144 304482 27985
rect 304650 27144 305218 27985
rect 305386 27144 305954 27985
rect 306122 27144 306690 27985
rect 306858 27144 307426 27985
rect 307594 27144 308162 27985
rect 308330 27144 308898 27985
rect 309066 27144 309634 27985
rect 309802 27144 310370 27985
rect 310538 27144 311106 27985
rect 311274 27144 311842 27985
rect 312010 27144 312578 27985
rect 312746 27144 313314 27985
rect 313482 27144 314050 27985
rect 314218 27144 314786 27985
rect 314954 27144 315522 27985
rect 315690 27144 316258 27985
rect 316426 27144 316994 27985
rect 317162 27144 317730 27985
rect 317898 27144 318466 27985
rect 318634 27144 319202 27985
rect 319370 27144 319938 27985
rect 320106 27144 320674 27985
rect 320842 27144 321410 27985
rect 321578 27144 322146 27985
rect 322314 27144 322882 27985
rect 323050 27144 323618 27985
rect 323786 27144 324354 27985
rect 324522 27144 325090 27985
rect 325258 27144 325826 27985
rect 325994 27144 326562 27985
rect 326730 27144 327298 27985
rect 327466 27144 328034 27985
rect 328202 27144 328770 27985
rect 328938 27144 329506 27985
rect 329674 27144 330242 27985
rect 330410 27144 330978 27985
rect 331146 27144 331714 27985
rect 331882 27144 332450 27985
rect 332618 27144 333186 27985
rect 333354 27144 333922 27985
rect 334090 27144 334658 27985
rect 334826 27144 335394 27985
rect 335562 27144 336130 27985
rect 336298 27144 336866 27985
rect 337034 27144 337602 27985
rect 337770 27144 338338 27985
rect 338506 27144 339074 27985
rect 339242 27144 339810 27985
rect 339978 27144 340546 27985
rect 340714 27144 341282 27985
rect 341450 27144 342018 27985
rect 342186 27144 342754 27985
rect 342922 27144 343490 27985
rect 343658 27144 344226 27985
rect 344394 27144 344962 27985
rect 345130 27144 345698 27985
rect 345866 27144 346434 27985
rect 346602 27144 347170 27985
rect 347338 27144 347906 27985
rect 348074 27144 348642 27985
rect 348810 27144 349378 27985
rect 349546 27144 350114 27985
rect 350282 27144 350850 27985
rect 351018 27144 351586 27985
rect 351754 27144 352322 27985
rect 352490 27144 353058 27985
rect 353226 27144 353794 27985
rect 353962 27144 354530 27985
rect 354698 27144 355266 27985
rect 355434 27144 356002 27985
rect 356170 27144 356738 27985
rect 356906 27144 357474 27985
rect 357642 27144 358210 27985
rect 358378 27144 358946 27985
rect 359114 27144 359682 27985
rect 359850 27144 360418 27985
rect 360586 27144 361154 27985
rect 361322 27144 361890 27985
rect 362058 27144 362626 27985
rect 362794 27144 363362 27985
rect 363530 27144 364098 27985
rect 364266 27144 364834 27985
rect 365002 27144 365570 27985
rect 365738 27144 366306 27985
rect 366474 27144 367042 27985
rect 367210 27144 367778 27985
rect 367946 27144 368514 27985
rect 368682 27144 369250 27985
rect 369418 27144 369986 27985
rect 370154 27144 370722 27985
rect 370890 27144 371458 27985
rect 371626 27144 372194 27985
rect 372362 27144 382334 27985
rect 5036 856 382334 27144
rect 5036 2 21306 856
rect 21474 2 21858 856
rect 22026 2 22410 856
rect 22578 2 22962 856
rect 23130 2 23514 856
rect 23682 2 24066 856
rect 24234 2 24618 856
rect 24786 2 25170 856
rect 25338 2 25722 856
rect 25890 2 26274 856
rect 26442 2 26826 856
rect 26994 2 27378 856
rect 27546 2 27930 856
rect 28098 2 28482 856
rect 28650 2 29034 856
rect 29202 2 29586 856
rect 29754 2 30138 856
rect 30306 2 30690 856
rect 30858 2 31242 856
rect 31410 2 31794 856
rect 31962 2 32346 856
rect 32514 2 32898 856
rect 33066 2 33450 856
rect 33618 2 34002 856
rect 34170 2 34554 856
rect 34722 2 35106 856
rect 35274 2 35658 856
rect 35826 2 36210 856
rect 36378 2 36762 856
rect 36930 2 37314 856
rect 37482 2 37866 856
rect 38034 2 38418 856
rect 38586 2 38970 856
rect 39138 2 39522 856
rect 39690 2 40074 856
rect 40242 2 40626 856
rect 40794 2 41178 856
rect 41346 2 41730 856
rect 41898 2 42282 856
rect 42450 2 42834 856
rect 43002 2 43386 856
rect 43554 2 43938 856
rect 44106 2 44490 856
rect 44658 2 45042 856
rect 45210 2 45594 856
rect 45762 2 46146 856
rect 46314 2 46698 856
rect 46866 2 47250 856
rect 47418 2 47802 856
rect 47970 2 48354 856
rect 48522 2 48906 856
rect 49074 2 49458 856
rect 49626 2 50010 856
rect 50178 2 50562 856
rect 50730 2 51114 856
rect 51282 2 51666 856
rect 51834 2 52218 856
rect 52386 2 52770 856
rect 52938 2 53322 856
rect 53490 2 53874 856
rect 54042 2 54426 856
rect 54594 2 54978 856
rect 55146 2 55530 856
rect 55698 2 56082 856
rect 56250 2 56634 856
rect 56802 2 57186 856
rect 57354 2 57738 856
rect 57906 2 58290 856
rect 58458 2 58842 856
rect 59010 2 59394 856
rect 59562 2 59946 856
rect 60114 2 60498 856
rect 60666 2 61050 856
rect 61218 2 61602 856
rect 61770 2 62154 856
rect 62322 2 62706 856
rect 62874 2 63258 856
rect 63426 2 63810 856
rect 63978 2 64362 856
rect 64530 2 64914 856
rect 65082 2 65466 856
rect 65634 2 66018 856
rect 66186 2 66570 856
rect 66738 2 67122 856
rect 67290 2 67674 856
rect 67842 2 68226 856
rect 68394 2 68778 856
rect 68946 2 69330 856
rect 69498 2 69882 856
rect 70050 2 70434 856
rect 70602 2 70986 856
rect 71154 2 71538 856
rect 71706 2 72090 856
rect 72258 2 72642 856
rect 72810 2 73194 856
rect 73362 2 73746 856
rect 73914 2 74298 856
rect 74466 2 74850 856
rect 75018 2 75402 856
rect 75570 2 75954 856
rect 76122 2 76506 856
rect 76674 2 77058 856
rect 77226 2 77610 856
rect 77778 2 78162 856
rect 78330 2 78714 856
rect 78882 2 79266 856
rect 79434 2 79818 856
rect 79986 2 80370 856
rect 80538 2 80922 856
rect 81090 2 81474 856
rect 81642 2 82026 856
rect 82194 2 82578 856
rect 82746 2 83130 856
rect 83298 2 83682 856
rect 83850 2 84234 856
rect 84402 2 84786 856
rect 84954 2 85338 856
rect 85506 2 85890 856
rect 86058 2 86442 856
rect 86610 2 86994 856
rect 87162 2 87546 856
rect 87714 2 88098 856
rect 88266 2 88650 856
rect 88818 2 89202 856
rect 89370 2 89754 856
rect 89922 2 90306 856
rect 90474 2 90858 856
rect 91026 2 91410 856
rect 91578 2 91962 856
rect 92130 2 92514 856
rect 92682 2 93066 856
rect 93234 2 93618 856
rect 93786 2 94170 856
rect 94338 2 94722 856
rect 94890 2 95274 856
rect 95442 2 95826 856
rect 95994 2 96378 856
rect 96546 2 96930 856
rect 97098 2 97482 856
rect 97650 2 98034 856
rect 98202 2 98586 856
rect 98754 2 99138 856
rect 99306 2 99690 856
rect 99858 2 100242 856
rect 100410 2 100794 856
rect 100962 2 101346 856
rect 101514 2 101898 856
rect 102066 2 102450 856
rect 102618 2 103002 856
rect 103170 2 103554 856
rect 103722 2 104106 856
rect 104274 2 104658 856
rect 104826 2 105210 856
rect 105378 2 105762 856
rect 105930 2 106314 856
rect 106482 2 106866 856
rect 107034 2 107418 856
rect 107586 2 107970 856
rect 108138 2 108522 856
rect 108690 2 109074 856
rect 109242 2 109626 856
rect 109794 2 110178 856
rect 110346 2 110730 856
rect 110898 2 111282 856
rect 111450 2 111834 856
rect 112002 2 112386 856
rect 112554 2 112938 856
rect 113106 2 113490 856
rect 113658 2 114042 856
rect 114210 2 114594 856
rect 114762 2 115146 856
rect 115314 2 115698 856
rect 115866 2 116250 856
rect 116418 2 116802 856
rect 116970 2 117354 856
rect 117522 2 117906 856
rect 118074 2 118458 856
rect 118626 2 119010 856
rect 119178 2 119562 856
rect 119730 2 120114 856
rect 120282 2 120666 856
rect 120834 2 121218 856
rect 121386 2 121770 856
rect 121938 2 122322 856
rect 122490 2 122874 856
rect 123042 2 123426 856
rect 123594 2 123978 856
rect 124146 2 124530 856
rect 124698 2 125082 856
rect 125250 2 125634 856
rect 125802 2 126186 856
rect 126354 2 126738 856
rect 126906 2 127290 856
rect 127458 2 127842 856
rect 128010 2 128394 856
rect 128562 2 128946 856
rect 129114 2 129498 856
rect 129666 2 130050 856
rect 130218 2 130602 856
rect 130770 2 131154 856
rect 131322 2 131706 856
rect 131874 2 132258 856
rect 132426 2 132810 856
rect 132978 2 133362 856
rect 133530 2 133914 856
rect 134082 2 134466 856
rect 134634 2 135018 856
rect 135186 2 135570 856
rect 135738 2 136122 856
rect 136290 2 136674 856
rect 136842 2 137226 856
rect 137394 2 137778 856
rect 137946 2 138330 856
rect 138498 2 138882 856
rect 139050 2 139434 856
rect 139602 2 139986 856
rect 140154 2 140538 856
rect 140706 2 141090 856
rect 141258 2 141642 856
rect 141810 2 142194 856
rect 142362 2 142746 856
rect 142914 2 143298 856
rect 143466 2 143850 856
rect 144018 2 144402 856
rect 144570 2 144954 856
rect 145122 2 145506 856
rect 145674 2 146058 856
rect 146226 2 146610 856
rect 146778 2 147162 856
rect 147330 2 147714 856
rect 147882 2 148266 856
rect 148434 2 148818 856
rect 148986 2 149370 856
rect 149538 2 149922 856
rect 150090 2 150474 856
rect 150642 2 151026 856
rect 151194 2 151578 856
rect 151746 2 152130 856
rect 152298 2 152682 856
rect 152850 2 153234 856
rect 153402 2 153786 856
rect 153954 2 154338 856
rect 154506 2 154890 856
rect 155058 2 155442 856
rect 155610 2 155994 856
rect 156162 2 156546 856
rect 156714 2 157098 856
rect 157266 2 157650 856
rect 157818 2 158202 856
rect 158370 2 158754 856
rect 158922 2 159306 856
rect 159474 2 159858 856
rect 160026 2 160410 856
rect 160578 2 160962 856
rect 161130 2 161514 856
rect 161682 2 162066 856
rect 162234 2 162618 856
rect 162786 2 163170 856
rect 163338 2 163722 856
rect 163890 2 164274 856
rect 164442 2 164826 856
rect 164994 2 165378 856
rect 165546 2 165930 856
rect 166098 2 166482 856
rect 166650 2 167034 856
rect 167202 2 167586 856
rect 167754 2 168138 856
rect 168306 2 168690 856
rect 168858 2 169242 856
rect 169410 2 169794 856
rect 169962 2 170346 856
rect 170514 2 170898 856
rect 171066 2 171450 856
rect 171618 2 172002 856
rect 172170 2 172554 856
rect 172722 2 173106 856
rect 173274 2 173658 856
rect 173826 2 174210 856
rect 174378 2 174762 856
rect 174930 2 175314 856
rect 175482 2 175866 856
rect 176034 2 176418 856
rect 176586 2 176970 856
rect 177138 2 177522 856
rect 177690 2 178074 856
rect 178242 2 178626 856
rect 178794 2 179178 856
rect 179346 2 179730 856
rect 179898 2 180282 856
rect 180450 2 180834 856
rect 181002 2 181386 856
rect 181554 2 181938 856
rect 182106 2 182490 856
rect 182658 2 183042 856
rect 183210 2 183594 856
rect 183762 2 184146 856
rect 184314 2 184698 856
rect 184866 2 185250 856
rect 185418 2 185802 856
rect 185970 2 186354 856
rect 186522 2 186906 856
rect 187074 2 187458 856
rect 187626 2 188010 856
rect 188178 2 188562 856
rect 188730 2 189114 856
rect 189282 2 189666 856
rect 189834 2 190218 856
rect 190386 2 190770 856
rect 190938 2 191322 856
rect 191490 2 191874 856
rect 192042 2 192426 856
rect 192594 2 192978 856
rect 193146 2 193530 856
rect 193698 2 194082 856
rect 194250 2 194634 856
rect 194802 2 195186 856
rect 195354 2 195738 856
rect 195906 2 196290 856
rect 196458 2 196842 856
rect 197010 2 197394 856
rect 197562 2 197946 856
rect 198114 2 198498 856
rect 198666 2 199050 856
rect 199218 2 199602 856
rect 199770 2 200154 856
rect 200322 2 200706 856
rect 200874 2 201258 856
rect 201426 2 201810 856
rect 201978 2 202362 856
rect 202530 2 202914 856
rect 203082 2 203466 856
rect 203634 2 204018 856
rect 204186 2 204570 856
rect 204738 2 205122 856
rect 205290 2 205674 856
rect 205842 2 206226 856
rect 206394 2 206778 856
rect 206946 2 207330 856
rect 207498 2 207882 856
rect 208050 2 208434 856
rect 208602 2 208986 856
rect 209154 2 209538 856
rect 209706 2 210090 856
rect 210258 2 210642 856
rect 210810 2 211194 856
rect 211362 2 211746 856
rect 211914 2 212298 856
rect 212466 2 212850 856
rect 213018 2 213402 856
rect 213570 2 213954 856
rect 214122 2 214506 856
rect 214674 2 215058 856
rect 215226 2 215610 856
rect 215778 2 216162 856
rect 216330 2 216714 856
rect 216882 2 217266 856
rect 217434 2 217818 856
rect 217986 2 218370 856
rect 218538 2 218922 856
rect 219090 2 219474 856
rect 219642 2 220026 856
rect 220194 2 220578 856
rect 220746 2 221130 856
rect 221298 2 221682 856
rect 221850 2 222234 856
rect 222402 2 222786 856
rect 222954 2 223338 856
rect 223506 2 223890 856
rect 224058 2 224442 856
rect 224610 2 224994 856
rect 225162 2 225546 856
rect 225714 2 226098 856
rect 226266 2 226650 856
rect 226818 2 227202 856
rect 227370 2 227754 856
rect 227922 2 228306 856
rect 228474 2 228858 856
rect 229026 2 229410 856
rect 229578 2 229962 856
rect 230130 2 230514 856
rect 230682 2 231066 856
rect 231234 2 231618 856
rect 231786 2 232170 856
rect 232338 2 232722 856
rect 232890 2 233274 856
rect 233442 2 233826 856
rect 233994 2 234378 856
rect 234546 2 234930 856
rect 235098 2 235482 856
rect 235650 2 236034 856
rect 236202 2 236586 856
rect 236754 2 237138 856
rect 237306 2 237690 856
rect 237858 2 238242 856
rect 238410 2 238794 856
rect 238962 2 239346 856
rect 239514 2 239898 856
rect 240066 2 240450 856
rect 240618 2 241002 856
rect 241170 2 241554 856
rect 241722 2 242106 856
rect 242274 2 242658 856
rect 242826 2 243210 856
rect 243378 2 243762 856
rect 243930 2 244314 856
rect 244482 2 244866 856
rect 245034 2 245418 856
rect 245586 2 245970 856
rect 246138 2 246522 856
rect 246690 2 247074 856
rect 247242 2 247626 856
rect 247794 2 248178 856
rect 248346 2 248730 856
rect 248898 2 249282 856
rect 249450 2 249834 856
rect 250002 2 250386 856
rect 250554 2 250938 856
rect 251106 2 251490 856
rect 251658 2 252042 856
rect 252210 2 252594 856
rect 252762 2 253146 856
rect 253314 2 253698 856
rect 253866 2 254250 856
rect 254418 2 254802 856
rect 254970 2 255354 856
rect 255522 2 255906 856
rect 256074 2 256458 856
rect 256626 2 257010 856
rect 257178 2 257562 856
rect 257730 2 258114 856
rect 258282 2 258666 856
rect 258834 2 259218 856
rect 259386 2 259770 856
rect 259938 2 260322 856
rect 260490 2 260874 856
rect 261042 2 261426 856
rect 261594 2 261978 856
rect 262146 2 262530 856
rect 262698 2 263082 856
rect 263250 2 263634 856
rect 263802 2 264186 856
rect 264354 2 264738 856
rect 264906 2 265290 856
rect 265458 2 265842 856
rect 266010 2 266394 856
rect 266562 2 266946 856
rect 267114 2 267498 856
rect 267666 2 268050 856
rect 268218 2 268602 856
rect 268770 2 269154 856
rect 269322 2 269706 856
rect 269874 2 270258 856
rect 270426 2 270810 856
rect 270978 2 271362 856
rect 271530 2 271914 856
rect 272082 2 272466 856
rect 272634 2 273018 856
rect 273186 2 273570 856
rect 273738 2 274122 856
rect 274290 2 274674 856
rect 274842 2 275226 856
rect 275394 2 275778 856
rect 275946 2 276330 856
rect 276498 2 276882 856
rect 277050 2 277434 856
rect 277602 2 277986 856
rect 278154 2 278538 856
rect 278706 2 279090 856
rect 279258 2 279642 856
rect 279810 2 280194 856
rect 280362 2 280746 856
rect 280914 2 281298 856
rect 281466 2 281850 856
rect 282018 2 282402 856
rect 282570 2 282954 856
rect 283122 2 283506 856
rect 283674 2 284058 856
rect 284226 2 284610 856
rect 284778 2 285162 856
rect 285330 2 285714 856
rect 285882 2 286266 856
rect 286434 2 286818 856
rect 286986 2 287370 856
rect 287538 2 287922 856
rect 288090 2 288474 856
rect 288642 2 289026 856
rect 289194 2 289578 856
rect 289746 2 290130 856
rect 290298 2 290682 856
rect 290850 2 291234 856
rect 291402 2 291786 856
rect 291954 2 292338 856
rect 292506 2 292890 856
rect 293058 2 293442 856
rect 293610 2 293994 856
rect 294162 2 294546 856
rect 294714 2 295098 856
rect 295266 2 295650 856
rect 295818 2 296202 856
rect 296370 2 296754 856
rect 296922 2 297306 856
rect 297474 2 297858 856
rect 298026 2 298410 856
rect 298578 2 298962 856
rect 299130 2 299514 856
rect 299682 2 300066 856
rect 300234 2 300618 856
rect 300786 2 301170 856
rect 301338 2 301722 856
rect 301890 2 302274 856
rect 302442 2 302826 856
rect 302994 2 303378 856
rect 303546 2 303930 856
rect 304098 2 304482 856
rect 304650 2 305034 856
rect 305202 2 305586 856
rect 305754 2 306138 856
rect 306306 2 306690 856
rect 306858 2 307242 856
rect 307410 2 307794 856
rect 307962 2 308346 856
rect 308514 2 308898 856
rect 309066 2 309450 856
rect 309618 2 310002 856
rect 310170 2 310554 856
rect 310722 2 311106 856
rect 311274 2 311658 856
rect 311826 2 312210 856
rect 312378 2 312762 856
rect 312930 2 313314 856
rect 313482 2 313866 856
rect 314034 2 314418 856
rect 314586 2 314970 856
rect 315138 2 315522 856
rect 315690 2 316074 856
rect 316242 2 316626 856
rect 316794 2 317178 856
rect 317346 2 317730 856
rect 317898 2 318282 856
rect 318450 2 318834 856
rect 319002 2 319386 856
rect 319554 2 319938 856
rect 320106 2 320490 856
rect 320658 2 321042 856
rect 321210 2 321594 856
rect 321762 2 322146 856
rect 322314 2 322698 856
rect 322866 2 323250 856
rect 323418 2 323802 856
rect 323970 2 324354 856
rect 324522 2 324906 856
rect 325074 2 325458 856
rect 325626 2 326010 856
rect 326178 2 326562 856
rect 326730 2 327114 856
rect 327282 2 327666 856
rect 327834 2 328218 856
rect 328386 2 328770 856
rect 328938 2 329322 856
rect 329490 2 329874 856
rect 330042 2 330426 856
rect 330594 2 330978 856
rect 331146 2 331530 856
rect 331698 2 332082 856
rect 332250 2 332634 856
rect 332802 2 333186 856
rect 333354 2 333738 856
rect 333906 2 334290 856
rect 334458 2 334842 856
rect 335010 2 335394 856
rect 335562 2 335946 856
rect 336114 2 336498 856
rect 336666 2 337050 856
rect 337218 2 337602 856
rect 337770 2 338154 856
rect 338322 2 338706 856
rect 338874 2 339258 856
rect 339426 2 339810 856
rect 339978 2 340362 856
rect 340530 2 340914 856
rect 341082 2 341466 856
rect 341634 2 342018 856
rect 342186 2 342570 856
rect 342738 2 343122 856
rect 343290 2 343674 856
rect 343842 2 344226 856
rect 344394 2 344778 856
rect 344946 2 345330 856
rect 345498 2 345882 856
rect 346050 2 346434 856
rect 346602 2 346986 856
rect 347154 2 347538 856
rect 347706 2 348090 856
rect 348258 2 348642 856
rect 348810 2 349194 856
rect 349362 2 349746 856
rect 349914 2 350298 856
rect 350466 2 350850 856
rect 351018 2 351402 856
rect 351570 2 351954 856
rect 352122 2 352506 856
rect 352674 2 353058 856
rect 353226 2 353610 856
rect 353778 2 354162 856
rect 354330 2 354714 856
rect 354882 2 355266 856
rect 355434 2 355818 856
rect 355986 2 356370 856
rect 356538 2 356922 856
rect 357090 2 357474 856
rect 357642 2 358026 856
rect 358194 2 358578 856
rect 358746 2 359130 856
rect 359298 2 359682 856
rect 359850 2 360234 856
rect 360402 2 360786 856
rect 360954 2 361338 856
rect 361506 2 361890 856
rect 362058 2 362442 856
rect 362610 2 382334 856
<< metal3 >>
rect 383200 26256 384400 26376
rect 383200 24352 384400 24472
rect 383200 22448 384400 22568
rect 383200 20544 384400 20664
rect 383200 18640 384400 18760
rect 383200 16736 384400 16856
rect 383200 14832 384400 14952
rect 383200 12928 384400 13048
rect 383200 11024 384400 11144
rect 383200 9120 384400 9240
rect 383200 7216 384400 7336
rect 383200 5312 384400 5432
rect 383200 3408 384400 3528
rect 383200 1504 384400 1624
<< obsm3 >>
rect 5026 26456 383200 27981
rect 5026 26176 383120 26456
rect 5026 24552 383200 26176
rect 5026 24272 383120 24552
rect 5026 22648 383200 24272
rect 5026 22368 383120 22648
rect 5026 20744 383200 22368
rect 5026 20464 383120 20744
rect 5026 18840 383200 20464
rect 5026 18560 383120 18840
rect 5026 16936 383200 18560
rect 5026 16656 383120 16936
rect 5026 15032 383200 16656
rect 5026 14752 383120 15032
rect 5026 13128 383200 14752
rect 5026 12848 383120 13128
rect 5026 11224 383200 12848
rect 5026 10944 383120 11224
rect 5026 9320 383200 10944
rect 5026 9040 383120 9320
rect 5026 7416 383200 9040
rect 5026 7136 383120 7416
rect 5026 5512 383200 7136
rect 5026 5232 383120 5512
rect 5026 3608 383200 5232
rect 5026 3328 383120 3608
rect 5026 1704 383200 3328
rect 5026 1424 383120 1704
rect 5026 35 383200 1424
<< metal4 >>
rect 5014 1040 5194 26704
rect 12394 1040 12574 26704
rect 20064 1040 20244 26704
rect 27444 1040 27624 26704
rect 35114 1040 35294 26704
rect 42494 1040 42674 26704
rect 50164 1040 50344 26704
rect 57544 1040 57724 26704
rect 65214 1040 65394 26704
rect 66854 1040 67034 26704
rect 71034 1040 71214 26704
rect 72594 1040 72774 26704
rect 76854 1040 77034 26704
rect 80264 1040 80444 26704
rect 81034 1040 81214 26704
rect 87644 1040 87824 26704
rect 95314 1040 95494 26704
rect 102694 1040 102874 26704
rect 110364 1040 110544 26704
rect 117744 1040 117924 26704
rect 125414 1040 125594 26704
rect 132794 1040 132974 26704
rect 140464 1040 140644 26704
rect 141284 1040 141464 26704
rect 147844 1040 148024 26704
rect 148664 1040 148844 26704
rect 155514 1040 155694 26704
rect 156334 1040 156514 26704
rect 162894 1040 163074 26704
rect 163714 1040 163894 26704
rect 170564 1040 170744 26704
rect 171384 1040 171564 26704
rect 177944 1040 178124 26704
rect 178764 1040 178944 26704
rect 185614 1040 185794 26704
rect 186434 1040 186614 26704
rect 192994 1040 193174 26704
rect 193814 1040 193994 26704
rect 200664 1040 200844 26704
rect 208044 1040 208224 26704
rect 215714 1040 215894 26704
rect 223094 1040 223274 26704
rect 230764 1040 230944 26704
rect 238144 1040 238324 26704
rect 245814 1040 245994 26704
rect 253194 1040 253374 26704
rect 255814 1040 255994 26704
rect 256614 1040 256794 26704
rect 260864 1040 261044 26704
rect 263194 1040 263374 26704
rect 263994 1040 264174 26704
rect 268244 1040 268424 26704
rect 270864 1040 271044 26704
rect 271664 1040 271844 26704
rect 275914 1040 276094 26704
rect 278244 1040 278424 26704
rect 279044 1040 279224 26704
rect 283294 1040 283474 26704
rect 290964 1040 291144 26704
rect 298344 1040 298524 26704
rect 306014 1040 306194 26704
rect 313394 1040 313574 26704
rect 321064 1040 321244 26704
rect 328444 1040 328624 26704
rect 336114 1040 336294 26704
rect 343494 1040 343674 26704
rect 351164 1040 351344 26704
rect 358544 1040 358724 26704
rect 366214 1040 366394 26704
rect 373594 1040 373774 26704
rect 381264 1040 381444 26704
<< obsm4 >>
rect 68323 26784 305749 27981
rect 68323 960 70954 26784
rect 71294 960 72514 26784
rect 72854 960 76774 26784
rect 77114 960 80184 26784
rect 80524 960 80954 26784
rect 81294 960 87564 26784
rect 87904 960 95234 26784
rect 95574 960 102614 26784
rect 102954 960 110284 26784
rect 110624 960 117664 26784
rect 118004 960 125334 26784
rect 125674 960 132714 26784
rect 133054 960 140384 26784
rect 140724 960 141204 26784
rect 141544 960 147764 26784
rect 148104 960 148584 26784
rect 148924 960 155434 26784
rect 155774 960 156254 26784
rect 156594 960 162814 26784
rect 163154 960 163634 26784
rect 163974 960 170484 26784
rect 170824 960 171304 26784
rect 171644 960 177864 26784
rect 178204 960 178684 26784
rect 179024 960 185534 26784
rect 185874 960 186354 26784
rect 186694 960 192914 26784
rect 193254 960 193734 26784
rect 194074 960 200584 26784
rect 200924 960 207964 26784
rect 208304 960 215634 26784
rect 215974 960 223014 26784
rect 223354 960 230684 26784
rect 231024 960 238064 26784
rect 238404 960 245734 26784
rect 246074 960 253114 26784
rect 253454 960 255734 26784
rect 256074 960 256534 26784
rect 256874 960 260784 26784
rect 261124 960 263114 26784
rect 263454 960 263914 26784
rect 264254 960 268164 26784
rect 268504 960 270784 26784
rect 271124 960 271584 26784
rect 271924 960 275834 26784
rect 276174 960 278164 26784
rect 278504 960 278964 26784
rect 279304 960 283214 26784
rect 283554 960 290884 26784
rect 291224 960 298264 26784
rect 298604 960 305749 26784
rect 68323 35 305749 960
<< labels >>
rlabel metal2 s 178130 -400 178186 800 6 caravel_clk
port 1 nsew signal input
rlabel metal3 s 383200 7216 384400 7336 6 caravel_clk2
port 2 nsew signal input
rlabel metal2 s 178682 -400 178738 800 6 caravel_rstn
port 3 nsew signal input
rlabel metal2 s 89626 27200 89682 28400 6 la_data_in_core[0]
port 4 nsew signal output
rlabel metal2 s 310426 27200 310482 28400 6 la_data_in_core[100]
port 5 nsew signal output
rlabel metal2 s 312634 27200 312690 28400 6 la_data_in_core[101]
port 6 nsew signal output
rlabel metal2 s 314842 27200 314898 28400 6 la_data_in_core[102]
port 7 nsew signal output
rlabel metal2 s 317050 27200 317106 28400 6 la_data_in_core[103]
port 8 nsew signal output
rlabel metal2 s 319258 27200 319314 28400 6 la_data_in_core[104]
port 9 nsew signal output
rlabel metal2 s 321466 27200 321522 28400 6 la_data_in_core[105]
port 10 nsew signal output
rlabel metal2 s 323674 27200 323730 28400 6 la_data_in_core[106]
port 11 nsew signal output
rlabel metal2 s 325882 27200 325938 28400 6 la_data_in_core[107]
port 12 nsew signal output
rlabel metal2 s 328090 27200 328146 28400 6 la_data_in_core[108]
port 13 nsew signal output
rlabel metal2 s 330298 27200 330354 28400 6 la_data_in_core[109]
port 14 nsew signal output
rlabel metal2 s 111706 27200 111762 28400 6 la_data_in_core[10]
port 15 nsew signal output
rlabel metal2 s 332506 27200 332562 28400 6 la_data_in_core[110]
port 16 nsew signal output
rlabel metal2 s 334714 27200 334770 28400 6 la_data_in_core[111]
port 17 nsew signal output
rlabel metal2 s 336922 27200 336978 28400 6 la_data_in_core[112]
port 18 nsew signal output
rlabel metal2 s 339130 27200 339186 28400 6 la_data_in_core[113]
port 19 nsew signal output
rlabel metal2 s 341338 27200 341394 28400 6 la_data_in_core[114]
port 20 nsew signal output
rlabel metal2 s 343546 27200 343602 28400 6 la_data_in_core[115]
port 21 nsew signal output
rlabel metal2 s 345754 27200 345810 28400 6 la_data_in_core[116]
port 22 nsew signal output
rlabel metal2 s 347962 27200 348018 28400 6 la_data_in_core[117]
port 23 nsew signal output
rlabel metal2 s 350170 27200 350226 28400 6 la_data_in_core[118]
port 24 nsew signal output
rlabel metal2 s 352378 27200 352434 28400 6 la_data_in_core[119]
port 25 nsew signal output
rlabel metal2 s 113914 27200 113970 28400 6 la_data_in_core[11]
port 26 nsew signal output
rlabel metal2 s 354586 27200 354642 28400 6 la_data_in_core[120]
port 27 nsew signal output
rlabel metal2 s 356794 27200 356850 28400 6 la_data_in_core[121]
port 28 nsew signal output
rlabel metal2 s 359002 27200 359058 28400 6 la_data_in_core[122]
port 29 nsew signal output
rlabel metal2 s 361210 27200 361266 28400 6 la_data_in_core[123]
port 30 nsew signal output
rlabel metal2 s 363418 27200 363474 28400 6 la_data_in_core[124]
port 31 nsew signal output
rlabel metal2 s 365626 27200 365682 28400 6 la_data_in_core[125]
port 32 nsew signal output
rlabel metal2 s 367834 27200 367890 28400 6 la_data_in_core[126]
port 33 nsew signal output
rlabel metal2 s 370042 27200 370098 28400 6 la_data_in_core[127]
port 34 nsew signal output
rlabel metal2 s 116122 27200 116178 28400 6 la_data_in_core[12]
port 35 nsew signal output
rlabel metal2 s 118330 27200 118386 28400 6 la_data_in_core[13]
port 36 nsew signal output
rlabel metal2 s 120538 27200 120594 28400 6 la_data_in_core[14]
port 37 nsew signal output
rlabel metal2 s 122746 27200 122802 28400 6 la_data_in_core[15]
port 38 nsew signal output
rlabel metal2 s 124954 27200 125010 28400 6 la_data_in_core[16]
port 39 nsew signal output
rlabel metal2 s 127162 27200 127218 28400 6 la_data_in_core[17]
port 40 nsew signal output
rlabel metal2 s 129370 27200 129426 28400 6 la_data_in_core[18]
port 41 nsew signal output
rlabel metal2 s 131578 27200 131634 28400 6 la_data_in_core[19]
port 42 nsew signal output
rlabel metal2 s 91834 27200 91890 28400 6 la_data_in_core[1]
port 43 nsew signal output
rlabel metal2 s 133786 27200 133842 28400 6 la_data_in_core[20]
port 44 nsew signal output
rlabel metal2 s 135994 27200 136050 28400 6 la_data_in_core[21]
port 45 nsew signal output
rlabel metal2 s 138202 27200 138258 28400 6 la_data_in_core[22]
port 46 nsew signal output
rlabel metal2 s 140410 27200 140466 28400 6 la_data_in_core[23]
port 47 nsew signal output
rlabel metal2 s 142618 27200 142674 28400 6 la_data_in_core[24]
port 48 nsew signal output
rlabel metal2 s 144826 27200 144882 28400 6 la_data_in_core[25]
port 49 nsew signal output
rlabel metal2 s 147034 27200 147090 28400 6 la_data_in_core[26]
port 50 nsew signal output
rlabel metal2 s 149242 27200 149298 28400 6 la_data_in_core[27]
port 51 nsew signal output
rlabel metal2 s 151450 27200 151506 28400 6 la_data_in_core[28]
port 52 nsew signal output
rlabel metal2 s 153658 27200 153714 28400 6 la_data_in_core[29]
port 53 nsew signal output
rlabel metal2 s 94042 27200 94098 28400 6 la_data_in_core[2]
port 54 nsew signal output
rlabel metal2 s 155866 27200 155922 28400 6 la_data_in_core[30]
port 55 nsew signal output
rlabel metal2 s 158074 27200 158130 28400 6 la_data_in_core[31]
port 56 nsew signal output
rlabel metal2 s 160282 27200 160338 28400 6 la_data_in_core[32]
port 57 nsew signal output
rlabel metal2 s 162490 27200 162546 28400 6 la_data_in_core[33]
port 58 nsew signal output
rlabel metal2 s 164698 27200 164754 28400 6 la_data_in_core[34]
port 59 nsew signal output
rlabel metal2 s 166906 27200 166962 28400 6 la_data_in_core[35]
port 60 nsew signal output
rlabel metal2 s 169114 27200 169170 28400 6 la_data_in_core[36]
port 61 nsew signal output
rlabel metal2 s 171322 27200 171378 28400 6 la_data_in_core[37]
port 62 nsew signal output
rlabel metal2 s 173530 27200 173586 28400 6 la_data_in_core[38]
port 63 nsew signal output
rlabel metal2 s 175738 27200 175794 28400 6 la_data_in_core[39]
port 64 nsew signal output
rlabel metal2 s 96250 27200 96306 28400 6 la_data_in_core[3]
port 65 nsew signal output
rlabel metal2 s 177946 27200 178002 28400 6 la_data_in_core[40]
port 66 nsew signal output
rlabel metal2 s 180154 27200 180210 28400 6 la_data_in_core[41]
port 67 nsew signal output
rlabel metal2 s 182362 27200 182418 28400 6 la_data_in_core[42]
port 68 nsew signal output
rlabel metal2 s 184570 27200 184626 28400 6 la_data_in_core[43]
port 69 nsew signal output
rlabel metal2 s 186778 27200 186834 28400 6 la_data_in_core[44]
port 70 nsew signal output
rlabel metal2 s 188986 27200 189042 28400 6 la_data_in_core[45]
port 71 nsew signal output
rlabel metal2 s 191194 27200 191250 28400 6 la_data_in_core[46]
port 72 nsew signal output
rlabel metal2 s 193402 27200 193458 28400 6 la_data_in_core[47]
port 73 nsew signal output
rlabel metal2 s 195610 27200 195666 28400 6 la_data_in_core[48]
port 74 nsew signal output
rlabel metal2 s 197818 27200 197874 28400 6 la_data_in_core[49]
port 75 nsew signal output
rlabel metal2 s 98458 27200 98514 28400 6 la_data_in_core[4]
port 76 nsew signal output
rlabel metal2 s 200026 27200 200082 28400 6 la_data_in_core[50]
port 77 nsew signal output
rlabel metal2 s 202234 27200 202290 28400 6 la_data_in_core[51]
port 78 nsew signal output
rlabel metal2 s 204442 27200 204498 28400 6 la_data_in_core[52]
port 79 nsew signal output
rlabel metal2 s 206650 27200 206706 28400 6 la_data_in_core[53]
port 80 nsew signal output
rlabel metal2 s 208858 27200 208914 28400 6 la_data_in_core[54]
port 81 nsew signal output
rlabel metal2 s 211066 27200 211122 28400 6 la_data_in_core[55]
port 82 nsew signal output
rlabel metal2 s 213274 27200 213330 28400 6 la_data_in_core[56]
port 83 nsew signal output
rlabel metal2 s 215482 27200 215538 28400 6 la_data_in_core[57]
port 84 nsew signal output
rlabel metal2 s 217690 27200 217746 28400 6 la_data_in_core[58]
port 85 nsew signal output
rlabel metal2 s 219898 27200 219954 28400 6 la_data_in_core[59]
port 86 nsew signal output
rlabel metal2 s 100666 27200 100722 28400 6 la_data_in_core[5]
port 87 nsew signal output
rlabel metal2 s 222106 27200 222162 28400 6 la_data_in_core[60]
port 88 nsew signal output
rlabel metal2 s 224314 27200 224370 28400 6 la_data_in_core[61]
port 89 nsew signal output
rlabel metal2 s 226522 27200 226578 28400 6 la_data_in_core[62]
port 90 nsew signal output
rlabel metal2 s 228730 27200 228786 28400 6 la_data_in_core[63]
port 91 nsew signal output
rlabel metal2 s 230938 27200 230994 28400 6 la_data_in_core[64]
port 92 nsew signal output
rlabel metal2 s 233146 27200 233202 28400 6 la_data_in_core[65]
port 93 nsew signal output
rlabel metal2 s 235354 27200 235410 28400 6 la_data_in_core[66]
port 94 nsew signal output
rlabel metal2 s 237562 27200 237618 28400 6 la_data_in_core[67]
port 95 nsew signal output
rlabel metal2 s 239770 27200 239826 28400 6 la_data_in_core[68]
port 96 nsew signal output
rlabel metal2 s 241978 27200 242034 28400 6 la_data_in_core[69]
port 97 nsew signal output
rlabel metal2 s 102874 27200 102930 28400 6 la_data_in_core[6]
port 98 nsew signal output
rlabel metal2 s 244186 27200 244242 28400 6 la_data_in_core[70]
port 99 nsew signal output
rlabel metal2 s 246394 27200 246450 28400 6 la_data_in_core[71]
port 100 nsew signal output
rlabel metal2 s 248602 27200 248658 28400 6 la_data_in_core[72]
port 101 nsew signal output
rlabel metal2 s 250810 27200 250866 28400 6 la_data_in_core[73]
port 102 nsew signal output
rlabel metal2 s 253018 27200 253074 28400 6 la_data_in_core[74]
port 103 nsew signal output
rlabel metal2 s 255226 27200 255282 28400 6 la_data_in_core[75]
port 104 nsew signal output
rlabel metal2 s 257434 27200 257490 28400 6 la_data_in_core[76]
port 105 nsew signal output
rlabel metal2 s 259642 27200 259698 28400 6 la_data_in_core[77]
port 106 nsew signal output
rlabel metal2 s 261850 27200 261906 28400 6 la_data_in_core[78]
port 107 nsew signal output
rlabel metal2 s 264058 27200 264114 28400 6 la_data_in_core[79]
port 108 nsew signal output
rlabel metal2 s 105082 27200 105138 28400 6 la_data_in_core[7]
port 109 nsew signal output
rlabel metal2 s 266266 27200 266322 28400 6 la_data_in_core[80]
port 110 nsew signal output
rlabel metal2 s 268474 27200 268530 28400 6 la_data_in_core[81]
port 111 nsew signal output
rlabel metal2 s 270682 27200 270738 28400 6 la_data_in_core[82]
port 112 nsew signal output
rlabel metal2 s 272890 27200 272946 28400 6 la_data_in_core[83]
port 113 nsew signal output
rlabel metal2 s 275098 27200 275154 28400 6 la_data_in_core[84]
port 114 nsew signal output
rlabel metal2 s 277306 27200 277362 28400 6 la_data_in_core[85]
port 115 nsew signal output
rlabel metal2 s 279514 27200 279570 28400 6 la_data_in_core[86]
port 116 nsew signal output
rlabel metal2 s 281722 27200 281778 28400 6 la_data_in_core[87]
port 117 nsew signal output
rlabel metal2 s 283930 27200 283986 28400 6 la_data_in_core[88]
port 118 nsew signal output
rlabel metal2 s 286138 27200 286194 28400 6 la_data_in_core[89]
port 119 nsew signal output
rlabel metal2 s 107290 27200 107346 28400 6 la_data_in_core[8]
port 120 nsew signal output
rlabel metal2 s 288346 27200 288402 28400 6 la_data_in_core[90]
port 121 nsew signal output
rlabel metal2 s 290554 27200 290610 28400 6 la_data_in_core[91]
port 122 nsew signal output
rlabel metal2 s 292762 27200 292818 28400 6 la_data_in_core[92]
port 123 nsew signal output
rlabel metal2 s 294970 27200 295026 28400 6 la_data_in_core[93]
port 124 nsew signal output
rlabel metal2 s 297178 27200 297234 28400 6 la_data_in_core[94]
port 125 nsew signal output
rlabel metal2 s 299386 27200 299442 28400 6 la_data_in_core[95]
port 126 nsew signal output
rlabel metal2 s 301594 27200 301650 28400 6 la_data_in_core[96]
port 127 nsew signal output
rlabel metal2 s 303802 27200 303858 28400 6 la_data_in_core[97]
port 128 nsew signal output
rlabel metal2 s 306010 27200 306066 28400 6 la_data_in_core[98]
port 129 nsew signal output
rlabel metal2 s 308218 27200 308274 28400 6 la_data_in_core[99]
port 130 nsew signal output
rlabel metal2 s 109498 27200 109554 28400 6 la_data_in_core[9]
port 131 nsew signal output
rlabel metal2 s 21362 -400 21418 800 6 la_data_in_mprj[0]
port 132 nsew signal output
rlabel metal2 s 243266 -400 243322 800 6 la_data_in_mprj[100]
port 133 nsew signal output
rlabel metal2 s 245474 -400 245530 800 6 la_data_in_mprj[101]
port 134 nsew signal output
rlabel metal2 s 247682 -400 247738 800 6 la_data_in_mprj[102]
port 135 nsew signal output
rlabel metal2 s 249890 -400 249946 800 6 la_data_in_mprj[103]
port 136 nsew signal output
rlabel metal2 s 252098 -400 252154 800 6 la_data_in_mprj[104]
port 137 nsew signal output
rlabel metal2 s 254306 -400 254362 800 6 la_data_in_mprj[105]
port 138 nsew signal output
rlabel metal2 s 256514 -400 256570 800 6 la_data_in_mprj[106]
port 139 nsew signal output
rlabel metal2 s 258722 -400 258778 800 6 la_data_in_mprj[107]
port 140 nsew signal output
rlabel metal2 s 260930 -400 260986 800 6 la_data_in_mprj[108]
port 141 nsew signal output
rlabel metal2 s 263138 -400 263194 800 6 la_data_in_mprj[109]
port 142 nsew signal output
rlabel metal2 s 43442 -400 43498 800 6 la_data_in_mprj[10]
port 143 nsew signal output
rlabel metal2 s 265346 -400 265402 800 6 la_data_in_mprj[110]
port 144 nsew signal output
rlabel metal2 s 267554 -400 267610 800 6 la_data_in_mprj[111]
port 145 nsew signal output
rlabel metal2 s 269762 -400 269818 800 6 la_data_in_mprj[112]
port 146 nsew signal output
rlabel metal2 s 271970 -400 272026 800 6 la_data_in_mprj[113]
port 147 nsew signal output
rlabel metal2 s 274178 -400 274234 800 6 la_data_in_mprj[114]
port 148 nsew signal output
rlabel metal2 s 276386 -400 276442 800 6 la_data_in_mprj[115]
port 149 nsew signal output
rlabel metal2 s 278594 -400 278650 800 6 la_data_in_mprj[116]
port 150 nsew signal output
rlabel metal2 s 280802 -400 280858 800 6 la_data_in_mprj[117]
port 151 nsew signal output
rlabel metal2 s 283010 -400 283066 800 6 la_data_in_mprj[118]
port 152 nsew signal output
rlabel metal2 s 285218 -400 285274 800 6 la_data_in_mprj[119]
port 153 nsew signal output
rlabel metal2 s 45650 -400 45706 800 6 la_data_in_mprj[11]
port 154 nsew signal output
rlabel metal2 s 287426 -400 287482 800 6 la_data_in_mprj[120]
port 155 nsew signal output
rlabel metal2 s 289634 -400 289690 800 6 la_data_in_mprj[121]
port 156 nsew signal output
rlabel metal2 s 291842 -400 291898 800 6 la_data_in_mprj[122]
port 157 nsew signal output
rlabel metal2 s 294050 -400 294106 800 6 la_data_in_mprj[123]
port 158 nsew signal output
rlabel metal2 s 296258 -400 296314 800 6 la_data_in_mprj[124]
port 159 nsew signal output
rlabel metal2 s 298466 -400 298522 800 6 la_data_in_mprj[125]
port 160 nsew signal output
rlabel metal2 s 300674 -400 300730 800 6 la_data_in_mprj[126]
port 161 nsew signal output
rlabel metal2 s 302882 -400 302938 800 6 la_data_in_mprj[127]
port 162 nsew signal output
rlabel metal2 s 47858 -400 47914 800 6 la_data_in_mprj[12]
port 163 nsew signal output
rlabel metal2 s 50066 -400 50122 800 6 la_data_in_mprj[13]
port 164 nsew signal output
rlabel metal2 s 52274 -400 52330 800 6 la_data_in_mprj[14]
port 165 nsew signal output
rlabel metal2 s 54482 -400 54538 800 6 la_data_in_mprj[15]
port 166 nsew signal output
rlabel metal2 s 56690 -400 56746 800 6 la_data_in_mprj[16]
port 167 nsew signal output
rlabel metal2 s 58898 -400 58954 800 6 la_data_in_mprj[17]
port 168 nsew signal output
rlabel metal2 s 61106 -400 61162 800 6 la_data_in_mprj[18]
port 169 nsew signal output
rlabel metal2 s 63314 -400 63370 800 6 la_data_in_mprj[19]
port 170 nsew signal output
rlabel metal2 s 23570 -400 23626 800 6 la_data_in_mprj[1]
port 171 nsew signal output
rlabel metal2 s 65522 -400 65578 800 6 la_data_in_mprj[20]
port 172 nsew signal output
rlabel metal2 s 67730 -400 67786 800 6 la_data_in_mprj[21]
port 173 nsew signal output
rlabel metal2 s 69938 -400 69994 800 6 la_data_in_mprj[22]
port 174 nsew signal output
rlabel metal2 s 72146 -400 72202 800 6 la_data_in_mprj[23]
port 175 nsew signal output
rlabel metal2 s 74354 -400 74410 800 6 la_data_in_mprj[24]
port 176 nsew signal output
rlabel metal2 s 76562 -400 76618 800 6 la_data_in_mprj[25]
port 177 nsew signal output
rlabel metal2 s 78770 -400 78826 800 6 la_data_in_mprj[26]
port 178 nsew signal output
rlabel metal2 s 80978 -400 81034 800 6 la_data_in_mprj[27]
port 179 nsew signal output
rlabel metal2 s 83186 -400 83242 800 6 la_data_in_mprj[28]
port 180 nsew signal output
rlabel metal2 s 85394 -400 85450 800 6 la_data_in_mprj[29]
port 181 nsew signal output
rlabel metal2 s 25778 -400 25834 800 6 la_data_in_mprj[2]
port 182 nsew signal output
rlabel metal2 s 87602 -400 87658 800 6 la_data_in_mprj[30]
port 183 nsew signal output
rlabel metal2 s 89810 -400 89866 800 6 la_data_in_mprj[31]
port 184 nsew signal output
rlabel metal2 s 92018 -400 92074 800 6 la_data_in_mprj[32]
port 185 nsew signal output
rlabel metal2 s 94226 -400 94282 800 6 la_data_in_mprj[33]
port 186 nsew signal output
rlabel metal2 s 96434 -400 96490 800 6 la_data_in_mprj[34]
port 187 nsew signal output
rlabel metal2 s 98642 -400 98698 800 6 la_data_in_mprj[35]
port 188 nsew signal output
rlabel metal2 s 100850 -400 100906 800 6 la_data_in_mprj[36]
port 189 nsew signal output
rlabel metal2 s 103058 -400 103114 800 6 la_data_in_mprj[37]
port 190 nsew signal output
rlabel metal2 s 105266 -400 105322 800 6 la_data_in_mprj[38]
port 191 nsew signal output
rlabel metal2 s 107474 -400 107530 800 6 la_data_in_mprj[39]
port 192 nsew signal output
rlabel metal2 s 27986 -400 28042 800 6 la_data_in_mprj[3]
port 193 nsew signal output
rlabel metal2 s 109682 -400 109738 800 6 la_data_in_mprj[40]
port 194 nsew signal output
rlabel metal2 s 111890 -400 111946 800 6 la_data_in_mprj[41]
port 195 nsew signal output
rlabel metal2 s 114098 -400 114154 800 6 la_data_in_mprj[42]
port 196 nsew signal output
rlabel metal2 s 116306 -400 116362 800 6 la_data_in_mprj[43]
port 197 nsew signal output
rlabel metal2 s 118514 -400 118570 800 6 la_data_in_mprj[44]
port 198 nsew signal output
rlabel metal2 s 120722 -400 120778 800 6 la_data_in_mprj[45]
port 199 nsew signal output
rlabel metal2 s 122930 -400 122986 800 6 la_data_in_mprj[46]
port 200 nsew signal output
rlabel metal2 s 125138 -400 125194 800 6 la_data_in_mprj[47]
port 201 nsew signal output
rlabel metal2 s 127346 -400 127402 800 6 la_data_in_mprj[48]
port 202 nsew signal output
rlabel metal2 s 129554 -400 129610 800 6 la_data_in_mprj[49]
port 203 nsew signal output
rlabel metal2 s 30194 -400 30250 800 6 la_data_in_mprj[4]
port 204 nsew signal output
rlabel metal2 s 131762 -400 131818 800 6 la_data_in_mprj[50]
port 205 nsew signal output
rlabel metal2 s 133970 -400 134026 800 6 la_data_in_mprj[51]
port 206 nsew signal output
rlabel metal2 s 136178 -400 136234 800 6 la_data_in_mprj[52]
port 207 nsew signal output
rlabel metal2 s 138386 -400 138442 800 6 la_data_in_mprj[53]
port 208 nsew signal output
rlabel metal2 s 140594 -400 140650 800 6 la_data_in_mprj[54]
port 209 nsew signal output
rlabel metal2 s 142802 -400 142858 800 6 la_data_in_mprj[55]
port 210 nsew signal output
rlabel metal2 s 145010 -400 145066 800 6 la_data_in_mprj[56]
port 211 nsew signal output
rlabel metal2 s 147218 -400 147274 800 6 la_data_in_mprj[57]
port 212 nsew signal output
rlabel metal2 s 149426 -400 149482 800 6 la_data_in_mprj[58]
port 213 nsew signal output
rlabel metal2 s 151634 -400 151690 800 6 la_data_in_mprj[59]
port 214 nsew signal output
rlabel metal2 s 32402 -400 32458 800 6 la_data_in_mprj[5]
port 215 nsew signal output
rlabel metal2 s 153842 -400 153898 800 6 la_data_in_mprj[60]
port 216 nsew signal output
rlabel metal2 s 156050 -400 156106 800 6 la_data_in_mprj[61]
port 217 nsew signal output
rlabel metal2 s 158258 -400 158314 800 6 la_data_in_mprj[62]
port 218 nsew signal output
rlabel metal2 s 160466 -400 160522 800 6 la_data_in_mprj[63]
port 219 nsew signal output
rlabel metal2 s 162674 -400 162730 800 6 la_data_in_mprj[64]
port 220 nsew signal output
rlabel metal2 s 164882 -400 164938 800 6 la_data_in_mprj[65]
port 221 nsew signal output
rlabel metal2 s 167090 -400 167146 800 6 la_data_in_mprj[66]
port 222 nsew signal output
rlabel metal2 s 169298 -400 169354 800 6 la_data_in_mprj[67]
port 223 nsew signal output
rlabel metal2 s 171506 -400 171562 800 6 la_data_in_mprj[68]
port 224 nsew signal output
rlabel metal2 s 173714 -400 173770 800 6 la_data_in_mprj[69]
port 225 nsew signal output
rlabel metal2 s 34610 -400 34666 800 6 la_data_in_mprj[6]
port 226 nsew signal output
rlabel metal2 s 175922 -400 175978 800 6 la_data_in_mprj[70]
port 227 nsew signal output
rlabel metal2 s 179234 -400 179290 800 6 la_data_in_mprj[71]
port 228 nsew signal output
rlabel metal2 s 181442 -400 181498 800 6 la_data_in_mprj[72]
port 229 nsew signal output
rlabel metal2 s 183650 -400 183706 800 6 la_data_in_mprj[73]
port 230 nsew signal output
rlabel metal2 s 185858 -400 185914 800 6 la_data_in_mprj[74]
port 231 nsew signal output
rlabel metal2 s 188066 -400 188122 800 6 la_data_in_mprj[75]
port 232 nsew signal output
rlabel metal2 s 190274 -400 190330 800 6 la_data_in_mprj[76]
port 233 nsew signal output
rlabel metal2 s 192482 -400 192538 800 6 la_data_in_mprj[77]
port 234 nsew signal output
rlabel metal2 s 194690 -400 194746 800 6 la_data_in_mprj[78]
port 235 nsew signal output
rlabel metal2 s 196898 -400 196954 800 6 la_data_in_mprj[79]
port 236 nsew signal output
rlabel metal2 s 36818 -400 36874 800 6 la_data_in_mprj[7]
port 237 nsew signal output
rlabel metal2 s 199106 -400 199162 800 6 la_data_in_mprj[80]
port 238 nsew signal output
rlabel metal2 s 201314 -400 201370 800 6 la_data_in_mprj[81]
port 239 nsew signal output
rlabel metal2 s 203522 -400 203578 800 6 la_data_in_mprj[82]
port 240 nsew signal output
rlabel metal2 s 205730 -400 205786 800 6 la_data_in_mprj[83]
port 241 nsew signal output
rlabel metal2 s 207938 -400 207994 800 6 la_data_in_mprj[84]
port 242 nsew signal output
rlabel metal2 s 210146 -400 210202 800 6 la_data_in_mprj[85]
port 243 nsew signal output
rlabel metal2 s 212354 -400 212410 800 6 la_data_in_mprj[86]
port 244 nsew signal output
rlabel metal2 s 214562 -400 214618 800 6 la_data_in_mprj[87]
port 245 nsew signal output
rlabel metal2 s 216770 -400 216826 800 6 la_data_in_mprj[88]
port 246 nsew signal output
rlabel metal2 s 218978 -400 219034 800 6 la_data_in_mprj[89]
port 247 nsew signal output
rlabel metal2 s 39026 -400 39082 800 6 la_data_in_mprj[8]
port 248 nsew signal output
rlabel metal2 s 221186 -400 221242 800 6 la_data_in_mprj[90]
port 249 nsew signal output
rlabel metal2 s 223394 -400 223450 800 6 la_data_in_mprj[91]
port 250 nsew signal output
rlabel metal2 s 225602 -400 225658 800 6 la_data_in_mprj[92]
port 251 nsew signal output
rlabel metal2 s 227810 -400 227866 800 6 la_data_in_mprj[93]
port 252 nsew signal output
rlabel metal2 s 230018 -400 230074 800 6 la_data_in_mprj[94]
port 253 nsew signal output
rlabel metal2 s 232226 -400 232282 800 6 la_data_in_mprj[95]
port 254 nsew signal output
rlabel metal2 s 234434 -400 234490 800 6 la_data_in_mprj[96]
port 255 nsew signal output
rlabel metal2 s 236642 -400 236698 800 6 la_data_in_mprj[97]
port 256 nsew signal output
rlabel metal2 s 238850 -400 238906 800 6 la_data_in_mprj[98]
port 257 nsew signal output
rlabel metal2 s 241058 -400 241114 800 6 la_data_in_mprj[99]
port 258 nsew signal output
rlabel metal2 s 41234 -400 41290 800 6 la_data_in_mprj[9]
port 259 nsew signal output
rlabel metal2 s 90362 27200 90418 28400 6 la_data_out_core[0]
port 260 nsew signal input
rlabel metal2 s 311162 27200 311218 28400 6 la_data_out_core[100]
port 261 nsew signal input
rlabel metal2 s 313370 27200 313426 28400 6 la_data_out_core[101]
port 262 nsew signal input
rlabel metal2 s 315578 27200 315634 28400 6 la_data_out_core[102]
port 263 nsew signal input
rlabel metal2 s 317786 27200 317842 28400 6 la_data_out_core[103]
port 264 nsew signal input
rlabel metal2 s 319994 27200 320050 28400 6 la_data_out_core[104]
port 265 nsew signal input
rlabel metal2 s 322202 27200 322258 28400 6 la_data_out_core[105]
port 266 nsew signal input
rlabel metal2 s 324410 27200 324466 28400 6 la_data_out_core[106]
port 267 nsew signal input
rlabel metal2 s 326618 27200 326674 28400 6 la_data_out_core[107]
port 268 nsew signal input
rlabel metal2 s 328826 27200 328882 28400 6 la_data_out_core[108]
port 269 nsew signal input
rlabel metal2 s 331034 27200 331090 28400 6 la_data_out_core[109]
port 270 nsew signal input
rlabel metal2 s 112442 27200 112498 28400 6 la_data_out_core[10]
port 271 nsew signal input
rlabel metal2 s 333242 27200 333298 28400 6 la_data_out_core[110]
port 272 nsew signal input
rlabel metal2 s 335450 27200 335506 28400 6 la_data_out_core[111]
port 273 nsew signal input
rlabel metal2 s 337658 27200 337714 28400 6 la_data_out_core[112]
port 274 nsew signal input
rlabel metal2 s 339866 27200 339922 28400 6 la_data_out_core[113]
port 275 nsew signal input
rlabel metal2 s 342074 27200 342130 28400 6 la_data_out_core[114]
port 276 nsew signal input
rlabel metal2 s 344282 27200 344338 28400 6 la_data_out_core[115]
port 277 nsew signal input
rlabel metal2 s 346490 27200 346546 28400 6 la_data_out_core[116]
port 278 nsew signal input
rlabel metal2 s 348698 27200 348754 28400 6 la_data_out_core[117]
port 279 nsew signal input
rlabel metal2 s 350906 27200 350962 28400 6 la_data_out_core[118]
port 280 nsew signal input
rlabel metal2 s 353114 27200 353170 28400 6 la_data_out_core[119]
port 281 nsew signal input
rlabel metal2 s 114650 27200 114706 28400 6 la_data_out_core[11]
port 282 nsew signal input
rlabel metal2 s 355322 27200 355378 28400 6 la_data_out_core[120]
port 283 nsew signal input
rlabel metal2 s 357530 27200 357586 28400 6 la_data_out_core[121]
port 284 nsew signal input
rlabel metal2 s 359738 27200 359794 28400 6 la_data_out_core[122]
port 285 nsew signal input
rlabel metal2 s 361946 27200 362002 28400 6 la_data_out_core[123]
port 286 nsew signal input
rlabel metal2 s 364154 27200 364210 28400 6 la_data_out_core[124]
port 287 nsew signal input
rlabel metal2 s 366362 27200 366418 28400 6 la_data_out_core[125]
port 288 nsew signal input
rlabel metal2 s 368570 27200 368626 28400 6 la_data_out_core[126]
port 289 nsew signal input
rlabel metal2 s 370778 27200 370834 28400 6 la_data_out_core[127]
port 290 nsew signal input
rlabel metal2 s 116858 27200 116914 28400 6 la_data_out_core[12]
port 291 nsew signal input
rlabel metal2 s 119066 27200 119122 28400 6 la_data_out_core[13]
port 292 nsew signal input
rlabel metal2 s 121274 27200 121330 28400 6 la_data_out_core[14]
port 293 nsew signal input
rlabel metal2 s 123482 27200 123538 28400 6 la_data_out_core[15]
port 294 nsew signal input
rlabel metal2 s 125690 27200 125746 28400 6 la_data_out_core[16]
port 295 nsew signal input
rlabel metal2 s 127898 27200 127954 28400 6 la_data_out_core[17]
port 296 nsew signal input
rlabel metal2 s 130106 27200 130162 28400 6 la_data_out_core[18]
port 297 nsew signal input
rlabel metal2 s 132314 27200 132370 28400 6 la_data_out_core[19]
port 298 nsew signal input
rlabel metal2 s 92570 27200 92626 28400 6 la_data_out_core[1]
port 299 nsew signal input
rlabel metal2 s 134522 27200 134578 28400 6 la_data_out_core[20]
port 300 nsew signal input
rlabel metal2 s 136730 27200 136786 28400 6 la_data_out_core[21]
port 301 nsew signal input
rlabel metal2 s 138938 27200 138994 28400 6 la_data_out_core[22]
port 302 nsew signal input
rlabel metal2 s 141146 27200 141202 28400 6 la_data_out_core[23]
port 303 nsew signal input
rlabel metal2 s 143354 27200 143410 28400 6 la_data_out_core[24]
port 304 nsew signal input
rlabel metal2 s 145562 27200 145618 28400 6 la_data_out_core[25]
port 305 nsew signal input
rlabel metal2 s 147770 27200 147826 28400 6 la_data_out_core[26]
port 306 nsew signal input
rlabel metal2 s 149978 27200 150034 28400 6 la_data_out_core[27]
port 307 nsew signal input
rlabel metal2 s 152186 27200 152242 28400 6 la_data_out_core[28]
port 308 nsew signal input
rlabel metal2 s 154394 27200 154450 28400 6 la_data_out_core[29]
port 309 nsew signal input
rlabel metal2 s 94778 27200 94834 28400 6 la_data_out_core[2]
port 310 nsew signal input
rlabel metal2 s 156602 27200 156658 28400 6 la_data_out_core[30]
port 311 nsew signal input
rlabel metal2 s 158810 27200 158866 28400 6 la_data_out_core[31]
port 312 nsew signal input
rlabel metal2 s 161018 27200 161074 28400 6 la_data_out_core[32]
port 313 nsew signal input
rlabel metal2 s 163226 27200 163282 28400 6 la_data_out_core[33]
port 314 nsew signal input
rlabel metal2 s 165434 27200 165490 28400 6 la_data_out_core[34]
port 315 nsew signal input
rlabel metal2 s 167642 27200 167698 28400 6 la_data_out_core[35]
port 316 nsew signal input
rlabel metal2 s 169850 27200 169906 28400 6 la_data_out_core[36]
port 317 nsew signal input
rlabel metal2 s 172058 27200 172114 28400 6 la_data_out_core[37]
port 318 nsew signal input
rlabel metal2 s 174266 27200 174322 28400 6 la_data_out_core[38]
port 319 nsew signal input
rlabel metal2 s 176474 27200 176530 28400 6 la_data_out_core[39]
port 320 nsew signal input
rlabel metal2 s 96986 27200 97042 28400 6 la_data_out_core[3]
port 321 nsew signal input
rlabel metal2 s 178682 27200 178738 28400 6 la_data_out_core[40]
port 322 nsew signal input
rlabel metal2 s 180890 27200 180946 28400 6 la_data_out_core[41]
port 323 nsew signal input
rlabel metal2 s 183098 27200 183154 28400 6 la_data_out_core[42]
port 324 nsew signal input
rlabel metal2 s 185306 27200 185362 28400 6 la_data_out_core[43]
port 325 nsew signal input
rlabel metal2 s 187514 27200 187570 28400 6 la_data_out_core[44]
port 326 nsew signal input
rlabel metal2 s 189722 27200 189778 28400 6 la_data_out_core[45]
port 327 nsew signal input
rlabel metal2 s 191930 27200 191986 28400 6 la_data_out_core[46]
port 328 nsew signal input
rlabel metal2 s 194138 27200 194194 28400 6 la_data_out_core[47]
port 329 nsew signal input
rlabel metal2 s 196346 27200 196402 28400 6 la_data_out_core[48]
port 330 nsew signal input
rlabel metal2 s 198554 27200 198610 28400 6 la_data_out_core[49]
port 331 nsew signal input
rlabel metal2 s 99194 27200 99250 28400 6 la_data_out_core[4]
port 332 nsew signal input
rlabel metal2 s 200762 27200 200818 28400 6 la_data_out_core[50]
port 333 nsew signal input
rlabel metal2 s 202970 27200 203026 28400 6 la_data_out_core[51]
port 334 nsew signal input
rlabel metal2 s 205178 27200 205234 28400 6 la_data_out_core[52]
port 335 nsew signal input
rlabel metal2 s 207386 27200 207442 28400 6 la_data_out_core[53]
port 336 nsew signal input
rlabel metal2 s 209594 27200 209650 28400 6 la_data_out_core[54]
port 337 nsew signal input
rlabel metal2 s 211802 27200 211858 28400 6 la_data_out_core[55]
port 338 nsew signal input
rlabel metal2 s 214010 27200 214066 28400 6 la_data_out_core[56]
port 339 nsew signal input
rlabel metal2 s 216218 27200 216274 28400 6 la_data_out_core[57]
port 340 nsew signal input
rlabel metal2 s 218426 27200 218482 28400 6 la_data_out_core[58]
port 341 nsew signal input
rlabel metal2 s 220634 27200 220690 28400 6 la_data_out_core[59]
port 342 nsew signal input
rlabel metal2 s 101402 27200 101458 28400 6 la_data_out_core[5]
port 343 nsew signal input
rlabel metal2 s 222842 27200 222898 28400 6 la_data_out_core[60]
port 344 nsew signal input
rlabel metal2 s 225050 27200 225106 28400 6 la_data_out_core[61]
port 345 nsew signal input
rlabel metal2 s 227258 27200 227314 28400 6 la_data_out_core[62]
port 346 nsew signal input
rlabel metal2 s 229466 27200 229522 28400 6 la_data_out_core[63]
port 347 nsew signal input
rlabel metal2 s 231674 27200 231730 28400 6 la_data_out_core[64]
port 348 nsew signal input
rlabel metal2 s 233882 27200 233938 28400 6 la_data_out_core[65]
port 349 nsew signal input
rlabel metal2 s 236090 27200 236146 28400 6 la_data_out_core[66]
port 350 nsew signal input
rlabel metal2 s 238298 27200 238354 28400 6 la_data_out_core[67]
port 351 nsew signal input
rlabel metal2 s 240506 27200 240562 28400 6 la_data_out_core[68]
port 352 nsew signal input
rlabel metal2 s 242714 27200 242770 28400 6 la_data_out_core[69]
port 353 nsew signal input
rlabel metal2 s 103610 27200 103666 28400 6 la_data_out_core[6]
port 354 nsew signal input
rlabel metal2 s 244922 27200 244978 28400 6 la_data_out_core[70]
port 355 nsew signal input
rlabel metal2 s 247130 27200 247186 28400 6 la_data_out_core[71]
port 356 nsew signal input
rlabel metal2 s 249338 27200 249394 28400 6 la_data_out_core[72]
port 357 nsew signal input
rlabel metal2 s 251546 27200 251602 28400 6 la_data_out_core[73]
port 358 nsew signal input
rlabel metal2 s 253754 27200 253810 28400 6 la_data_out_core[74]
port 359 nsew signal input
rlabel metal2 s 255962 27200 256018 28400 6 la_data_out_core[75]
port 360 nsew signal input
rlabel metal2 s 258170 27200 258226 28400 6 la_data_out_core[76]
port 361 nsew signal input
rlabel metal2 s 260378 27200 260434 28400 6 la_data_out_core[77]
port 362 nsew signal input
rlabel metal2 s 262586 27200 262642 28400 6 la_data_out_core[78]
port 363 nsew signal input
rlabel metal2 s 264794 27200 264850 28400 6 la_data_out_core[79]
port 364 nsew signal input
rlabel metal2 s 105818 27200 105874 28400 6 la_data_out_core[7]
port 365 nsew signal input
rlabel metal2 s 267002 27200 267058 28400 6 la_data_out_core[80]
port 366 nsew signal input
rlabel metal2 s 269210 27200 269266 28400 6 la_data_out_core[81]
port 367 nsew signal input
rlabel metal2 s 271418 27200 271474 28400 6 la_data_out_core[82]
port 368 nsew signal input
rlabel metal2 s 273626 27200 273682 28400 6 la_data_out_core[83]
port 369 nsew signal input
rlabel metal2 s 275834 27200 275890 28400 6 la_data_out_core[84]
port 370 nsew signal input
rlabel metal2 s 278042 27200 278098 28400 6 la_data_out_core[85]
port 371 nsew signal input
rlabel metal2 s 280250 27200 280306 28400 6 la_data_out_core[86]
port 372 nsew signal input
rlabel metal2 s 282458 27200 282514 28400 6 la_data_out_core[87]
port 373 nsew signal input
rlabel metal2 s 284666 27200 284722 28400 6 la_data_out_core[88]
port 374 nsew signal input
rlabel metal2 s 286874 27200 286930 28400 6 la_data_out_core[89]
port 375 nsew signal input
rlabel metal2 s 108026 27200 108082 28400 6 la_data_out_core[8]
port 376 nsew signal input
rlabel metal2 s 289082 27200 289138 28400 6 la_data_out_core[90]
port 377 nsew signal input
rlabel metal2 s 291290 27200 291346 28400 6 la_data_out_core[91]
port 378 nsew signal input
rlabel metal2 s 293498 27200 293554 28400 6 la_data_out_core[92]
port 379 nsew signal input
rlabel metal2 s 295706 27200 295762 28400 6 la_data_out_core[93]
port 380 nsew signal input
rlabel metal2 s 297914 27200 297970 28400 6 la_data_out_core[94]
port 381 nsew signal input
rlabel metal2 s 300122 27200 300178 28400 6 la_data_out_core[95]
port 382 nsew signal input
rlabel metal2 s 302330 27200 302386 28400 6 la_data_out_core[96]
port 383 nsew signal input
rlabel metal2 s 304538 27200 304594 28400 6 la_data_out_core[97]
port 384 nsew signal input
rlabel metal2 s 306746 27200 306802 28400 6 la_data_out_core[98]
port 385 nsew signal input
rlabel metal2 s 308954 27200 309010 28400 6 la_data_out_core[99]
port 386 nsew signal input
rlabel metal2 s 110234 27200 110290 28400 6 la_data_out_core[9]
port 387 nsew signal input
rlabel metal2 s 21914 -400 21970 800 6 la_data_out_mprj[0]
port 388 nsew signal input
rlabel metal2 s 243818 -400 243874 800 6 la_data_out_mprj[100]
port 389 nsew signal input
rlabel metal2 s 246026 -400 246082 800 6 la_data_out_mprj[101]
port 390 nsew signal input
rlabel metal2 s 248234 -400 248290 800 6 la_data_out_mprj[102]
port 391 nsew signal input
rlabel metal2 s 250442 -400 250498 800 6 la_data_out_mprj[103]
port 392 nsew signal input
rlabel metal2 s 252650 -400 252706 800 6 la_data_out_mprj[104]
port 393 nsew signal input
rlabel metal2 s 254858 -400 254914 800 6 la_data_out_mprj[105]
port 394 nsew signal input
rlabel metal2 s 257066 -400 257122 800 6 la_data_out_mprj[106]
port 395 nsew signal input
rlabel metal2 s 259274 -400 259330 800 6 la_data_out_mprj[107]
port 396 nsew signal input
rlabel metal2 s 261482 -400 261538 800 6 la_data_out_mprj[108]
port 397 nsew signal input
rlabel metal2 s 263690 -400 263746 800 6 la_data_out_mprj[109]
port 398 nsew signal input
rlabel metal2 s 43994 -400 44050 800 6 la_data_out_mprj[10]
port 399 nsew signal input
rlabel metal2 s 265898 -400 265954 800 6 la_data_out_mprj[110]
port 400 nsew signal input
rlabel metal2 s 268106 -400 268162 800 6 la_data_out_mprj[111]
port 401 nsew signal input
rlabel metal2 s 270314 -400 270370 800 6 la_data_out_mprj[112]
port 402 nsew signal input
rlabel metal2 s 272522 -400 272578 800 6 la_data_out_mprj[113]
port 403 nsew signal input
rlabel metal2 s 274730 -400 274786 800 6 la_data_out_mprj[114]
port 404 nsew signal input
rlabel metal2 s 276938 -400 276994 800 6 la_data_out_mprj[115]
port 405 nsew signal input
rlabel metal2 s 279146 -400 279202 800 6 la_data_out_mprj[116]
port 406 nsew signal input
rlabel metal2 s 281354 -400 281410 800 6 la_data_out_mprj[117]
port 407 nsew signal input
rlabel metal2 s 283562 -400 283618 800 6 la_data_out_mprj[118]
port 408 nsew signal input
rlabel metal2 s 285770 -400 285826 800 6 la_data_out_mprj[119]
port 409 nsew signal input
rlabel metal2 s 46202 -400 46258 800 6 la_data_out_mprj[11]
port 410 nsew signal input
rlabel metal2 s 287978 -400 288034 800 6 la_data_out_mprj[120]
port 411 nsew signal input
rlabel metal2 s 290186 -400 290242 800 6 la_data_out_mprj[121]
port 412 nsew signal input
rlabel metal2 s 292394 -400 292450 800 6 la_data_out_mprj[122]
port 413 nsew signal input
rlabel metal2 s 294602 -400 294658 800 6 la_data_out_mprj[123]
port 414 nsew signal input
rlabel metal2 s 296810 -400 296866 800 6 la_data_out_mprj[124]
port 415 nsew signal input
rlabel metal2 s 299018 -400 299074 800 6 la_data_out_mprj[125]
port 416 nsew signal input
rlabel metal2 s 301226 -400 301282 800 6 la_data_out_mprj[126]
port 417 nsew signal input
rlabel metal2 s 303434 -400 303490 800 6 la_data_out_mprj[127]
port 418 nsew signal input
rlabel metal2 s 48410 -400 48466 800 6 la_data_out_mprj[12]
port 419 nsew signal input
rlabel metal2 s 50618 -400 50674 800 6 la_data_out_mprj[13]
port 420 nsew signal input
rlabel metal2 s 52826 -400 52882 800 6 la_data_out_mprj[14]
port 421 nsew signal input
rlabel metal2 s 55034 -400 55090 800 6 la_data_out_mprj[15]
port 422 nsew signal input
rlabel metal2 s 57242 -400 57298 800 6 la_data_out_mprj[16]
port 423 nsew signal input
rlabel metal2 s 59450 -400 59506 800 6 la_data_out_mprj[17]
port 424 nsew signal input
rlabel metal2 s 61658 -400 61714 800 6 la_data_out_mprj[18]
port 425 nsew signal input
rlabel metal2 s 63866 -400 63922 800 6 la_data_out_mprj[19]
port 426 nsew signal input
rlabel metal2 s 24122 -400 24178 800 6 la_data_out_mprj[1]
port 427 nsew signal input
rlabel metal2 s 66074 -400 66130 800 6 la_data_out_mprj[20]
port 428 nsew signal input
rlabel metal2 s 68282 -400 68338 800 6 la_data_out_mprj[21]
port 429 nsew signal input
rlabel metal2 s 70490 -400 70546 800 6 la_data_out_mprj[22]
port 430 nsew signal input
rlabel metal2 s 72698 -400 72754 800 6 la_data_out_mprj[23]
port 431 nsew signal input
rlabel metal2 s 74906 -400 74962 800 6 la_data_out_mprj[24]
port 432 nsew signal input
rlabel metal2 s 77114 -400 77170 800 6 la_data_out_mprj[25]
port 433 nsew signal input
rlabel metal2 s 79322 -400 79378 800 6 la_data_out_mprj[26]
port 434 nsew signal input
rlabel metal2 s 81530 -400 81586 800 6 la_data_out_mprj[27]
port 435 nsew signal input
rlabel metal2 s 83738 -400 83794 800 6 la_data_out_mprj[28]
port 436 nsew signal input
rlabel metal2 s 85946 -400 86002 800 6 la_data_out_mprj[29]
port 437 nsew signal input
rlabel metal2 s 26330 -400 26386 800 6 la_data_out_mprj[2]
port 438 nsew signal input
rlabel metal2 s 88154 -400 88210 800 6 la_data_out_mprj[30]
port 439 nsew signal input
rlabel metal2 s 90362 -400 90418 800 6 la_data_out_mprj[31]
port 440 nsew signal input
rlabel metal2 s 92570 -400 92626 800 6 la_data_out_mprj[32]
port 441 nsew signal input
rlabel metal2 s 94778 -400 94834 800 6 la_data_out_mprj[33]
port 442 nsew signal input
rlabel metal2 s 96986 -400 97042 800 6 la_data_out_mprj[34]
port 443 nsew signal input
rlabel metal2 s 99194 -400 99250 800 6 la_data_out_mprj[35]
port 444 nsew signal input
rlabel metal2 s 101402 -400 101458 800 6 la_data_out_mprj[36]
port 445 nsew signal input
rlabel metal2 s 103610 -400 103666 800 6 la_data_out_mprj[37]
port 446 nsew signal input
rlabel metal2 s 105818 -400 105874 800 6 la_data_out_mprj[38]
port 447 nsew signal input
rlabel metal2 s 108026 -400 108082 800 6 la_data_out_mprj[39]
port 448 nsew signal input
rlabel metal2 s 28538 -400 28594 800 6 la_data_out_mprj[3]
port 449 nsew signal input
rlabel metal2 s 110234 -400 110290 800 6 la_data_out_mprj[40]
port 450 nsew signal input
rlabel metal2 s 112442 -400 112498 800 6 la_data_out_mprj[41]
port 451 nsew signal input
rlabel metal2 s 114650 -400 114706 800 6 la_data_out_mprj[42]
port 452 nsew signal input
rlabel metal2 s 116858 -400 116914 800 6 la_data_out_mprj[43]
port 453 nsew signal input
rlabel metal2 s 119066 -400 119122 800 6 la_data_out_mprj[44]
port 454 nsew signal input
rlabel metal2 s 121274 -400 121330 800 6 la_data_out_mprj[45]
port 455 nsew signal input
rlabel metal2 s 123482 -400 123538 800 6 la_data_out_mprj[46]
port 456 nsew signal input
rlabel metal2 s 125690 -400 125746 800 6 la_data_out_mprj[47]
port 457 nsew signal input
rlabel metal2 s 127898 -400 127954 800 6 la_data_out_mprj[48]
port 458 nsew signal input
rlabel metal2 s 130106 -400 130162 800 6 la_data_out_mprj[49]
port 459 nsew signal input
rlabel metal2 s 30746 -400 30802 800 6 la_data_out_mprj[4]
port 460 nsew signal input
rlabel metal2 s 132314 -400 132370 800 6 la_data_out_mprj[50]
port 461 nsew signal input
rlabel metal2 s 134522 -400 134578 800 6 la_data_out_mprj[51]
port 462 nsew signal input
rlabel metal2 s 136730 -400 136786 800 6 la_data_out_mprj[52]
port 463 nsew signal input
rlabel metal2 s 138938 -400 138994 800 6 la_data_out_mprj[53]
port 464 nsew signal input
rlabel metal2 s 141146 -400 141202 800 6 la_data_out_mprj[54]
port 465 nsew signal input
rlabel metal2 s 143354 -400 143410 800 6 la_data_out_mprj[55]
port 466 nsew signal input
rlabel metal2 s 145562 -400 145618 800 6 la_data_out_mprj[56]
port 467 nsew signal input
rlabel metal2 s 147770 -400 147826 800 6 la_data_out_mprj[57]
port 468 nsew signal input
rlabel metal2 s 149978 -400 150034 800 6 la_data_out_mprj[58]
port 469 nsew signal input
rlabel metal2 s 152186 -400 152242 800 6 la_data_out_mprj[59]
port 470 nsew signal input
rlabel metal2 s 32954 -400 33010 800 6 la_data_out_mprj[5]
port 471 nsew signal input
rlabel metal2 s 154394 -400 154450 800 6 la_data_out_mprj[60]
port 472 nsew signal input
rlabel metal2 s 156602 -400 156658 800 6 la_data_out_mprj[61]
port 473 nsew signal input
rlabel metal2 s 158810 -400 158866 800 6 la_data_out_mprj[62]
port 474 nsew signal input
rlabel metal2 s 161018 -400 161074 800 6 la_data_out_mprj[63]
port 475 nsew signal input
rlabel metal2 s 163226 -400 163282 800 6 la_data_out_mprj[64]
port 476 nsew signal input
rlabel metal2 s 165434 -400 165490 800 6 la_data_out_mprj[65]
port 477 nsew signal input
rlabel metal2 s 167642 -400 167698 800 6 la_data_out_mprj[66]
port 478 nsew signal input
rlabel metal2 s 169850 -400 169906 800 6 la_data_out_mprj[67]
port 479 nsew signal input
rlabel metal2 s 172058 -400 172114 800 6 la_data_out_mprj[68]
port 480 nsew signal input
rlabel metal2 s 174266 -400 174322 800 6 la_data_out_mprj[69]
port 481 nsew signal input
rlabel metal2 s 35162 -400 35218 800 6 la_data_out_mprj[6]
port 482 nsew signal input
rlabel metal2 s 176474 -400 176530 800 6 la_data_out_mprj[70]
port 483 nsew signal input
rlabel metal2 s 179786 -400 179842 800 6 la_data_out_mprj[71]
port 484 nsew signal input
rlabel metal2 s 181994 -400 182050 800 6 la_data_out_mprj[72]
port 485 nsew signal input
rlabel metal2 s 184202 -400 184258 800 6 la_data_out_mprj[73]
port 486 nsew signal input
rlabel metal2 s 186410 -400 186466 800 6 la_data_out_mprj[74]
port 487 nsew signal input
rlabel metal2 s 188618 -400 188674 800 6 la_data_out_mprj[75]
port 488 nsew signal input
rlabel metal2 s 190826 -400 190882 800 6 la_data_out_mprj[76]
port 489 nsew signal input
rlabel metal2 s 193034 -400 193090 800 6 la_data_out_mprj[77]
port 490 nsew signal input
rlabel metal2 s 195242 -400 195298 800 6 la_data_out_mprj[78]
port 491 nsew signal input
rlabel metal2 s 197450 -400 197506 800 6 la_data_out_mprj[79]
port 492 nsew signal input
rlabel metal2 s 37370 -400 37426 800 6 la_data_out_mprj[7]
port 493 nsew signal input
rlabel metal2 s 199658 -400 199714 800 6 la_data_out_mprj[80]
port 494 nsew signal input
rlabel metal2 s 201866 -400 201922 800 6 la_data_out_mprj[81]
port 495 nsew signal input
rlabel metal2 s 204074 -400 204130 800 6 la_data_out_mprj[82]
port 496 nsew signal input
rlabel metal2 s 206282 -400 206338 800 6 la_data_out_mprj[83]
port 497 nsew signal input
rlabel metal2 s 208490 -400 208546 800 6 la_data_out_mprj[84]
port 498 nsew signal input
rlabel metal2 s 210698 -400 210754 800 6 la_data_out_mprj[85]
port 499 nsew signal input
rlabel metal2 s 212906 -400 212962 800 6 la_data_out_mprj[86]
port 500 nsew signal input
rlabel metal2 s 215114 -400 215170 800 6 la_data_out_mprj[87]
port 501 nsew signal input
rlabel metal2 s 217322 -400 217378 800 6 la_data_out_mprj[88]
port 502 nsew signal input
rlabel metal2 s 219530 -400 219586 800 6 la_data_out_mprj[89]
port 503 nsew signal input
rlabel metal2 s 39578 -400 39634 800 6 la_data_out_mprj[8]
port 504 nsew signal input
rlabel metal2 s 221738 -400 221794 800 6 la_data_out_mprj[90]
port 505 nsew signal input
rlabel metal2 s 223946 -400 224002 800 6 la_data_out_mprj[91]
port 506 nsew signal input
rlabel metal2 s 226154 -400 226210 800 6 la_data_out_mprj[92]
port 507 nsew signal input
rlabel metal2 s 228362 -400 228418 800 6 la_data_out_mprj[93]
port 508 nsew signal input
rlabel metal2 s 230570 -400 230626 800 6 la_data_out_mprj[94]
port 509 nsew signal input
rlabel metal2 s 232778 -400 232834 800 6 la_data_out_mprj[95]
port 510 nsew signal input
rlabel metal2 s 234986 -400 235042 800 6 la_data_out_mprj[96]
port 511 nsew signal input
rlabel metal2 s 237194 -400 237250 800 6 la_data_out_mprj[97]
port 512 nsew signal input
rlabel metal2 s 239402 -400 239458 800 6 la_data_out_mprj[98]
port 513 nsew signal input
rlabel metal2 s 241610 -400 241666 800 6 la_data_out_mprj[99]
port 514 nsew signal input
rlabel metal2 s 41786 -400 41842 800 6 la_data_out_mprj[9]
port 515 nsew signal input
rlabel metal2 s 22466 -400 22522 800 6 la_iena_mprj[0]
port 516 nsew signal input
rlabel metal2 s 244370 -400 244426 800 6 la_iena_mprj[100]
port 517 nsew signal input
rlabel metal2 s 246578 -400 246634 800 6 la_iena_mprj[101]
port 518 nsew signal input
rlabel metal2 s 248786 -400 248842 800 6 la_iena_mprj[102]
port 519 nsew signal input
rlabel metal2 s 250994 -400 251050 800 6 la_iena_mprj[103]
port 520 nsew signal input
rlabel metal2 s 253202 -400 253258 800 6 la_iena_mprj[104]
port 521 nsew signal input
rlabel metal2 s 255410 -400 255466 800 6 la_iena_mprj[105]
port 522 nsew signal input
rlabel metal2 s 257618 -400 257674 800 6 la_iena_mprj[106]
port 523 nsew signal input
rlabel metal2 s 259826 -400 259882 800 6 la_iena_mprj[107]
port 524 nsew signal input
rlabel metal2 s 262034 -400 262090 800 6 la_iena_mprj[108]
port 525 nsew signal input
rlabel metal2 s 264242 -400 264298 800 6 la_iena_mprj[109]
port 526 nsew signal input
rlabel metal2 s 44546 -400 44602 800 6 la_iena_mprj[10]
port 527 nsew signal input
rlabel metal2 s 266450 -400 266506 800 6 la_iena_mprj[110]
port 528 nsew signal input
rlabel metal2 s 268658 -400 268714 800 6 la_iena_mprj[111]
port 529 nsew signal input
rlabel metal2 s 270866 -400 270922 800 6 la_iena_mprj[112]
port 530 nsew signal input
rlabel metal2 s 273074 -400 273130 800 6 la_iena_mprj[113]
port 531 nsew signal input
rlabel metal2 s 275282 -400 275338 800 6 la_iena_mprj[114]
port 532 nsew signal input
rlabel metal2 s 277490 -400 277546 800 6 la_iena_mprj[115]
port 533 nsew signal input
rlabel metal2 s 279698 -400 279754 800 6 la_iena_mprj[116]
port 534 nsew signal input
rlabel metal2 s 281906 -400 281962 800 6 la_iena_mprj[117]
port 535 nsew signal input
rlabel metal2 s 284114 -400 284170 800 6 la_iena_mprj[118]
port 536 nsew signal input
rlabel metal2 s 286322 -400 286378 800 6 la_iena_mprj[119]
port 537 nsew signal input
rlabel metal2 s 46754 -400 46810 800 6 la_iena_mprj[11]
port 538 nsew signal input
rlabel metal2 s 288530 -400 288586 800 6 la_iena_mprj[120]
port 539 nsew signal input
rlabel metal2 s 290738 -400 290794 800 6 la_iena_mprj[121]
port 540 nsew signal input
rlabel metal2 s 292946 -400 293002 800 6 la_iena_mprj[122]
port 541 nsew signal input
rlabel metal2 s 295154 -400 295210 800 6 la_iena_mprj[123]
port 542 nsew signal input
rlabel metal2 s 297362 -400 297418 800 6 la_iena_mprj[124]
port 543 nsew signal input
rlabel metal2 s 299570 -400 299626 800 6 la_iena_mprj[125]
port 544 nsew signal input
rlabel metal2 s 301778 -400 301834 800 6 la_iena_mprj[126]
port 545 nsew signal input
rlabel metal2 s 303986 -400 304042 800 6 la_iena_mprj[127]
port 546 nsew signal input
rlabel metal2 s 48962 -400 49018 800 6 la_iena_mprj[12]
port 547 nsew signal input
rlabel metal2 s 51170 -400 51226 800 6 la_iena_mprj[13]
port 548 nsew signal input
rlabel metal2 s 53378 -400 53434 800 6 la_iena_mprj[14]
port 549 nsew signal input
rlabel metal2 s 55586 -400 55642 800 6 la_iena_mprj[15]
port 550 nsew signal input
rlabel metal2 s 57794 -400 57850 800 6 la_iena_mprj[16]
port 551 nsew signal input
rlabel metal2 s 60002 -400 60058 800 6 la_iena_mprj[17]
port 552 nsew signal input
rlabel metal2 s 62210 -400 62266 800 6 la_iena_mprj[18]
port 553 nsew signal input
rlabel metal2 s 64418 -400 64474 800 6 la_iena_mprj[19]
port 554 nsew signal input
rlabel metal2 s 24674 -400 24730 800 6 la_iena_mprj[1]
port 555 nsew signal input
rlabel metal2 s 66626 -400 66682 800 6 la_iena_mprj[20]
port 556 nsew signal input
rlabel metal2 s 68834 -400 68890 800 6 la_iena_mprj[21]
port 557 nsew signal input
rlabel metal2 s 71042 -400 71098 800 6 la_iena_mprj[22]
port 558 nsew signal input
rlabel metal2 s 73250 -400 73306 800 6 la_iena_mprj[23]
port 559 nsew signal input
rlabel metal2 s 75458 -400 75514 800 6 la_iena_mprj[24]
port 560 nsew signal input
rlabel metal2 s 77666 -400 77722 800 6 la_iena_mprj[25]
port 561 nsew signal input
rlabel metal2 s 79874 -400 79930 800 6 la_iena_mprj[26]
port 562 nsew signal input
rlabel metal2 s 82082 -400 82138 800 6 la_iena_mprj[27]
port 563 nsew signal input
rlabel metal2 s 84290 -400 84346 800 6 la_iena_mprj[28]
port 564 nsew signal input
rlabel metal2 s 86498 -400 86554 800 6 la_iena_mprj[29]
port 565 nsew signal input
rlabel metal2 s 26882 -400 26938 800 6 la_iena_mprj[2]
port 566 nsew signal input
rlabel metal2 s 88706 -400 88762 800 6 la_iena_mprj[30]
port 567 nsew signal input
rlabel metal2 s 90914 -400 90970 800 6 la_iena_mprj[31]
port 568 nsew signal input
rlabel metal2 s 93122 -400 93178 800 6 la_iena_mprj[32]
port 569 nsew signal input
rlabel metal2 s 95330 -400 95386 800 6 la_iena_mprj[33]
port 570 nsew signal input
rlabel metal2 s 97538 -400 97594 800 6 la_iena_mprj[34]
port 571 nsew signal input
rlabel metal2 s 99746 -400 99802 800 6 la_iena_mprj[35]
port 572 nsew signal input
rlabel metal2 s 101954 -400 102010 800 6 la_iena_mprj[36]
port 573 nsew signal input
rlabel metal2 s 104162 -400 104218 800 6 la_iena_mprj[37]
port 574 nsew signal input
rlabel metal2 s 106370 -400 106426 800 6 la_iena_mprj[38]
port 575 nsew signal input
rlabel metal2 s 108578 -400 108634 800 6 la_iena_mprj[39]
port 576 nsew signal input
rlabel metal2 s 29090 -400 29146 800 6 la_iena_mprj[3]
port 577 nsew signal input
rlabel metal2 s 110786 -400 110842 800 6 la_iena_mprj[40]
port 578 nsew signal input
rlabel metal2 s 112994 -400 113050 800 6 la_iena_mprj[41]
port 579 nsew signal input
rlabel metal2 s 115202 -400 115258 800 6 la_iena_mprj[42]
port 580 nsew signal input
rlabel metal2 s 117410 -400 117466 800 6 la_iena_mprj[43]
port 581 nsew signal input
rlabel metal2 s 119618 -400 119674 800 6 la_iena_mprj[44]
port 582 nsew signal input
rlabel metal2 s 121826 -400 121882 800 6 la_iena_mprj[45]
port 583 nsew signal input
rlabel metal2 s 124034 -400 124090 800 6 la_iena_mprj[46]
port 584 nsew signal input
rlabel metal2 s 126242 -400 126298 800 6 la_iena_mprj[47]
port 585 nsew signal input
rlabel metal2 s 128450 -400 128506 800 6 la_iena_mprj[48]
port 586 nsew signal input
rlabel metal2 s 130658 -400 130714 800 6 la_iena_mprj[49]
port 587 nsew signal input
rlabel metal2 s 31298 -400 31354 800 6 la_iena_mprj[4]
port 588 nsew signal input
rlabel metal2 s 132866 -400 132922 800 6 la_iena_mprj[50]
port 589 nsew signal input
rlabel metal2 s 135074 -400 135130 800 6 la_iena_mprj[51]
port 590 nsew signal input
rlabel metal2 s 137282 -400 137338 800 6 la_iena_mprj[52]
port 591 nsew signal input
rlabel metal2 s 139490 -400 139546 800 6 la_iena_mprj[53]
port 592 nsew signal input
rlabel metal2 s 141698 -400 141754 800 6 la_iena_mprj[54]
port 593 nsew signal input
rlabel metal2 s 143906 -400 143962 800 6 la_iena_mprj[55]
port 594 nsew signal input
rlabel metal2 s 146114 -400 146170 800 6 la_iena_mprj[56]
port 595 nsew signal input
rlabel metal2 s 148322 -400 148378 800 6 la_iena_mprj[57]
port 596 nsew signal input
rlabel metal2 s 150530 -400 150586 800 6 la_iena_mprj[58]
port 597 nsew signal input
rlabel metal2 s 152738 -400 152794 800 6 la_iena_mprj[59]
port 598 nsew signal input
rlabel metal2 s 33506 -400 33562 800 6 la_iena_mprj[5]
port 599 nsew signal input
rlabel metal2 s 154946 -400 155002 800 6 la_iena_mprj[60]
port 600 nsew signal input
rlabel metal2 s 157154 -400 157210 800 6 la_iena_mprj[61]
port 601 nsew signal input
rlabel metal2 s 159362 -400 159418 800 6 la_iena_mprj[62]
port 602 nsew signal input
rlabel metal2 s 161570 -400 161626 800 6 la_iena_mprj[63]
port 603 nsew signal input
rlabel metal2 s 163778 -400 163834 800 6 la_iena_mprj[64]
port 604 nsew signal input
rlabel metal2 s 165986 -400 166042 800 6 la_iena_mprj[65]
port 605 nsew signal input
rlabel metal2 s 168194 -400 168250 800 6 la_iena_mprj[66]
port 606 nsew signal input
rlabel metal2 s 170402 -400 170458 800 6 la_iena_mprj[67]
port 607 nsew signal input
rlabel metal2 s 172610 -400 172666 800 6 la_iena_mprj[68]
port 608 nsew signal input
rlabel metal2 s 174818 -400 174874 800 6 la_iena_mprj[69]
port 609 nsew signal input
rlabel metal2 s 35714 -400 35770 800 6 la_iena_mprj[6]
port 610 nsew signal input
rlabel metal2 s 177026 -400 177082 800 6 la_iena_mprj[70]
port 611 nsew signal input
rlabel metal2 s 180338 -400 180394 800 6 la_iena_mprj[71]
port 612 nsew signal input
rlabel metal2 s 182546 -400 182602 800 6 la_iena_mprj[72]
port 613 nsew signal input
rlabel metal2 s 184754 -400 184810 800 6 la_iena_mprj[73]
port 614 nsew signal input
rlabel metal2 s 186962 -400 187018 800 6 la_iena_mprj[74]
port 615 nsew signal input
rlabel metal2 s 189170 -400 189226 800 6 la_iena_mprj[75]
port 616 nsew signal input
rlabel metal2 s 191378 -400 191434 800 6 la_iena_mprj[76]
port 617 nsew signal input
rlabel metal2 s 193586 -400 193642 800 6 la_iena_mprj[77]
port 618 nsew signal input
rlabel metal2 s 195794 -400 195850 800 6 la_iena_mprj[78]
port 619 nsew signal input
rlabel metal2 s 198002 -400 198058 800 6 la_iena_mprj[79]
port 620 nsew signal input
rlabel metal2 s 37922 -400 37978 800 6 la_iena_mprj[7]
port 621 nsew signal input
rlabel metal2 s 200210 -400 200266 800 6 la_iena_mprj[80]
port 622 nsew signal input
rlabel metal2 s 202418 -400 202474 800 6 la_iena_mprj[81]
port 623 nsew signal input
rlabel metal2 s 204626 -400 204682 800 6 la_iena_mprj[82]
port 624 nsew signal input
rlabel metal2 s 206834 -400 206890 800 6 la_iena_mprj[83]
port 625 nsew signal input
rlabel metal2 s 209042 -400 209098 800 6 la_iena_mprj[84]
port 626 nsew signal input
rlabel metal2 s 211250 -400 211306 800 6 la_iena_mprj[85]
port 627 nsew signal input
rlabel metal2 s 213458 -400 213514 800 6 la_iena_mprj[86]
port 628 nsew signal input
rlabel metal2 s 215666 -400 215722 800 6 la_iena_mprj[87]
port 629 nsew signal input
rlabel metal2 s 217874 -400 217930 800 6 la_iena_mprj[88]
port 630 nsew signal input
rlabel metal2 s 220082 -400 220138 800 6 la_iena_mprj[89]
port 631 nsew signal input
rlabel metal2 s 40130 -400 40186 800 6 la_iena_mprj[8]
port 632 nsew signal input
rlabel metal2 s 222290 -400 222346 800 6 la_iena_mprj[90]
port 633 nsew signal input
rlabel metal2 s 224498 -400 224554 800 6 la_iena_mprj[91]
port 634 nsew signal input
rlabel metal2 s 226706 -400 226762 800 6 la_iena_mprj[92]
port 635 nsew signal input
rlabel metal2 s 228914 -400 228970 800 6 la_iena_mprj[93]
port 636 nsew signal input
rlabel metal2 s 231122 -400 231178 800 6 la_iena_mprj[94]
port 637 nsew signal input
rlabel metal2 s 233330 -400 233386 800 6 la_iena_mprj[95]
port 638 nsew signal input
rlabel metal2 s 235538 -400 235594 800 6 la_iena_mprj[96]
port 639 nsew signal input
rlabel metal2 s 237746 -400 237802 800 6 la_iena_mprj[97]
port 640 nsew signal input
rlabel metal2 s 239954 -400 240010 800 6 la_iena_mprj[98]
port 641 nsew signal input
rlabel metal2 s 242162 -400 242218 800 6 la_iena_mprj[99]
port 642 nsew signal input
rlabel metal2 s 42338 -400 42394 800 6 la_iena_mprj[9]
port 643 nsew signal input
rlabel metal2 s 91098 27200 91154 28400 6 la_oenb_core[0]
port 644 nsew signal output
rlabel metal2 s 311898 27200 311954 28400 6 la_oenb_core[100]
port 645 nsew signal output
rlabel metal2 s 314106 27200 314162 28400 6 la_oenb_core[101]
port 646 nsew signal output
rlabel metal2 s 316314 27200 316370 28400 6 la_oenb_core[102]
port 647 nsew signal output
rlabel metal2 s 318522 27200 318578 28400 6 la_oenb_core[103]
port 648 nsew signal output
rlabel metal2 s 320730 27200 320786 28400 6 la_oenb_core[104]
port 649 nsew signal output
rlabel metal2 s 322938 27200 322994 28400 6 la_oenb_core[105]
port 650 nsew signal output
rlabel metal2 s 325146 27200 325202 28400 6 la_oenb_core[106]
port 651 nsew signal output
rlabel metal2 s 327354 27200 327410 28400 6 la_oenb_core[107]
port 652 nsew signal output
rlabel metal2 s 329562 27200 329618 28400 6 la_oenb_core[108]
port 653 nsew signal output
rlabel metal2 s 331770 27200 331826 28400 6 la_oenb_core[109]
port 654 nsew signal output
rlabel metal2 s 113178 27200 113234 28400 6 la_oenb_core[10]
port 655 nsew signal output
rlabel metal2 s 333978 27200 334034 28400 6 la_oenb_core[110]
port 656 nsew signal output
rlabel metal2 s 336186 27200 336242 28400 6 la_oenb_core[111]
port 657 nsew signal output
rlabel metal2 s 338394 27200 338450 28400 6 la_oenb_core[112]
port 658 nsew signal output
rlabel metal2 s 340602 27200 340658 28400 6 la_oenb_core[113]
port 659 nsew signal output
rlabel metal2 s 342810 27200 342866 28400 6 la_oenb_core[114]
port 660 nsew signal output
rlabel metal2 s 345018 27200 345074 28400 6 la_oenb_core[115]
port 661 nsew signal output
rlabel metal2 s 347226 27200 347282 28400 6 la_oenb_core[116]
port 662 nsew signal output
rlabel metal2 s 349434 27200 349490 28400 6 la_oenb_core[117]
port 663 nsew signal output
rlabel metal2 s 351642 27200 351698 28400 6 la_oenb_core[118]
port 664 nsew signal output
rlabel metal2 s 353850 27200 353906 28400 6 la_oenb_core[119]
port 665 nsew signal output
rlabel metal2 s 115386 27200 115442 28400 6 la_oenb_core[11]
port 666 nsew signal output
rlabel metal2 s 356058 27200 356114 28400 6 la_oenb_core[120]
port 667 nsew signal output
rlabel metal2 s 358266 27200 358322 28400 6 la_oenb_core[121]
port 668 nsew signal output
rlabel metal2 s 360474 27200 360530 28400 6 la_oenb_core[122]
port 669 nsew signal output
rlabel metal2 s 362682 27200 362738 28400 6 la_oenb_core[123]
port 670 nsew signal output
rlabel metal2 s 364890 27200 364946 28400 6 la_oenb_core[124]
port 671 nsew signal output
rlabel metal2 s 367098 27200 367154 28400 6 la_oenb_core[125]
port 672 nsew signal output
rlabel metal2 s 369306 27200 369362 28400 6 la_oenb_core[126]
port 673 nsew signal output
rlabel metal2 s 371514 27200 371570 28400 6 la_oenb_core[127]
port 674 nsew signal output
rlabel metal2 s 117594 27200 117650 28400 6 la_oenb_core[12]
port 675 nsew signal output
rlabel metal2 s 119802 27200 119858 28400 6 la_oenb_core[13]
port 676 nsew signal output
rlabel metal2 s 122010 27200 122066 28400 6 la_oenb_core[14]
port 677 nsew signal output
rlabel metal2 s 124218 27200 124274 28400 6 la_oenb_core[15]
port 678 nsew signal output
rlabel metal2 s 126426 27200 126482 28400 6 la_oenb_core[16]
port 679 nsew signal output
rlabel metal2 s 128634 27200 128690 28400 6 la_oenb_core[17]
port 680 nsew signal output
rlabel metal2 s 130842 27200 130898 28400 6 la_oenb_core[18]
port 681 nsew signal output
rlabel metal2 s 133050 27200 133106 28400 6 la_oenb_core[19]
port 682 nsew signal output
rlabel metal2 s 93306 27200 93362 28400 6 la_oenb_core[1]
port 683 nsew signal output
rlabel metal2 s 135258 27200 135314 28400 6 la_oenb_core[20]
port 684 nsew signal output
rlabel metal2 s 137466 27200 137522 28400 6 la_oenb_core[21]
port 685 nsew signal output
rlabel metal2 s 139674 27200 139730 28400 6 la_oenb_core[22]
port 686 nsew signal output
rlabel metal2 s 141882 27200 141938 28400 6 la_oenb_core[23]
port 687 nsew signal output
rlabel metal2 s 144090 27200 144146 28400 6 la_oenb_core[24]
port 688 nsew signal output
rlabel metal2 s 146298 27200 146354 28400 6 la_oenb_core[25]
port 689 nsew signal output
rlabel metal2 s 148506 27200 148562 28400 6 la_oenb_core[26]
port 690 nsew signal output
rlabel metal2 s 150714 27200 150770 28400 6 la_oenb_core[27]
port 691 nsew signal output
rlabel metal2 s 152922 27200 152978 28400 6 la_oenb_core[28]
port 692 nsew signal output
rlabel metal2 s 155130 27200 155186 28400 6 la_oenb_core[29]
port 693 nsew signal output
rlabel metal2 s 95514 27200 95570 28400 6 la_oenb_core[2]
port 694 nsew signal output
rlabel metal2 s 157338 27200 157394 28400 6 la_oenb_core[30]
port 695 nsew signal output
rlabel metal2 s 159546 27200 159602 28400 6 la_oenb_core[31]
port 696 nsew signal output
rlabel metal2 s 161754 27200 161810 28400 6 la_oenb_core[32]
port 697 nsew signal output
rlabel metal2 s 163962 27200 164018 28400 6 la_oenb_core[33]
port 698 nsew signal output
rlabel metal2 s 166170 27200 166226 28400 6 la_oenb_core[34]
port 699 nsew signal output
rlabel metal2 s 168378 27200 168434 28400 6 la_oenb_core[35]
port 700 nsew signal output
rlabel metal2 s 170586 27200 170642 28400 6 la_oenb_core[36]
port 701 nsew signal output
rlabel metal2 s 172794 27200 172850 28400 6 la_oenb_core[37]
port 702 nsew signal output
rlabel metal2 s 175002 27200 175058 28400 6 la_oenb_core[38]
port 703 nsew signal output
rlabel metal2 s 177210 27200 177266 28400 6 la_oenb_core[39]
port 704 nsew signal output
rlabel metal2 s 97722 27200 97778 28400 6 la_oenb_core[3]
port 705 nsew signal output
rlabel metal2 s 179418 27200 179474 28400 6 la_oenb_core[40]
port 706 nsew signal output
rlabel metal2 s 181626 27200 181682 28400 6 la_oenb_core[41]
port 707 nsew signal output
rlabel metal2 s 183834 27200 183890 28400 6 la_oenb_core[42]
port 708 nsew signal output
rlabel metal2 s 186042 27200 186098 28400 6 la_oenb_core[43]
port 709 nsew signal output
rlabel metal2 s 188250 27200 188306 28400 6 la_oenb_core[44]
port 710 nsew signal output
rlabel metal2 s 190458 27200 190514 28400 6 la_oenb_core[45]
port 711 nsew signal output
rlabel metal2 s 192666 27200 192722 28400 6 la_oenb_core[46]
port 712 nsew signal output
rlabel metal2 s 194874 27200 194930 28400 6 la_oenb_core[47]
port 713 nsew signal output
rlabel metal2 s 197082 27200 197138 28400 6 la_oenb_core[48]
port 714 nsew signal output
rlabel metal2 s 199290 27200 199346 28400 6 la_oenb_core[49]
port 715 nsew signal output
rlabel metal2 s 99930 27200 99986 28400 6 la_oenb_core[4]
port 716 nsew signal output
rlabel metal2 s 201498 27200 201554 28400 6 la_oenb_core[50]
port 717 nsew signal output
rlabel metal2 s 203706 27200 203762 28400 6 la_oenb_core[51]
port 718 nsew signal output
rlabel metal2 s 205914 27200 205970 28400 6 la_oenb_core[52]
port 719 nsew signal output
rlabel metal2 s 208122 27200 208178 28400 6 la_oenb_core[53]
port 720 nsew signal output
rlabel metal2 s 210330 27200 210386 28400 6 la_oenb_core[54]
port 721 nsew signal output
rlabel metal2 s 212538 27200 212594 28400 6 la_oenb_core[55]
port 722 nsew signal output
rlabel metal2 s 214746 27200 214802 28400 6 la_oenb_core[56]
port 723 nsew signal output
rlabel metal2 s 216954 27200 217010 28400 6 la_oenb_core[57]
port 724 nsew signal output
rlabel metal2 s 219162 27200 219218 28400 6 la_oenb_core[58]
port 725 nsew signal output
rlabel metal2 s 221370 27200 221426 28400 6 la_oenb_core[59]
port 726 nsew signal output
rlabel metal2 s 102138 27200 102194 28400 6 la_oenb_core[5]
port 727 nsew signal output
rlabel metal2 s 223578 27200 223634 28400 6 la_oenb_core[60]
port 728 nsew signal output
rlabel metal2 s 225786 27200 225842 28400 6 la_oenb_core[61]
port 729 nsew signal output
rlabel metal2 s 227994 27200 228050 28400 6 la_oenb_core[62]
port 730 nsew signal output
rlabel metal2 s 230202 27200 230258 28400 6 la_oenb_core[63]
port 731 nsew signal output
rlabel metal2 s 232410 27200 232466 28400 6 la_oenb_core[64]
port 732 nsew signal output
rlabel metal2 s 234618 27200 234674 28400 6 la_oenb_core[65]
port 733 nsew signal output
rlabel metal2 s 236826 27200 236882 28400 6 la_oenb_core[66]
port 734 nsew signal output
rlabel metal2 s 239034 27200 239090 28400 6 la_oenb_core[67]
port 735 nsew signal output
rlabel metal2 s 241242 27200 241298 28400 6 la_oenb_core[68]
port 736 nsew signal output
rlabel metal2 s 243450 27200 243506 28400 6 la_oenb_core[69]
port 737 nsew signal output
rlabel metal2 s 104346 27200 104402 28400 6 la_oenb_core[6]
port 738 nsew signal output
rlabel metal2 s 245658 27200 245714 28400 6 la_oenb_core[70]
port 739 nsew signal output
rlabel metal2 s 247866 27200 247922 28400 6 la_oenb_core[71]
port 740 nsew signal output
rlabel metal2 s 250074 27200 250130 28400 6 la_oenb_core[72]
port 741 nsew signal output
rlabel metal2 s 252282 27200 252338 28400 6 la_oenb_core[73]
port 742 nsew signal output
rlabel metal2 s 254490 27200 254546 28400 6 la_oenb_core[74]
port 743 nsew signal output
rlabel metal2 s 256698 27200 256754 28400 6 la_oenb_core[75]
port 744 nsew signal output
rlabel metal2 s 258906 27200 258962 28400 6 la_oenb_core[76]
port 745 nsew signal output
rlabel metal2 s 261114 27200 261170 28400 6 la_oenb_core[77]
port 746 nsew signal output
rlabel metal2 s 263322 27200 263378 28400 6 la_oenb_core[78]
port 747 nsew signal output
rlabel metal2 s 265530 27200 265586 28400 6 la_oenb_core[79]
port 748 nsew signal output
rlabel metal2 s 106554 27200 106610 28400 6 la_oenb_core[7]
port 749 nsew signal output
rlabel metal2 s 267738 27200 267794 28400 6 la_oenb_core[80]
port 750 nsew signal output
rlabel metal2 s 269946 27200 270002 28400 6 la_oenb_core[81]
port 751 nsew signal output
rlabel metal2 s 272154 27200 272210 28400 6 la_oenb_core[82]
port 752 nsew signal output
rlabel metal2 s 274362 27200 274418 28400 6 la_oenb_core[83]
port 753 nsew signal output
rlabel metal2 s 276570 27200 276626 28400 6 la_oenb_core[84]
port 754 nsew signal output
rlabel metal2 s 278778 27200 278834 28400 6 la_oenb_core[85]
port 755 nsew signal output
rlabel metal2 s 280986 27200 281042 28400 6 la_oenb_core[86]
port 756 nsew signal output
rlabel metal2 s 283194 27200 283250 28400 6 la_oenb_core[87]
port 757 nsew signal output
rlabel metal2 s 285402 27200 285458 28400 6 la_oenb_core[88]
port 758 nsew signal output
rlabel metal2 s 287610 27200 287666 28400 6 la_oenb_core[89]
port 759 nsew signal output
rlabel metal2 s 108762 27200 108818 28400 6 la_oenb_core[8]
port 760 nsew signal output
rlabel metal2 s 289818 27200 289874 28400 6 la_oenb_core[90]
port 761 nsew signal output
rlabel metal2 s 292026 27200 292082 28400 6 la_oenb_core[91]
port 762 nsew signal output
rlabel metal2 s 294234 27200 294290 28400 6 la_oenb_core[92]
port 763 nsew signal output
rlabel metal2 s 296442 27200 296498 28400 6 la_oenb_core[93]
port 764 nsew signal output
rlabel metal2 s 298650 27200 298706 28400 6 la_oenb_core[94]
port 765 nsew signal output
rlabel metal2 s 300858 27200 300914 28400 6 la_oenb_core[95]
port 766 nsew signal output
rlabel metal2 s 303066 27200 303122 28400 6 la_oenb_core[96]
port 767 nsew signal output
rlabel metal2 s 305274 27200 305330 28400 6 la_oenb_core[97]
port 768 nsew signal output
rlabel metal2 s 307482 27200 307538 28400 6 la_oenb_core[98]
port 769 nsew signal output
rlabel metal2 s 309690 27200 309746 28400 6 la_oenb_core[99]
port 770 nsew signal output
rlabel metal2 s 110970 27200 111026 28400 6 la_oenb_core[9]
port 771 nsew signal output
rlabel metal2 s 23018 -400 23074 800 6 la_oenb_mprj[0]
port 772 nsew signal input
rlabel metal2 s 244922 -400 244978 800 6 la_oenb_mprj[100]
port 773 nsew signal input
rlabel metal2 s 247130 -400 247186 800 6 la_oenb_mprj[101]
port 774 nsew signal input
rlabel metal2 s 249338 -400 249394 800 6 la_oenb_mprj[102]
port 775 nsew signal input
rlabel metal2 s 251546 -400 251602 800 6 la_oenb_mprj[103]
port 776 nsew signal input
rlabel metal2 s 253754 -400 253810 800 6 la_oenb_mprj[104]
port 777 nsew signal input
rlabel metal2 s 255962 -400 256018 800 6 la_oenb_mprj[105]
port 778 nsew signal input
rlabel metal2 s 258170 -400 258226 800 6 la_oenb_mprj[106]
port 779 nsew signal input
rlabel metal2 s 260378 -400 260434 800 6 la_oenb_mprj[107]
port 780 nsew signal input
rlabel metal2 s 262586 -400 262642 800 6 la_oenb_mprj[108]
port 781 nsew signal input
rlabel metal2 s 264794 -400 264850 800 6 la_oenb_mprj[109]
port 782 nsew signal input
rlabel metal2 s 45098 -400 45154 800 6 la_oenb_mprj[10]
port 783 nsew signal input
rlabel metal2 s 267002 -400 267058 800 6 la_oenb_mprj[110]
port 784 nsew signal input
rlabel metal2 s 269210 -400 269266 800 6 la_oenb_mprj[111]
port 785 nsew signal input
rlabel metal2 s 271418 -400 271474 800 6 la_oenb_mprj[112]
port 786 nsew signal input
rlabel metal2 s 273626 -400 273682 800 6 la_oenb_mprj[113]
port 787 nsew signal input
rlabel metal2 s 275834 -400 275890 800 6 la_oenb_mprj[114]
port 788 nsew signal input
rlabel metal2 s 278042 -400 278098 800 6 la_oenb_mprj[115]
port 789 nsew signal input
rlabel metal2 s 280250 -400 280306 800 6 la_oenb_mprj[116]
port 790 nsew signal input
rlabel metal2 s 282458 -400 282514 800 6 la_oenb_mprj[117]
port 791 nsew signal input
rlabel metal2 s 284666 -400 284722 800 6 la_oenb_mprj[118]
port 792 nsew signal input
rlabel metal2 s 286874 -400 286930 800 6 la_oenb_mprj[119]
port 793 nsew signal input
rlabel metal2 s 47306 -400 47362 800 6 la_oenb_mprj[11]
port 794 nsew signal input
rlabel metal2 s 289082 -400 289138 800 6 la_oenb_mprj[120]
port 795 nsew signal input
rlabel metal2 s 291290 -400 291346 800 6 la_oenb_mprj[121]
port 796 nsew signal input
rlabel metal2 s 293498 -400 293554 800 6 la_oenb_mprj[122]
port 797 nsew signal input
rlabel metal2 s 295706 -400 295762 800 6 la_oenb_mprj[123]
port 798 nsew signal input
rlabel metal2 s 297914 -400 297970 800 6 la_oenb_mprj[124]
port 799 nsew signal input
rlabel metal2 s 300122 -400 300178 800 6 la_oenb_mprj[125]
port 800 nsew signal input
rlabel metal2 s 302330 -400 302386 800 6 la_oenb_mprj[126]
port 801 nsew signal input
rlabel metal2 s 304538 -400 304594 800 6 la_oenb_mprj[127]
port 802 nsew signal input
rlabel metal2 s 49514 -400 49570 800 6 la_oenb_mprj[12]
port 803 nsew signal input
rlabel metal2 s 51722 -400 51778 800 6 la_oenb_mprj[13]
port 804 nsew signal input
rlabel metal2 s 53930 -400 53986 800 6 la_oenb_mprj[14]
port 805 nsew signal input
rlabel metal2 s 56138 -400 56194 800 6 la_oenb_mprj[15]
port 806 nsew signal input
rlabel metal2 s 58346 -400 58402 800 6 la_oenb_mprj[16]
port 807 nsew signal input
rlabel metal2 s 60554 -400 60610 800 6 la_oenb_mprj[17]
port 808 nsew signal input
rlabel metal2 s 62762 -400 62818 800 6 la_oenb_mprj[18]
port 809 nsew signal input
rlabel metal2 s 64970 -400 65026 800 6 la_oenb_mprj[19]
port 810 nsew signal input
rlabel metal2 s 25226 -400 25282 800 6 la_oenb_mprj[1]
port 811 nsew signal input
rlabel metal2 s 67178 -400 67234 800 6 la_oenb_mprj[20]
port 812 nsew signal input
rlabel metal2 s 69386 -400 69442 800 6 la_oenb_mprj[21]
port 813 nsew signal input
rlabel metal2 s 71594 -400 71650 800 6 la_oenb_mprj[22]
port 814 nsew signal input
rlabel metal2 s 73802 -400 73858 800 6 la_oenb_mprj[23]
port 815 nsew signal input
rlabel metal2 s 76010 -400 76066 800 6 la_oenb_mprj[24]
port 816 nsew signal input
rlabel metal2 s 78218 -400 78274 800 6 la_oenb_mprj[25]
port 817 nsew signal input
rlabel metal2 s 80426 -400 80482 800 6 la_oenb_mprj[26]
port 818 nsew signal input
rlabel metal2 s 82634 -400 82690 800 6 la_oenb_mprj[27]
port 819 nsew signal input
rlabel metal2 s 84842 -400 84898 800 6 la_oenb_mprj[28]
port 820 nsew signal input
rlabel metal2 s 87050 -400 87106 800 6 la_oenb_mprj[29]
port 821 nsew signal input
rlabel metal2 s 27434 -400 27490 800 6 la_oenb_mprj[2]
port 822 nsew signal input
rlabel metal2 s 89258 -400 89314 800 6 la_oenb_mprj[30]
port 823 nsew signal input
rlabel metal2 s 91466 -400 91522 800 6 la_oenb_mprj[31]
port 824 nsew signal input
rlabel metal2 s 93674 -400 93730 800 6 la_oenb_mprj[32]
port 825 nsew signal input
rlabel metal2 s 95882 -400 95938 800 6 la_oenb_mprj[33]
port 826 nsew signal input
rlabel metal2 s 98090 -400 98146 800 6 la_oenb_mprj[34]
port 827 nsew signal input
rlabel metal2 s 100298 -400 100354 800 6 la_oenb_mprj[35]
port 828 nsew signal input
rlabel metal2 s 102506 -400 102562 800 6 la_oenb_mprj[36]
port 829 nsew signal input
rlabel metal2 s 104714 -400 104770 800 6 la_oenb_mprj[37]
port 830 nsew signal input
rlabel metal2 s 106922 -400 106978 800 6 la_oenb_mprj[38]
port 831 nsew signal input
rlabel metal2 s 109130 -400 109186 800 6 la_oenb_mprj[39]
port 832 nsew signal input
rlabel metal2 s 29642 -400 29698 800 6 la_oenb_mprj[3]
port 833 nsew signal input
rlabel metal2 s 111338 -400 111394 800 6 la_oenb_mprj[40]
port 834 nsew signal input
rlabel metal2 s 113546 -400 113602 800 6 la_oenb_mprj[41]
port 835 nsew signal input
rlabel metal2 s 115754 -400 115810 800 6 la_oenb_mprj[42]
port 836 nsew signal input
rlabel metal2 s 117962 -400 118018 800 6 la_oenb_mprj[43]
port 837 nsew signal input
rlabel metal2 s 120170 -400 120226 800 6 la_oenb_mprj[44]
port 838 nsew signal input
rlabel metal2 s 122378 -400 122434 800 6 la_oenb_mprj[45]
port 839 nsew signal input
rlabel metal2 s 124586 -400 124642 800 6 la_oenb_mprj[46]
port 840 nsew signal input
rlabel metal2 s 126794 -400 126850 800 6 la_oenb_mprj[47]
port 841 nsew signal input
rlabel metal2 s 129002 -400 129058 800 6 la_oenb_mprj[48]
port 842 nsew signal input
rlabel metal2 s 131210 -400 131266 800 6 la_oenb_mprj[49]
port 843 nsew signal input
rlabel metal2 s 31850 -400 31906 800 6 la_oenb_mprj[4]
port 844 nsew signal input
rlabel metal2 s 133418 -400 133474 800 6 la_oenb_mprj[50]
port 845 nsew signal input
rlabel metal2 s 135626 -400 135682 800 6 la_oenb_mprj[51]
port 846 nsew signal input
rlabel metal2 s 137834 -400 137890 800 6 la_oenb_mprj[52]
port 847 nsew signal input
rlabel metal2 s 140042 -400 140098 800 6 la_oenb_mprj[53]
port 848 nsew signal input
rlabel metal2 s 142250 -400 142306 800 6 la_oenb_mprj[54]
port 849 nsew signal input
rlabel metal2 s 144458 -400 144514 800 6 la_oenb_mprj[55]
port 850 nsew signal input
rlabel metal2 s 146666 -400 146722 800 6 la_oenb_mprj[56]
port 851 nsew signal input
rlabel metal2 s 148874 -400 148930 800 6 la_oenb_mprj[57]
port 852 nsew signal input
rlabel metal2 s 151082 -400 151138 800 6 la_oenb_mprj[58]
port 853 nsew signal input
rlabel metal2 s 153290 -400 153346 800 6 la_oenb_mprj[59]
port 854 nsew signal input
rlabel metal2 s 34058 -400 34114 800 6 la_oenb_mprj[5]
port 855 nsew signal input
rlabel metal2 s 155498 -400 155554 800 6 la_oenb_mprj[60]
port 856 nsew signal input
rlabel metal2 s 157706 -400 157762 800 6 la_oenb_mprj[61]
port 857 nsew signal input
rlabel metal2 s 159914 -400 159970 800 6 la_oenb_mprj[62]
port 858 nsew signal input
rlabel metal2 s 162122 -400 162178 800 6 la_oenb_mprj[63]
port 859 nsew signal input
rlabel metal2 s 164330 -400 164386 800 6 la_oenb_mprj[64]
port 860 nsew signal input
rlabel metal2 s 166538 -400 166594 800 6 la_oenb_mprj[65]
port 861 nsew signal input
rlabel metal2 s 168746 -400 168802 800 6 la_oenb_mprj[66]
port 862 nsew signal input
rlabel metal2 s 170954 -400 171010 800 6 la_oenb_mprj[67]
port 863 nsew signal input
rlabel metal2 s 173162 -400 173218 800 6 la_oenb_mprj[68]
port 864 nsew signal input
rlabel metal2 s 175370 -400 175426 800 6 la_oenb_mprj[69]
port 865 nsew signal input
rlabel metal2 s 36266 -400 36322 800 6 la_oenb_mprj[6]
port 866 nsew signal input
rlabel metal2 s 177578 -400 177634 800 6 la_oenb_mprj[70]
port 867 nsew signal input
rlabel metal2 s 180890 -400 180946 800 6 la_oenb_mprj[71]
port 868 nsew signal input
rlabel metal2 s 183098 -400 183154 800 6 la_oenb_mprj[72]
port 869 nsew signal input
rlabel metal2 s 185306 -400 185362 800 6 la_oenb_mprj[73]
port 870 nsew signal input
rlabel metal2 s 187514 -400 187570 800 6 la_oenb_mprj[74]
port 871 nsew signal input
rlabel metal2 s 189722 -400 189778 800 6 la_oenb_mprj[75]
port 872 nsew signal input
rlabel metal2 s 191930 -400 191986 800 6 la_oenb_mprj[76]
port 873 nsew signal input
rlabel metal2 s 194138 -400 194194 800 6 la_oenb_mprj[77]
port 874 nsew signal input
rlabel metal2 s 196346 -400 196402 800 6 la_oenb_mprj[78]
port 875 nsew signal input
rlabel metal2 s 198554 -400 198610 800 6 la_oenb_mprj[79]
port 876 nsew signal input
rlabel metal2 s 38474 -400 38530 800 6 la_oenb_mprj[7]
port 877 nsew signal input
rlabel metal2 s 200762 -400 200818 800 6 la_oenb_mprj[80]
port 878 nsew signal input
rlabel metal2 s 202970 -400 203026 800 6 la_oenb_mprj[81]
port 879 nsew signal input
rlabel metal2 s 205178 -400 205234 800 6 la_oenb_mprj[82]
port 880 nsew signal input
rlabel metal2 s 207386 -400 207442 800 6 la_oenb_mprj[83]
port 881 nsew signal input
rlabel metal2 s 209594 -400 209650 800 6 la_oenb_mprj[84]
port 882 nsew signal input
rlabel metal2 s 211802 -400 211858 800 6 la_oenb_mprj[85]
port 883 nsew signal input
rlabel metal2 s 214010 -400 214066 800 6 la_oenb_mprj[86]
port 884 nsew signal input
rlabel metal2 s 216218 -400 216274 800 6 la_oenb_mprj[87]
port 885 nsew signal input
rlabel metal2 s 218426 -400 218482 800 6 la_oenb_mprj[88]
port 886 nsew signal input
rlabel metal2 s 220634 -400 220690 800 6 la_oenb_mprj[89]
port 887 nsew signal input
rlabel metal2 s 40682 -400 40738 800 6 la_oenb_mprj[8]
port 888 nsew signal input
rlabel metal2 s 222842 -400 222898 800 6 la_oenb_mprj[90]
port 889 nsew signal input
rlabel metal2 s 225050 -400 225106 800 6 la_oenb_mprj[91]
port 890 nsew signal input
rlabel metal2 s 227258 -400 227314 800 6 la_oenb_mprj[92]
port 891 nsew signal input
rlabel metal2 s 229466 -400 229522 800 6 la_oenb_mprj[93]
port 892 nsew signal input
rlabel metal2 s 231674 -400 231730 800 6 la_oenb_mprj[94]
port 893 nsew signal input
rlabel metal2 s 233882 -400 233938 800 6 la_oenb_mprj[95]
port 894 nsew signal input
rlabel metal2 s 236090 -400 236146 800 6 la_oenb_mprj[96]
port 895 nsew signal input
rlabel metal2 s 238298 -400 238354 800 6 la_oenb_mprj[97]
port 896 nsew signal input
rlabel metal2 s 240506 -400 240562 800 6 la_oenb_mprj[98]
port 897 nsew signal input
rlabel metal2 s 242714 -400 242770 800 6 la_oenb_mprj[99]
port 898 nsew signal input
rlabel metal2 s 42890 -400 42946 800 6 la_oenb_mprj[9]
port 899 nsew signal input
rlabel metal2 s 305090 -400 305146 800 6 mprj_ack_i_core
port 900 nsew signal output
rlabel metal2 s 13082 27200 13138 28400 6 mprj_ack_i_user
port 901 nsew signal input
rlabel metal2 s 307298 -400 307354 800 6 mprj_adr_o_core[0]
port 902 nsew signal input
rlabel metal2 s 326066 -400 326122 800 6 mprj_adr_o_core[10]
port 903 nsew signal input
rlabel metal2 s 327722 -400 327778 800 6 mprj_adr_o_core[11]
port 904 nsew signal input
rlabel metal2 s 329378 -400 329434 800 6 mprj_adr_o_core[12]
port 905 nsew signal input
rlabel metal2 s 331034 -400 331090 800 6 mprj_adr_o_core[13]
port 906 nsew signal input
rlabel metal2 s 332690 -400 332746 800 6 mprj_adr_o_core[14]
port 907 nsew signal input
rlabel metal2 s 334346 -400 334402 800 6 mprj_adr_o_core[15]
port 908 nsew signal input
rlabel metal2 s 336002 -400 336058 800 6 mprj_adr_o_core[16]
port 909 nsew signal input
rlabel metal2 s 337658 -400 337714 800 6 mprj_adr_o_core[17]
port 910 nsew signal input
rlabel metal2 s 339314 -400 339370 800 6 mprj_adr_o_core[18]
port 911 nsew signal input
rlabel metal2 s 340970 -400 341026 800 6 mprj_adr_o_core[19]
port 912 nsew signal input
rlabel metal2 s 309506 -400 309562 800 6 mprj_adr_o_core[1]
port 913 nsew signal input
rlabel metal2 s 342626 -400 342682 800 6 mprj_adr_o_core[20]
port 914 nsew signal input
rlabel metal2 s 344282 -400 344338 800 6 mprj_adr_o_core[21]
port 915 nsew signal input
rlabel metal2 s 345938 -400 345994 800 6 mprj_adr_o_core[22]
port 916 nsew signal input
rlabel metal2 s 347594 -400 347650 800 6 mprj_adr_o_core[23]
port 917 nsew signal input
rlabel metal2 s 349250 -400 349306 800 6 mprj_adr_o_core[24]
port 918 nsew signal input
rlabel metal2 s 350906 -400 350962 800 6 mprj_adr_o_core[25]
port 919 nsew signal input
rlabel metal2 s 352562 -400 352618 800 6 mprj_adr_o_core[26]
port 920 nsew signal input
rlabel metal2 s 354218 -400 354274 800 6 mprj_adr_o_core[27]
port 921 nsew signal input
rlabel metal2 s 355874 -400 355930 800 6 mprj_adr_o_core[28]
port 922 nsew signal input
rlabel metal2 s 357530 -400 357586 800 6 mprj_adr_o_core[29]
port 923 nsew signal input
rlabel metal2 s 311714 -400 311770 800 6 mprj_adr_o_core[2]
port 924 nsew signal input
rlabel metal2 s 359186 -400 359242 800 6 mprj_adr_o_core[30]
port 925 nsew signal input
rlabel metal2 s 360842 -400 360898 800 6 mprj_adr_o_core[31]
port 926 nsew signal input
rlabel metal2 s 313922 -400 313978 800 6 mprj_adr_o_core[3]
port 927 nsew signal input
rlabel metal2 s 316130 -400 316186 800 6 mprj_adr_o_core[4]
port 928 nsew signal input
rlabel metal2 s 317786 -400 317842 800 6 mprj_adr_o_core[5]
port 929 nsew signal input
rlabel metal2 s 319442 -400 319498 800 6 mprj_adr_o_core[6]
port 930 nsew signal input
rlabel metal2 s 321098 -400 321154 800 6 mprj_adr_o_core[7]
port 931 nsew signal input
rlabel metal2 s 322754 -400 322810 800 6 mprj_adr_o_core[8]
port 932 nsew signal input
rlabel metal2 s 324410 -400 324466 800 6 mprj_adr_o_core[9]
port 933 nsew signal input
rlabel metal2 s 16026 27200 16082 28400 6 mprj_adr_o_user[0]
port 934 nsew signal output
rlabel metal2 s 41050 27200 41106 28400 6 mprj_adr_o_user[10]
port 935 nsew signal output
rlabel metal2 s 43258 27200 43314 28400 6 mprj_adr_o_user[11]
port 936 nsew signal output
rlabel metal2 s 45466 27200 45522 28400 6 mprj_adr_o_user[12]
port 937 nsew signal output
rlabel metal2 s 47674 27200 47730 28400 6 mprj_adr_o_user[13]
port 938 nsew signal output
rlabel metal2 s 49882 27200 49938 28400 6 mprj_adr_o_user[14]
port 939 nsew signal output
rlabel metal2 s 52090 27200 52146 28400 6 mprj_adr_o_user[15]
port 940 nsew signal output
rlabel metal2 s 54298 27200 54354 28400 6 mprj_adr_o_user[16]
port 941 nsew signal output
rlabel metal2 s 56506 27200 56562 28400 6 mprj_adr_o_user[17]
port 942 nsew signal output
rlabel metal2 s 58714 27200 58770 28400 6 mprj_adr_o_user[18]
port 943 nsew signal output
rlabel metal2 s 60922 27200 60978 28400 6 mprj_adr_o_user[19]
port 944 nsew signal output
rlabel metal2 s 18970 27200 19026 28400 6 mprj_adr_o_user[1]
port 945 nsew signal output
rlabel metal2 s 63130 27200 63186 28400 6 mprj_adr_o_user[20]
port 946 nsew signal output
rlabel metal2 s 65338 27200 65394 28400 6 mprj_adr_o_user[21]
port 947 nsew signal output
rlabel metal2 s 67546 27200 67602 28400 6 mprj_adr_o_user[22]
port 948 nsew signal output
rlabel metal2 s 69754 27200 69810 28400 6 mprj_adr_o_user[23]
port 949 nsew signal output
rlabel metal2 s 71962 27200 72018 28400 6 mprj_adr_o_user[24]
port 950 nsew signal output
rlabel metal2 s 74170 27200 74226 28400 6 mprj_adr_o_user[25]
port 951 nsew signal output
rlabel metal2 s 76378 27200 76434 28400 6 mprj_adr_o_user[26]
port 952 nsew signal output
rlabel metal2 s 78586 27200 78642 28400 6 mprj_adr_o_user[27]
port 953 nsew signal output
rlabel metal2 s 80794 27200 80850 28400 6 mprj_adr_o_user[28]
port 954 nsew signal output
rlabel metal2 s 83002 27200 83058 28400 6 mprj_adr_o_user[29]
port 955 nsew signal output
rlabel metal2 s 21914 27200 21970 28400 6 mprj_adr_o_user[2]
port 956 nsew signal output
rlabel metal2 s 85210 27200 85266 28400 6 mprj_adr_o_user[30]
port 957 nsew signal output
rlabel metal2 s 87418 27200 87474 28400 6 mprj_adr_o_user[31]
port 958 nsew signal output
rlabel metal2 s 24858 27200 24914 28400 6 mprj_adr_o_user[3]
port 959 nsew signal output
rlabel metal2 s 27802 27200 27858 28400 6 mprj_adr_o_user[4]
port 960 nsew signal output
rlabel metal2 s 30010 27200 30066 28400 6 mprj_adr_o_user[5]
port 961 nsew signal output
rlabel metal2 s 32218 27200 32274 28400 6 mprj_adr_o_user[6]
port 962 nsew signal output
rlabel metal2 s 34426 27200 34482 28400 6 mprj_adr_o_user[7]
port 963 nsew signal output
rlabel metal2 s 36634 27200 36690 28400 6 mprj_adr_o_user[8]
port 964 nsew signal output
rlabel metal2 s 38842 27200 38898 28400 6 mprj_adr_o_user[9]
port 965 nsew signal output
rlabel metal2 s 305642 -400 305698 800 6 mprj_cyc_o_core
port 966 nsew signal input
rlabel metal2 s 13818 27200 13874 28400 6 mprj_cyc_o_user
port 967 nsew signal output
rlabel metal2 s 307850 -400 307906 800 6 mprj_dat_i_core[0]
port 968 nsew signal output
rlabel metal2 s 326618 -400 326674 800 6 mprj_dat_i_core[10]
port 969 nsew signal output
rlabel metal2 s 328274 -400 328330 800 6 mprj_dat_i_core[11]
port 970 nsew signal output
rlabel metal2 s 329930 -400 329986 800 6 mprj_dat_i_core[12]
port 971 nsew signal output
rlabel metal2 s 331586 -400 331642 800 6 mprj_dat_i_core[13]
port 972 nsew signal output
rlabel metal2 s 333242 -400 333298 800 6 mprj_dat_i_core[14]
port 973 nsew signal output
rlabel metal2 s 334898 -400 334954 800 6 mprj_dat_i_core[15]
port 974 nsew signal output
rlabel metal2 s 336554 -400 336610 800 6 mprj_dat_i_core[16]
port 975 nsew signal output
rlabel metal2 s 338210 -400 338266 800 6 mprj_dat_i_core[17]
port 976 nsew signal output
rlabel metal2 s 339866 -400 339922 800 6 mprj_dat_i_core[18]
port 977 nsew signal output
rlabel metal2 s 341522 -400 341578 800 6 mprj_dat_i_core[19]
port 978 nsew signal output
rlabel metal2 s 310058 -400 310114 800 6 mprj_dat_i_core[1]
port 979 nsew signal output
rlabel metal2 s 343178 -400 343234 800 6 mprj_dat_i_core[20]
port 980 nsew signal output
rlabel metal2 s 344834 -400 344890 800 6 mprj_dat_i_core[21]
port 981 nsew signal output
rlabel metal2 s 346490 -400 346546 800 6 mprj_dat_i_core[22]
port 982 nsew signal output
rlabel metal2 s 348146 -400 348202 800 6 mprj_dat_i_core[23]
port 983 nsew signal output
rlabel metal2 s 349802 -400 349858 800 6 mprj_dat_i_core[24]
port 984 nsew signal output
rlabel metal2 s 351458 -400 351514 800 6 mprj_dat_i_core[25]
port 985 nsew signal output
rlabel metal2 s 353114 -400 353170 800 6 mprj_dat_i_core[26]
port 986 nsew signal output
rlabel metal2 s 354770 -400 354826 800 6 mprj_dat_i_core[27]
port 987 nsew signal output
rlabel metal2 s 356426 -400 356482 800 6 mprj_dat_i_core[28]
port 988 nsew signal output
rlabel metal2 s 358082 -400 358138 800 6 mprj_dat_i_core[29]
port 989 nsew signal output
rlabel metal2 s 312266 -400 312322 800 6 mprj_dat_i_core[2]
port 990 nsew signal output
rlabel metal2 s 359738 -400 359794 800 6 mprj_dat_i_core[30]
port 991 nsew signal output
rlabel metal2 s 361394 -400 361450 800 6 mprj_dat_i_core[31]
port 992 nsew signal output
rlabel metal2 s 314474 -400 314530 800 6 mprj_dat_i_core[3]
port 993 nsew signal output
rlabel metal2 s 316682 -400 316738 800 6 mprj_dat_i_core[4]
port 994 nsew signal output
rlabel metal2 s 318338 -400 318394 800 6 mprj_dat_i_core[5]
port 995 nsew signal output
rlabel metal2 s 319994 -400 320050 800 6 mprj_dat_i_core[6]
port 996 nsew signal output
rlabel metal2 s 321650 -400 321706 800 6 mprj_dat_i_core[7]
port 997 nsew signal output
rlabel metal2 s 323306 -400 323362 800 6 mprj_dat_i_core[8]
port 998 nsew signal output
rlabel metal2 s 324962 -400 325018 800 6 mprj_dat_i_core[9]
port 999 nsew signal output
rlabel metal2 s 16762 27200 16818 28400 6 mprj_dat_i_user[0]
port 1000 nsew signal input
rlabel metal2 s 41786 27200 41842 28400 6 mprj_dat_i_user[10]
port 1001 nsew signal input
rlabel metal2 s 43994 27200 44050 28400 6 mprj_dat_i_user[11]
port 1002 nsew signal input
rlabel metal2 s 46202 27200 46258 28400 6 mprj_dat_i_user[12]
port 1003 nsew signal input
rlabel metal2 s 48410 27200 48466 28400 6 mprj_dat_i_user[13]
port 1004 nsew signal input
rlabel metal2 s 50618 27200 50674 28400 6 mprj_dat_i_user[14]
port 1005 nsew signal input
rlabel metal2 s 52826 27200 52882 28400 6 mprj_dat_i_user[15]
port 1006 nsew signal input
rlabel metal2 s 55034 27200 55090 28400 6 mprj_dat_i_user[16]
port 1007 nsew signal input
rlabel metal2 s 57242 27200 57298 28400 6 mprj_dat_i_user[17]
port 1008 nsew signal input
rlabel metal2 s 59450 27200 59506 28400 6 mprj_dat_i_user[18]
port 1009 nsew signal input
rlabel metal2 s 61658 27200 61714 28400 6 mprj_dat_i_user[19]
port 1010 nsew signal input
rlabel metal2 s 19706 27200 19762 28400 6 mprj_dat_i_user[1]
port 1011 nsew signal input
rlabel metal2 s 63866 27200 63922 28400 6 mprj_dat_i_user[20]
port 1012 nsew signal input
rlabel metal2 s 66074 27200 66130 28400 6 mprj_dat_i_user[21]
port 1013 nsew signal input
rlabel metal2 s 68282 27200 68338 28400 6 mprj_dat_i_user[22]
port 1014 nsew signal input
rlabel metal2 s 70490 27200 70546 28400 6 mprj_dat_i_user[23]
port 1015 nsew signal input
rlabel metal2 s 72698 27200 72754 28400 6 mprj_dat_i_user[24]
port 1016 nsew signal input
rlabel metal2 s 74906 27200 74962 28400 6 mprj_dat_i_user[25]
port 1017 nsew signal input
rlabel metal2 s 77114 27200 77170 28400 6 mprj_dat_i_user[26]
port 1018 nsew signal input
rlabel metal2 s 79322 27200 79378 28400 6 mprj_dat_i_user[27]
port 1019 nsew signal input
rlabel metal2 s 81530 27200 81586 28400 6 mprj_dat_i_user[28]
port 1020 nsew signal input
rlabel metal2 s 83738 27200 83794 28400 6 mprj_dat_i_user[29]
port 1021 nsew signal input
rlabel metal2 s 22650 27200 22706 28400 6 mprj_dat_i_user[2]
port 1022 nsew signal input
rlabel metal2 s 85946 27200 86002 28400 6 mprj_dat_i_user[30]
port 1023 nsew signal input
rlabel metal2 s 88154 27200 88210 28400 6 mprj_dat_i_user[31]
port 1024 nsew signal input
rlabel metal2 s 25594 27200 25650 28400 6 mprj_dat_i_user[3]
port 1025 nsew signal input
rlabel metal2 s 28538 27200 28594 28400 6 mprj_dat_i_user[4]
port 1026 nsew signal input
rlabel metal2 s 30746 27200 30802 28400 6 mprj_dat_i_user[5]
port 1027 nsew signal input
rlabel metal2 s 32954 27200 33010 28400 6 mprj_dat_i_user[6]
port 1028 nsew signal input
rlabel metal2 s 35162 27200 35218 28400 6 mprj_dat_i_user[7]
port 1029 nsew signal input
rlabel metal2 s 37370 27200 37426 28400 6 mprj_dat_i_user[8]
port 1030 nsew signal input
rlabel metal2 s 39578 27200 39634 28400 6 mprj_dat_i_user[9]
port 1031 nsew signal input
rlabel metal2 s 308402 -400 308458 800 6 mprj_dat_o_core[0]
port 1032 nsew signal input
rlabel metal2 s 327170 -400 327226 800 6 mprj_dat_o_core[10]
port 1033 nsew signal input
rlabel metal2 s 328826 -400 328882 800 6 mprj_dat_o_core[11]
port 1034 nsew signal input
rlabel metal2 s 330482 -400 330538 800 6 mprj_dat_o_core[12]
port 1035 nsew signal input
rlabel metal2 s 332138 -400 332194 800 6 mprj_dat_o_core[13]
port 1036 nsew signal input
rlabel metal2 s 333794 -400 333850 800 6 mprj_dat_o_core[14]
port 1037 nsew signal input
rlabel metal2 s 335450 -400 335506 800 6 mprj_dat_o_core[15]
port 1038 nsew signal input
rlabel metal2 s 337106 -400 337162 800 6 mprj_dat_o_core[16]
port 1039 nsew signal input
rlabel metal2 s 338762 -400 338818 800 6 mprj_dat_o_core[17]
port 1040 nsew signal input
rlabel metal2 s 340418 -400 340474 800 6 mprj_dat_o_core[18]
port 1041 nsew signal input
rlabel metal2 s 342074 -400 342130 800 6 mprj_dat_o_core[19]
port 1042 nsew signal input
rlabel metal2 s 310610 -400 310666 800 6 mprj_dat_o_core[1]
port 1043 nsew signal input
rlabel metal2 s 343730 -400 343786 800 6 mprj_dat_o_core[20]
port 1044 nsew signal input
rlabel metal2 s 345386 -400 345442 800 6 mprj_dat_o_core[21]
port 1045 nsew signal input
rlabel metal2 s 347042 -400 347098 800 6 mprj_dat_o_core[22]
port 1046 nsew signal input
rlabel metal2 s 348698 -400 348754 800 6 mprj_dat_o_core[23]
port 1047 nsew signal input
rlabel metal2 s 350354 -400 350410 800 6 mprj_dat_o_core[24]
port 1048 nsew signal input
rlabel metal2 s 352010 -400 352066 800 6 mprj_dat_o_core[25]
port 1049 nsew signal input
rlabel metal2 s 353666 -400 353722 800 6 mprj_dat_o_core[26]
port 1050 nsew signal input
rlabel metal2 s 355322 -400 355378 800 6 mprj_dat_o_core[27]
port 1051 nsew signal input
rlabel metal2 s 356978 -400 357034 800 6 mprj_dat_o_core[28]
port 1052 nsew signal input
rlabel metal2 s 358634 -400 358690 800 6 mprj_dat_o_core[29]
port 1053 nsew signal input
rlabel metal2 s 312818 -400 312874 800 6 mprj_dat_o_core[2]
port 1054 nsew signal input
rlabel metal2 s 360290 -400 360346 800 6 mprj_dat_o_core[30]
port 1055 nsew signal input
rlabel metal2 s 361946 -400 362002 800 6 mprj_dat_o_core[31]
port 1056 nsew signal input
rlabel metal2 s 315026 -400 315082 800 6 mprj_dat_o_core[3]
port 1057 nsew signal input
rlabel metal2 s 317234 -400 317290 800 6 mprj_dat_o_core[4]
port 1058 nsew signal input
rlabel metal2 s 318890 -400 318946 800 6 mprj_dat_o_core[5]
port 1059 nsew signal input
rlabel metal2 s 320546 -400 320602 800 6 mprj_dat_o_core[6]
port 1060 nsew signal input
rlabel metal2 s 322202 -400 322258 800 6 mprj_dat_o_core[7]
port 1061 nsew signal input
rlabel metal2 s 323858 -400 323914 800 6 mprj_dat_o_core[8]
port 1062 nsew signal input
rlabel metal2 s 325514 -400 325570 800 6 mprj_dat_o_core[9]
port 1063 nsew signal input
rlabel metal2 s 17498 27200 17554 28400 6 mprj_dat_o_user[0]
port 1064 nsew signal output
rlabel metal2 s 42522 27200 42578 28400 6 mprj_dat_o_user[10]
port 1065 nsew signal output
rlabel metal2 s 44730 27200 44786 28400 6 mprj_dat_o_user[11]
port 1066 nsew signal output
rlabel metal2 s 46938 27200 46994 28400 6 mprj_dat_o_user[12]
port 1067 nsew signal output
rlabel metal2 s 49146 27200 49202 28400 6 mprj_dat_o_user[13]
port 1068 nsew signal output
rlabel metal2 s 51354 27200 51410 28400 6 mprj_dat_o_user[14]
port 1069 nsew signal output
rlabel metal2 s 53562 27200 53618 28400 6 mprj_dat_o_user[15]
port 1070 nsew signal output
rlabel metal2 s 55770 27200 55826 28400 6 mprj_dat_o_user[16]
port 1071 nsew signal output
rlabel metal2 s 57978 27200 58034 28400 6 mprj_dat_o_user[17]
port 1072 nsew signal output
rlabel metal2 s 60186 27200 60242 28400 6 mprj_dat_o_user[18]
port 1073 nsew signal output
rlabel metal2 s 62394 27200 62450 28400 6 mprj_dat_o_user[19]
port 1074 nsew signal output
rlabel metal2 s 20442 27200 20498 28400 6 mprj_dat_o_user[1]
port 1075 nsew signal output
rlabel metal2 s 64602 27200 64658 28400 6 mprj_dat_o_user[20]
port 1076 nsew signal output
rlabel metal2 s 66810 27200 66866 28400 6 mprj_dat_o_user[21]
port 1077 nsew signal output
rlabel metal2 s 69018 27200 69074 28400 6 mprj_dat_o_user[22]
port 1078 nsew signal output
rlabel metal2 s 71226 27200 71282 28400 6 mprj_dat_o_user[23]
port 1079 nsew signal output
rlabel metal2 s 73434 27200 73490 28400 6 mprj_dat_o_user[24]
port 1080 nsew signal output
rlabel metal2 s 75642 27200 75698 28400 6 mprj_dat_o_user[25]
port 1081 nsew signal output
rlabel metal2 s 77850 27200 77906 28400 6 mprj_dat_o_user[26]
port 1082 nsew signal output
rlabel metal2 s 80058 27200 80114 28400 6 mprj_dat_o_user[27]
port 1083 nsew signal output
rlabel metal2 s 82266 27200 82322 28400 6 mprj_dat_o_user[28]
port 1084 nsew signal output
rlabel metal2 s 84474 27200 84530 28400 6 mprj_dat_o_user[29]
port 1085 nsew signal output
rlabel metal2 s 23386 27200 23442 28400 6 mprj_dat_o_user[2]
port 1086 nsew signal output
rlabel metal2 s 86682 27200 86738 28400 6 mprj_dat_o_user[30]
port 1087 nsew signal output
rlabel metal2 s 88890 27200 88946 28400 6 mprj_dat_o_user[31]
port 1088 nsew signal output
rlabel metal2 s 26330 27200 26386 28400 6 mprj_dat_o_user[3]
port 1089 nsew signal output
rlabel metal2 s 29274 27200 29330 28400 6 mprj_dat_o_user[4]
port 1090 nsew signal output
rlabel metal2 s 31482 27200 31538 28400 6 mprj_dat_o_user[5]
port 1091 nsew signal output
rlabel metal2 s 33690 27200 33746 28400 6 mprj_dat_o_user[6]
port 1092 nsew signal output
rlabel metal2 s 35898 27200 35954 28400 6 mprj_dat_o_user[7]
port 1093 nsew signal output
rlabel metal2 s 38106 27200 38162 28400 6 mprj_dat_o_user[8]
port 1094 nsew signal output
rlabel metal2 s 40314 27200 40370 28400 6 mprj_dat_o_user[9]
port 1095 nsew signal output
rlabel metal2 s 362498 -400 362554 800 6 mprj_iena_wb
port 1096 nsew signal input
rlabel metal2 s 308954 -400 309010 800 6 mprj_sel_o_core[0]
port 1097 nsew signal input
rlabel metal2 s 311162 -400 311218 800 6 mprj_sel_o_core[1]
port 1098 nsew signal input
rlabel metal2 s 313370 -400 313426 800 6 mprj_sel_o_core[2]
port 1099 nsew signal input
rlabel metal2 s 315578 -400 315634 800 6 mprj_sel_o_core[3]
port 1100 nsew signal input
rlabel metal2 s 18234 27200 18290 28400 6 mprj_sel_o_user[0]
port 1101 nsew signal output
rlabel metal2 s 21178 27200 21234 28400 6 mprj_sel_o_user[1]
port 1102 nsew signal output
rlabel metal2 s 24122 27200 24178 28400 6 mprj_sel_o_user[2]
port 1103 nsew signal output
rlabel metal2 s 27066 27200 27122 28400 6 mprj_sel_o_user[3]
port 1104 nsew signal output
rlabel metal2 s 306194 -400 306250 800 6 mprj_stb_o_core
port 1105 nsew signal input
rlabel metal2 s 14554 27200 14610 28400 6 mprj_stb_o_user
port 1106 nsew signal output
rlabel metal2 s 306746 -400 306802 800 6 mprj_we_o_core
port 1107 nsew signal input
rlabel metal2 s 15290 27200 15346 28400 6 mprj_we_o_user
port 1108 nsew signal output
rlabel metal3 s 383200 9120 384400 9240 6 user1_vcc_powergood
port 1109 nsew signal output
rlabel metal3 s 383200 11024 384400 11144 6 user1_vdd_powergood
port 1110 nsew signal output
rlabel metal3 s 383200 12928 384400 13048 6 user2_vcc_powergood
port 1111 nsew signal output
rlabel metal3 s 383200 14832 384400 14952 6 user2_vdd_powergood
port 1112 nsew signal output
rlabel metal2 s 11610 27200 11666 28400 6 user_clock
port 1113 nsew signal output
rlabel metal2 s 372250 27200 372306 28400 6 user_clock2
port 1114 nsew signal output
rlabel metal3 s 383200 16736 384400 16856 6 user_irq[0]
port 1115 nsew signal output
rlabel metal3 s 383200 18640 384400 18760 6 user_irq[1]
port 1116 nsew signal output
rlabel metal3 s 383200 20544 384400 20664 6 user_irq[2]
port 1117 nsew signal output
rlabel metal3 s 383200 1504 384400 1624 6 user_irq_core[0]
port 1118 nsew signal input
rlabel metal3 s 383200 3408 384400 3528 6 user_irq_core[1]
port 1119 nsew signal input
rlabel metal3 s 383200 5312 384400 5432 6 user_irq_core[2]
port 1120 nsew signal input
rlabel metal3 s 383200 22448 384400 22568 6 user_irq_ena[0]
port 1121 nsew signal input
rlabel metal3 s 383200 24352 384400 24472 6 user_irq_ena[1]
port 1122 nsew signal input
rlabel metal3 s 383200 26256 384400 26376 6 user_irq_ena[2]
port 1123 nsew signal input
rlabel metal2 s 12346 27200 12402 28400 6 user_reset
port 1124 nsew signal output
rlabel metal4 s 5014 1040 5194 26704 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 20064 1040 20244 26704 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 35114 1040 35294 26704 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 50164 1040 50344 26704 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 65214 1040 65394 26704 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 80264 1040 80444 26704 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 95314 1040 95494 26704 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 110364 1040 110544 26704 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 125414 1040 125594 26704 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 140464 1040 140644 26704 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 155514 1040 155694 26704 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 170564 1040 170744 26704 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 185614 1040 185794 26704 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 200664 1040 200844 26704 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 215714 1040 215894 26704 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 230764 1040 230944 26704 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 245814 1040 245994 26704 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 260864 1040 261044 26704 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 275914 1040 276094 26704 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 290964 1040 291144 26704 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 306014 1040 306194 26704 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 321064 1040 321244 26704 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 336114 1040 336294 26704 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 351164 1040 351344 26704 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 366214 1040 366394 26704 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 381264 1040 381444 26704 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 141284 1040 141464 26704 6 vccd1
port 1126 nsew power bidirectional
rlabel metal4 s 156334 1040 156514 26704 6 vccd1
port 1126 nsew power bidirectional
rlabel metal4 s 171384 1040 171564 26704 6 vccd1
port 1126 nsew power bidirectional
rlabel metal4 s 186434 1040 186614 26704 6 vccd1
port 1126 nsew power bidirectional
rlabel metal4 s 66854 1040 67034 26704 6 vccd2
port 1127 nsew power bidirectional
rlabel metal4 s 76854 1040 77034 26704 6 vccd2
port 1127 nsew power bidirectional
rlabel metal4 s 255814 1040 255994 26704 6 vdda1
port 1128 nsew power bidirectional
rlabel metal4 s 270864 1040 271044 26704 6 vdda1
port 1128 nsew power bidirectional
rlabel metal4 s 256614 1040 256794 26704 6 vdda2
port 1129 nsew power bidirectional
rlabel metal4 s 271664 1040 271844 26704 6 vdda2
port 1129 nsew power bidirectional
rlabel metal4 s 263194 1040 263374 26704 6 vssa1
port 1130 nsew ground bidirectional
rlabel metal4 s 278244 1040 278424 26704 6 vssa1
port 1130 nsew ground bidirectional
rlabel metal4 s 263994 1040 264174 26704 6 vssa2
port 1131 nsew ground bidirectional
rlabel metal4 s 279044 1040 279224 26704 6 vssa2
port 1131 nsew ground bidirectional
rlabel metal4 s 12394 1040 12574 26704 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 27444 1040 27624 26704 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 42494 1040 42674 26704 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 57544 1040 57724 26704 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 72594 1040 72774 26704 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 87644 1040 87824 26704 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 102694 1040 102874 26704 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 117744 1040 117924 26704 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 132794 1040 132974 26704 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 147844 1040 148024 26704 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 162894 1040 163074 26704 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 177944 1040 178124 26704 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 192994 1040 193174 26704 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 208044 1040 208224 26704 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 223094 1040 223274 26704 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 238144 1040 238324 26704 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 253194 1040 253374 26704 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 268244 1040 268424 26704 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 283294 1040 283474 26704 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 298344 1040 298524 26704 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 313394 1040 313574 26704 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 328444 1040 328624 26704 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 343494 1040 343674 26704 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 358544 1040 358724 26704 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 373594 1040 373774 26704 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 148664 1040 148844 26704 6 vssd1
port 1133 nsew ground bidirectional
rlabel metal4 s 163714 1040 163894 26704 6 vssd1
port 1133 nsew ground bidirectional
rlabel metal4 s 178764 1040 178944 26704 6 vssd1
port 1133 nsew ground bidirectional
rlabel metal4 s 193814 1040 193994 26704 6 vssd1
port 1133 nsew ground bidirectional
rlabel metal4 s 71034 1040 71214 26704 6 vssd2
port 1134 nsew ground bidirectional
rlabel metal4 s 81034 1040 81214 26704 6 vssd2
port 1134 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 384000 28000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 17673590
string GDS_FILE /home/hosni/caravel_sky130/caravel/openlane/mgmt_protect/runs/23_02_07_02_42/results/signoff/mgmt_protect.magic.gds
string GDS_START 723546
<< end >>

