* NGSPICE file created from caravel_openframe.ext - technology: sky130A

.subckt sky130_fd_io__com_ctl_ls_octl VCC_IO VPB OUT_H_N OUT_H IN RST_H SET_H HLD_H_N
+ a_992_934# a_181_1305# a_n17_1379#
X0 a_361_1391# a_181_1305# a_128_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X1 VCC_IO a_130_181# OUT_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X2 a_128_1391# a_181_1305# a_361_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X3 a_n17_1379# a_634_829# a_128_1391# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 a_128_1391# a_634_829# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.15
X5 a_361_1391# HLD_H_N a_130_181# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.6
X6 a_634_829# a_992_934# a_181_1305# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.25
X7 a_361_1391# a_181_1305# a_128_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X8 a_n17_1379# a_634_829# a_128_1391# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9 OUT_H_N a_65_861# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X10 a_n17_1379# a_992_934# a_724_1391# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11 a_128_1391# a_634_829# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 a_724_1391# a_992_934# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13 a_65_861# HLD_H_N a_957_1391# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X14 OUT_H a_130_181# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.28 pd=2.56 as=0.14 ps=1.28 w=1 l=0.6
X15 a_n17_1379# a_992_934# a_724_1391# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X16 a_65_861# a_130_181# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.199 ps=2.03 w=0.75 l=0.5
X17 a_724_1391# a_992_934# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X18 a_n17_1379# a_65_861# a_130_181# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.199 ps=2.03 w=0.75 l=1
X19 a_181_1305# IN a_992_934# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.25
X20 a_957_1391# a_181_1305# a_724_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X21 a_n17_1379# IN a_992_934# a_n17_1379# sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.25
X22 a_n17_1379# a_65_861# OUT_H_N a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.6
X23 a_130_181# a_65_861# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.199 ps=2.03 w=0.75 l=0.5
X24 a_724_1391# a_181_1305# a_957_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X25 a_957_1391# a_181_1305# a_724_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X26 a_65_861# a_130_181# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.105 ps=1.03 w=0.75 l=1
X27 a_634_829# a_992_934# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8 ad=0.28 pd=2.56 as=0.14 ps=1.28 w=1 l=0.25
X28 a_130_181# SET_H a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X29 a_724_1391# a_181_1305# a_957_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X30 a_n17_1379# RST_H a_65_861# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X31 a_128_1391# a_181_1305# a_361_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
.ends

.subckt sky130_fd_io__gpiov2_octl DM_H[1] DM_H[0] DM_H[2] DM_H_N[0] DM_H_N[1] DM_H_N[2]
+ PUEN_2OR1_H PDEN_H_N[1] PDEN_H_N[0] SLOW SLOW_H VCC_IO a_n8755_2384# a_n9051_2020#
+ w_n9346_2317# a_n9227_2020# a_n9283_2046# a_5840_3586# m1_n8913_3102# VPWR a_n8875_2020#
+ a_4338_3622# a_3924_6676# a_n8931_2384# a_4514_3388# SLOW_H_N VGND a_5813_4576#
+ HLD_I_H_N OD_H
Xsky130_fd_io__com_ctl_ls_octl_0 VCC_IO VPWR SLOW_H_N SLOW_H SLOW OD_H VGND HLD_I_H_N
+ m2_5755_2254# VPWR VGND sky130_fd_io__com_ctl_ls_octl
X0 a_4667_4619# a_3966_4619# a_4491_4619# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X1 a_5720_3560# a_5315_3924# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X2 VCC_IO DM_H[2] a_3933_3414# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X3 a_4282_3414# DM_H[2] VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X4 VCC_IO DM_H_N[0] a_4520_6066# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X5 a_3871_7368# a_3924_6676# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X6 a_n8755_2384# a_n9280_2384# a_n8755_2046# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X7 a_n9107_2384# a_n9227_2020# a_n9280_2384# w_n9346_2317# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X8 a_4634_3414# a_4514_3388# a_4458_3414# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X9 a_4872_6702# DM_H_N[2] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X10 VCC_IO DM_H[2] a_3966_4619# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X11 a_4996_5728# a_4520_6066# PUEN_2OR1_H VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.185 ps=1.93 w=0.7 l=0.6
X12 VCC_IO a_4347_7368# a_5651_5728# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X13 VCC_IO a_5052_5702# PUEN_2OR1_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X14 a_5488_3924# DM_H_N[1] a_5315_3924# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X15 a_5813_4576# a_5693_4550# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X16 VCC_IO a_5720_3560# a_5840_3586# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X17 VCC_IO DM_H[0] a_5052_5702# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X18 a_4282_3816# DM_H[2] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X19 VCC_IO DM_H_N[0] a_5175_7368# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X20 a_4634_3816# a_3933_3414# a_4458_3414# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X21 a_4491_4619# a_4371_4587# a_4315_4619# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X22 a_5513_4576# a_3871_7368# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.6
X23 PDEN_H_N[1] a_5651_6702# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X24 a_5315_3924# DM_H_N[1] VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.196 ps=1.96 w=0.7 l=0.6
X25 VCC_IO DM_H[1] a_4667_4619# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X26 a_n8931_2384# a_n9051_2020# a_n9107_2384# w_n9346_2317# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X27 a_4044_6066# DM_H_N[1] a_3871_6066# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X28 a_n8755_2046# a_n8875_2020# a_n9283_2046# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X29 PDEN_H_N[0] a_5651_5728# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X30 a_4520_6066# a_3871_6066# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X31 a_4347_7368# DM_H[0] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X32 a_n8931_2384# a_n9280_2384# a_n8755_2384# w_n9346_2317# sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X33 VCC_IO a_4458_3414# a_5488_3924# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X34 a_5513_4576# a_3871_7368# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.185 ps=1.93 w=0.7 l=0.6
X35 a_4371_4587# DM_H[1] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X36 VGND a_4458_3414# a_5315_3924# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X37 VCC_IO a_5693_4550# a_5813_4576# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X38 a_4338_3622# DM_H[0] VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X39 PUEN_2OR1_H a_4520_6066# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X40 VGND PUEN_2OR1_H a_4044_7368# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X41 PDEN_H_N[1] a_5651_6702# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X42 a_5348_7368# a_4872_6702# a_5175_7368# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.185 ps=1.93 w=0.7 l=0.6
X43 VCC_IO DM_H_N[0] a_4520_6066# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X44 VGND a_5651_6702# PDEN_H_N[1] VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X45 VCC_IO DM_H[1] a_4347_7368# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X46 VCC_IO DM_H_N[1] a_4872_6702# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X47 a_n8755_2384# a_n8875_2020# a_n8931_2384# w_n9346_2317# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X48 a_5840_3586# a_5720_3560# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X49 a_4458_3414# a_4338_3622# a_4282_3816# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X50 a_4315_5349# DM_H[2] VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X51 VCC_IO a_5175_7368# a_5651_6702# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X52 VCC_IO a_4347_7368# a_5651_5728# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X53 a_4338_3622# DM_H[0] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X54 VGND a_5693_4550# a_5813_4576# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X55 a_4667_5349# a_4371_4587# a_4491_4619# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X56 VGND DM_H_N[2] a_3871_6066# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X57 a_5813_4576# a_5693_4550# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X58 a_5840_3586# a_5720_3560# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X59 a_5348_5728# a_4491_4619# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X60 VGND a_5651_5728# PDEN_H_N[0] VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X61 VGND a_3933_3414# a_4634_3414# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X62 a_4315_4619# DM_H[2] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X63 a_5693_4550# a_5513_4576# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X64 a_4667_4619# a_3966_4619# a_4491_4619# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X65 PDEN_H_N[0] a_5651_5728# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X66 a_4044_6066# DM_H_N[1] a_3871_6066# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X67 VGND DM_H_N[0] a_5348_7368# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X68 a_3871_7368# a_3924_6676# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X69 a_4872_6702# DM_H_N[2] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X70 VCC_IO a_5720_3560# a_5840_3586# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X71 a_4282_3816# DM_H[2] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X72 VCC_IO DM_H[0] a_4634_3816# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X73 VCC_IO PUEN_2OR1_H a_3871_7368# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X74 a_4634_3816# a_3933_3414# a_4458_3414# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X75 a_5813_4576# a_5693_4550# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.185 ps=1.93 w=0.7 l=0.6
X76 a_4491_4619# DM_H[1] a_4315_5349# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X77 a_n9280_2384# a_n9227_2020# a_n9283_2046# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.196 ps=1.96 w=0.7 l=0.6
X78 VGND a_3966_4619# a_4667_5349# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X79 VGND a_5052_5702# a_4996_5728# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X80 a_5175_7368# a_4872_6702# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X81 VGND a_5720_3560# a_5840_3586# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X82 VCC_IO a_5651_6702# PDEN_H_N[1] VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X83 a_n8931_2384# a_n9280_2384# a_n8755_2384# w_n9346_2317# sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X84 a_5052_5702# DM_H[0] a_5348_5728# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X85 VGND DM_H[2] a_3933_3414# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.185 ps=1.93 w=0.7 l=0.6
X86 a_4491_4619# a_4371_4587# a_4315_4619# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X87 a_5720_3560# a_5315_3924# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X88 VCC_IO DM_H[1] a_4667_4619# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X89 a_4520_7368# DM_H[0] a_4347_7368# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.185 ps=1.93 w=0.7 l=0.6
X90 VCC_IO DM_H[2] a_3966_4619# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X91 PUEN_2OR1_H a_4520_6066# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X92 VCC_IO DM_H[2] a_3933_3414# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X93 VCC_IO DM_H_N[2] a_4044_6066# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X94 a_n9283_2046# a_n9051_2020# a_n9280_2384# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X95 a_4371_4587# DM_H[1] VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X96 a_5052_5702# a_4491_4619# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X97 a_4520_5728# a_3871_6066# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.185 ps=1.93 w=0.7 l=0.6
X98 VCC_IO a_5651_5728# PDEN_H_N[0] VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X99 VCC_IO DM_H_N[0] a_5175_7368# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X100 a_n8755_2384# a_n8875_2020# a_n8931_2384# w_n9346_2317# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X101 a_5488_3924# DM_H_N[1] a_5315_3924# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X102 a_4371_4587# DM_H[1] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X103 a_n9107_2384# a_n9227_2020# a_n9280_2384# w_n9346_2317# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X104 VGND DM_H[1] a_4520_7368# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X105 a_4872_6702# DM_H_N[1] a_4872_7368# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X106 VGND a_5175_7368# a_5651_6702# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.185 ps=1.93 w=0.7 l=0.6
X107 a_5693_4550# a_5513_4576# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X108 PDEN_H_N[0] a_5651_5728# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X109 PDEN_H_N[1] a_5651_6702# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X110 a_4338_3622# DM_H[0] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X111 VCC_IO a_5052_5702# PUEN_2OR1_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X112 a_4347_7368# DM_H[0] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X113 a_4520_6066# DM_H_N[0] a_4520_5728# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X114 VCC_IO DM_H[0] a_5052_5702# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X115 a_5513_4576# a_3871_7368# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.6
X116 VGND a_4347_7368# a_5651_5728# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.185 ps=1.93 w=0.7 l=0.6
X117 VCC_IO a_4458_3414# a_5488_3924# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X118 a_n8931_2384# a_n9051_2020# a_n9107_2384# w_n9346_2317# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X119 a_4044_7368# a_3924_6676# a_3871_7368# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.185 ps=1.93 w=0.7 l=0.6
X120 a_4872_7368# DM_H_N[2] VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X121 a_5693_4550# a_5513_4576# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X122 VCC_IO DM_H[0] a_4634_3816# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X123 a_4458_3414# DM_H[0] a_4282_3414# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X124 a_4520_6066# a_3871_6066# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X125 VCC_IO DM_H[1] a_4347_7368# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X126 a_3871_6066# DM_H_N[1] VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.196 ps=1.96 w=0.7 l=0.6
X127 VCC_IO DM_H_N[1] a_4872_6702# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X128 VCC_IO a_5175_7368# a_5651_6702# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X129 VCC_IO DM_H_N[2] a_4044_6066# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X130 VCC_IO PUEN_2OR1_H a_3871_7368# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X131 a_5052_5702# a_4491_4619# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X132 a_5720_3560# a_5315_3924# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X133 a_5840_3586# a_5720_3560# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X134 VCC_IO a_5693_4550# a_5813_4576# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X135 a_5175_7368# a_4872_6702# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X136 VCC_IO a_5651_5728# PDEN_H_N[0] VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X137 a_4458_3414# a_4338_3622# a_4282_3816# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X138 VCC_IO a_5651_6702# PDEN_H_N[1] VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X139 a_4315_4619# DM_H[2] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X140 VGND DM_H[2] a_3966_4619# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.185 ps=1.93 w=0.7 l=0.6
.ends

.subckt sky130_fd_io__gpio_dat_ls_1v2 IN OUT_H_N RST_H SET_H HLD_H_N VCC_IO VGND OUT_H
+ VPWR_KA
X0 a_2251_36# a_2251_2228# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.25
X1 a_28_633# SET_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X2 a_1720_1202# HLD_H_N a_28_14# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=10.5 as=1.33 ps=10.5 w=5 l=0.5
X3 a_1251_128# VPWR_KA a_1484_128# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X4 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.9
X5 a_2080_128# a_2251_2228# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X6 a_1484_128# VPWR_KA a_1251_128# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X7 VGND a_2251_2228# a_2080_128# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X8 a_1484_128# a_2251_36# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X9 VGND a_2251_36# a_1484_128# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X10 VPWR_KA a_2251_2228# a_2251_36# VPWR_KA sky130_fd_pr__pfet_01v8_hvt ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.25
X11 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.9
X12 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.9
X13 a_1251_128# VPWR_KA a_1484_128# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X14 a_28_633# a_28_14# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.5
X15 VGND IN a_2251_2228# VGND sky130_fd_pr__nfet_01v8 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.25
X16 OUT_H a_28_633# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.5
X17 a_1484_128# a_2251_36# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X18 a_2080_128# a_2251_2228# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X19 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.9
X20 a_1251_128# VPWR_KA a_1484_128# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X21 a_1484_128# VPWR_KA a_1251_128# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X22 VGND a_2251_36# a_1484_128# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X23 a_1484_128# a_2251_36# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X24 VGND a_28_633# OUT_H VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.6
X25 VGND a_2251_2228# a_2080_128# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X26 a_2251_2228# IN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.25
X27 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.9
X28 a_1484_128# VPWR_KA a_1251_128# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X29 VGND a_2251_36# a_1484_128# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X30 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.9
X31 a_2251_2228# IN VPWR_KA VPWR_KA sky130_fd_pr__pfet_01v8_hvt ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.25
X32 VGND a_28_633# a_28_14# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.185 ps=1.93 w=0.7 l=0.6
X33 a_2080_128# a_2251_2228# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X34 a_1484_128# VPWR_KA a_1251_128# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X35 VGND a_2251_36# a_1484_128# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X36 VGND a_2251_2228# a_2251_36# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.25
X37 a_28_633# a_28_14# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X38 VGND a_2251_2228# a_2080_128# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X39 a_28_14# a_28_633# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.5
X40 a_1251_128# VPWR_KA a_1484_128# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X41 a_1251_128# HLD_H_N a_28_633# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.6 as=1.33 ps=10.5 w=5 l=0.5
X42 VCC_IO a_28_14# OUT_H_N VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X43 a_1484_128# a_2251_36# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X44 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.9
X45 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.9
X46 VGND RST_H a_28_14# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X47 OUT_H_N a_28_14# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.28 pd=2.56 as=0.14 ps=1.28 w=1 l=0.6
X48 a_2080_128# a_2251_2228# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X49 VGND a_2251_2228# a_2080_128# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_io__gpio_dat_lsv2 IN OUT_H_N RST_H SET_H HLD_H_N VCC_IO VGND OUT_H
+ VPWR_KA a_28_14#
X0 a_2251_36# a_2251_2228# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.25
X1 a_28_633# SET_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X2 a_1720_1202# HLD_H_N a_28_14# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=10.5 as=1.33 ps=10.5 w=5 l=0.5
X3 a_1251_128# VPWR_KA a_1484_128# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X4 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.9
X5 a_2080_128# a_2251_2228# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X6 a_1484_128# VPWR_KA a_1251_128# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X7 VGND a_2251_2228# a_2080_128# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X8 a_1484_128# a_2251_36# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X9 VGND a_2251_36# a_1484_128# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X10 VPWR_KA a_2251_2228# a_2251_36# VPWR_KA sky130_fd_pr__pfet_01v8_hvt ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.25
X11 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.9
X12 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.9
X13 a_1251_128# VPWR_KA a_1484_128# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X14 a_28_633# a_28_14# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.5
X15 VGND IN a_2251_2228# VGND sky130_fd_pr__nfet_01v8 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.25
X16 OUT_H a_28_633# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.5
X17 a_1484_128# a_2251_36# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X18 a_2080_128# a_2251_2228# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X19 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.9
X20 a_1251_128# VPWR_KA a_1484_128# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X21 a_1484_128# VPWR_KA a_1251_128# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X22 VGND a_2251_36# a_1484_128# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X23 a_1484_128# a_2251_36# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X24 VGND a_28_633# OUT_H VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.6
X25 VGND a_2251_2228# a_2080_128# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X26 a_2251_2228# IN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.25
X27 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.9
X28 a_1484_128# VPWR_KA a_1251_128# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X29 VGND a_2251_36# a_1484_128# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X30 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.9
X31 a_2251_2228# IN VPWR_KA VPWR_KA sky130_fd_pr__pfet_01v8_hvt ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.25
X32 VGND a_28_633# a_28_14# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.185 ps=1.93 w=0.7 l=0.6
X33 a_2080_128# a_2251_2228# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X34 a_1484_128# VPWR_KA a_1251_128# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X35 VGND a_2251_36# a_1484_128# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X36 VGND a_2251_2228# a_2251_36# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.25
X37 a_28_633# a_28_14# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X38 VGND a_2251_2228# a_2080_128# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X39 a_28_14# a_28_633# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.5
X40 a_1251_128# VPWR_KA a_1484_128# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X41 a_1251_128# HLD_H_N a_28_633# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.6 as=1.33 ps=10.5 w=5 l=0.5
X42 VCC_IO a_28_14# OUT_H_N VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X43 a_1484_128# a_2251_36# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X44 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.9
X45 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.9
X46 VGND RST_H a_28_14# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X47 OUT_H_N a_28_14# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.28 pd=2.56 as=0.14 ps=1.28 w=1 l=0.6
X48 a_2080_128# a_2251_2228# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X49 VGND a_2251_2228# a_2080_128# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_io__com_cclat PU_DIS_H PD_DIS_H VGND OE_H_N DRVHI_H VCC_IO DRVLO_H_N
X0 a_947_1193# DRVLO_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.5
X1 VCC_IO a_505_1193# a_3417_1193# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.6
X2 VCC_IO a_505_1193# a_3417_1193# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.6
X3 a_3417_1193# DRVHI_H a_4762_1193# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X4 a_4762_1193# DRVHI_H a_3417_1193# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X5 VGND DRVHI_H a_2361_1095# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X6 VCC_IO PU_DIS_H a_638_279# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.5
X7 VCC_IO a_2361_1095# DRVLO_H_N VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X8 DRVLO_H_N a_2361_1095# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X9 DRVHI_H a_947_1193# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X10 a_2361_1095# DRVHI_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X11 VCC_IO a_947_1193# DRVHI_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X12 DRVLO_H_N a_2361_1095# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X13 VCC_IO a_2361_1095# DRVLO_H_N VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X14 DRVHI_H a_947_1193# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.5
X15 VCC_IO a_947_1193# DRVHI_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X16 VGND PU_DIS_H a_638_279# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X17 a_4762_1193# DRVHI_H a_3417_1193# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X18 a_2361_1095# PD_DIS_H a_4762_1193# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X19 VGND PD_DIS_H a_2361_1095# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X20 a_505_1193# a_176_279# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.5
X21 VCC_IO a_638_279# a_947_1193# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X22 a_3417_1193# DRVHI_H a_4762_1193# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.5
X23 a_2361_1095# PD_DIS_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X24 VGND a_947_1193# DRVHI_H VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X25 DRVLO_H_N a_2361_1095# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X26 VGND a_947_1193# DRVHI_H VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X27 a_987_279# a_176_279# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X28 DRVHI_H a_947_1193# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X29 a_4762_1193# PD_DIS_H a_2361_1095# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X30 DRVHI_H a_947_1193# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X31 VCC_IO OE_H_N a_176_279# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.5
X32 a_3417_1193# a_505_1193# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.6
X33 a_2361_1095# PD_DIS_H a_4762_1193# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X34 a_987_279# DRVLO_H_N a_1628_279# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X35 VGND a_2361_1095# DRVLO_H_N VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X36 DRVHI_H a_947_1193# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X37 a_947_1193# a_176_279# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X38 VGND OE_H_N a_176_279# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X39 VCC_IO a_947_1193# DRVHI_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X40 VCC_IO a_2361_1095# DRVLO_H_N VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X41 DRVLO_H_N a_2361_1095# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X42 VCC_IO a_505_1193# a_3417_1193# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.6
X43 DRVHI_H a_947_1193# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X44 VCC_IO a_505_1193# a_3417_1193# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.6
X45 a_4762_1193# PD_DIS_H a_2361_1095# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.5
X46 VGND a_176_279# a_987_279# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X47 VGND a_947_1193# DRVHI_H VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X48 a_947_1193# a_638_279# a_1628_279# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X49 VGND a_2361_1095# DRVLO_H_N VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X50 DRVLO_H_N a_2361_1095# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X51 a_1628_279# DRVLO_H_N a_987_279# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X52 a_3417_1193# a_505_1193# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.6
X53 a_505_1193# a_176_279# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X54 DRVLO_H_N a_2361_1095# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X55 VGND a_505_1193# a_2361_1095# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X56 a_3417_1193# a_505_1193# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.6
X57 VGND a_176_279# a_987_279# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X58 a_3417_1193# a_505_1193# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.6
X59 VGND a_2361_1095# DRVLO_H_N VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X60 a_2361_1095# a_505_1193# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X61 a_987_279# a_176_279# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X62 a_1628_279# a_638_279# a_947_1193# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
.ends

.subckt sky130_fd_io__com_opath_datoev2 OE_H DRVLO_H_N VCC_IO HLD_I_OVR_H a_5565_99#
+ OUT OE_N sky130_fd_io__com_cclat_0/PD_DIS_H VPWR_KA DRVHI_H li_5565_99# sky130_fd_io__gpio_dat_ls_1v2_0/SET_H
+ VGND OD_H
Xsky130_fd_io__gpio_dat_ls_1v2_0 OUT sky130_fd_io__com_cclat_0/PU_DIS_H VGND sky130_fd_io__gpio_dat_ls_1v2_0/SET_H
+ HLD_I_OVR_H VCC_IO VGND sky130_fd_io__com_cclat_0/PD_DIS_H VPWR_KA sky130_fd_io__gpio_dat_ls_1v2
Xsky130_fd_io__gpio_dat_lsv2_0 OE_N OE_H VGND OD_H HLD_I_OVR_H VCC_IO VGND sky130_fd_io__com_cclat_0/OE_H_N
+ VPWR_KA a_28_1762# sky130_fd_io__gpio_dat_lsv2
Xsky130_fd_io__com_cclat_0 sky130_fd_io__com_cclat_0/PU_DIS_H sky130_fd_io__com_cclat_0/PD_DIS_H
+ VGND sky130_fd_io__com_cclat_0/OE_H_N DRVHI_H VCC_IO DRVLO_H_N sky130_fd_io__com_cclat
.ends

.subckt sky130_fd_io__com_pdpredrvr_weakv2 DRVLO_H_N PDEN_H_N VGND_IO VCC_IO PD_H
X0 PD_H DRVLO_H_N a_73_866# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X1 a_73_866# PDEN_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X2 PD_H PDEN_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X3 VGND_IO DRVLO_H_N PD_H VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X4 VCC_IO PDEN_H_N a_73_866# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
.ends

.subckt sky130_fd_io__gpiov2_octl_mux SEL_H_N A_H Y_H B_H SEL_H a_1266_1185# w_1191_2415#
X0 Y_H SEL_H A_H a_1266_1185# sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X1 A_H SEL_H_N Y_H w_1191_2415# sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.5
X2 Y_H SEL_H B_H w_1191_2415# sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X3 B_H SEL_H_N Y_H a_1266_1185# sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.5
.ends

.subckt sky130_fd_io__gpiov2_pdpredrvr_strong sky130_fd_io__gpiov2_octl_mux_0/SEL_H
+ sky130_fd_io__gpiov2_octl_mux_0/B_H sky130_fd_io__gpiov2_octl_mux_0/SEL_H_N sky130_fd_io__gpiov2_octl_mux_0/w_1191_2415#
+ sky130_fd_io__gpiov2_octl_mux_0/A_H sky130_fd_io__gpiov2_octl_mux_0/Y_H VSUBS
Xsky130_fd_io__gpiov2_octl_mux_0 sky130_fd_io__gpiov2_octl_mux_0/SEL_H_N sky130_fd_io__gpiov2_octl_mux_0/A_H
+ sky130_fd_io__gpiov2_octl_mux_0/Y_H sky130_fd_io__gpiov2_octl_mux_0/B_H sky130_fd_io__gpiov2_octl_mux_0/SEL_H
+ VSUBS sky130_fd_io__gpiov2_octl_mux_0/w_1191_2415# sky130_fd_io__gpiov2_octl_mux
.ends

.subckt sky130_fd_io__feascom_pupredrvr_nbiasv2 EN_H EN_H_N VGND_IO DRVHI_H NBIAS
+ PUEN_H VCC_IO PU_H_N a_261_220# a_2821_220# a_2874_118# a_1772_220#
X0 VCC_IO DRVHI_H a_207_1014# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.192 pd=1.38 as=0.14 ps=1.28 w=1 l=0.5
X1 VCC_IO a_250_1898# a_1507_1397# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.8
X2 VGND_IO a_261_220# a_261_220# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X3 a_1507_1397# a_250_1898# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.8
X4 a_261_220# a_261_220# VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X5 a_1672_194# a_207_1014# VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.5
X6 NBIAS a_250_1898# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.192 ps=1.38 w=1 l=0.8
X7 a_250_1898# a_562_1898# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X8 VGND_IO a_1672_194# a_1772_220# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
R0 a_562_1898# m1_2838_1831# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R1 m1_1014_127# NBIAS sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X9 VCC_IO a_250_1898# a_2874_118# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.5
X10 NBIAS NBIAS a_261_220# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
R2 m1_1014_800# NBIAS sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X11 VGND_IO a_1672_194# a_1772_220# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
R3 m1_575_1252# EN_H sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X12 VCC_IO DRVHI_H a_562_1898# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.185 pd=1.51 as=0.14 ps=1.28 w=1 l=0.5
X13 a_261_220# a_261_220# VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
R4 m1_2838_1794# a_620_1263# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R5 m1_612_1252# a_620_1263# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X14 a_250_1898# DRVHI_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.5
X15 VGND_IO DRVHI_H a_207_1014# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.324 pd=2.02 as=0.265 ps=2.53 w=1 l=0.6
X16 VGND_IO a_207_1014# NBIAS VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X17 VGND_IO a_250_1898# a_1004_990# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=4
X18 NBIAS NBIAS a_261_220# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
R6 m1_1409_1332# NBIAS sky130_fd_pr__res_generic_m1 w=0.23 l=10m
X19 VCC_IO a_250_1898# NBIAS VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.8
X20 a_2874_118# a_250_1898# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.04 ps=5.51 w=5 l=0.5
X21 a_583_914# EN_H VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.203 pd=1.77 as=0.324 ps=2.02 w=1.5 l=0.5
X22 a_2821_220# a_2874_118# a_2874_118# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
R7 m1_1608_646# a_1772_220# sky130_fd_pr__res_generic_m1 w=0.23 l=10m
X23 a_1772_220# a_1672_194# VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X24 NBIAS a_250_1898# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.8
X25 a_207_1014# DRVHI_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.5
X26 a_250_1898# a_562_1898# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
R8 m1_2596_1928# a_2421_2014# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X27 a_261_220# NBIAS NBIAS VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X28 NBIAS EN_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X29 VCC_IO a_250_1898# a_1507_1397# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.8
X30 VCC_IO a_562_1898# a_250_1898# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=1.04 pd=5.51 as=0.42 ps=3.28 w=3 l=0.5
X31 a_1772_220# a_1672_194# VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X32 a_2821_220# a_2821_220# a_1672_194# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.5
R9 m1_2596_1928# a_250_1898# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R10 m1_702_1715# PU_H_N sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R11 m1_1409_1332# a_1507_1397# sky130_fd_pr__res_generic_m1 w=0.23 l=10m
X33 a_1507_1397# a_250_1898# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.8
R12 m1_1046_126# a_261_220# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X34 VCC_IO EN_H a_250_1898# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.5
X35 a_562_1898# PUEN_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.5
X36 a_2421_2014# PU_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.185 ps=1.51 w=0.42 l=8
X37 a_737_914# a_620_1263# a_583_914# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.203 pd=1.77 as=0.203 ps=1.77 w=1.5 l=0.5
R13 a_620_1263# m1_702_1715# sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R14 m1_1014_800# a_1004_990# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X38 VCC_IO a_250_1898# NBIAS VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.8
X39 a_261_220# NBIAS NBIAS VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.5
X40 VGND_IO a_261_220# a_261_220# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
R15 m1_1608_646# a_261_220# sky130_fd_pr__res_generic_m1 w=0.23 l=10m
X41 VCC_IO a_562_1898# a_250_1898# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X42 a_250_1898# DRVHI_H a_737_914# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.203 ps=1.77 w=1.5 l=0.5
X43 a_1672_194# a_2821_220# a_2821_220# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X44 a_562_1898# a_620_1263# a_620_1263# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.5
X45 a_1672_194# VCC_IO VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=8
X46 a_2874_118# a_2874_118# a_2821_220# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
.ends

.subckt sky130_fd_io__gpiov2_pupredrvr_strong_nd2 DRVHI_H PUEN_H EN_FAST[0] EN_FAST[1]
+ EN_FAST[2] EN_FAST[3] VGND_IO VCC_IO PU_H_N a_158_632#
R0 PU_H_N m1_1184_866# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X0 VCC_IO DRVHI_H PU_H_N VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.6
X1 a_311_632# DRVHI_H a_158_632# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.157 pd=1.71 as=0.398 ps=3.53 w=1.5 l=0.5
X2 VGND_IO EN_FAST[3] a_311_632# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.157 ps=1.71 w=1.5 l=1
R1 m1_1184_866# a_158_632# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X3 PU_H_N DRVHI_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.6
X4 PU_H_N PUEN_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.6
X5 VCC_IO DRVHI_H PU_H_N VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.6
R2 a_1008_2434# PU_H_N sky130_fd_pr__res_generic_po w=0.33 l=4
X6 a_158_632# DRVHI_H a_809_1060# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.165 ps=1.72 w=1.5 l=0.5
R3 a_1008_2434# a_158_632# sky130_fd_pr__res_generic_po w=0.33 l=11
X7 a_809_632# EN_FAST[2] VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.165 pd=1.72 as=0.21 ps=1.78 w=1.5 l=1
X8 a_158_632# DRVHI_H a_809_632# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.165 ps=1.72 w=1.5 l=0.5
X9 a_311_1060# DRVHI_H a_158_632# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.157 pd=1.71 as=0.398 ps=3.53 w=1.5 l=0.5
X10 VGND_IO EN_FAST[0] a_311_1060# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.157 ps=1.71 w=1.5 l=1
X11 PU_H_N DRVHI_H a_158_109# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.111 ps=1.37 w=0.42 l=4
X12 VGND_IO PUEN_H a_158_109# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.111 ps=1.37 w=0.42 l=4
X13 a_809_1060# EN_FAST[1] VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.165 pd=1.72 as=0.21 ps=1.78 w=1.5 l=1
.ends

.subckt sky130_fd_io__gpiov2_pupredrvr_strong_nd2_a DRVHI_H PUEN_H EN_FAST[0] EN_FAST[1]
+ EN_FAST[2] EN_FAST[3] VGND_IO VCC_IO PU_H_N a_353_606# a_609_606#
R0 PU_H_N m1_1184_866# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X0 VCC_IO DRVHI_H PU_H_N VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.6
X1 a_311_632# DRVHI_H a_158_632# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.157 pd=1.71 as=0.398 ps=3.53 w=1.5 l=0.5
X2 VGND_IO a_353_606# a_311_632# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.157 ps=1.71 w=1.5 l=1
X3 VGND_IO PUEN_H a_158_199# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.111 ps=1.37 w=0.42 l=4
R1 m1_1184_866# a_158_632# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X4 PU_H_N DRVHI_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.6
X5 PU_H_N PUEN_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.6
X6 VCC_IO DRVHI_H PU_H_N VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.6
R2 a_1008_2434# PU_H_N sky130_fd_pr__res_generic_po w=0.33 l=4
X7 a_158_632# DRVHI_H a_809_1060# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.165 ps=1.72 w=1.5 l=0.5
R3 a_1008_2434# a_158_632# sky130_fd_pr__res_generic_po w=0.33 l=11
X8 a_809_632# a_609_606# VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.165 pd=1.72 as=0.21 ps=1.78 w=1.5 l=1
X9 a_158_632# DRVHI_H a_809_632# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.165 ps=1.72 w=1.5 l=0.5
X10 a_311_1060# DRVHI_H a_158_632# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.157 pd=1.71 as=0.398 ps=3.53 w=1.5 l=0.5
X11 VGND_IO EN_FAST[0] a_311_1060# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.157 ps=1.71 w=1.5 l=1
X12 PU_H_N DRVHI_H a_158_199# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.111 ps=1.37 w=0.42 l=4
X13 a_809_1060# EN_FAST[1] VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.165 pd=1.72 as=0.21 ps=1.78 w=1.5 l=1
.ends

.subckt sky130_fd_io__gpio_pupredrvr_strongv2 VCC_IO PU_H_N[3] PU_H_N[2] SLOW_H_N
+ sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_1772_220# sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/a_158_632#
+ sky130_fd_io__feascom_pupredrvr_nbiasv2_0/NBIAS sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_261_220#
+ sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2821_220# PUEN_H DRVHI_H sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2874_118#
+ VSUBS
Xsky130_fd_io__feascom_pupredrvr_nbiasv2_0 sky130_fd_io__feascom_pupredrvr_nbiasv2_0/EN_H
+ sky130_fd_io__feascom_pupredrvr_nbiasv2_0/EN_H_N VSUBS DRVHI_H sky130_fd_io__feascom_pupredrvr_nbiasv2_0/NBIAS
+ PUEN_H VCC_IO PU_H_N[2] sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_261_220# sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2821_220#
+ sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2874_118# sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_1772_220#
+ sky130_fd_io__feascom_pupredrvr_nbiasv2
Xsky130_fd_io__gpiov2_pupredrvr_strong_nd2_0 DRVHI_H PUEN_H sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/EN_FAST[0]
+ sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/EN_FAST[1] sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/EN_FAST[2]
+ sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/EN_FAST[3] VSUBS VCC_IO PU_H_N[3] sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/a_158_632#
+ sky130_fd_io__gpiov2_pupredrvr_strong_nd2
Xsky130_fd_io__gpiov2_pupredrvr_strong_nd2_a_0 DRVHI_H PUEN_H sky130_fd_io__gpiov2_pupredrvr_strong_nd2_a_0/EN_FAST[3]
+ sky130_fd_io__gpiov2_pupredrvr_strong_nd2_a_0/EN_FAST[3] sky130_fd_io__gpiov2_pupredrvr_strong_nd2_a_0/EN_FAST[3]
+ sky130_fd_io__gpiov2_pupredrvr_strong_nd2_a_0/EN_FAST[3] VSUBS VCC_IO PU_H_N[2]
+ sky130_fd_io__gpiov2_pupredrvr_strong_nd2_a_0/EN_FAST[3] sky130_fd_io__gpiov2_pupredrvr_strong_nd2_a_0/EN_FAST[3]
+ sky130_fd_io__gpiov2_pupredrvr_strong_nd2_a
R0 m1_6556_1365# sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/EN_FAST[0] sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R1 m1_6555_1273# VSUBS sky130_fd_pr__res_generic_m1 w=0.65 l=10m
X0 VCC_IO PUEN_H sky130_fd_io__feascom_pupredrvr_nbiasv2_0/EN_H_N VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
R2 sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/EN_FAST[1] m1_6299_1273# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R3 VSUBS m1_6266_605# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R4 m1_5759_509# sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/EN_FAST[3] sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X1 sky130_fd_io__feascom_pupredrvr_nbiasv2_0/EN_H_N SLOW_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
R5 m1_4777_1326# sky130_fd_io__gpiov2_pupredrvr_strong_nd2_a_0/EN_FAST[3] sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R6 m1_5786_421# sky130_fd_io__feascom_pupredrvr_nbiasv2_0/NBIAS sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R7 m1_4655_1468# sky130_fd_io__gpiov2_pupredrvr_strong_nd2_a_0/EN_FAST[3] sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R8 m1_6266_568# sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/EN_FAST[2] sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R9 sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/EN_FAST[3] m1_5786_421# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R10 sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/EN_FAST[3] m1_6300_1402# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
X2 sky130_fd_io__feascom_pupredrvr_nbiasv2_0/EN_H sky130_fd_io__feascom_pupredrvr_nbiasv2_0/EN_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
R11 sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/EN_FAST[2] m1_6265_477# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R12 m1_5722_509# sky130_fd_io__feascom_pupredrvr_nbiasv2_0/EN_H sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R13 m1_6299_1273# VSUBS sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R14 m1_6300_1365# sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/EN_FAST[1] sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R15 sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/EN_FAST[0] m1_6555_1273# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R16 m1_6265_477# sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/EN_FAST[3] sky130_fd_pr__res_generic_m1 w=0.65 l=10m
X3 VSUBS PUEN_H a_483_1179# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X4 a_483_1179# SLOW_H_N sky130_fd_io__feascom_pupredrvr_nbiasv2_0/EN_H_N VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X5 sky130_fd_io__feascom_pupredrvr_nbiasv2_0/EN_H sky130_fd_io__feascom_pupredrvr_nbiasv2_0/EN_H_N VSUBS VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
R17 m1_4740_1326# sky130_fd_io__feascom_pupredrvr_nbiasv2_0/EN_H sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R18 sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/EN_FAST[3] m1_6556_1402# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R19 m1_4655_1468# sky130_fd_io__feascom_pupredrvr_nbiasv2_0/NBIAS sky130_fd_pr__res_generic_m1 w=0.26 l=10m
.ends

.subckt sky130_fd_io__gpiov2_obpredrvr sky130_fd_io__gpio_pupredrvr_strongv2_0/SLOW_H_N
+ sky130_fd_io__com_pdpredrvr_weakv2_0/PDEN_H_N sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_261_220#
+ sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/SEL_H_N
+ sky130_fd_io__com_pdpredrvr_weakv2_0/VCC_IO sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2821_220#
+ sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2874_118#
+ sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/A_H sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/Y_H
+ sky130_fd_io__gpio_pupredrvr_strongv2_0/PUEN_H sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/SEL_H
+ sky130_fd_io__com_pdpredrvr_weakv2_0/PD_H sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_1772_220#
+ sky130_fd_io__gpio_pupredrvr_strongv2_0/DRVHI_H sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/a_158_632#
+ sky130_fd_io__gpio_pupredrvr_strongv2_0/PU_H_N[2] sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/w_1191_2415#
+ sky130_fd_io__gpio_pupredrvr_strongv2_0/PU_H_N[3] sky130_fd_io__com_pdpredrvr_weakv2_0/DRVLO_H_N
+ sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/B_H sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/NBIAS
+ VSUBS sky130_fd_io__gpio_pupredrvr_strongv2_0/VCC_IO
Xsky130_fd_io__com_pdpredrvr_weakv2_0 sky130_fd_io__com_pdpredrvr_weakv2_0/DRVLO_H_N
+ sky130_fd_io__com_pdpredrvr_weakv2_0/PDEN_H_N VSUBS sky130_fd_io__com_pdpredrvr_weakv2_0/VCC_IO
+ sky130_fd_io__com_pdpredrvr_weakv2_0/PD_H sky130_fd_io__com_pdpredrvr_weakv2
Xsky130_fd_io__gpiov2_pdpredrvr_strong_0 sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/SEL_H
+ sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/B_H sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/SEL_H_N
+ sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/w_1191_2415#
+ sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/A_H sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/Y_H
+ VSUBS sky130_fd_io__gpiov2_pdpredrvr_strong
Xsky130_fd_io__gpio_pupredrvr_strongv2_0 sky130_fd_io__gpio_pupredrvr_strongv2_0/VCC_IO
+ sky130_fd_io__gpio_pupredrvr_strongv2_0/PU_H_N[3] sky130_fd_io__gpio_pupredrvr_strongv2_0/PU_H_N[2]
+ sky130_fd_io__gpio_pupredrvr_strongv2_0/SLOW_H_N sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_1772_220#
+ sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/a_158_632#
+ sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/NBIAS
+ sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_261_220#
+ sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2821_220#
+ sky130_fd_io__gpio_pupredrvr_strongv2_0/PUEN_H sky130_fd_io__gpio_pupredrvr_strongv2_0/DRVHI_H
+ sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2874_118#
+ VSUBS sky130_fd_io__gpio_pupredrvr_strongv2
.ends

.subckt sky130_fd_io__gpiov2_octl_dat VPWR_KA SLOW HLD_I_OVR_H OD_H SLOW_H_N DRVHI_H
+ PU_H_N[2] PU_H_N[1] PU_H_N[0] PD_H[1] PD_H[0] PD_H[4] PD_H[3] PD_H[2] a_1106_3203#
+ a_3125_3203# a_4416_3253# sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/NBIAS
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_261_220#
+ a_n433_1745# a_8354_4056# sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2821_220#
+ DM_H[0] sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/Y_H
+ DM_H[1] DM_H_N[0] DM_H_N[1] DM_H[2] DM_H_N[2] a_1415_3203# sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2874_118#
+ OE_N sky130_fd_io__com_opath_datoev2_0/li_5565_99# a_9656_1708# sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/a_158_632#
+ HLD_I_H_N a_1528_3203# a_2205_3177# VGND_IO VPWR sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_1772_220#
+ OUT VCC_IO PU_H_N[3] VGND
Xsky130_fd_io__gpiov2_octl_0 DM_H[1] DM_H[0] DM_H[2] DM_H_N[0] DM_H_N[1] DM_H_N[2]
+ sky130_fd_io__gpiov2_octl_0/PUEN_2OR1_H sky130_fd_io__gpiov2_octl_0/PDEN_H_N[1]
+ sky130_fd_io__gpiov2_octl_0/PDEN_H_N[0] SLOW sky130_fd_io__gpiov2_octl_0/SLOW_H
+ VCC_IO sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/SEL_H_N
+ DM_H[1] VCC_IO DM_H[0] VGND a_7799_1681# VCC_IO VPWR DM_H[2] a_13335_4479# VCC_IO
+ VCC_IO a_13335_4479# SLOW_H_N VGND sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/PUEN_H
+ HLD_I_H_N OD_H sky130_fd_io__gpiov2_octl
Xsky130_fd_io__com_opath_datoev2_0 sky130_fd_io__com_opath_datoev2_0/OE_H DRVLO_H_N
+ VCC_IO HLD_I_OVR_H VGND OUT OE_N sky130_fd_io__com_opath_datoev2_0/sky130_fd_io__com_cclat_0/PD_DIS_H
+ VPWR_KA DRVHI_H sky130_fd_io__com_opath_datoev2_0/li_5565_99# OD_H VGND OD_H sky130_fd_io__com_opath_datoev2
Xsky130_fd_io__gpiov2_obpredrvr_0 SLOW_H_N sky130_fd_io__gpiov2_octl_0/PDEN_H_N[0]
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_261_220#
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/SEL_H_N
+ VCC_IO sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2821_220#
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2874_118#
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/A_H
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/Y_H
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/PUEN_H
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/SEL_H
+ PD_H[0] sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_1772_220#
+ DRVHI_H sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/a_158_632#
+ PU_H_N[2] VCC_IO PU_H_N[3] DRVLO_H_N DRVLO_H_N sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/NBIAS
+ VGND_IO VCC_IO sky130_fd_io__gpiov2_obpredrvr
X0 PD_H[4] DRVLO_H_N a_12137_3347# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=1
X1 VCC_IO a_n461_1863# a_10398_443# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.5
X2 VCC_IO sky130_fd_io__gpiov2_octl_0/PDEN_H_N[1] a_8876_944# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X3 a_8354_4056# PD_H[4] a_8354_3203# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.111 ps=1.37 w=0.42 l=4
X4 a_3125_3203# a_1415_3203# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X5 a_1528_3203# a_2205_3177# a_2205_3177# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.5
X6 a_1415_3203# a_1528_3203# a_1528_3203# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X7 VCC_IO a_1415_3203# a_3125_3203# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X8 VCC_IO DRVLO_H_N a_1159_3105# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.5
X9 VGND_IO a_7610_2597# a_1106_3203# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=1
R0 m1_10510_2769# a_7462_4229# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X10 PU_H_N[0] a_7799_1681# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.6
X11 a_2205_3177# a_2205_3177# a_1528_3203# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X12 a_1528_3203# a_1528_3203# a_1415_3203# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X13 VGND_IO a_7799_1681# a_7743_1707# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X14 VCC_IO a_4416_3253# a_4416_3253# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X15 a_11758_843# sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/Y_H PD_H[3] VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=2
X16 VCC_IO DRVHI_H PU_H_N[1] VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X17 sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/SEL_H sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/SEL_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.6
X18 a_1106_3203# a_1106_3203# a_4416_3253# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X19 a_4416_3253# a_4416_3253# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X20 PD_H[3] sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/Y_H VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
R1 m1_10378_2704# m1_10351_2626# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R2 m1_8330_3159# a_7610_2597# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
X21 VCC_IO a_n461_1863# a_9290_3718# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X22 VGND PD_H[4] sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/A_H VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.111 ps=1.37 w=0.42 l=0.5
X23 a_1415_3203# a_1159_3105# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.5
R3 m1_10312_2627# a_1106_3203# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X24 PD_H[3] sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/Y_H a_11053_559# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.5
X25 a_7161_3177# sky130_fd_io__gpiov2_octl_0/PDEN_H_N[1] VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.335 ps=2.67 w=1 l=0.6
R4 m1_8994_2542# a_7512_2477# sky130_fd_pr__res_generic_m1 w=2.5 l=10m
X26 a_n408_4001# sky130_fd_io__gpiov2_octl_0/SLOW_H a_n112_4027# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
R5 m1_7727_3684# a_7462_4229# sky130_fd_pr__res_generic_m1 w=0.64 l=10m
X27 VCC_IO DRVHI_H PU_H_N[1] VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X28 VCC_IO a_7610_2597# a_8026_3203# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.111 ps=1.37 w=0.42 l=4
X29 a_7462_4229# a_7161_3177# VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.21 ps=1.42 w=1 l=0.6
X30 a_9290_3718# a_1106_3203# a_9882_3718# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
R6 a_7462_4229# m1_10378_2741# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R7 a_8354_3203# m1_8330_3159# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R8 m1_10312_2627# m1_10351_2626# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R9 m1_10523_1531# VCC_IO sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X31 a_10564_1155# a_11085_1123# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X32 a_n408_1837# sky130_fd_io__gpiov2_octl_0/SLOW_H a_n112_1863# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
R10 m1_9138_2849# a_1106_3203# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X33 a_8876_944# sky130_fd_io__gpiov2_octl_0/PDEN_H_N[1] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X34 VCC_IO sky130_fd_io__gpiov2_octl_0/SLOW_H a_n408_1837# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X35 VCC_IO a_n461_4027# a_9935_2938# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.63 pd=3.42 as=0.42 ps=3.28 w=3 l=0.6
X36 a_4416_3253# a_1106_3203# a_1106_3203# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.5
X37 a_1106_3203# a_1106_3203# a_4416_3253# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X38 a_7512_2477# sky130_fd_io__gpiov2_octl_0/PDEN_H_N[1] VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X39 a_11053_559# a_10919_675# a_10398_443# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.5
X40 a_1106_3203# a_1106_3203# a_4416_3253# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
R11 a_11085_1123# m1_10523_1531# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X41 a_4416_3253# a_1106_3203# a_1106_3203# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X42 PD_H[2] DRVLO_H_N a_10194_3718# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.5
X43 a_9656_1708# DRVHI_H PU_H_N[1] VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X44 a_3125_3203# a_1415_3203# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X45 a_12137_3347# DRVLO_H_N PD_H[4] VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=1
X46 a_1159_3105# DRVLO_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.5
X47 VGND a_n408_4001# a_n461_4027# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.185 ps=1.93 w=0.7 l=0.6
X48 PD_H[3] sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/Y_H VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X49 VCC_IO sky130_fd_io__gpiov2_octl_0/SLOW_H a_n408_4001# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X50 VGND_IO a_7610_2597# a_9179_2770# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=1
X51 PD_H[3] sky130_fd_io__gpiov2_octl_0/PDEN_H_N[1] VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
R12 m1_10547_2769# a_10919_675# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X52 VCC_IO a_1415_3203# a_3125_3203# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X53 a_7613_3603# a_7462_4229# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.315 pd=3.21 as=0.795 ps=6.53 w=3 l=0.5
X54 a_3125_3203# a_1415_3203# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.5
X55 sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/SEL_H sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/SEL_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.6
X56 a_10873_1155# sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/Y_H PD_H[3] VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X57 VGND a_n408_1837# a_n461_1863# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.185 ps=1.93 w=0.7 l=0.6
X58 VCC_IO a_1159_3105# a_1106_3203# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.5
X59 PD_H[2] DRVLO_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X60 VCC_IO a_n408_1837# a_n461_1863# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X61 PD_H[3] sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/Y_H a_10564_1155# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.398 ps=3.53 w=1.5 l=0.5
X62 PD_H[4] sky130_fd_io__gpiov2_octl_0/PDEN_H_N[1] VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X63 a_11862_3305# sky130_fd_io__gpiov2_octl_0/PDEN_H_N[1] a_11009_3305# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.111 ps=1.37 w=0.42 l=4
X64 a_8876_944# DRVLO_H_N PD_H[1] VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.5
R13 m1_4181_3684# a_4416_3253# sky130_fd_pr__res_generic_m1 w=0.23 l=10m
X65 a_7755_3603# a_7638_3476# a_7613_3603# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.315 pd=3.21 as=0.315 ps=3.21 w=3 l=0.5
X66 PD_H[2] DRVLO_H_N a_9882_3718# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X67 VCC_IO PD_H[4] sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/A_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.5
X68 sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/SEL_H sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/SEL_H_N VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.185 ps=1.93 w=0.7 l=0.6
X69 a_11009_3305# DRVLO_H_N PD_H[2] VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.111 ps=1.37 w=0.42 l=4
X70 a_9656_1708# sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/PUEN_H VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X71 a_n112_4027# sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/SEL_H_N VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
R14 m1_7764_3684# a_7638_3476# sky130_fd_pr__res_generic_m1 w=0.64 l=10m
X72 VGND_IO sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/Y_H PD_H[3] VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X73 VCC_IO sky130_fd_io__gpiov2_octl_0/SLOW_H a_n408_1837# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X74 a_7610_2597# DRVLO_H_N a_7755_3603# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.315 ps=3.21 w=3 l=0.5
R15 m1_5837_4210# a_1106_3203# sky130_fd_pr__res_generic_m1 w=0.23 l=10m
X75 VGND_IO sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/Y_H PD_H[3] VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X76 a_9179_2770# a_7610_2597# VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=1
X77 VGND_IO DRVLO_H_N PD_H[2] VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X78 VGND_IO a_n461_4027# a_7161_3177# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.42 as=0.14 ps=1.28 w=1 l=0.6
X79 a_n112_1863# sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/SEL_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X80 a_n408_1837# sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/SEL_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X81 VCC_IO a_n408_4001# a_n461_4027# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
R16 m1_9138_2849# a_9179_2770# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X82 VGND_IO sky130_fd_io__gpiov2_octl_0/PDEN_H_N[1] PD_H[2] VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X83 a_4416_3253# a_4416_3253# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X84 a_8354_4056# PD_H[4] VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.111 ps=1.37 w=0.42 l=4
X85 a_1106_3203# a_7610_2597# VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=1
X86 a_4416_3253# a_1106_3203# a_1106_3203# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X87 a_1106_3203# a_1106_3203# a_4416_3253# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.5
X88 a_10194_3718# DRVLO_H_N PD_H[2] VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X89 PU_H_N[1] sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/PUEN_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.5
X90 a_1528_3203# a_2205_3177# a_2205_3177# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X91 a_7638_3476# a_7638_3476# a_7512_2477# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.5
X92 a_1415_3203# a_1528_3203# a_1528_3203# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.5
X93 VGND_IO sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/PUEN_H a_9656_1708# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X94 a_2205_3177# a_2205_3177# a_1528_3203# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X95 a_1106_3203# a_7161_3177# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.5
X96 PU_H_N[0] DRVHI_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.6
X97 VGND_IO sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/Y_H PD_H[3] VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X98 VCC_IO a_4416_3253# a_4416_3253# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X99 VCC_IO a_4416_3253# a_4416_3253# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
R17 m1_10375_2471# a_1106_3203# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R18 m1_4181_3684# a_3125_3203# sky130_fd_pr__res_generic_m1 w=0.23 l=10m
X100 a_4416_3253# a_4416_3253# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X101 a_9290_3718# a_n461_1863# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X102 VCC_IO sky130_fd_io__gpiov2_octl_0/PDEN_H_N[1] a_11009_3747# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.111 ps=1.37 w=0.42 l=4
X103 PU_H_N[1] DRVHI_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
R19 m1_8014_3310# a_8026_3203# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
X104 a_n408_4001# sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/SEL_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X105 VCC_IO a_n408_1837# a_n461_1863# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X106 VCC_IO sky130_fd_io__gpiov2_octl_0/SLOW_H a_n408_4001# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X107 VGND_IO DRVLO_H_N a_7512_2477# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
R20 m1_10375_2471# a_10919_675# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X108 VCC_IO a_1106_3203# a_12137_3347# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.111 ps=1.37 w=0.42 l=1
R21 m1_9297_3844# PD_H[4] sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X109 PD_H[3] sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/Y_H a_10849_843# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=2
X110 VCC_IO VGND_IO a_1415_3203# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.111 ps=1.37 w=0.42 l=8
X111 VGND_IO sky130_fd_io__gpiov2_octl_0/PDEN_H_N[1] PD_H[3] VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
R22 a_1106_3203# m1_8014_3310# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
X112 a_7610_2597# a_7512_2477# VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=10.5 as=1.33 ps=10.5 w=5 l=0.6
X113 a_10398_443# a_n461_1863# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.5
X114 a_4416_3253# a_1106_3203# a_1106_3203# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
R23 m1_9297_3844# a_7638_3476# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X115 a_10398_443# a_11085_1123# a_11053_559# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.5
X116 a_n408_1837# sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/SEL_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X117 VGND_IO DRVLO_H_N a_1159_3105# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
R24 m1_5874_4210# a_4416_3253# sky130_fd_pr__res_generic_m1 w=0.23 l=10m
X118 VCC_IO DRVHI_H PU_H_N[0] VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.6
X119 VGND_IO DRVLO_H_N PD_H[4] VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X120 PD_H[2] a_n461_1863# VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X121 VGND_IO DRVLO_H_N a_7610_2597# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X122 PD_H[1] sky130_fd_io__gpiov2_octl_0/PDEN_H_N[1] VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X123 a_11862_3305# sky130_fd_io__gpiov2_octl_0/PDEN_H_N[1] a_9290_3718# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.111 ps=1.37 w=0.42 l=4
X124 a_4416_3253# a_4416_3253# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.5
X125 VCC_IO a_1415_3203# a_3125_3203# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X126 VCC_IO a_1415_3203# a_3125_3203# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.5
X127 a_9290_3718# a_n461_1863# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.5
X128 a_3125_3203# a_1415_3203# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X129 a_11053_559# sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/Y_H PD_H[3] VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.5
X130 a_9935_2938# sky130_fd_io__gpiov2_octl_0/PDEN_H_N[1] a_7161_3177# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=1 ps=6.67 w=3 l=0.6
X131 VCC_IO a_n408_4001# a_n461_4027# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X132 a_1528_3203# a_1528_3203# a_1415_3203# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
R25 m1_10778_2548# a_11085_1123# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X133 VCC_IO a_10919_675# a_10873_1155# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X134 a_7462_4229# a_7161_3177# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.63 ps=3.42 w=3 l=0.6
X135 a_10398_443# sky130_fd_io__gpiov2_octl_0/PDEN_H_N[1] a_11758_843# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=2
X136 VCC_IO a_4416_3253# a_4416_3253# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X137 a_10194_3718# a_1106_3203# a_9290_3718# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.5
X138 PU_H_N[1] DRVHI_H a_9656_1708# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X139 PD_H[1] DRVLO_H_N a_8876_944# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X140 a_7610_2597# a_7462_4229# VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X141 VGND_IO DRVLO_H_N PD_H[1] VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X142 PD_H[4] DRVLO_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X143 a_7743_1707# DRVHI_H PU_H_N[0] VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
R26 a_7638_3476# m1_8994_2579# sky130_fd_pr__res_generic_m1 w=2.5 l=10m
X144 a_2205_3177# a_7610_2597# VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=10.5 as=1.33 ps=10.5 w=5 l=0.6
X145 a_9882_3718# DRVLO_H_N PD_H[2] VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X146 VCC_IO sky130_fd_io__gpiov2_octl_0/PDEN_H_N[1] a_10849_843# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.111 ps=1.37 w=0.42 l=4
R27 a_10919_675# m1_10778_2585# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X147 PD_H[4] DRVLO_H_N a_11009_3747# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.111 ps=1.37 w=0.42 l=4
X148 a_n408_4001# sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/SEL_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
.ends

.subckt sky130_fd_io__com_res_weak_bentbigres a_419_6804# a_419_8054# a_n256_8772#
+ a_419_8146# a_n258_6046# a_419_9396# a_n2_6046#
R0 a_n256_8772# a_n258_6046# sky130_fd_pr__res_generic_po w=0.8 l=12
R1 a_419_9396# a_419_8146# sky130_fd_pr__res_generic_po w=0.8 l=6
R2 a_n258_6046# a_n2_6046# sky130_fd_pr__res_generic_po w=0.8 l=50
R3 a_419_8054# a_419_6804# sky130_fd_pr__res_generic_po w=0.8 l=6
.ends

.subckt sky130_fd_io__com_res_weak RA RB sky130_fd_io__com_res_weak_bentbigres_0/a_n258_6046#
+ li_n135_8054# a_n160_10423# li_n135_6820# a_n160_9488#
Xsky130_fd_io__com_res_weak_bentbigres_0 li_n135_6820# li_n135_8054# li_n135_6820#
+ li_n135_8054# sky130_fd_io__com_res_weak_bentbigres_0/a_n258_6046# a_n160_9488#
+ RA sky130_fd_io__com_res_weak_bentbigres
R0 a_n160_10423# a_n160_9838# sky130_fd_pr__res_generic_po w=0.8 l=1.5
R1 a_n160_9838# a_n160_9488# sky130_fd_pr__res_generic_po w=0.8 l=1.5
R2 a_n160_10423# m1_n147_10115# sky130_fd_pr__res_generic_m1 w=0.66 l=10m
R3 a_n160_9488# m1_n147_8777# sky130_fd_pr__res_generic_m1 w=0.66 l=10m
R4 a_n160_10423# m1_532_10115# sky130_fd_pr__res_generic_m1 w=0.66 l=10m
R5 a_517_9818# m1_532_9534# sky130_fd_pr__res_generic_m1 w=0.66 l=10m
R6 m1_n147_8777# li_n135_8054# sky130_fd_pr__res_generic_m1 w=0.66 l=10m
R7 m1_n147_10115# a_n160_9838# sky130_fd_pr__res_generic_m1 w=0.66 l=10m
R8 m1_532_10115# a_517_9818# sky130_fd_pr__res_generic_m1 w=0.66 l=10m
R9 a_517_9818# RB sky130_fd_pr__res_generic_po w=0.8 l=1.5
R10 m1_532_9534# RB sky130_fd_pr__res_generic_m1 w=0.66 l=10m
R11 a_n160_9838# m1_n147_9555# sky130_fd_pr__res_generic_m1 w=0.66 l=10m
R12 li_n135_8054# m1_n146_7735# sky130_fd_pr__res_generic_m1 w=0.66 l=10m
R13 a_n160_10423# a_517_9818# sky130_fd_pr__res_generic_po w=0.8 l=1.5
R14 m1_n147_9555# a_n160_9488# sky130_fd_pr__res_generic_m1 w=0.66 l=10m
R15 m1_n146_7434# li_n135_6820# sky130_fd_pr__res_generic_m1 w=0.66 l=10m
.ends

.subckt sky130_fd_io__pfet_con_diff_wo_abt_270v2 w_415_600# a_2303_1380# a_13777_1380#
+ a_8817_1380# a_4287_1380# a_7263_1380# a_12223_1380# a_9247_1380# a_2865_1380# a_5841_1380#
+ a_4849_1380# a_10801_1380# a_14135_1380# a_1311_1380# a_12785_1380# a_7825_1380#
+ a_3295_1380# a_9809_1380# a_1001_1552# a_6271_1380# a_5279_1380# a_11231_1380# a_10239_1380#
+ a_8255_1380# a_1873_1380# a_13215_1380# a_3857_1380# a_11793_1380# a_881_1380# a_6833_1380#
X0 a_1001_1552# a_13777_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.97 pd=6.19 as=3.78 ps=11.5 w=5 l=0.6
X1 a_1001_1552# a_4849_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X2 a_1001_1552# a_8817_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X3 w_415_600# a_10239_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X4 a_1001_1552# a_1873_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X5 w_415_600# a_3295_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X6 w_415_600# a_14135_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=4.3 pd=11.7 as=2.97 ps=6.19 w=5 l=0.6
X7 a_1001_1552# a_5841_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X8 w_415_600# a_2303_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X9 w_415_600# a_7263_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X10 a_1001_1552# a_4849_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X11 w_415_600# a_11231_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X12 a_1001_1552# a_12785_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X13 w_415_600# a_10239_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X14 a_1001_1552# a_8817_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X15 w_415_600# a_3295_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X16 w_415_600# a_2303_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X17 w_415_600# a_7263_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X18 a_1001_1552# a_12785_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X19 a_1001_1552# a_3857_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X20 a_1001_1552# a_7825_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X21 w_415_600# a_13215_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X22 w_415_600# a_1311_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X23 w_415_600# a_6271_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X24 a_1001_1552# a_3857_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X25 w_415_600# a_5279_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X26 a_1001_1552# a_11793_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X27 a_1001_1552# a_7825_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X28 w_415_600# a_9247_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X29 a_1001_1552# a_10801_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X30 w_415_600# a_13215_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X31 w_415_600# a_1311_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X32 w_415_600# a_6271_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X33 a_1001_1552# a_881_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=4.32 ps=11.7 w=5 l=0.6
X34 a_1001_1552# a_2865_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X35 w_415_600# a_5279_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X36 a_1001_1552# a_11793_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X37 a_1001_1552# a_10801_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X38 a_1001_1552# a_6833_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X39 w_415_600# a_9247_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X40 w_415_600# a_12223_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X41 a_1001_1552# a_881_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=4.32 ps=11.7 w=5 l=0.6
X42 a_1001_1552# a_9809_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X43 a_1001_1552# a_2865_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X44 w_415_600# a_4287_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X45 a_1001_1552# a_6833_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X46 w_415_600# a_8255_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X47 w_415_600# a_12223_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X48 a_1001_1552# a_13777_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.97 pd=6.19 as=3.78 ps=11.5 w=5 l=0.6
X49 a_1001_1552# a_9809_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X50 a_1001_1552# a_1873_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X51 w_415_600# a_4287_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X52 w_415_600# a_14135_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=4.3 pd=11.7 as=2.97 ps=6.19 w=5 l=0.6
X53 w_415_600# a_8255_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X54 a_1001_1552# a_5841_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X55 w_415_600# a_11231_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
.ends

.subckt sky130_fd_io__gpio_pudrvr_strongv2 PU_H_N[3] PU_H_N[2] VCC_IO m1_1330_n459#
+ TIE_HI_ESD m1_6027_281# m1_3418_50# VNB a_14575_n157# m1_6652_281# m1_3028_333#
+ PAD m1_14880_n614# li_9083_n155#
Xsky130_fd_io__pfet_con_diff_wo_abt_270v2_0 VCC_IO PU_H_N[2] m1_14229_1478# m1_8837_1478#
+ PU_H_N[3] PU_H_N[3] m1_11745_1478# m1_8837_1478# PU_H_N[2] PU_H_N[3] PU_H_N[3] m1_10391_1478#
+ m1_14229_1478# PU_H_N[2] PU_H_N[2] PU_H_N[3] PU_H_N[2] m1_10391_1478# PAD PU_H_N[3]
+ PU_H_N[3] m1_11745_1478# m1_10391_1478# m1_8837_1478# PU_H_N[2] m1_13667_1478# PU_H_N[3]
+ m1_11745_1478# PU_H_N[2] PU_H_N[3] sky130_fd_io__pfet_con_diff_wo_abt_270v2
R0 m1_14229_1478# m2_14532_958# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R1 m1_13667_1478# m2_13593_958# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R2 m2_12849_n185# PU_H_N[2] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R3 m1_8837_1478# m2_10673_n208# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R4 m1_10391_1478# m2_10945_92# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R5 m2_11422_n209# PU_H_N[2] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R6 m1_13667_1478# m2_14075_958# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R7 m2_10673_n208# PU_H_N[2] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R8 m2_10197_n209# TIE_HI_ESD sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R9 m1_11745_1478# m2_12608_116# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R10 m2_10945_n209# TIE_HI_ESD sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R11 m1_10391_1478# m2_11422_92# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R12 m1_11745_1478# m2_12849_116# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R13 m2_12608_n185# PU_H_N[3] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R14 m2_14769_657# PU_H_N[2] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R15 m2_11186_n208# PU_H_N[3] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R16 m2_13837_658# PU_H_N[3] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R17 TIE_HI_ESD a_14575_n157# sky130_fd_pr__res_generic_po w=0.5 l=10.2
R18 m2_14286_658# TIE_HI_ESD sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R19 m1_8837_1478# m2_10197_92# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R20 m1_8837_1478# m2_10439_92# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R21 m2_14532_657# PU_H_N[3] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R22 m1_10391_1478# m2_11186_n208# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R23 m2_13593_657# TIE_HI_ESD sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R24 m1_13667_1478# m2_13837_658# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R25 m1_14229_1478# m2_14769_958# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R26 m1_11745_1478# m2_12365_n184# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R27 m2_10439_n209# PU_H_N[3] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R28 m2_12365_n184# TIE_HI_ESD sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R29 m1_14229_1478# m2_14286_658# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R30 m2_14075_657# PU_H_N[2] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
.ends

.subckt sky130_fd_io__nfet_con_diff_wo_abt_270v2 VCC_IO VSSIO PAD a_10282_1285# a_5322_1285#
+ a_12266_1285# a_7306_1285# a_3900_1285# a_2908_1285# a_5884_1285# a_14178_1285#
+ a_10844_1285# a_1354_1285# a_7868_1285# a_12828_1285# a_8860_1285# a_13820_1285#
+ a_4330_1285# a_3338_1285# a_11274_1285# a_6314_1285# a_8298_1285# a_13258_1285#
+ a_9290_1285# a_1916_1285# a_4892_1285# a_6876_1285# a_924_1285# a_11836_1285# a_2346_1285#
+ a_9852_1285#
X0 VSSIO a_5322_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X1 PAD a_9852_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X2 VSSIO a_11274_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X3 PAD a_10844_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X4 PAD a_6876_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X5 VSSIO a_2346_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X6 PAD a_1916_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X7 VSSIO a_12266_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X8 VSSIO a_6314_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X9 PAD a_11836_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X10 VSSIO a_9290_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X11 PAD a_4892_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X12 VSSIO a_10282_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X13 VSSIO a_4330_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X14 PAD a_3900_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X15 PAD a_8860_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X16 VSSIO a_3338_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X17 VSSIO a_8298_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X18 PAD a_924_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.42 ps=11.4 w=5 l=0.6
X19 VSSIO a_7306_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X20 PAD a_13820_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=2.97 pd=6.19 as=3.78 ps=11.5 w=5 l=0.6
X21 PAD a_2908_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X22 PAD a_7868_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X23 VSSIO a_13258_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X24 PAD a_12828_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X25 VSSIO a_14178_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.42 pd=11.4 as=2.97 ps=6.19 w=5 l=0.6
X26 VSSIO a_1354_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X27 PAD a_5884_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X28 VSSIO a_11274_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X29 VSSIO a_5322_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X30 PAD a_9852_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X31 PAD a_10844_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X32 VSSIO a_2346_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X33 PAD a_6876_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X34 VSSIO a_6314_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X35 PAD a_1916_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X36 VSSIO a_12266_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X37 PAD a_11836_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X38 PAD a_4892_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X39 VSSIO a_4330_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X40 VSSIO a_9290_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X41 PAD a_8860_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X42 VSSIO a_10282_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X43 PAD a_924_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.42 ps=11.4 w=5 l=0.6
X44 PAD a_3900_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X45 VSSIO a_3338_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X46 VSSIO a_8298_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X47 PAD a_2908_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X48 PAD a_7868_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X49 VSSIO a_13258_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X50 VSSIO a_7306_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X51 PAD a_13820_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=2.97 pd=6.19 as=3.78 ps=11.5 w=5 l=0.6
X52 PAD a_12828_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X53 VSSIO a_1354_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X54 VSSIO a_14178_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.42 pd=11.4 as=2.97 ps=6.19 w=5 l=0.6
X55 PAD a_5884_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
.ends

.subckt sky130_fd_io__gpiov2_pddrvr_strong sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_3338_1285#
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_4330_1285# sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_10282_1285#
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_6314_1285# sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_12266_1285#
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_8298_1285# sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_9290_1285#
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_1916_1285# sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/VSSIO
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_4892_1285# sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/VCC_IO
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_10844_1285# sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/PAD
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_6876_1285# sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_14178_1285#
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_2346_1285# sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_12828_1285#
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_13820_1285# sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_924_1285#
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_9852_1285# sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_5322_1285#
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_11274_1285# sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_7306_1285#
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_13258_1285# sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_3900_1285#
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_2908_1285# sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_5884_1285#
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_1354_1285# sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_7868_1285#
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_11836_1285# sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_8860_1285#
Xsky130_fd_io__nfet_con_diff_wo_abt_270v2_0 sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/VCC_IO
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/VSSIO sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/PAD
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_10282_1285# sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_5322_1285#
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_12266_1285# sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_7306_1285#
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_3900_1285# sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_2908_1285#
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_5884_1285# sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_14178_1285#
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_10844_1285# sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_1354_1285#
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_7868_1285# sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_12828_1285#
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_8860_1285# sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_13820_1285#
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_4330_1285# sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_3338_1285#
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_11274_1285# sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_6314_1285#
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_8298_1285# sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_13258_1285#
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_9290_1285# sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_1916_1285#
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_4892_1285# sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_6876_1285#
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_924_1285# sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_11836_1285#
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_2346_1285# sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_9852_1285#
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2
.ends

.subckt sky130_fd_io__com_pudrvr_weakv2 PU_H_N PAD w_258_n30# a_756_297#
X0 PAD PU_H_N w_258_n30# w_258_n30# sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X1 PAD PU_H_N w_258_n30# w_258_n30# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X2 w_258_n30# PU_H_N a_756_297# w_258_n30# sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X3 w_258_n30# PU_H_N a_756_297# w_258_n30# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X4 w_258_n30# PU_H_N PAD w_258_n30# sky130_fd_pr__pfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.5
X5 w_258_n30# PU_H_N PAD w_258_n30# sky130_fd_pr__pfet_g5v0d10v5 ad=1.86 pd=14.5 as=0.98 ps=7.28 w=7 l=0.5
X6 a_756_297# PU_H_N w_258_n30# w_258_n30# sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.5
X7 a_756_297# PU_H_N w_258_n30# w_258_n30# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.86 ps=14.5 w=7 l=0.5
.ends

.subckt sky130_fd_io__res250_sub_small a_10_2# a_2142_2#
R0 a_10_2# a_2142_2# sky130_fd_pr__res_generic_po w=2 l=10.1
.ends

.subckt sky130_fd_io__res250only_small PAD ROUT
Xsky130_fd_io__res250_sub_small_0 PAD ROUT sky130_fd_io__res250_sub_small
.ends

.subckt sky130_fd_io__gpio_pddrvr_weakv2 PD_H PAD dw_n122_84# w_168_168#
X0 w_168_168# PD_H PAD w_168_168# sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=10.5 as=1.33 ps=10.5 w=5 l=0.6
X1 w_168_168# PD_H PAD w_168_168# sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=10.5 as=1.33 ps=10.5 w=5 l=0.6
X2 w_168_168# PD_H PAD w_168_168# sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=10.5 as=1.33 ps=10.5 w=5 l=0.6
X3 w_168_168# PD_H PAD w_168_168# sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=10.5 as=1.33 ps=10.5 w=5 l=0.6
X4 w_168_168# PD_H PAD w_168_168# sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=10.5 as=1.33 ps=10.5 w=5 l=0.6
X5 w_168_168# PD_H PAD w_168_168# sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=10.5 as=1.33 ps=10.5 w=5 l=0.6
.ends

.subckt sky130_fd_io__gpio_odrvr_subv2 VGND PD_H[0] PD_H[2] PD_H[1] PD_H[3] TIE_LO_ESD
+ FORCE_HI_H_N FORCE_LO_H FORCE_LOVOL_H PU_H_N[0] PU_H_N[1] PU_H_N[2] PU_H_N[3] VSSIO_AMX
+ VGND_IO TIE_HI_ESD w_588_14893# m3_6107_13425# w_n915_9930# li_5884_n9263# m2_8191_n10933#
+ sky130_fd_io__gpiov2_pddrvr_strong_0/sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/VSSIO
+ sky130_fd_io__gpio_pudrvr_strongv2_0/m1_14880_n614# sky130_fd_io__gpio_pudrvr_strongv2_0/li_9083_n155#
+ m1_2782_13727# PAD w_5497_14893# VCC_IO
Xsky130_fd_io__com_res_weak_0 sky130_fd_io__com_res_weak_0/RA sky130_fd_io__com_res_weak_0/RB
+ sky130_fd_io__com_res_weak_0/sky130_fd_io__com_res_weak_bentbigres_0/a_n258_6046#
+ sky130_fd_io__com_res_weak_0/li_n135_8054# sky130_fd_io__com_res_weak_0/a_n160_10423#
+ sky130_fd_io__com_res_weak_0/li_n135_6820# sky130_fd_io__com_res_weak_0/a_n160_9488#
+ sky130_fd_io__com_res_weak
Xsky130_fd_io__gpio_pudrvr_strongv2_0 PU_H_N[3] PU_H_N[2] VCC_IO VCC_IO TIE_HI_ESD
+ VCC_IO PU_H_N[0] VGND VCC_IO VCC_IO VCC_IO PAD sky130_fd_io__gpio_pudrvr_strongv2_0/m1_14880_n614#
+ sky130_fd_io__gpio_pudrvr_strongv2_0/li_9083_n155# sky130_fd_io__gpio_pudrvr_strongv2
Xsky130_fd_io__gpiov2_pddrvr_strong_0 m1_11278_13727# m1_9854_13727# PD_H[3] m1_8317_13727#
+ m1_2782_13727# PD_H[2] PD_H[3] m1_12832_13727# sky130_fd_io__gpiov2_pddrvr_strong_0/sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/VSSIO
+ m1_9854_13727# VCC_IO PD_H[3] PAD m1_8317_13727# m1_870_13727# m1_12832_13727# m1_2220_13727#
+ m1_870_13727# m1_12832_13727# PD_H[3] m1_9854_13727# PD_H[3] m1_7742_13727# m1_870_13727#
+ m1_11278_13727# m1_11278_13727# m1_8317_13727# m1_12832_13727# PD_H[2] PD_H[3] PD_H[2]
+ sky130_fd_io__gpiov2_pddrvr_strong
Xsky130_fd_io__com_pudrvr_weakv2_0 PU_H_N[0] sky130_fd_io__com_res_weak_0/RA VCC_IO
+ sky130_fd_io__com_res_weak_0/RA sky130_fd_io__com_pudrvr_weakv2
Xsky130_fd_io__res250only_small_0 PAD sky130_fd_io__com_res_weak_0/RB sky130_fd_io__res250only_small
Xsky130_fd_io__gpio_pddrvr_weakv2_0 PD_H[0] sky130_fd_io__com_res_weak_0/RA VCC_IO
+ w_5497_14893# sky130_fd_io__gpio_pddrvr_weakv2
R0 a_10314_7886# sky130_fd_io__com_res_weak_0/RB sky130_fd_pr__res_generic_po w=2 l=2
R1 TIE_LO_ESD m2_1933_16117# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R2 m2_982_15816# m1_870_13727# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R3 PD_H[2] m2_10071_16117# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R4 m2_12848_15816# m1_12832_13727# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R5 a_9612_7886# a_10314_7886# sky130_fd_pr__res_generic_po w=2 l=3
X0 VCC_IO PU_H_N[1] a_782_15260# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=1.86 pd=14.5 as=0.98 ps=7.28 w=7 l=0.5
R6 TIE_LO_ESD m2_9451_16117# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R7 PD_H[3] m2_7318_15817# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R8 m2_13278_15816# m1_12832_13727# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
X1 a_782_15260# PD_H[1] w_588_14893# w_588_14893# sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=10.5 as=1.33 ps=10.5 w=5 l=0.6
X2 a_782_15260# PU_H_N[1] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.86 ps=14.5 w=7 l=0.5
R9 TIE_LO_ESD m2_499_16117# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R10 PD_H[2] m2_6889_16117# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R11 m2_11414_15816# m1_11278_13727# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R12 TIE_LO_ESD m2_10931_16117# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
X3 a_782_15260# PD_H[1] w_588_14893# w_588_14893# sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=10.5 as=1.33 ps=10.5 w=5 l=0.6
X4 a_782_15260# PD_H[1] w_588_14893# w_588_14893# sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=10.5 as=1.33 ps=10.5 w=5 l=0.6
R13 m2_1933_15816# m1_2220_13727# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R14 m2_10071_15816# m1_9854_13727# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R15 m2_9451_15816# m1_8317_13727# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R16 PD_H[3] m2_1650_16117# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R17 m2_7318_15817# m1_7742_13727# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R18 PD_H[2] m2_1345_15817# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R19 m2_499_15816# m1_870_13727# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R20 m2_6889_15816# m1_7742_13727# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
X5 a_782_15260# PU_H_N[1] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.86 ps=14.5 w=7 l=0.5
R21 m2_10931_15816# m1_9854_13727# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R22 m1_9882_7996# a_10314_7886# sky130_fd_pr__res_generic_m1 w=1.32 l=10m
R23 PD_H[3] m2_9020_15817# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R24 TIE_LO_ESD m2_13707_15817# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R25 m2_1650_15816# m1_2220_13727# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R26 PD_H[2] m2_8591_16117# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R27 PD_H[3] m2_740_15817# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R28 m1_9882_7996# a_9612_7886# sky130_fd_pr__res_generic_m1 w=1.32 l=10m
R29 m2_1345_15817# m1_2220_13727# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
X6 a_782_15260# PU_H_N[1] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
R30 PD_H[3] m2_10500_15817# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R31 PD_H[3] m2_11843_15817# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R32 m2_13707_15817# m1_12832_13727# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
X7 VCC_IO PU_H_N[1] a_782_15260# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
R33 m2_9020_15817# m1_8317_13727# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R34 m2_8591_15816# m1_8317_13727# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R35 TIE_LO_ESD m2_12274_16117# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R36 m2_740_15817# m1_870_13727# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R37 TIE_LO_ESD m2_7749_16117# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R38 m2_10500_15817# m1_9854_13727# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R39 m2_11843_15817# m1_11278_13727# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
X8 a_782_15260# PD_H[1] w_588_14893# w_588_14893# sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=10.5 as=1.33 ps=10.5 w=5 l=0.6
X9 VCC_IO PU_H_N[1] a_782_15260# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=1.86 pd=14.5 as=0.98 ps=7.28 w=7 l=0.5
X10 a_782_15260# PU_H_N[1] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
R40 PD_H[2] m2_982_16117# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R41 PD_H[2] m2_12848_16117# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R42 m2_12274_15816# m1_11278_13727# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
X11 VCC_IO PU_H_N[1] a_782_15260# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
R43 a_782_15260# a_9612_7886# sky130_fd_pr__res_generic_po w=2 l=5
R44 PD_H[3] m2_13278_16117# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R45 TIE_LO_ESD VGND_IO sky130_fd_pr__res_generic_po w=0.5 l=10.2
R46 m2_7749_15816# m1_7742_13727# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R47 PD_H[2] m2_11414_16117# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
.ends

.subckt sky130_fd_io__gpio_odrvrv2 PAD PD_H[0] PD_H[1] PD_H[2] PD_H[3] PU_H_N[0] PU_H_N[1]
+ PU_H_N[2] PU_H_N[3] TIE_HI_ESD FORCE_HI_H_N FORCE_LO_H VSSIO_AMX w_n915_9930# FORCE_LOVOL_H
+ sky130_fd_io__gpio_odrvr_subv2_0/m3_6107_13425# TIE_LO_ESD w_5497_14893# sky130_fd_io__gpio_odrvr_subv2_0/li_5884_n9263#
+ sky130_fd_io__gpio_odrvr_subv2_0/m2_8191_n10933# w_588_14893# sky130_fd_io__gpio_odrvr_subv2_0/sky130_fd_io__gpio_pudrvr_strongv2_0/li_9083_n155#
+ sky130_fd_io__gpio_odrvr_subv2_0/sky130_fd_io__gpio_pudrvr_strongv2_0/m1_14880_n614#
+ sky130_fd_io__gpio_odrvr_subv2_0/m1_2782_13727# VGND VCC_IO VGND_IO
Xsky130_fd_io__gpio_odrvr_subv2_0 VGND PD_H[0] PD_H[2] PD_H[1] PD_H[3] TIE_LO_ESD
+ FORCE_HI_H_N FORCE_LO_H FORCE_LOVOL_H PU_H_N[0] PU_H_N[1] PU_H_N[2] PU_H_N[3] VSSIO_AMX
+ VGND_IO TIE_HI_ESD w_588_14893# sky130_fd_io__gpio_odrvr_subv2_0/m3_6107_13425#
+ w_n915_9930# sky130_fd_io__gpio_odrvr_subv2_0/li_5884_n9263# sky130_fd_io__gpio_odrvr_subv2_0/m2_8191_n10933#
+ VGND_IO sky130_fd_io__gpio_odrvr_subv2_0/sky130_fd_io__gpio_pudrvr_strongv2_0/m1_14880_n614#
+ sky130_fd_io__gpio_odrvr_subv2_0/sky130_fd_io__gpio_pudrvr_strongv2_0/li_9083_n155#
+ sky130_fd_io__gpio_odrvr_subv2_0/m1_2782_13727# PAD w_5497_14893# VCC_IO sky130_fd_io__gpio_odrvr_subv2
.ends

.subckt sky130_fd_io__gpio_opathv2 HLD_I_OVR_H HLD_I_H_N OD_H SLOW VPWR TIE_HI_ESD
+ sky130_fd_io__gpiov2_octl_dat_0/a_1528_3203# sky130_fd_io__gpiov2_octl_dat_0/a_2205_3177#
+ sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/a_158_632#
+ sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/Y_H
+ DM_H[0] DM_H_N[0] sky130_fd_io__gpiov2_octl_dat_0/a_1106_3203# DM_H[2] DM_H_N[1]
+ m1_4747_14860# sky130_fd_io__gpio_odrvrv2_0/sky130_fd_io__gpio_odrvr_subv2_0/sky130_fd_io__gpio_pudrvr_strongv2_0/li_9083_n155#
+ TIE_LO_ESD sky130_fd_io__gpiov2_octl_dat_0/a_3125_3203# sky130_fd_io__gpiov2_octl_dat_0/a_4416_3253#
+ sky130_fd_io__gpio_odrvrv2_0/PU_H_N[2] m2_2157_n626# sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2821_220#
+ m1_5007_14796# DM_H[1] PAD sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2874_118#
+ sky130_fd_io__gpiov2_octl_dat_0/a_8354_4056# w_5597_30124# DM_H_N[2] sky130_fd_io__gpiov2_octl_dat_0/a_1415_3203#
+ VSSIO_AMX sky130_fd_io__gpio_odrvrv2_0/sky130_fd_io__gpio_odrvr_subv2_0/m3_6107_13425#
+ sky130_fd_io__gpiov2_octl_dat_0/a_9656_1708# VGND_IO OE_N OUT w_688_30124# VPWR_KA
+ VCC_IO sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/NBIAS
+ VGND sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_1772_220#
+ sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_261_220#
Xsky130_fd_io__gpiov2_octl_dat_0 VPWR_KA SLOW HLD_I_OVR_H OD_H sky130_fd_io__gpiov2_octl_dat_0/SLOW_H_N
+ sky130_fd_io__gpiov2_octl_dat_0/DRVHI_H sky130_fd_io__gpio_odrvrv2_0/PU_H_N[2] sky130_fd_io__gpio_odrvrv2_0/PU_H_N[1]
+ sky130_fd_io__gpio_odrvrv2_0/PU_H_N[0] sky130_fd_io__gpio_odrvrv2_0/PD_H[1] sky130_fd_io__gpio_odrvrv2_0/PD_H[0]
+ sky130_fd_io__gpiov2_octl_dat_0/PD_H[4] sky130_fd_io__gpio_odrvrv2_0/PD_H[3] sky130_fd_io__gpio_odrvrv2_0/PD_H[2]
+ sky130_fd_io__gpiov2_octl_dat_0/a_1106_3203# sky130_fd_io__gpiov2_octl_dat_0/a_3125_3203#
+ sky130_fd_io__gpiov2_octl_dat_0/a_4416_3253# sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/NBIAS
+ sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_261_220#
+ VGND sky130_fd_io__gpiov2_octl_dat_0/a_8354_4056# sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2821_220#
+ DM_H[0] sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/Y_H
+ DM_H[1] DM_H_N[0] DM_H_N[1] DM_H[2] DM_H_N[2] sky130_fd_io__gpiov2_octl_dat_0/a_1415_3203#
+ sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2874_118#
+ OE_N VGND sky130_fd_io__gpiov2_octl_dat_0/a_9656_1708# sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/a_158_632#
+ HLD_I_H_N sky130_fd_io__gpiov2_octl_dat_0/a_1528_3203# sky130_fd_io__gpiov2_octl_dat_0/a_2205_3177#
+ VGND_IO VPWR sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_1772_220#
+ OUT VCC_IO sky130_fd_io__gpio_odrvrv2_0/PU_H_N[3] VGND sky130_fd_io__gpiov2_octl_dat
Xsky130_fd_io__gpio_odrvrv2_0 PAD sky130_fd_io__gpio_odrvrv2_0/PD_H[0] sky130_fd_io__gpio_odrvrv2_0/PD_H[1]
+ sky130_fd_io__gpio_odrvrv2_0/PD_H[2] sky130_fd_io__gpio_odrvrv2_0/PD_H[3] sky130_fd_io__gpio_odrvrv2_0/PU_H_N[0]
+ sky130_fd_io__gpio_odrvrv2_0/PU_H_N[1] sky130_fd_io__gpio_odrvrv2_0/PU_H_N[2] sky130_fd_io__gpio_odrvrv2_0/PU_H_N[3]
+ TIE_HI_ESD VSSIO_AMX VSSIO_AMX VSSIO_AMX w_n815_25161# VSSIO_AMX sky130_fd_io__gpio_odrvrv2_0/sky130_fd_io__gpio_odrvr_subv2_0/m3_6107_13425#
+ TIE_LO_ESD w_5597_30124# VGND VGND w_688_30124# sky130_fd_io__gpio_odrvrv2_0/sky130_fd_io__gpio_odrvr_subv2_0/sky130_fd_io__gpio_pudrvr_strongv2_0/li_9083_n155#
+ sky130_fd_io__gpio_odrvrv2_0/PU_H_N[1] sky130_fd_io__gpiov2_octl_dat_0/PD_H[4] VGND
+ VCC_IO VGND_IO sky130_fd_io__gpio_odrvrv2
.ends

.subckt sky130_fd_io__amux_switch_1v2b AMUXBUS_HV PG_AMX_VDDA_H_N NG_AMX_VPMP_H NG_PAD_VPMP_H
+ PAD_HV_P0 PAD_HV_P1 PG_PAD_VDDIOQ_H_N PAD_HV_N0 PAD_HV_N1 VDDA VSSD PAD_HV_N2 VDDIO
+ PAD_HV_N3 w_7010_315# w_3919_213#
X0 PAD_HV_N0 NG_PAD_VPMP_H w_3919_213# w_3919_213# sky130_fd_pr__nfet_g5v0d10v5 ad=1.23 pd=7.35 as=0.98 ps=7.28 w=7 l=0.5
X1 AMUXBUS_HV NG_AMX_VPMP_H w_3919_213# w_3919_213# sky130_fd_pr__nfet_g5v0d10v5 ad=1.23 pd=7.35 as=0.98 ps=7.28 w=7 l=0.5
X2 PAD_HV_N1 NG_PAD_VPMP_H w_3919_213# w_3919_213# sky130_fd_pr__nfet_g5v0d10v5 ad=1.23 pd=7.35 as=0.98 ps=7.28 w=7 l=0.5
X3 w_3919_213# PG_PAD_VDDIOQ_H_N PAD_HV_P0 VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.23 ps=7.35 w=7 l=0.5
X4 w_7010_315# NG_PAD_VPMP_H PAD_HV_N2 w_7010_315# sky130_fd_pr__nfet_g5v0d10v5 ad=1.23 pd=7.35 as=0.98 ps=7.28 w=7 l=0.5
X5 AMUXBUS_HV PG_AMX_VDDA_H_N w_3919_213# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.23 ps=7.35 w=7 l=0.5
X6 w_3919_213# PG_AMX_VDDA_H_N AMUXBUS_HV VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1.23 pd=7.35 as=0.98 ps=7.28 w=7 l=0.5
X7 w_3919_213# NG_PAD_VPMP_H PAD_HV_N1 w_3919_213# sky130_fd_pr__nfet_g5v0d10v5 ad=1.96 pd=14.6 as=1.23 ps=7.35 w=7 l=0.5
X8 PAD_HV_N2 NG_PAD_VPMP_H w_7010_315# w_7010_315# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.23 ps=7.35 w=7 l=0.5
X9 w_3919_213# NG_AMX_VPMP_H AMUXBUS_HV w_3919_213# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.23 ps=7.35 w=7 l=0.5
X10 w_3919_213# PG_AMX_VDDA_H_N AMUXBUS_HV VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1.23 pd=7.35 as=1.96 ps=14.6 w=7 l=0.5
X11 w_3919_213# NG_PAD_VPMP_H PAD_HV_N0 w_3919_213# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=2.2 ps=14.6 w=7 l=0.5
X12 w_7010_315# NG_AMX_VPMP_H AMUXBUS_HV w_7010_315# sky130_fd_pr__nfet_g5v0d10v5 ad=1.23 pd=7.35 as=0.98 ps=7.28 w=7 l=0.5
X13 w_7010_315# NG_PAD_VPMP_H PAD_HV_N3 w_7010_315# sky130_fd_pr__nfet_g5v0d10v5 ad=1.23 pd=7.35 as=0.98 ps=7.28 w=7 l=0.5
X14 w_3919_213# NG_PAD_VPMP_H PAD_HV_N1 w_3919_213# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.23 ps=7.35 w=7 l=0.5
X15 AMUXBUS_HV NG_AMX_VPMP_H w_3919_213# w_3919_213# sky130_fd_pr__nfet_g5v0d10v5 ad=1.23 pd=7.35 as=0.98 ps=7.28 w=7 l=0.5
X16 AMUXBUS_HV NG_AMX_VPMP_H w_3919_213# w_3919_213# sky130_fd_pr__nfet_g5v0d10v5 ad=2.2 pd=14.6 as=0.98 ps=7.28 w=7 l=0.5
X17 w_3919_213# PG_PAD_VDDIOQ_H_N PAD_HV_P0 VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=2.2 ps=14.6 w=7 l=0.5
X18 w_7010_315# NG_AMX_VPMP_H AMUXBUS_HV w_7010_315# sky130_fd_pr__nfet_g5v0d10v5 ad=1.23 pd=7.35 as=0.98 ps=7.28 w=7 l=0.5
X19 AMUXBUS_HV PG_AMX_VDDA_H_N w_3919_213# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.23 ps=7.35 w=7 l=0.5
X20 PAD_HV_N3 NG_PAD_VPMP_H w_7010_315# w_7010_315# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.23 ps=7.35 w=7 l=0.5
X21 AMUXBUS_HV NG_AMX_VPMP_H w_3919_213# w_3919_213# sky130_fd_pr__nfet_g5v0d10v5 ad=1.23 pd=7.35 as=1.96 ps=14.6 w=7 l=0.5
X22 PAD_HV_P1 PG_PAD_VDDIOQ_H_N w_3919_213# VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=2.2 pd=14.6 as=0.98 ps=7.28 w=7 l=0.5
X23 PAD_HV_P1 PG_PAD_VDDIOQ_H_N w_3919_213# VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=1.23 pd=7.35 as=0.98 ps=7.28 w=7 l=0.5
X24 PAD_HV_N2 NG_PAD_VPMP_H w_7010_315# w_7010_315# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=2.2 ps=14.6 w=7 l=0.5
X25 AMUXBUS_HV NG_AMX_VPMP_H w_7010_315# w_7010_315# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.23 ps=7.35 w=7 l=0.5
X26 PAD_HV_N3 NG_PAD_VPMP_H w_7010_315# w_7010_315# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.23 ps=7.35 w=7 l=0.5
X27 w_3919_213# NG_AMX_VPMP_H AMUXBUS_HV w_3919_213# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.23 ps=7.35 w=7 l=0.5
X28 PAD_HV_N1 NG_PAD_VPMP_H w_3919_213# w_3919_213# sky130_fd_pr__nfet_g5v0d10v5 ad=1.23 pd=7.35 as=0.98 ps=7.28 w=7 l=0.5
X29 w_7010_315# NG_PAD_VPMP_H PAD_HV_N2 w_7010_315# sky130_fd_pr__nfet_g5v0d10v5 ad=1.23 pd=7.35 as=0.98 ps=7.28 w=7 l=0.5
X30 w_7010_315# NG_AMX_VPMP_H AMUXBUS_HV w_7010_315# sky130_fd_pr__nfet_g5v0d10v5 ad=2.2 pd=14.6 as=0.98 ps=7.28 w=7 l=0.5
X31 w_7010_315# NG_AMX_VPMP_H AMUXBUS_HV w_7010_315# sky130_fd_pr__nfet_g5v0d10v5 ad=1.23 pd=7.35 as=1.96 ps=14.6 w=7 l=0.5
X32 w_3919_213# PG_PAD_VDDIOQ_H_N PAD_HV_P1 VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.23 ps=7.35 w=7 l=0.5
X33 w_3919_213# PG_AMX_VDDA_H_N AMUXBUS_HV VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=2.2 pd=14.6 as=0.98 ps=7.28 w=7 l=0.5
X34 PAD_HV_P0 PG_PAD_VDDIOQ_H_N w_3919_213# VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=1.23 pd=7.35 as=0.98 ps=7.28 w=7 l=0.5
X35 w_3919_213# NG_AMX_VPMP_H AMUXBUS_HV w_3919_213# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.23 ps=7.35 w=7 l=0.5
X36 w_3919_213# NG_PAD_VPMP_H PAD_HV_N0 w_3919_213# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.23 ps=7.35 w=7 l=0.5
X37 AMUXBUS_HV NG_AMX_VPMP_H w_7010_315# w_7010_315# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.23 ps=7.35 w=7 l=0.5
X38 AMUXBUS_HV NG_AMX_VPMP_H w_7010_315# w_7010_315# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.23 ps=7.35 w=7 l=0.5
X39 w_7010_315# NG_PAD_VPMP_H PAD_HV_N3 w_7010_315# sky130_fd_pr__nfet_g5v0d10v5 ad=2.2 pd=14.6 as=0.98 ps=7.28 w=7 l=0.5
.ends

.subckt sky130_fd_io__res75only_small PAD ROUT
R0 PAD ROUT sky130_fd_pr__res_generic_po w=2 l=3.15
.ends

.subckt sky130_fd_io__inv_1 VNB VPB VPWR VGND Y A
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.83 as=0.386 ps=2.93 w=1.12 l=0.15
X1 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.211 pd=2.05 as=0.263 ps=2.19 w=0.74 l=0.15
.ends

.subckt sky130_fd_io__nor2_1 VNB VPB VPWR VGND B Y A
X0 a_116_368# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.151 pd=1.39 as=0.33 ps=2.83 w=1.12 l=0.15
X1 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=1.02 as=0.211 ps=2.05 w=0.74 l=0.15
X2 Y B a_116_368# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.83 as=0.151 ps=1.39 w=1.12 l=0.15
X3 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.211 pd=2.05 as=0.104 ps=1.02 w=0.74 l=0.15
.ends

.subckt sky130_fd_io__nand2_1 VNB VPB VPWR VGND B Y A
X0 a_117_74# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0888 pd=0.98 as=0.211 ps=2.05 w=0.74 l=0.15
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.319 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X2 Y A a_117_74# VNB sky130_fd_pr__nfet_01v8 ad=0.211 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.168 pd=1.42 as=0.319 ps=2.81 w=1.12 l=0.15
.ends

.subckt sky130_fd_io__gpiov2_amux_decoder sky130_fd_io__inv_1_8/A sky130_fd_io__inv_1_0/Y
+ sky130_fd_io__inv_1_11/A sky130_fd_io__inv_1_2/Y sky130_fd_io__inv_1_13/A sky130_fd_io__nor2_1_0/Y
+ sky130_fd_io__inv_1_4/Y sky130_fd_io__nand2_1_0/Y sky130_fd_io__inv_1_1/A sky130_fd_io__nor2_1_2/Y
+ sky130_fd_io__nand2_1_2/Y sky130_fd_io__inv_1_6/Y sky130_fd_io__inv_1_3/A sky130_fd_io__nor2_1_1/B
+ sky130_fd_io__inv_1_8/Y sky130_fd_io__nand2_1_1/B sky130_fd_io__nor2_1_1/A sky130_fd_io__inv_1_11/Y
+ sky130_fd_io__inv_1_5/A sky130_fd_io__nand2_1_1/A sky130_fd_io__nor2_1_3/B sky130_fd_io__nor2_1_3/A
+ sky130_fd_io__tap_1_2/VGND sky130_fd_io__inv_1_13/Y sky130_fd_io__nand2_1_3/B sky130_fd_io__inv_1_7/A
+ sky130_fd_io__inv_1_10/A sky130_fd_io__nand2_1_3/A sky130_fd_io__inv_1_1/Y sky130_fd_io__inv_1_12/A
+ sky130_fd_io__inv_1_9/A sky130_fd_io__inv_1_8/VGND sky130_fd_io__inv_1_3/Y sky130_fd_io__inv_1_14/A
+ sky130_fd_io__inv_1_0/A sky130_fd_io__nor2_1_1/Y sky130_fd_io__nand2_1_1/Y sky130_fd_io__inv_1_5/Y
+ sky130_fd_io__nor2_1_0/B sky130_fd_io__nor2_1_3/Y sky130_fd_io__inv_1_2/A sky130_fd_io__nor2_1_0/A
+ sky130_fd_io__inv_1_7/Y sky130_fd_io__nand2_1_3/Y sky130_fd_io__inv_1_10/Y sky130_fd_io__nand2_1_0/B
+ sky130_fd_io__tap_1_2/VPB sky130_fd_io__inv_1_4/A sky130_fd_io__nand2_1_0/A sky130_fd_io__nor2_1_2/B
+ sky130_fd_io__inv_1_9/Y sky130_fd_io__nor2_1_2/A sky130_fd_io__inv_1_12/Y sky130_fd_io__inv_1_6/A
+ sky130_fd_io__nand2_1_2/B sky130_fd_io__nand2_1_2/A sky130_fd_io__tap_1_2/VPWR sky130_fd_io__tap_1_1/VGND
+ VSUBS sky130_fd_io__inv_1_14/Y
Xsky130_fd_io__inv_1_10 VSUBS sky130_fd_io__tap_1_2/VPB sky130_fd_io__tap_1_2/VPWR
+ sky130_fd_io__tap_1_2/VGND sky130_fd_io__inv_1_10/Y sky130_fd_io__inv_1_10/A sky130_fd_io__inv_1
Xsky130_fd_io__inv_1_11 VSUBS sky130_fd_io__tap_1_2/VPB sky130_fd_io__tap_1_2/VPWR
+ sky130_fd_io__tap_1_2/VGND sky130_fd_io__inv_1_11/Y sky130_fd_io__inv_1_11/A sky130_fd_io__inv_1
Xsky130_fd_io__inv_1_12 VSUBS sky130_fd_io__tap_1_2/VPB sky130_fd_io__tap_1_2/VPWR
+ sky130_fd_io__inv_1_8/VGND sky130_fd_io__inv_1_12/Y sky130_fd_io__inv_1_12/A sky130_fd_io__inv_1
Xsky130_fd_io__inv_1_13 VSUBS sky130_fd_io__tap_1_2/VPB sky130_fd_io__tap_1_2/VPWR
+ sky130_fd_io__inv_1_8/VGND sky130_fd_io__inv_1_13/Y sky130_fd_io__inv_1_13/A sky130_fd_io__inv_1
Xsky130_fd_io__inv_1_14 VSUBS sky130_fd_io__tap_1_2/VPB sky130_fd_io__tap_1_2/VPWR
+ sky130_fd_io__tap_1_1/VGND sky130_fd_io__inv_1_14/Y sky130_fd_io__inv_1_14/A sky130_fd_io__inv_1
Xsky130_fd_io__inv_1_0 VSUBS sky130_fd_io__tap_1_2/VPB sky130_fd_io__tap_1_2/VPWR
+ sky130_fd_io__tap_1_1/VGND sky130_fd_io__inv_1_0/Y sky130_fd_io__inv_1_0/A sky130_fd_io__inv_1
Xsky130_fd_io__inv_1_1 VSUBS sky130_fd_io__tap_1_2/VPB sky130_fd_io__tap_1_2/VPWR
+ sky130_fd_io__tap_1_1/VGND sky130_fd_io__inv_1_1/Y sky130_fd_io__inv_1_1/A sky130_fd_io__inv_1
Xsky130_fd_io__inv_1_2 VSUBS sky130_fd_io__tap_1_2/VPB sky130_fd_io__tap_1_2/VPWR
+ sky130_fd_io__tap_1_1/VGND sky130_fd_io__inv_1_2/Y sky130_fd_io__inv_1_2/A sky130_fd_io__inv_1
Xsky130_fd_io__inv_1_3 VSUBS sky130_fd_io__tap_1_2/VPB sky130_fd_io__tap_1_2/VPWR
+ sky130_fd_io__tap_1_1/VGND sky130_fd_io__inv_1_3/Y sky130_fd_io__inv_1_3/A sky130_fd_io__inv_1
Xsky130_fd_io__inv_1_4 VSUBS sky130_fd_io__tap_1_2/VPB sky130_fd_io__tap_1_2/VPWR
+ sky130_fd_io__tap_1_1/VGND sky130_fd_io__inv_1_4/Y sky130_fd_io__inv_1_4/A sky130_fd_io__inv_1
Xsky130_fd_io__inv_1_5 VSUBS sky130_fd_io__tap_1_2/VPB sky130_fd_io__tap_1_2/VPWR
+ sky130_fd_io__tap_1_2/VGND sky130_fd_io__inv_1_5/Y sky130_fd_io__inv_1_5/A sky130_fd_io__inv_1
Xsky130_fd_io__inv_1_6 VSUBS sky130_fd_io__tap_1_2/VPB sky130_fd_io__tap_1_2/VPWR
+ sky130_fd_io__tap_1_1/VGND sky130_fd_io__inv_1_6/Y sky130_fd_io__inv_1_6/A sky130_fd_io__inv_1
Xsky130_fd_io__nor2_1_0 VSUBS sky130_fd_io__tap_1_2/VPB sky130_fd_io__tap_1_2/VPWR
+ sky130_fd_io__tap_1_1/VGND sky130_fd_io__nor2_1_0/B sky130_fd_io__nor2_1_0/Y sky130_fd_io__nor2_1_0/A
+ sky130_fd_io__nor2_1
Xsky130_fd_io__inv_1_7 VSUBS sky130_fd_io__tap_1_2/VPB sky130_fd_io__tap_1_2/VPWR
+ sky130_fd_io__tap_1_2/VGND sky130_fd_io__inv_1_7/Y sky130_fd_io__inv_1_7/A sky130_fd_io__inv_1
Xsky130_fd_io__nor2_1_2 VSUBS sky130_fd_io__tap_1_2/VPB sky130_fd_io__tap_1_2/VPWR
+ sky130_fd_io__tap_1_1/VGND sky130_fd_io__nor2_1_2/B sky130_fd_io__nor2_1_2/Y sky130_fd_io__nor2_1_2/A
+ sky130_fd_io__nor2_1
Xsky130_fd_io__nor2_1_1 VSUBS sky130_fd_io__tap_1_2/VPB sky130_fd_io__tap_1_2/VPWR
+ sky130_fd_io__tap_1_1/VGND sky130_fd_io__nor2_1_1/B sky130_fd_io__nor2_1_1/Y sky130_fd_io__nor2_1_1/A
+ sky130_fd_io__nor2_1
Xsky130_fd_io__nor2_1_3 VSUBS sky130_fd_io__tap_1_2/VPB sky130_fd_io__tap_1_2/VPWR
+ sky130_fd_io__tap_1_1/VGND sky130_fd_io__nor2_1_3/B sky130_fd_io__nor2_1_3/Y sky130_fd_io__nor2_1_3/A
+ sky130_fd_io__nor2_1
Xsky130_fd_io__inv_1_8 VSUBS sky130_fd_io__tap_1_2/VPB sky130_fd_io__tap_1_2/VPWR
+ sky130_fd_io__inv_1_8/VGND sky130_fd_io__inv_1_8/Y sky130_fd_io__inv_1_8/A sky130_fd_io__inv_1
Xsky130_fd_io__inv_1_9 VSUBS sky130_fd_io__tap_1_2/VPB sky130_fd_io__tap_1_2/VPWR
+ sky130_fd_io__tap_1_2/VGND sky130_fd_io__inv_1_9/Y sky130_fd_io__inv_1_9/A sky130_fd_io__inv_1
Xsky130_fd_io__nand2_1_0 VSUBS sky130_fd_io__tap_1_2/VPB sky130_fd_io__tap_1_2/VPWR
+ sky130_fd_io__tap_1_2/VGND sky130_fd_io__nand2_1_0/B sky130_fd_io__nand2_1_0/Y sky130_fd_io__nand2_1_0/A
+ sky130_fd_io__nand2_1
Xsky130_fd_io__nand2_1_1 VSUBS sky130_fd_io__tap_1_2/VPB sky130_fd_io__tap_1_2/VPWR
+ sky130_fd_io__inv_1_8/VGND sky130_fd_io__nand2_1_1/B sky130_fd_io__nand2_1_1/Y sky130_fd_io__nand2_1_1/A
+ sky130_fd_io__nand2_1
Xsky130_fd_io__nand2_1_2 VSUBS sky130_fd_io__tap_1_2/VPB sky130_fd_io__tap_1_2/VPWR
+ sky130_fd_io__tap_1_2/VGND sky130_fd_io__nand2_1_2/B sky130_fd_io__nand2_1_2/Y sky130_fd_io__nand2_1_2/A
+ sky130_fd_io__nand2_1
Xsky130_fd_io__nand2_1_3 VSUBS sky130_fd_io__tap_1_2/VPB sky130_fd_io__tap_1_2/VPWR
+ sky130_fd_io__tap_1_2/VGND sky130_fd_io__nand2_1_3/B sky130_fd_io__nand2_1_3/Y sky130_fd_io__nand2_1_3/A
+ sky130_fd_io__nand2_1
.ends

.subckt sky130_fd_io__gpiov2_amux_ctl_logic sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_4/A
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_9/Y sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_2/Y
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_6/A sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_1/Y
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_1/B sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_0/Y
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_8/A sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_1/A
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_3/Y sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_11/Y
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_0/B sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_3/B
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_0/A sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_2/Y
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_3/A sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_13/Y
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_2/B sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_10/A
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_4/Y sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_2/A
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_1/A sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_12/A
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_6/Y sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_3/A
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_14/A sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_8/Y
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_1/Y sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_5/A
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_0/Y sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_0/B
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_3/Y sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__tap_1_0/VPWR
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_8/VGND sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_10/Y
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_7/A sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_0/A
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_2/Y sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_1/Y
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_2/B sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_9/A
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_2/A sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_12/Y
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_1/B sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_1/A
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_3/Y sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_14/Y
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_0/A sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__tap_1_2/VPB
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_11/A sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_3/B
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_5/Y sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__tap_1_0/VPB
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__tap_1_2/VPWR sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__tap_1_0/VGND
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_3/A sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_2/A
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__tap_1_1/VGND VSUBS sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_13/A
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_7/Y sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_0/Y
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__tap_1_2/VGND
Xsky130_fd_io__gpiov2_amux_decoder_0 sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_8/A
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_0/Y sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_11/A
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_2/Y sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_13/A
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_0/Y sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_4/Y
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_0/Y sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_1/A
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_2/Y sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_2/Y
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_6/Y sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_3/A
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_1/B sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_8/Y
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_1/B sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_1/A
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_11/Y sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_5/A
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_1/A sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_3/B
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_3/A sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__tap_1_2/VGND
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_13/Y sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_3/B
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_7/A sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_10/A
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_3/A sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_1/Y
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_12/A sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_9/A
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_8/VGND sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_3/Y
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_14/A sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_0/A
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_1/Y sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_1/Y
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_5/Y sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_0/B
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_3/Y sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_2/A
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_0/A sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_7/Y
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_3/Y sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_10/Y
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_0/B sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__tap_1_2/VPB
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_4/A sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_0/A
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_2/B sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_9/Y
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_2/A sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_12/Y
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_6/A sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_2/B
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_2/A sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__tap_1_2/VPWR
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__tap_1_1/VGND VSUBS sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_14/Y
+ sky130_fd_io__gpiov2_amux_decoder
.ends

.subckt sky130_fd_io__gpiov2_amux sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_0/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_9/Y
+ sky130_fd_io__amux_switch_1v2b_0/PAD_HV_P0 sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_3/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_13/Y
+ sky130_fd_io__res75only_small_0/ROUT sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_6/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_10/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_2/Y
+ sky130_fd_io__amux_switch_1v2b_1/PAD_HV_N3 sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_0/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_8/A
+ sky130_fd_io__amux_switch_1v2b_1/PAD_HV_N2 sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_12/A
+ sky130_fd_io__amux_switch_1v2b_1/PG_AMX_VDDA_H_N sky130_fd_io__amux_switch_1v2b_1/PAD_HV_N1
+ sky130_fd_io__res75only_small_7/ROUT sky130_fd_io__amux_switch_1v2b_0/NG_PAD_VPMP_H
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_2/Y
+ sky130_fd_io__amux_switch_1v2b_1/PAD_HV_N0 sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_1/B
+ sky130_fd_io__amux_switch_1v2b_0/NG_AMX_VPMP_H sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_1/A
+ sky130_fd_io__amux_switch_1v2b_1/PAD_HV_P1 sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_14/A
+ sky130_fd_io__amux_switch_1v2b_1/PAD_HV_P0 sky130_fd_io__res75only_small_13/PAD
+ sky130_fd_io__res75only_small_4/ROUT sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_1/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_3/B
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_4/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_3/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_1/A
+ w_11765_4495# sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_3/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_0/B
+ sky130_fd_io__amux_switch_1v2b_0/PG_AMX_VDDA_H_N sky130_fd_io__res75only_small_2/PAD
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_6/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_0/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_10/Y
+ sky130_fd_io__amux_switch_1v2b_1/PG_PAD_VDDIOQ_H_N sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_3/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_2/B
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_8/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_2/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_12/Y
+ w_11765_6609# sky130_fd_io__amux_switch_1v2b_1/VDDA sky130_fd_io__res75only_small_8/ROUT
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_5/A
+ sky130_fd_io__res75only_small_9/PAD sky130_fd_io__amux_switch_1v2b_1/NG_PAD_VPMP_H
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_1/Y
+ sky130_fd_io__res75only_small_13/ROUT sky130_fd_io__res75only_small_5/ROUT sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_14/Y
+ sky130_fd_io__amux_switch_1v2b_1/NG_AMX_VPMP_H sky130_fd_io__res75only_small_1/PAD
+ sky130_fd_io__res75only_small_8/PAD sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_7/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_11/A
+ sky130_fd_io__res75only_small_10/ROUT sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_3/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_0/B
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_1/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_9/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_0/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_13/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_0/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__tap_1_0/VPWR
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__tap_1_2/VGND
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_2/B
+ sky130_fd_io__res75only_small_0/PAD sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_3/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_2/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_0/A
+ sky130_fd_io__amux_switch_1v2b_0/PG_PAD_VDDIOQ_H_N sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__tap_1_1/VGND
+ sky130_fd_io__res75only_small_9/ROUT w_8674_6609# sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_2/Y
+ sky130_fd_io__amux_switch_1v2b_0/AMUXBUS_HV sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_5/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__tap_1_0/VPB
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_2/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__tap_1_2/VPWR
+ sky130_fd_io__amux_switch_1v2b_0/PAD_HV_N3 sky130_fd_io__res75only_small_6/ROUT
+ sky130_fd_io__res75only_small_7/PAD sky130_fd_io__amux_switch_1v2b_1/AMUXBUS_HV
+ sky130_fd_io__amux_switch_1v2b_0/PAD_HV_N2 sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_1/B
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_7/Y
+ sky130_fd_io__amux_switch_1v2b_0/PAD_HV_N1 sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_1/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_11/Y
+ w_8674_4393# sky130_fd_io__res75only_small_3/ROUT sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__tap_1_2/VPB
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__tap_1_0/VGND
+ sky130_fd_io__amux_switch_1v2b_0/PAD_HV_N0 sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_4/A
+ sky130_fd_io__amux_switch_1v2b_0/VDDIO sky130_fd_io__res75only_small_5/PAD sky130_fd_io__amux_switch_1v2b_0/PAD_HV_P1
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_3/B
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_8/VGND
+ VSUBS sky130_fd_io__amux_switch_1v2b_1/VDDIO
Xsky130_fd_io__amux_switch_1v2b_0 sky130_fd_io__amux_switch_1v2b_0/AMUXBUS_HV sky130_fd_io__amux_switch_1v2b_0/PG_AMX_VDDA_H_N
+ sky130_fd_io__amux_switch_1v2b_0/NG_AMX_VPMP_H sky130_fd_io__amux_switch_1v2b_0/NG_PAD_VPMP_H
+ sky130_fd_io__amux_switch_1v2b_0/PAD_HV_P0 sky130_fd_io__amux_switch_1v2b_0/PAD_HV_P1
+ sky130_fd_io__amux_switch_1v2b_0/PG_PAD_VDDIOQ_H_N sky130_fd_io__amux_switch_1v2b_0/PAD_HV_N0
+ sky130_fd_io__amux_switch_1v2b_0/PAD_HV_N1 sky130_fd_io__amux_switch_1v2b_1/VDDA
+ VSUBS sky130_fd_io__amux_switch_1v2b_0/PAD_HV_N2 sky130_fd_io__amux_switch_1v2b_0/VDDIO
+ sky130_fd_io__amux_switch_1v2b_0/PAD_HV_N3 w_11765_6609# w_8674_6609# sky130_fd_io__amux_switch_1v2b
Xsky130_fd_io__amux_switch_1v2b_1 sky130_fd_io__amux_switch_1v2b_1/AMUXBUS_HV sky130_fd_io__amux_switch_1v2b_1/PG_AMX_VDDA_H_N
+ sky130_fd_io__amux_switch_1v2b_1/NG_AMX_VPMP_H sky130_fd_io__amux_switch_1v2b_1/NG_PAD_VPMP_H
+ sky130_fd_io__amux_switch_1v2b_1/PAD_HV_P0 sky130_fd_io__amux_switch_1v2b_1/PAD_HV_P1
+ sky130_fd_io__amux_switch_1v2b_1/PG_PAD_VDDIOQ_H_N sky130_fd_io__amux_switch_1v2b_1/PAD_HV_N0
+ sky130_fd_io__amux_switch_1v2b_1/PAD_HV_N1 sky130_fd_io__amux_switch_1v2b_1/VDDA
+ VSUBS sky130_fd_io__amux_switch_1v2b_1/PAD_HV_N2 sky130_fd_io__amux_switch_1v2b_1/VDDIO
+ sky130_fd_io__amux_switch_1v2b_1/PAD_HV_N3 w_11765_4495# w_8674_4393# sky130_fd_io__amux_switch_1v2b
Xsky130_fd_io__res75only_small_10 sky130_fd_io__res75only_small_10/PAD sky130_fd_io__res75only_small_10/ROUT
+ sky130_fd_io__res75only_small
Xsky130_fd_io__res75only_small_11 sky130_fd_io__res75only_small_2/PAD sky130_fd_io__res75only_small_10/PAD
+ sky130_fd_io__res75only_small
Xsky130_fd_io__res75only_small_13 sky130_fd_io__res75only_small_13/PAD sky130_fd_io__res75only_small_13/ROUT
+ sky130_fd_io__res75only_small
Xsky130_fd_io__res75only_small_12 sky130_fd_io__res75only_small_1/PAD sky130_fd_io__res75only_small_13/PAD
+ sky130_fd_io__res75only_small
Xsky130_fd_io__res75only_small_0 sky130_fd_io__res75only_small_0/PAD sky130_fd_io__res75only_small_0/ROUT
+ sky130_fd_io__res75only_small
Xsky130_fd_io__res75only_small_1 sky130_fd_io__res75only_small_1/PAD sky130_fd_io__res75only_small_3/PAD
+ sky130_fd_io__res75only_small
Xsky130_fd_io__res75only_small_2 sky130_fd_io__res75only_small_2/PAD sky130_fd_io__res75only_small_0/PAD
+ sky130_fd_io__res75only_small
Xsky130_fd_io__res75only_small_3 sky130_fd_io__res75only_small_3/PAD sky130_fd_io__res75only_small_3/ROUT
+ sky130_fd_io__res75only_small
Xsky130_fd_io__res75only_small_4 sky130_fd_io__res75only_small_5/PAD sky130_fd_io__res75only_small_4/ROUT
+ sky130_fd_io__res75only_small
Xsky130_fd_io__gpiov2_amux_ctl_logic_0 sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_4/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_9/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_2/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_6/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_1/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_1/B
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_0/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_8/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_1/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_3/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_11/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_0/B
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_3/B
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_0/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_2/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_3/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_13/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_2/B
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_10/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_4/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_2/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_1/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_12/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_6/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_3/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_14/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_8/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_1/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_5/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_0/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_0/B
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_3/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__tap_1_0/VPWR
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_8/VGND
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_10/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_7/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_0/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_2/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_1/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_2/B
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_9/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_2/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_12/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_1/B
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_1/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_3/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_14/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_0/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__tap_1_2/VPB
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_11/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_3/B
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_5/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__tap_1_0/VPB
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__tap_1_2/VPWR
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__tap_1_0/VGND
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_3/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_2/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__tap_1_1/VGND
+ VSUBS sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_13/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_7/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_0/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__tap_1_2/VGND
+ sky130_fd_io__gpiov2_amux_ctl_logic
Xsky130_fd_io__res75only_small_5 sky130_fd_io__res75only_small_5/PAD sky130_fd_io__res75only_small_5/ROUT
+ sky130_fd_io__res75only_small
Xsky130_fd_io__res75only_small_6 sky130_fd_io__res75only_small_8/PAD sky130_fd_io__res75only_small_6/ROUT
+ sky130_fd_io__res75only_small
Xsky130_fd_io__res75only_small_7 sky130_fd_io__res75only_small_7/PAD sky130_fd_io__res75only_small_7/ROUT
+ sky130_fd_io__res75only_small
Xsky130_fd_io__res75only_small_8 sky130_fd_io__res75only_small_8/PAD sky130_fd_io__res75only_small_8/ROUT
+ sky130_fd_io__res75only_small
Xsky130_fd_io__res75only_small_9 sky130_fd_io__res75only_small_9/PAD sky130_fd_io__res75only_small_9/ROUT
+ sky130_fd_io__res75only_small
.ends

.subckt sky130_fd_io__gpiov2_ipath_hvls OUT OUT_B MODE_NORMAL_N IN_VCCHIB INB_VCCHIB
+ IN_VDDIO MODE_VCCHIB_N MODE_NORMAL MODE_VCCHIB VDDIO_Q VSSD
X0 a_1290_2876# MODE_VCCHIB_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.5
X1 VSSD OUT_B OUT VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.5
X2 a_1752_1955# a_1175_2172# OUT_B VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X3 a_602_2876# IN_VCCHIB a_1930_201# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.5
X4 VDDIO_Q OUT_B OUT VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.5
X5 a_1930_201# MODE_VCCHIB VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X6 VDDIO_Q OUT_B OUT VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.5
X7 a_621_2778# MODE_VCCHIB_N VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.5
X8 a_2024_2876# MODE_NORMAL_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X9 OUT OUT_B VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X10 VDDIO_Q MODE_VCCHIB_N a_1290_2876# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X11 a_1930_201# IN_VCCHIB a_602_2876# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X12 a_621_2778# INB_VCCHIB a_881_201# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X13 a_881_201# MODE_VCCHIB VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X14 OUT OUT_B VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X15 VSSD MODE_VCCHIB a_1752_1955# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X16 VSSD MODE_VCCHIB a_1930_201# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X17 VSSD MODE_VCCHIB a_1930_201# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.5
X18 a_621_2778# a_602_2876# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X19 VSSD OUT_B OUT VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.5
X20 a_1290_2876# a_1175_2172# OUT_B VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X21 VDDIO_Q MODE_NORMAL_N a_2024_2876# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.5
X22 a_1752_2267# MODE_NORMAL VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X23 a_881_201# MODE_VCCHIB VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.5
X24 a_881_201# INB_VCCHIB a_621_2778# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X25 a_1175_2172# a_602_2876# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.398 ps=3.53 w=1.5 l=0.5
X26 VDDIO_Q MODE_NORMAL a_2911_2876# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.5
X27 VDDIO_Q OUT_B OUT VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X28 VSSD MODE_VCCHIB a_881_201# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X29 VDDIO_Q a_621_2778# a_602_2876# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.398 ps=3.53 w=1.5 l=0.5
X30 a_2024_2876# IN_VDDIO OUT_B VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.5
X31 OUT_B a_1175_2172# a_1290_2876# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.5
X32 OUT_B IN_VDDIO a_1752_2267# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.5
X33 VSSD MODE_VCCHIB a_881_201# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X34 a_881_201# INB_VCCHIB a_621_2778# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X35 a_602_2876# IN_VCCHIB a_1930_201# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X36 a_2911_2876# MODE_VCCHIB OUT_B VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.5
X37 OUT OUT_B VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X38 a_1930_201# MODE_VCCHIB VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X39 OUT_B IN_VDDIO a_2024_2876# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X40 a_1175_2172# a_602_2876# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.398 ps=3.53 w=1.5 l=0.5
.ends

.subckt sky130_fd_io__gpiov2_vcchib_in_buf IN_H MODE_VCCHIB_LV_N VCCHIB VSSD OUT OUT_N
X0 VCCHIB MODE_VCCHIB_LV_N a_612_2476# VCCHIB sky130_fd_pr__pfet_01v8 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.25
X1 VSSD VSSD VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=4.58 ps=36.7 w=1 l=0.8
X2 a_612_2476# MODE_VCCHIB_LV_N VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.25
X3 VCCHIB MODE_VCCHIB_LV_N a_612_2476# VCCHIB sky130_fd_pr__pfet_01v8 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.25
X4 OUT OUT_N VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.25
X5 a_538_595# a_591_563# a_751_595# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.8
X6 a_446_3055# MODE_VCCHIB_LV_N VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.25
X7 VCCHIB a_446_3055# OUT_N VCCHIB sky130_fd_pr__pfet_01v8 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.25
X8 VSSD a_446_3055# OUT_N VSSD sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.25
X9 VSSD OUT_N OUT VSSD sky130_fd_pr__nfet_01v8 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.25
X10 a_751_595# IN_H VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.8
X11 a_751_595# a_591_563# a_538_595# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.8
X12 VCCHIB MODE_VCCHIB_LV_N a_612_3332# VCCHIB sky130_fd_pr__pfet_01v8 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.25
X13 VSSD MODE_VCCHIB_LV_N a_446_3055# VSSD sky130_fd_pr__nfet_01v8 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.25
X14 a_446_3055# a_591_563# a_612_3332# VCCHIB sky130_fd_pr__pfet_01v8 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.25
X15 a_612_3332# a_591_563# a_446_3055# VCCHIB sky130_fd_pr__pfet_01v8 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.25
X16 a_446_3055# a_591_563# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.25
X17 a_751_595# a_591_563# a_538_595# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.8
X18 VSSD OUT_N OUT VSSD sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.25
X19 VSSD IN_H a_751_595# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X20 a_751_595# IN_H a_591_563# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X21 a_591_563# IN_H a_612_2476# VCCHIB sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.8
X22 a_591_563# IN_H a_751_595# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.8
X23 a_538_595# MODE_VCCHIB_LV_N VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.25
X24 VSSD VSSD VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=10.5 as=0 ps=0 w=5 l=0.8
X25 a_612_2476# IN_H a_591_563# VCCHIB sky130_fd_pr__pfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.8
X26 VSSD a_591_563# a_446_3055# VSSD sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.25
X27 OUT OUT_N VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.25
.ends

.subckt sky130_fd_io__gpiov2_in_buf OUT OUT_N MODE_NORMAL_N IN_H IN_VT VTRIP_SEL_H
+ VTRIP_SEL_H_N VDDIO_Q VSSD m1_n467_n748#
X0 a_1761_1865# a_973_1767# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X1 a_249_n802# IN_H VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X2 a_2073_1865# a_36_n802# a_249_n802# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.8
X3 VSSD a_36_n802# a_2651_1865# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.5
X4 VDDIO_Q VDDIO_Q VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=1.33 pd=10.5 as=11.5 ps=89.5 w=5 l=0.8
X5 a_249_n802# IN_H VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X6 VDDIO_Q MODE_NORMAL_N a_219_1865# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.5
X7 a_249_n802# IN_H a_36_n802# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X8 a_219_1865# MODE_NORMAL_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.5
X9 a_3531_2403# MODE_NORMAL_N a_3358_2403# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X10 a_36_n802# IN_H a_249_n802# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X11 VSSD VSSD VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=10.5 as=15.1 ps=118 w=5 l=0.8
X12 a_3358_2403# MODE_NORMAL_N VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.196 ps=1.96 w=0.7 l=0.6
X13 a_2385_1865# MODE_NORMAL_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.5
X14 a_36_n802# IN_H a_219_1865# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.8
X15 VDDIO_Q MODE_NORMAL_N a_2073_1865# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X16 VDDIO_Q VTRIP_SEL_H a_3531_2403# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X17 a_249_n802# a_36_n802# a_2073_1865# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.8
X18 VSSD VTRIP_SEL_H a_3358_2403# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X19 a_917_1865# a_973_1767# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.5
X20 VSSD IN_H a_249_n802# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X21 VDDIO_Q a_2651_1865# OUT_N VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.5
X22 OUT OUT_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.5
X23 VSSD IN_H a_249_n802# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X24 a_973_1767# a_3358_2403# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X25 a_2651_1865# a_36_n802# a_2385_1865# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.5
X26 VDDIO_Q a_973_1767# a_1761_1865# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X27 a_2073_1865# MODE_NORMAL_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X28 a_973_1767# a_3358_2403# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X29 a_249_n802# IN_H a_36_n802# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X30 a_2651_1865# MODE_NORMAL_N VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X31 a_249_n802# IN_H a_36_n802# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.8
X32 a_36_n802# IN_H a_249_n802# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X33 a_1761_1865# a_36_n802# a_249_n802# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X34 a_249_n802# a_36_n802# a_1761_1865# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.8
X35 a_2073_1865# a_36_n802# a_249_n802# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.8
X36 a_249_n802# a_36_n802# a_2073_1865# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.8
X37 a_249_n802# IN_H VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X38 a_3531_2403# MODE_NORMAL_N a_3358_2403# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X39 VSSD IN_VT a_249_n802# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X40 VSSD IN_H a_249_n802# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=10.5 as=1.33 ps=10.5 w=5 l=0.8
X41 VSSD VTRIP_SEL_H_N IN_VT VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=1
X42 VDDIO_Q VTRIP_SEL_H a_3531_2403# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X43 VSSD VSSD VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=10.5 as=0 ps=0 w=5 l=0.8
X44 VDDIO_Q a_973_1767# a_917_1865# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X45 a_249_n802# a_36_n802# a_1761_1865# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X46 a_917_1865# IN_H a_36_n802# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X47 a_973_1767# a_3358_2403# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X48 a_1761_1865# a_36_n802# a_249_n802# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X49 VSSD MODE_NORMAL_N a_2651_1865# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X50 a_2651_1865# a_36_n802# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X51 VSSD a_2651_1865# OUT_N VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.5
X52 OUT OUT_N VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.5
.ends

.subckt sky130_fd_io__gpiov2_ipath_lvls IN_VCCHIB IN_VDDIO MODE_NORMAL_LV MODE_NORMAL_LV_N
+ MODE_VCCHIB_LV MODE_VCCHIB_LV_N VCCHIB VSSD OUT OUT_B a_323_2354#
X0 VSSD OUT_B OUT VSSD sky130_fd_pr__nfet_01v8 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.25
X1 VCCHIB MODE_NORMAL_LV_N a_436_2754# VCCHIB sky130_fd_pr__pfet_01v8 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.25
X2 VCCHIB MODE_VCCHIB_LV_N a_1504_2754# VCCHIB sky130_fd_pr__pfet_01v8 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.25
X3 a_823_n317# MODE_NORMAL_LV VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.25
X4 a_1679_n317# IN_VCCHIB OUT_B VSSD sky130_fd_pr__nfet_01v8 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.25
X5 OUT OUT_B VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.25
X6 a_114_2354# IN_VDDIO VCCHIB VCCHIB sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.5
X7 a_1504_2754# IN_VCCHIB OUT_B VCCHIB sky130_fd_pr__pfet_01v8 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.25
X8 a_323_2354# a_114_2354# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.25
X9 a_436_2754# MODE_NORMAL_LV_N VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.25
X10 OUT_B a_323_2354# a_436_2754# VCCHIB sky130_fd_pr__pfet_01v8 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.25
X11 VCCHIB OUT_B OUT VCCHIB sky130_fd_pr__pfet_01v8 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.25
X12 VCCHIB MODE_NORMAL_LV a_114_2354# VCCHIB sky130_fd_pr__pfet_01v8 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.25
X13 VCCHIB OUT_B OUT VCCHIB sky130_fd_pr__pfet_01v8 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.25
X14 a_823_n317# a_323_2354# OUT_B VSSD sky130_fd_pr__nfet_01v8 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.25
X15 a_1679_n317# MODE_VCCHIB_LV VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.25
X16 a_2141_2754# MODE_NORMAL_LV OUT_B VCCHIB sky130_fd_pr__pfet_01v8 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.25
X17 a_1504_2754# MODE_VCCHIB_LV_N VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.25
X18 VSSD MODE_NORMAL_LV a_823_n317# VSSD sky130_fd_pr__nfet_01v8 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.25
X19 VSSD MODE_VCCHIB_LV a_1679_n317# VSSD sky130_fd_pr__nfet_01v8 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.25
X20 a_316_n17# IN_VDDIO a_114_2354# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.398 ps=3.53 w=1.5 l=0.5
X21 VCCHIB MODE_VCCHIB_LV a_2141_2754# VCCHIB sky130_fd_pr__pfet_01v8 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.25
X22 VCCHIB IN_VDDIO a_114_2354# VCCHIB sky130_fd_pr__pfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.5
X23 OUT_B IN_VCCHIB a_1504_2754# VCCHIB sky130_fd_pr__pfet_01v8 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.25
X24 VSSD MODE_NORMAL_LV a_316_n17# VSSD sky130_fd_pr__nfet_01v8 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.25
X25 OUT OUT_B VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.25
X26 a_436_2754# a_323_2354# OUT_B VCCHIB sky130_fd_pr__pfet_01v8 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.25
X27 a_323_2354# a_114_2354# VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.25
X28 OUT OUT_B VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.25
X29 OUT_B a_323_2354# a_823_n317# VSSD sky130_fd_pr__nfet_01v8 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.25
X30 OUT_B IN_VCCHIB a_1679_n317# VSSD sky130_fd_pr__nfet_01v8 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.25
.ends

.subckt sky130_fd_io__gpiov2_inbuf_lvinv_x1 IN VGND VPWR OUT
X0 VPWR IN OUT VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.25
X1 VGND IN OUT VGND sky130_fd_pr__nfet_01v8 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.25
.ends

.subckt sky130_fd_io__gpiov2_ibuf_se VTRIP_SEL_H_N VCCHIB ENABLE_VDDIO_LV MODE_NORMAL_N
+ IBUFMUX_OUT IN_VT IN_H VTRIP_SEL_H MODE_VCCHIB_N sky130_fd_io__gpiov2_in_buf_0/m1_n467_n748#
+ VDDIO_Q VSSD sky130_fd_io__gpiov2_ipath_lvls_0/a_323_2354# IBUFMUX_OUT_H
Xsky130_fd_io__gpiov2_ipath_hvls_0 IBUFMUX_OUT_H sky130_fd_io__gpiov2_ipath_hvls_0/OUT_B
+ MODE_NORMAL_N sky130_fd_io__gpiov2_vcchib_in_buf_0/OUT sky130_fd_io__gpiov2_vcchib_in_buf_0/OUT_N
+ sky130_fd_io__gpiov2_in_buf_0/OUT MODE_VCCHIB_N sky130_fd_io__gpiov2_ipath_hvls_0/MODE_NORMAL
+ sky130_fd_io__gpiov2_ipath_hvls_0/MODE_VCCHIB VDDIO_Q VSSD sky130_fd_io__gpiov2_ipath_hvls
Xsky130_fd_io__gpiov2_vcchib_in_buf_0 IN_H sky130_fd_io__gpiov2_inbuf_lvinv_x1_1/IN
+ VCCHIB VSSD sky130_fd_io__gpiov2_vcchib_in_buf_0/OUT sky130_fd_io__gpiov2_vcchib_in_buf_0/OUT_N
+ sky130_fd_io__gpiov2_vcchib_in_buf
Xsky130_fd_io__gpiov2_in_buf_0 sky130_fd_io__gpiov2_in_buf_0/OUT sky130_fd_io__gpiov2_in_buf_0/OUT_N
+ MODE_NORMAL_N IN_H IN_VT VTRIP_SEL_H VTRIP_SEL_H_N VDDIO_Q VSSD sky130_fd_io__gpiov2_in_buf_0/m1_n467_n748#
+ sky130_fd_io__gpiov2_in_buf
Xsky130_fd_io__gpiov2_ipath_lvls_0 sky130_fd_io__gpiov2_vcchib_in_buf_0/OUT sky130_fd_io__gpiov2_in_buf_0/OUT
+ sky130_fd_io__gpiov2_inbuf_lvinv_x1_0/OUT sky130_fd_io__gpiov2_inbuf_lvinv_x1_0/IN
+ sky130_fd_io__gpiov2_inbuf_lvinv_x1_1/OUT sky130_fd_io__gpiov2_inbuf_lvinv_x1_1/IN
+ VCCHIB VSSD IBUFMUX_OUT sky130_fd_io__gpiov2_ipath_lvls_0/OUT_B sky130_fd_io__gpiov2_ipath_lvls_0/a_323_2354#
+ sky130_fd_io__gpiov2_ipath_lvls
Xsky130_fd_io__gpiov2_inbuf_lvinv_x1_0 sky130_fd_io__gpiov2_inbuf_lvinv_x1_0/IN VSSD
+ VCCHIB sky130_fd_io__gpiov2_inbuf_lvinv_x1_0/OUT sky130_fd_io__gpiov2_inbuf_lvinv_x1
Xsky130_fd_io__gpiov2_inbuf_lvinv_x1_1 sky130_fd_io__gpiov2_inbuf_lvinv_x1_1/IN VSSD
+ VCCHIB sky130_fd_io__gpiov2_inbuf_lvinv_x1_1/OUT sky130_fd_io__gpiov2_inbuf_lvinv_x1
X0 VCCHIB ENABLE_VDDIO_LV sky130_fd_io__gpiov2_inbuf_lvinv_x1_1/IN VCCHIB sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X1 VCCHIB sky130_fd_io__gpiov2_ipath_hvls_0/MODE_NORMAL sky130_fd_io__gpiov2_inbuf_lvinv_x1_0/IN VCCHIB sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X2 VSSD MODE_NORMAL_N sky130_fd_io__gpiov2_ipath_hvls_0/MODE_NORMAL VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.185 ps=1.93 w=0.7 l=0.6
X3 sky130_fd_io__gpiov2_inbuf_lvinv_x1_1/IN sky130_fd_io__gpiov2_ipath_hvls_0/MODE_VCCHIB VCCHIB VCCHIB sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X4 sky130_fd_io__gpiov2_inbuf_lvinv_x1_0/IN ENABLE_VDDIO_LV VCCHIB VCCHIB sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X5 sky130_fd_io__gpiov2_ipath_hvls_0/MODE_VCCHIB MODE_VCCHIB_N VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X6 VDDIO_Q MODE_NORMAL_N sky130_fd_io__gpiov2_ipath_hvls_0/MODE_NORMAL VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X7 VCCHIB ENABLE_VDDIO_LV sky130_fd_io__gpiov2_inbuf_lvinv_x1_1/IN VCCHIB sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X8 VCCHIB sky130_fd_io__gpiov2_ipath_hvls_0/MODE_NORMAL sky130_fd_io__gpiov2_inbuf_lvinv_x1_0/IN VCCHIB sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X9 sky130_fd_io__gpiov2_ipath_hvls_0/MODE_VCCHIB MODE_VCCHIB_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X10 sky130_fd_io__gpiov2_inbuf_lvinv_x1_1/IN sky130_fd_io__gpiov2_ipath_hvls_0/MODE_VCCHIB VCCHIB VCCHIB sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X11 sky130_fd_io__gpiov2_inbuf_lvinv_x1_0/IN ENABLE_VDDIO_LV VCCHIB VCCHIB sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X12 VDDIO_Q MODE_NORMAL_N sky130_fd_io__gpiov2_ipath_hvls_0/MODE_NORMAL VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X13 sky130_fd_io__gpiov2_ipath_hvls_0/MODE_VCCHIB MODE_VCCHIB_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X14 VSSD ENABLE_VDDIO_LV a_10411_1726# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X15 sky130_fd_io__gpiov2_inbuf_lvinv_x1_0/IN sky130_fd_io__gpiov2_ipath_hvls_0/MODE_NORMAL a_10763_1726# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X16 a_10411_1726# sky130_fd_io__gpiov2_ipath_hvls_0/MODE_VCCHIB sky130_fd_io__gpiov2_inbuf_lvinv_x1_1/IN VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.185 ps=1.93 w=0.7 l=0.6
X17 a_10763_1726# ENABLE_VDDIO_LV VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
.ends

.subckt sky130_fd_io__signal_5_sym_hv_local_5term GATE NWELLRING VGND NBODY IN m1_204_67#
X0 IN GATE VGND NBODY sky130_fd_pr__esd_nfet_g5v0d10v5 ad=3.73 pd=11.4 as=3.73 ps=11.4 w=5.75 l=0.6
R0 NBODY m1_534_67# sky130_fd_pr__res_generic_m1 w=0.02 l=5m
R1 NWELLRING m1_204_67# sky130_fd_pr__res_generic_m1 w=0.02 l=5m
.ends

.subckt sky130_fd_io__gpiov2_buf_localesd VTRIP_SEL_H OUT_VT VDDIO_Q OUT_H IN_H VSSD
Xsky130_fd_io__signal_5_sym_hv_local_5term_0 VSSD VDDIO_Q VSSD VSSD OUT_H VDDIO_Q
+ sky130_fd_io__signal_5_sym_hv_local_5term
Xsky130_fd_io__signal_5_sym_hv_local_5term_1 VSSD VDDIO_Q OUT_H VSSD VDDIO_Q VDDIO_Q
+ sky130_fd_io__signal_5_sym_hv_local_5term
Xsky130_fd_io__res250only_small_0 IN_H OUT_H sky130_fd_io__res250only_small
X0 OUT_H VTRIP_SEL_H OUT_VT VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=1
.ends

.subckt sky130_fd_io__gpiov2_ipath ENABLE_VDDIO_LV OUT_H VCCHIB DM_H_N[1] DM_H_N[0]
+ DM_H_N[2] INP_DIS_H_N IB_MODE_SEL_H IB_MODE_SEL_H_N VTRIP_SEL_H_N PAD OUT VSSD MODE_VCCHIB_N
+ m1_2058_35701# VDDIO_Q
Xsky130_fd_io__gpiov2_ibuf_se_0 sky130_fd_io__gpiov2_ibuf_se_0/VTRIP_SEL_H_N VCCHIB
+ ENABLE_VDDIO_LV sky130_fd_io__gpiov2_ibuf_se_0/MODE_NORMAL_N OUT sky130_fd_io__gpiov2_ibuf_se_0/IN_VT
+ sky130_fd_io__gpiov2_ibuf_se_0/IN_H sky130_fd_io__gpiov2_ibuf_se_0/VTRIP_SEL_H MODE_VCCHIB_N
+ PAD VDDIO_Q VSSD m2_15184_37210# OUT_H sky130_fd_io__gpiov2_ibuf_se
Xsky130_fd_io__gpiov2_buf_localesd_0 sky130_fd_io__gpiov2_ibuf_se_0/VTRIP_SEL_H sky130_fd_io__gpiov2_ibuf_se_0/IN_VT
+ VDDIO_Q sky130_fd_io__gpiov2_ibuf_se_0/IN_H PAD VSSD sky130_fd_io__gpiov2_buf_localesd
X0 VDDIO_Q a_9920_140# sky130_fd_io__gpiov2_ibuf_se_0/MODE_NORMAL_N VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X1 VDDIO_Q DM_H_N[2] a_10749_140# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X2 a_10749_140# a_11211_140# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X3 VSSD a_9920_140# a_9864_832# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X4 VSSD DM_H_N[2] a_11331_832# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X5 a_11331_832# a_11211_140# a_10749_140# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.185 ps=1.93 w=0.7 l=0.6
X6 VDDIO_Q sky130_fd_io__gpiov2_ibuf_se_0/VTRIP_SEL_H sky130_fd_io__gpiov2_ibuf_se_0/VTRIP_SEL_H_N VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X7 a_9399_166# VTRIP_SEL_H_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X8 a_10573_140# a_10749_140# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X9 VDDIO_Q a_10573_140# a_9920_140# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X10 a_11211_140# a_11563_140# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X11 VSSD a_10573_140# a_9920_140# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.185 ps=1.93 w=0.7 l=0.6
X12 a_11211_140# a_11563_140# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X13 sky130_fd_io__gpiov2_ibuf_se_0/VTRIP_SEL_H sky130_fd_io__gpiov2_ibuf_se_0/MODE_NORMAL_N a_9399_166# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X14 VDDIO_Q INP_DIS_H_N a_10573_140# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X15 MODE_VCCHIB_N a_9920_140# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X16 VDDIO_Q sky130_fd_io__gpiov2_ibuf_se_0/VTRIP_SEL_H sky130_fd_io__gpiov2_ibuf_se_0/VTRIP_SEL_H_N VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X17 a_9399_166# VTRIP_SEL_H_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X18 a_10573_140# a_10749_140# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X19 VSSD sky130_fd_io__gpiov2_ibuf_se_0/VTRIP_SEL_H sky130_fd_io__gpiov2_ibuf_se_0/VTRIP_SEL_H_N VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.185 ps=1.93 w=0.7 l=0.6
X20 sky130_fd_io__gpiov2_ibuf_se_0/VTRIP_SEL_H VTRIP_SEL_H_N VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X21 a_10869_832# a_10749_140# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X22 sky130_fd_io__gpiov2_ibuf_se_0/MODE_NORMAL_N IB_MODE_SEL_H_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X23 VDDIO_Q DM_H_N[1] a_11563_140# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X24 a_11563_140# DM_H_N[0] VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X25 VDDIO_Q IB_MODE_SEL_H MODE_VCCHIB_N VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X26 sky130_fd_io__gpiov2_ibuf_se_0/VTRIP_SEL_H sky130_fd_io__gpiov2_ibuf_se_0/MODE_NORMAL_N a_9399_166# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X27 VDDIO_Q INP_DIS_H_N a_10573_140# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X28 VSSD sky130_fd_io__gpiov2_ibuf_se_0/MODE_NORMAL_N sky130_fd_io__gpiov2_ibuf_se_0/VTRIP_SEL_H VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.196 pd=1.96 as=0.098 ps=0.98 w=0.7 l=0.6
X29 a_10573_140# INP_DIS_H_N a_10869_832# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X30 VDDIO_Q a_9920_140# sky130_fd_io__gpiov2_ibuf_se_0/MODE_NORMAL_N VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X31 VDDIO_Q DM_H_N[2] a_10749_140# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X32 MODE_VCCHIB_N a_9920_140# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X33 a_10749_140# a_11211_140# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X34 a_10216_832# a_9920_140# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X35 sky130_fd_io__gpiov2_ibuf_se_0/MODE_NORMAL_N IB_MODE_SEL_H_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X36 VDDIO_Q DM_H_N[1] a_11563_140# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X37 a_9864_832# IB_MODE_SEL_H_N sky130_fd_io__gpiov2_ibuf_se_0/MODE_NORMAL_N VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.185 ps=1.93 w=0.7 l=0.6
X38 VDDIO_Q a_10573_140# a_9920_140# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X39 VSSD DM_H_N[1] a_11969_832# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X40 VDDIO_Q IB_MODE_SEL_H MODE_VCCHIB_N VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X41 a_11563_140# DM_H_N[0] VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X42 a_11211_140# a_11563_140# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X43 a_11969_832# DM_H_N[0] a_11563_140# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.185 ps=1.93 w=0.7 l=0.6
X44 MODE_VCCHIB_N IB_MODE_SEL_H a_10216_832# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
.ends

.subckt sky130_fd_io__com_ctl_ls_en_1_v2 DM[1] VCC_IO VPB OUT_H_N OUT_H RST_H SET_H
+ VPWR HLD_H_N a_1150_n777# w_1114_n948# a_1762_n1276# a_n17_1379#
X0 a_361_1391# VPWR a_128_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X1 VCC_IO a_130_181# OUT_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X2 a_128_1391# VPWR a_361_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X3 a_n17_1379# a_634_829# a_128_1391# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 a_128_1391# a_634_829# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.15
X5 a_361_1391# HLD_H_N a_130_181# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.6
X6 a_361_1391# VPWR a_128_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X7 a_n17_1379# a_634_829# a_128_1391# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8 OUT_H_N a_65_861# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X9 a_n17_1379# a_992_934# a_724_1391# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10 a_1150_n777# DM[1] a_992_934# w_1114_n948# sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.25
X11 a_128_1391# a_634_829# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 a_724_1391# a_992_934# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13 a_65_861# HLD_H_N a_957_1391# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X14 OUT_H a_130_181# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.28 pd=2.56 as=0.14 ps=1.28 w=1 l=0.6
X15 a_n17_1379# a_992_934# a_724_1391# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X16 a_65_861# a_130_181# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.199 ps=2.03 w=0.75 l=0.5
X17 a_724_1391# a_992_934# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X18 a_n17_1379# a_65_861# a_130_181# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.199 ps=2.03 w=0.75 l=1
X19 a_634_829# a_992_934# a_1150_n777# w_1114_n948# sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.25
X20 a_957_1391# VPWR a_724_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X21 a_n17_1379# a_65_861# OUT_H_N a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.6
X22 a_130_181# a_65_861# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.199 ps=2.03 w=0.75 l=0.5
X23 a_724_1391# VPWR a_957_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X24 a_957_1391# VPWR a_724_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X25 a_65_861# a_130_181# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.105 ps=1.03 w=0.75 l=1
X26 a_130_181# SET_H a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X27 a_1762_n1276# DM[1] a_992_934# a_n17_1379# sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.25
X28 a_724_1391# VPWR a_957_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X29 a_n17_1379# RST_H a_65_861# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X30 a_634_829# a_992_934# a_1762_n1276# a_n17_1379# sky130_fd_pr__nfet_01v8 ad=0.28 pd=2.56 as=0.14 ps=1.28 w=1 l=0.25
X31 a_128_1391# VPWR a_361_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
.ends

.subckt sky130_fd_io__com_ctl_ls_v2 VCC_IO VPB OUT_H_N OUT_H IN RST_H SET_H VPWR HLD_H_N
+ a_n17_1379#
X0 a_361_1391# VPWR a_128_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X1 VCC_IO a_130_181# OUT_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X2 a_128_1391# VPWR a_361_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X3 a_n17_1379# a_634_829# a_128_1391# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 a_128_1391# a_634_829# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.15
X5 a_361_1391# HLD_H_N a_130_181# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.6
X6 a_634_829# a_992_934# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.25
X7 a_361_1391# VPWR a_128_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X8 a_n17_1379# a_634_829# a_128_1391# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9 OUT_H_N a_65_861# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X10 a_n17_1379# a_992_934# a_724_1391# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11 a_128_1391# a_634_829# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 a_724_1391# a_992_934# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13 a_65_861# HLD_H_N a_957_1391# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X14 OUT_H a_130_181# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.28 pd=2.56 as=0.14 ps=1.28 w=1 l=0.6
X15 a_n17_1379# a_992_934# a_724_1391# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X16 a_65_861# a_130_181# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.199 ps=2.03 w=0.75 l=0.5
X17 a_724_1391# a_992_934# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X18 a_n17_1379# a_65_861# a_130_181# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.199 ps=2.03 w=0.75 l=1
X19 VPWR IN a_992_934# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.25
X20 a_957_1391# VPWR a_724_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X21 a_n17_1379# IN a_992_934# a_n17_1379# sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.25
X22 a_n17_1379# a_65_861# OUT_H_N a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.6
X23 a_130_181# a_65_861# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.199 ps=2.03 w=0.75 l=0.5
X24 a_724_1391# VPWR a_957_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X25 a_957_1391# VPWR a_724_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X26 a_65_861# a_130_181# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.105 ps=1.03 w=0.75 l=1
X27 a_634_829# a_992_934# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8 ad=0.28 pd=2.56 as=0.14 ps=1.28 w=1 l=0.25
X28 a_130_181# SET_H a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X29 a_724_1391# VPWR a_957_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X30 a_n17_1379# RST_H a_65_861# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X31 a_128_1391# VPWR a_361_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
.ends

.subckt sky130_fd_io__com_ctl_lsv2 SET_H HLD_H_N VGND OUT_H OUT_H_N RST_H VPWR VCC_IO
+ m1_5675_1428# w_5775_333# w_4727_n1281# m1_5585_1428# IN
X0 a_4739_1530# HLD_H_N a_4700_968# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X1 OUT_H a_4739_1530# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X2 OUT_H_N a_4793_n866# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X3 a_4700_638# VPWR a_4933_638# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.9
X4 VGND SET_H a_4739_1530# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X5 VGND a_4739_1530# OUT_H VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X6 VCC_IO a_4793_n866# a_4739_1530# w_4727_n1281# sky130_fd_pr__pfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.199 ps=2.03 w=0.75 l=0.5
X7 a_4700_968# VPWR a_4933_968# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.9
X8 a_4933_968# a_4944_2840# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9 a_4793_n866# RST_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X10 VGND IN a_4944_2496# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.25
X11 a_4933_968# a_4944_2840# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 a_4933_638# VPWR a_4700_638# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X13 a_4933_638# HLD_H_N a_4793_n866# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X14 a_4933_968# VPWR a_4700_968# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X15 a_4700_968# VPWR a_4933_968# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X16 VCC_IO a_4793_n866# OUT_H_N VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X17 VGND a_4944_2840# a_4933_968# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X18 VGND a_4944_2496# a_4700_638# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X19 VGND a_4944_2496# a_4700_638# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X20 a_4944_2840# a_4944_2496# VPWR w_5775_333# sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.25
X21 a_4933_638# VPWR a_4700_638# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.9
X22 VCC_IO a_4739_1530# a_4793_n866# w_4727_n1281# sky130_fd_pr__pfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.199 ps=2.03 w=0.75 l=0.5
X23 a_4739_1530# a_4793_n866# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.199 ps=2.03 w=0.75 l=1
X24 a_4933_638# VPWR a_4700_638# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X25 a_4944_2840# a_4944_2496# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.25
X26 VGND a_4944_2840# a_4933_968# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X27 a_4793_n866# a_4739_1530# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.199 ps=2.03 w=0.75 l=1
X28 a_4933_968# VPWR a_4700_968# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.9
X29 VPWR IN a_4944_2496# w_5775_333# sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.25
X30 a_4700_638# a_4944_2496# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X31 a_4700_638# a_4944_2496# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
.ends

.subckt sky130_fd_io__com_ctl_ls_1v2 VCC_IO VPB OUT_H_N OUT_H IN RST_H SET_H VPWR
+ HLD_H_N a_n17_1379#
X0 a_361_1391# VPWR a_128_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X1 VCC_IO a_130_181# OUT_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X2 a_128_1391# VPWR a_361_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X3 a_n17_1379# a_634_829# a_128_1391# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 a_128_1391# a_634_829# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.15
X5 a_361_1391# HLD_H_N a_130_181# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.6
X6 a_634_829# a_992_934# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.25
X7 a_361_1391# VPWR a_128_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X8 a_n17_1379# a_634_829# a_128_1391# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9 OUT_H_N a_65_861# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X10 a_n17_1379# a_992_934# a_724_1391# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11 a_128_1391# a_634_829# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 a_724_1391# a_992_934# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13 a_65_861# HLD_H_N a_957_1391# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X14 OUT_H a_130_181# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.28 pd=2.56 as=0.14 ps=1.28 w=1 l=0.6
X15 a_n17_1379# a_992_934# a_724_1391# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X16 a_65_861# a_130_181# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.199 ps=2.03 w=0.75 l=0.5
X17 a_724_1391# a_992_934# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X18 a_n17_1379# a_65_861# a_130_181# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.199 ps=2.03 w=0.75 l=1
X19 VPWR IN a_992_934# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.25
X20 a_957_1391# VPWR a_724_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X21 a_n17_1379# IN a_992_934# a_n17_1379# sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.25
X22 a_n17_1379# a_65_861# OUT_H_N a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.6
X23 a_130_181# a_65_861# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.199 ps=2.03 w=0.75 l=0.5
X24 a_724_1391# VPWR a_957_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X25 a_957_1391# VPWR a_724_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X26 a_65_861# a_130_181# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.105 ps=1.03 w=0.75 l=1
X27 a_634_829# a_992_934# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8 ad=0.28 pd=2.56 as=0.14 ps=1.28 w=1 l=0.25
X28 a_130_181# SET_H a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X29 a_724_1391# VPWR a_957_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X30 a_n17_1379# RST_H a_65_861# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X31 a_128_1391# VPWR a_361_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
.ends

.subckt sky130_fd_io__gpiov2_ctl_lsbank VTRIP_SEL_H VTRIP_SEL INP_DIS INP_DIS_H DM[0]
+ DM_H[0] DM[2] DM_H[2] DM_H_N[2] VCC_IO STARTUP_ST_H STARTUP_RST_H OD_I_H IB_MODE_SEL_H_N
+ IB_MODE_SEL sky130_fd_io__com_ctl_ls_en_1_v2_0/a_1762_n1276# sky130_fd_io__com_ctl_lsv2_0/VCC_IO
+ DM_H[1] INP_DIS_H_N w_15552_2653# m1_2266_545# DM_H_N[1] DM[1] DM_H_N[0] VTRIP_SEL_H_N
+ HLD_I_H_N IB_MODE_SEL_H VPWR VGND
Xsky130_fd_io__com_ctl_ls_en_1_v2_0 DM[1] VCC_IO VPWR DM_H_N[1] DM_H[1] sky130_fd_io__com_ctl_ls_en_1_v2_0/RST_H
+ sky130_fd_io__com_ctl_ls_en_1_v2_0/SET_H VPWR HLD_I_H_N VPWR VPWR sky130_fd_io__com_ctl_ls_en_1_v2_0/a_1762_n1276#
+ VGND sky130_fd_io__com_ctl_ls_en_1_v2
Xsky130_fd_io__com_ctl_ls_v2_0 VCC_IO VPWR DM_H_N[2] DM_H[2] DM[2] sky130_fd_io__com_ctl_ls_v2_0/RST_H
+ sky130_fd_io__com_ctl_ls_v2_0/SET_H VPWR HLD_I_H_N VGND sky130_fd_io__com_ctl_ls_v2
Xsky130_fd_io__com_ctl_ls_v2_1 VCC_IO VPWR INP_DIS_H_N INP_DIS_H INP_DIS sky130_fd_io__com_ctl_ls_v2_1/RST_H
+ sky130_fd_io__com_ctl_ls_v2_1/SET_H VPWR HLD_I_H_N VGND sky130_fd_io__com_ctl_ls_v2
Xsky130_fd_io__com_ctl_ls_v2_2 VCC_IO VPWR DM_H_N[0] DM_H[0] DM[0] sky130_fd_io__com_ctl_ls_v2_2/RST_H
+ sky130_fd_io__com_ctl_ls_v2_2/SET_H VPWR HLD_I_H_N VGND sky130_fd_io__com_ctl_ls_v2
Xsky130_fd_io__com_ctl_lsv2_0 sky130_fd_io__com_ctl_lsv2_0/SET_H HLD_I_H_N VGND IB_MODE_SEL_H
+ IB_MODE_SEL_H_N sky130_fd_io__com_ctl_lsv2_0/RST_H VPWR sky130_fd_io__com_ctl_lsv2_0/VCC_IO
+ VGND VPWR w_15552_2653# VGND IB_MODE_SEL sky130_fd_io__com_ctl_lsv2
Xsky130_fd_io__com_ctl_ls_1v2_0 VCC_IO VPWR VTRIP_SEL_H_N VTRIP_SEL_H VTRIP_SEL sky130_fd_io__com_ctl_ls_1v2_0/RST_H
+ sky130_fd_io__com_ctl_ls_1v2_0/SET_H VPWR HLD_I_H_N VGND sky130_fd_io__com_ctl_ls_1v2
R0 sky130_fd_io__com_ctl_ls_en_1_v2_0/SET_H m1_2266_320# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R1 m1_14183_362# sky130_fd_io__com_ctl_ls_1v2_0/RST_H sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R2 m1_6620_334# STARTUP_ST_H sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R3 m2_15089_329# sky130_fd_io__com_ctl_lsv2_0/SET_H sky130_fd_pr__res_generic_m2 w=0.26 l=10m
R4 STARTUP_RST_H m1_6420_507# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R5 m1_5875_412# STARTUP_RST_H sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R6 m1_6148_320# STARTUP_ST_H sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R7 m1_10303_506# sky130_fd_io__com_ctl_ls_v2_0/SET_H sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R8 sky130_fd_io__com_ctl_ls_v2_1/RST_H m1_6620_334# sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R9 m1_14183_362# OD_I_H sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R10 sky130_fd_io__com_ctl_ls_v2_2/SET_H m1_6148_320# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R11 OD_I_H m1_10303_543# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R12 m1_10029_412# OD_I_H sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R13 m2_15027_104# sky130_fd_io__com_ctl_lsv2_0/SET_H sky130_fd_pr__res_generic_m2 w=0.26 l=10m
R14 m1_6707_412# sky130_fd_io__com_ctl_ls_v2_1/RST_H sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R15 m1_6421_319# STARTUP_ST_H sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R16 m1_14456_624# sky130_fd_io__com_ctl_ls_1v2_0/SET_H sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R17 m1_5955_333# STARTUP_ST_H sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R18 m1_14457_430# OD_I_H sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R19 m2_14799_410# OD_I_H sky130_fd_pr__res_generic_m2 w=0.26 l=10m
R20 sky130_fd_io__com_ctl_ls_v2_1/SET_H m1_6421_356# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R21 m2_14799_410# sky130_fd_io__com_ctl_lsv2_0/RST_H sky130_fd_pr__res_generic_m2 w=0.26 l=10m
R22 VGND m2_15089_329# sky130_fd_pr__res_generic_m2 w=0.26 l=10m
R23 VGND m1_14456_624# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R24 sky130_fd_io__com_ctl_ls_v2_2/RST_H m1_5955_370# sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R25 sky130_fd_io__com_ctl_ls_1v2_0/SET_H m1_14457_467# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R26 m1_10109_333# VGND sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R27 m1_10302_320# VGND sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R28 m1_2553_412# m1_2266_545# sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R29 sky130_fd_io__com_ctl_ls_v2_0/RST_H m1_10109_370# sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R30 sky130_fd_io__com_ctl_ls_v2_0/SET_H m1_10302_320# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R31 m1_2267_506# sky130_fd_io__com_ctl_ls_en_1_v2_0/SET_H sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R32 m1_14263_617# sky130_fd_io__com_ctl_ls_1v2_0/RST_H sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R33 m1_2467_333# VGND sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R34 m1_2266_545# m1_2267_543# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R35 VGND m1_14263_654# sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R36 sky130_fd_io__com_ctl_ls_en_1_v2_0/RST_H m1_2467_370# sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R37 m1_6149_506# sky130_fd_io__com_ctl_ls_v2_2/SET_H sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R38 m1_14911_509# sky130_fd_io__com_ctl_lsv2_0/RST_H sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R39 m1_10029_412# sky130_fd_io__com_ctl_ls_v2_0/RST_H sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R40 m2_14990_104# OD_I_H sky130_fd_pr__res_generic_m2 w=0.26 l=10m
R41 STARTUP_RST_H m1_6149_543# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R42 m1_2553_412# sky130_fd_io__com_ctl_ls_en_1_v2_0/RST_H sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R43 VGND m1_14911_546# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R44 m1_2266_320# VGND sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R45 m1_6744_412# STARTUP_RST_H sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R46 m1_5875_412# sky130_fd_io__com_ctl_ls_v2_2/RST_H sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R47 m1_6420_507# sky130_fd_io__com_ctl_ls_v2_1/SET_H sky130_fd_pr__res_generic_m1 w=0.26 l=10m
.ends

.subckt sky130_fd_io__com_ctl_ls VCC_IO VPB OUT_H_N OUT_H IN RST_H SET_H VPWR HLD_H_N
+ a_n17_1379#
X0 a_361_1391# VPWR a_128_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X1 VCC_IO a_130_181# OUT_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X2 a_128_1391# VPWR a_361_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X3 a_n17_1379# a_634_829# a_128_1391# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 a_128_1391# a_634_829# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.15
X5 a_361_1391# HLD_H_N a_130_181# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.6
X6 a_634_829# a_992_934# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.25
X7 a_361_1391# VPWR a_128_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X8 a_n17_1379# a_634_829# a_128_1391# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9 OUT_H_N a_65_861# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X10 a_n17_1379# a_992_934# a_724_1391# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11 a_128_1391# a_634_829# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 a_724_1391# a_992_934# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13 a_65_861# HLD_H_N a_957_1391# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X14 OUT_H a_130_181# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.28 pd=2.56 as=0.14 ps=1.28 w=1 l=0.6
X15 a_n17_1379# a_992_934# a_724_1391# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X16 a_65_861# a_130_181# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.199 ps=2.03 w=0.75 l=0.5
X17 a_724_1391# a_992_934# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X18 a_n17_1379# a_65_861# a_130_181# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.199 ps=2.03 w=0.75 l=1
X19 VPWR IN a_992_934# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.25
X20 a_957_1391# VPWR a_724_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X21 a_n17_1379# IN a_992_934# a_n17_1379# sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.25
X22 a_n17_1379# a_65_861# OUT_H_N a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.6
X23 a_130_181# a_65_861# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.199 ps=2.03 w=0.75 l=0.5
X24 a_724_1391# VPWR a_957_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X25 a_957_1391# VPWR a_724_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X26 a_65_861# a_130_181# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.105 ps=1.03 w=0.75 l=1
X27 a_634_829# a_992_934# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8 ad=0.28 pd=2.56 as=0.14 ps=1.28 w=1 l=0.25
X28 a_130_181# SET_H a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X29 a_724_1391# VPWR a_957_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X30 a_n17_1379# RST_H a_65_861# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X31 a_128_1391# VPWR a_361_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
.ends

.subckt sky130_fd_io__com_ctl_hldv2 HLD_OVR VCC_IO VGND HLD_I_H_N OD_I_H VPWR HLD_I_H
+ sky130_fd_io__com_ctl_ls_0/VCC_IO sky130_fd_io__com_ctl_ls_0/VPB a_8218_3918# a_3023_3554#
+ m2_3556_4143# m1_3684_4201# a_2671_3554# m2_3665_4182#
Xsky130_fd_io__com_ctl_ls_0 sky130_fd_io__com_ctl_ls_0/VCC_IO sky130_fd_io__com_ctl_ls_0/VPB
+ sky130_fd_io__com_ctl_ls_0/OUT_H_N sky130_fd_io__com_ctl_ls_0/OUT_H HLD_OVR sky130_fd_io__com_ctl_ls_0/RST_H
+ VGND VPWR sky130_fd_io__com_ctl_ls_0/HLD_H_N VGND sky130_fd_io__com_ctl_ls
X0 a_2967_3580# a_2671_3554# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X1 sky130_fd_io__com_ctl_ls_0/HLD_H_N a_2967_3918# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.6
X2 a_3743_3580# sky130_fd_io__com_ctl_ls_0/HLD_H_N VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.185 ps=1.93 w=0.7 l=0.6
X3 VCC_IO sky130_fd_io__com_ctl_ls_0/HLD_H_N a_3743_3580# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X4 VGND a_3743_3580# a_4447_3580# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X5 a_4447_3580# a_3743_3580# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X6 VCC_IO a_3743_3580# a_4447_3580# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X7 a_5855_3580# a_3743_3580# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X8 VCC_IO a_3743_3580# a_4447_3580# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X9 a_5855_3580# a_3743_3580# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X10 a_5855_3580# a_3743_3580# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X11 VCC_IO a_3743_3580# a_5855_3580# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X12 VCC_IO sky130_fd_io__com_ctl_ls_0/RST_H a_7214_3580# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X13 OD_I_H a_7214_3580# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X14 VCC_IO a_7214_3580# OD_I_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X15 VCC_IO OD_I_H a_8391_3918# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X16 VGND a_2671_3554# sky130_fd_io__com_ctl_ls_0/RST_H VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.185 ps=1.93 w=0.7 l=0.6
X17 VCC_IO a_3023_3554# a_2967_3918# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X18 VGND sky130_fd_io__com_ctl_ls_0/HLD_H_N a_3743_3580# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X19 a_4447_3580# a_3743_3580# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X20 a_4447_3580# a_3743_3580# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X21 VCC_IO a_3743_3580# a_5855_3580# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X22 a_5855_3580# a_3743_3580# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X23 VCC_IO a_3743_3580# a_5855_3580# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X24 VCC_IO a_3743_3580# a_5855_3580# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X25 OD_I_H a_7214_3580# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X26 a_8391_3918# a_8271_3554# a_8218_3918# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X27 VCC_IO a_7214_3580# OD_I_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X28 a_8743_3918# sky130_fd_io__com_ctl_ls_0/HLD_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X29 a_2967_3918# a_2671_3554# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X30 a_3743_3580# sky130_fd_io__com_ctl_ls_0/HLD_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X31 a_3743_3580# sky130_fd_io__com_ctl_ls_0/HLD_H_N VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X32 a_4447_3580# a_3743_3580# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X33 VCC_IO a_3743_3580# a_4447_3580# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
R0 HLD_I_H a_3743_3580# sky130_fd_pr__res_generic_m1 w=0.23 l=10m
X34 VCC_IO a_3743_3580# a_4447_3580# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X35 a_8271_3554# sky130_fd_io__com_ctl_ls_0/OUT_H a_8743_3918# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X36 VCC_IO a_2671_3554# sky130_fd_io__com_ctl_ls_0/RST_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X37 a_5855_3580# a_3743_3580# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X38 VGND a_3743_3580# a_4447_3580# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X39 a_5855_3580# a_3743_3580# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X40 sky130_fd_io__com_ctl_ls_0/HLD_H_N a_2967_3918# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.6
X41 VCC_IO sky130_fd_io__com_ctl_ls_0/HLD_H_N a_3743_3580# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X42 VGND sky130_fd_io__com_ctl_ls_0/RST_H a_7214_3580# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.185 ps=1.93 w=0.7 l=0.6
X43 VGND a_7214_3580# OD_I_H VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X44 VCC_IO sky130_fd_io__com_ctl_ls_0/HLD_H_N a_3743_3580# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X45 VGND OD_I_H a_8218_3918# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X46 a_4447_3580# a_3743_3580# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X47 VCC_IO a_3743_3580# a_4447_3580# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X48 a_5855_3580# a_3743_3580# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X49 VCC_IO a_3743_3580# a_5855_3580# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X50 OD_I_H a_7214_3580# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X51 a_2967_3918# a_3023_3554# a_2967_3580# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X52 a_4447_3580# a_3743_3580# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X53 VGND a_3743_3580# a_5855_3580# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X54 VGND a_3743_3580# a_5855_3580# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X55 OD_I_H a_7214_3580# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X56 a_3743_3580# sky130_fd_io__com_ctl_ls_0/HLD_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X57 a_8218_3918# a_8271_3554# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.196 ps=1.96 w=0.7 l=0.6
X58 a_4447_3580# a_3743_3580# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X59 a_8271_3554# sky130_fd_io__com_ctl_ls_0/HLD_H_N VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
R1 a_4447_3580# HLD_I_H_N sky130_fd_pr__res_generic_m1 w=0.23 l=0.025
X60 VCC_IO a_3743_3580# a_5855_3580# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X61 a_5855_3580# a_3743_3580# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
R2 HLD_I_H_N a_5855_3580# sky130_fd_pr__res_generic_m1 w=0.23 l=0.025
X62 VCC_IO a_7214_3580# OD_I_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X63 a_4447_3580# a_3743_3580# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X64 VGND a_3743_3580# a_4447_3580# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X65 VCC_IO a_3743_3580# a_4447_3580# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X66 a_5855_3580# a_3743_3580# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X67 a_2967_3918# a_2671_3554# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X68 a_5855_3580# a_3743_3580# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X69 VCC_IO sky130_fd_io__com_ctl_ls_0/RST_H a_7214_3580# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X70 a_3743_3580# sky130_fd_io__com_ctl_ls_0/HLD_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X71 VCC_IO a_7214_3580# OD_I_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X72 VGND sky130_fd_io__com_ctl_ls_0/OUT_H a_8271_3554# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.196 pd=1.96 as=0.098 ps=0.98 w=0.7 l=0.6
X73 VCC_IO a_3743_3580# a_4447_3580# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X74 VCC_IO OD_I_H a_8391_3918# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X75 VCC_IO a_3023_3554# a_2967_3918# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X76 sky130_fd_io__com_ctl_ls_0/HLD_H_N a_2967_3918# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.185 ps=1.93 w=0.7 l=0.6
X77 VGND sky130_fd_io__com_ctl_ls_0/HLD_H_N a_3743_3580# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X78 a_4447_3580# a_3743_3580# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X79 VGND a_3743_3580# a_4447_3580# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X80 a_4447_3580# a_3743_3580# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X81 a_5855_3580# a_3743_3580# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X82 VCC_IO a_2671_3554# sky130_fd_io__com_ctl_ls_0/RST_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X83 VCC_IO a_3743_3580# a_5855_3580# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X84 VGND a_3743_3580# a_5855_3580# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X85 VCC_IO sky130_fd_io__com_ctl_ls_0/HLD_H_N a_3743_3580# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X86 VCC_IO a_3743_3580# a_5855_3580# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X87 OD_I_H a_7214_3580# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X88 OD_I_H a_7214_3580# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X89 a_8391_3918# a_8271_3554# a_8218_3918# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X90 a_8743_3918# sky130_fd_io__com_ctl_ls_0/HLD_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X91 a_4447_3580# a_3743_3580# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X92 a_4447_3580# a_3743_3580# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X93 VCC_IO a_3743_3580# a_4447_3580# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X94 a_5855_3580# a_3743_3580# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X95 VGND a_3743_3580# a_5855_3580# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X96 VGND a_7214_3580# OD_I_H VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X97 a_3743_3580# sky130_fd_io__com_ctl_ls_0/HLD_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X98 a_8271_3554# sky130_fd_io__com_ctl_ls_0/OUT_H a_8743_3918# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
.ends

.subckt sky130_fd_io__gpiov2_ctl DM[0] VTRIP_SEL_H_N DM[2] DM_H[0] DM_H[2] DM_H_N[1]
+ INP_DIS INP_DIS_H_N HLD_OVR VTRIP_SEL VTRIP_SEL_H OD_I_H INP_STARTUP_EN_H IB_MODE_SEL_H_N
+ IB_MODE_SEL ENABLE_INP_H HLD_H_N HLD_I_OVR_H ENABLE_H DM[1] a_11799_3638# li_18199_5031#
+ DM_H_N[0] IB_MODE_SEL_H sky130_fd_io__gpiov2_ctl_lsbank_0/sky130_fd_io__com_ctl_ls_en_1_v2_0/a_1762_n1276#
+ DM_H_N[2] DM_H[1] HLD_I_H_N VPWR sky130_fd_io__com_ctl_hldv2_0/HLD_I_H VGND VCC_IO
Xsky130_fd_io__gpiov2_ctl_lsbank_0 VTRIP_SEL_H VTRIP_SEL INP_DIS sky130_fd_io__gpiov2_ctl_lsbank_0/INP_DIS_H
+ DM[0] DM_H[0] DM[2] DM_H[2] DM_H_N[2] VCC_IO INP_STARTUP_EN_H sky130_fd_io__gpiov2_ctl_lsbank_0/STARTUP_RST_H
+ OD_I_H IB_MODE_SEL_H_N IB_MODE_SEL sky130_fd_io__gpiov2_ctl_lsbank_0/sky130_fd_io__com_ctl_ls_en_1_v2_0/a_1762_n1276#
+ VCC_IO DM_H[1] INP_DIS_H_N VCC_IO OD_I_H DM_H_N[1] DM[1] DM_H_N[0] VTRIP_SEL_H_N
+ HLD_I_H_N IB_MODE_SEL_H VPWR VGND sky130_fd_io__gpiov2_ctl_lsbank
Xsky130_fd_io__com_ctl_hldv2_0 HLD_OVR VCC_IO VGND HLD_I_H_N OD_I_H VPWR sky130_fd_io__com_ctl_hldv2_0/HLD_I_H
+ VCC_IO VPWR HLD_I_OVR_H HLD_H_N OD_I_H OD_I_H ENABLE_H OD_I_H sky130_fd_io__com_ctl_hldv2
X0 INP_STARTUP_EN_H a_11094_4330# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X1 VCC_IO ENABLE_INP_H a_11919_3664# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X2 a_11919_3664# a_11799_3638# sky130_fd_io__gpiov2_ctl_lsbank_0/STARTUP_RST_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X3 sky130_fd_io__gpiov2_ctl_lsbank_0/STARTUP_RST_H a_11799_3638# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.196 ps=1.96 w=0.7 l=0.6
X4 VCC_IO ENABLE_INP_H a_11919_3664# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X5 a_11094_4330# ENABLE_INP_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X6 VGND ENABLE_INP_H sky130_fd_io__gpiov2_ctl_lsbank_0/STARTUP_RST_H VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X7 VCC_IO OD_I_H a_11094_4330# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X8 INP_STARTUP_EN_H a_11094_4330# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X9 a_11094_4330# ENABLE_INP_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X10 a_11267_4330# ENABLE_INP_H a_11094_4330# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.185 ps=1.93 w=0.7 l=0.6
X11 VCC_IO OD_I_H a_11094_4330# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X12 a_11919_3664# a_11799_3638# sky130_fd_io__gpiov2_ctl_lsbank_0/STARTUP_RST_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X13 VGND OD_I_H a_11267_4330# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X14 INP_STARTUP_EN_H a_11094_4330# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
.ends

.subckt sky130_fd_io__top_gpiov2 VSSIO_Q PAD_A_NOESD_H ANALOG_POL ENABLE_VDDIO IN_H
+ IN DM[0] DM[1] DM[2] HLD_OVR INP_DIS ENABLE_VDDA_H VTRIP_SEL OE_N OUT SLOW TIE_LO_ESD
+ PAD_A_ESD_0_H ANALOG_SEL ENABLE_INP_H PAD_A_ESD_1_H TIE_HI_ESD ENABLE_H IB_MODE_SEL
+ ENABLE_VSWITCH_H ANALOG_EN sky130_fd_io__overlay_gpiov2_m4_0/sky130_fd_io__top_gpio_pad_0/b_1500_19531#
+ w_9674_16869# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/PG_AMX_VDDA_H_N
+ w_12765_16869# w_12765_14755# w_9674_14653# HLD_H_N VDDIO_Q VSWITCH VSSA VCCHIB
+ VDDIO PAD VDDA AMUXBUS_B VCCD AMUXBUS_A VSSIO VSSD
Xsky130_fd_io__gpio_opathv2_0 sky130_fd_io__gpiov2_ctl_0/HLD_I_OVR_H sky130_fd_io__gpiov2_ctl_0/HLD_I_H_N
+ sky130_fd_io__gpiov2_ctl_0/OD_I_H SLOW VCCD TIE_HI_ESD li_3442_6400# li_3302_6400#
+ li_7854_5377# sky130_fd_io__gpio_opathv2_0/sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/Y_H
+ sky130_fd_io__gpiov2_ctl_0/DM_H[0] sky130_fd_io__gpiov2_ctl_0/DM_H_N[0] li_7943_6398#
+ sky130_fd_io__gpiov2_ctl_0/DM_H[2] sky130_fd_io__gpiov2_ctl_0/DM_H_N[1] VSSD PAD
+ TIE_LO_ESD li_4745_6400# li_7636_6398# sky130_fd_io__gpio_opathv2_0/sky130_fd_io__gpio_odrvrv2_0/PU_H_N[2]
+ sky130_fd_io__gpiov2_ctl_0/VTRIP_SEL_H_N li_5278_5352# VSSD sky130_fd_io__gpiov2_ctl_0/DM_H[1]
+ PAD li_5245_3919# li_9062_7268# VSSIO sky130_fd_io__gpiov2_ctl_0/DM_H_N[2] li_2678_6400#
+ VDDA VSSIO li_10974_4971# VSSIO OE_N OUT VSSIO VCCHIB VDDIO sky130_fd_io__gpio_opathv2_0/sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/NBIAS
+ VSSD li_3958_5352# li_3334_5352# sky130_fd_io__gpio_opathv2
Xsky130_fd_io__gpiov2_amux_0 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_0/B
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_9/Y
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_13/ROUT sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_6/Y
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_13/Y
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_0/ROUT ANALOG_EN ANALOG_POL
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_3/B
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_10/ROUT sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_0/Y
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_8/A
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_10/ROUT sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_13/Y
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/PG_AMX_VDDA_H_N sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_3/ROUT
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_7/ROUT sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/NG_PAD_VPMP_H
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_2/Y
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_3/ROUT sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_1/B
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/NG_AMX_VPMP_H sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_13/Y
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_0/ROUT sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_2/Y
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_13/ROUT PAD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_4/ROUT
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_1/Y
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_3/Y
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_4/Y
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_11/Y
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_5/Y
+ w_12765_14755# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_3/Y
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_0/B
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/PG_AMX_VDDA_H_N PAD
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_6/Y
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_6/Y
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_11/A
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/PG_PAD_VDDIOQ_H_N sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_4/Y
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_2/B
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_8/Y
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_6/Y
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_12/Y
+ w_12765_16869# VDDA sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_8/ROUT
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_5/A
+ VSSA sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/NG_PAD_VPMP_H
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_2/B
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_13/ROUT sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_5/ROUT
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_14/Y
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/NG_AMX_VPMP_H PAD VSSA
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_7/A
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_11/A
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_10/ROUT sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_1/B
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_12/Y
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_1/Y
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_9/A
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_1/B
+ ANALOG_SEL sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_2/A
+ VCCD VSSD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_4/Y
+ PAD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_3/Y
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_11/A
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_7/Y
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/PG_PAD_VDDIOQ_H_N VSSD
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_9/ROUT w_9674_16869# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_2/Y
+ AMUXBUS_A sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_5/Y
+ VCCD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_2/A
+ VCCD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_10/ROUT sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_6/ROUT
+ VSSA AMUXBUS_B sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_10/ROUT
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_1/B
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_7/Y
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_3/ROUT sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_6/Y
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_11/Y
+ w_9674_14653# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_3/ROUT VCCD
+ VSSD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_3/ROUT OUT VDDIO_Q
+ PAD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_0/ROUT sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_3/B
+ VSSD VSSD VDDIO_Q sky130_fd_io__gpiov2_amux
Xsky130_fd_io__res75only_small_0 PAD_A_ESD_1_H sky130_fd_io__res75only_small_1/PAD
+ sky130_fd_io__res75only_small
Xsky130_fd_io__res75only_small_1 sky130_fd_io__res75only_small_1/PAD PAD sky130_fd_io__res75only_small
Xsky130_fd_io__res75only_small_2 PAD_A_ESD_0_H sky130_fd_io__res75only_small_3/PAD
+ sky130_fd_io__res75only_small
Xsky130_fd_io__res75only_small_3 sky130_fd_io__res75only_small_3/PAD PAD sky130_fd_io__res75only_small
Xsky130_fd_io__gpiov2_ipath_0 ENABLE_VDDIO IN_H VCCHIB sky130_fd_io__gpiov2_ctl_0/DM_H_N[1]
+ sky130_fd_io__gpiov2_ctl_0/DM_H_N[0] sky130_fd_io__gpiov2_ctl_0/DM_H_N[2] sky130_fd_io__gpiov2_ctl_0/INP_DIS_H_N
+ sky130_fd_io__gpiov2_ctl_0/IB_MODE_SEL_H sky130_fd_io__gpiov2_ctl_0/IB_MODE_SEL_H_N
+ sky130_fd_io__gpiov2_ctl_0/VTRIP_SEL_H_N PAD IN VSSD sky130_fd_io__gpiov2_ipath_0/MODE_VCCHIB_N
+ VDDIO VDDIO_Q sky130_fd_io__gpiov2_ipath
Xsky130_fd_io__gpiov2_ctl_0 DM[0] sky130_fd_io__gpiov2_ctl_0/VTRIP_SEL_H_N DM[2] sky130_fd_io__gpiov2_ctl_0/DM_H[0]
+ sky130_fd_io__gpiov2_ctl_0/DM_H[2] sky130_fd_io__gpiov2_ctl_0/DM_H_N[1] INP_DIS
+ sky130_fd_io__gpiov2_ctl_0/INP_DIS_H_N HLD_OVR VTRIP_SEL sky130_fd_io__gpiov2_ctl_0/VTRIP_SEL_H
+ sky130_fd_io__gpiov2_ctl_0/OD_I_H sky130_fd_io__gpiov2_ctl_0/INP_STARTUP_EN_H sky130_fd_io__gpiov2_ctl_0/IB_MODE_SEL_H_N
+ IB_MODE_SEL ENABLE_INP_H HLD_H_N sky130_fd_io__gpiov2_ctl_0/HLD_I_OVR_H ENABLE_H
+ DM[1] ENABLE_H PAD sky130_fd_io__gpiov2_ctl_0/DM_H_N[0] sky130_fd_io__gpiov2_ctl_0/IB_MODE_SEL_H
+ VSSD sky130_fd_io__gpiov2_ctl_0/DM_H_N[2] sky130_fd_io__gpiov2_ctl_0/DM_H[1] sky130_fd_io__gpiov2_ctl_0/HLD_I_H_N
+ VCCD sky130_fd_io__gpiov2_ctl_0/sky130_fd_io__com_ctl_hldv2_0/HLD_I_H VSSD VDDIO_Q
+ sky130_fd_io__gpiov2_ctl
X0 a_3218_11709# a_282_14802# a_1024_11940# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X1 VSWITCH a_1225_14186# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/NG_AMX_VPMP_H VSWITCH sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X2 a_13902_2778# VCCD a_14397_2496# VSSD sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X3 VSSIO_Q a_387_12076# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_5/ROUT VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.6 as=0.7 ps=5.28 w=5 l=0.5
X4 a_14053_2496# VCCD a_14092_2778# VSSD sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X5 a_8765_11461# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/PG_AMX_VDDA_H_N VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X6 a_7015_11461# a_6895_11435# VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X7 a_382_14828# a_231_9686# a_497_17084# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X8 VCCD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_14/Y a_6895_11435# VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X9 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/NG_AMX_VPMP_H a_478_17182# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.5
X10 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_5/ROUT a_2250_17651# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=2.1 pd=15.3 as=4.2 ps=30.6 w=15 l=0.5
X11 a_14092_2778# a_13902_2778# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.199 ps=2.03 w=0.75 l=0.5
X12 VCCD a_6895_11435# a_7015_11461# VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X13 a_3462_14827# a_3642_14801# a_620_18182# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X14 a_10924_13064# a_334_12102# a_10768_13064# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X15 a_10350_10272# VCCD a_10583_10272# VSSD sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X16 VSSA a_377_12820# a_2162_14426# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X17 VSSA a_478_17182# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/NG_AMX_VPMP_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.5
X18 VSSD a_231_9686# a_178_9778# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.398 ps=3.53 w=1.5 l=0.5
X19 a_9877_11799# a_8765_11461# a_8067_11435# VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X20 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/NG_PAD_VPMP_H a_1225_12852# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.6
X21 a_10768_13064# a_2250_17651# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_9/A VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.5
X22 a_2159_13760# a_689_12820# a_1024_12357# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X23 VCCD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_5/A a_12443_12112# VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.155 pd=1.37 as=0.14 ps=1.28 w=1 l=0.6
X24 a_9406_11799# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/NG_PAD_VPMP_H VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X25 VDDA a_184_18182# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/PG_AMX_VDDA_H_N VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.5
X26 a_8699_10272# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_9/A VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X27 VSWITCH a_1024_12357# a_387_12076# VSWITCH sky130_fd_pr__pfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.105 ps=1.03 w=0.75 l=2
X28 VCCD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_1/Y sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_5/A VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X29 a_324_14186# a_689_12820# a_789_14186# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X30 a_620_17850# a_178_9778# a_2080_14827# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.5
X31 VDDA a_497_17084# a_229_14828# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=1
X32 a_10406_10767# a_7173_10183# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X33 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/PG_AMX_VDDA_H_N a_184_18182# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.5
X34 a_1072_12852# VCCD a_593_13378# VSSA sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X35 w_12765_16869# sky130_fd_io__gpiov2_ctl_0/sky130_fd_io__com_ctl_hldv2_0/HLD_I_H VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.118 pd=1.4 as=0.118 ps=1.4 w=0.42 l=0.5
X36 a_789_14186# a_689_12820# a_324_14186# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X37 VSSA a_478_17182# a_184_18182# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.5
R0 PAD PAD_A_NOESD_H sky130_fd_pr__res_generic_m3 w=1.07 l=0.035
X38 w_9674_14653# a_6367_11435# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_6/ROUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.84 pd=6.56 as=0.84 ps=6.56 w=3 l=0.5
X39 a_620_18182# a_184_18182# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=1
X40 a_1079_9778# a_282_14802# a_926_9778# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.398 ps=3.53 w=1.5 l=0.5
X41 a_6367_11435# a_6543_11435# VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X42 a_1225_14186# a_689_12820# a_1072_14186# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.398 ps=3.53 w=1.5 l=0.5
X43 a_11173_10272# VCCD a_10940_10272# VSSD sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X44 a_9067_10698# VCCD a_8699_10272# VSSD sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X45 a_2250_17651# a_7173_10183# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X46 VSSIO_Q a_387_12076# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_5/ROUT VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X47 VSSD ANALOG_EN a_13816_1289# VSSD sky130_fd_pr__nfet_01v8 ad=0.263 pd=2.19 as=0.211 ps=2.05 w=0.74 l=0.15
X48 a_3218_11709# ENABLE_VSWITCH_H VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.5
X49 a_1077_11842# a_1024_11940# VSWITCH VSWITCH sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=1
X50 VSSA VSSA a_387_12076# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X51 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/NG_PAD_VPMP_H a_1225_14186# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.6
X52 VSSD a_6895_11435# a_7015_11461# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X53 VDDA ENABLE_VDDA_H a_195_17182# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X54 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_7/A a_11131_11430# VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.155 ps=1.37 w=0.42 l=0.5
X55 a_643_12102# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/NG_PAD_VPMP_H VSWITCH VSWITCH sky130_fd_pr__pfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X56 a_8067_11435# a_8765_11461# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.196 ps=1.96 w=0.7 l=0.6
X57 a_229_14828# a_282_14802# a_382_14828# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X58 a_2749_13760# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_0/Y VSSA VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X59 a_7367_11461# a_7015_11461# VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X60 w_9674_14653# sky130_fd_io__gpiov2_ctl_0/sky130_fd_io__com_ctl_hldv2_0/HLD_I_H VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.118 pd=1.4 as=0.118 ps=1.4 w=0.42 l=0.5
X61 a_593_13760# VCCD a_1072_14186# VSSA sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X62 a_2982_13760# a_689_12820# a_2162_14426# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.398 ps=3.53 w=1.5 l=0.5
X63 a_6895_11435# a_7539_11435# VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X64 VSWITCH a_387_12076# a_334_12102# VSWITCH sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.398 ps=3.53 w=1.5 l=0.5
X65 a_643_12102# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/NG_PAD_VPMP_H VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.105 ps=1.03 w=0.75 l=0.5
X66 a_14092_2778# VCCD a_14053_2496# VSSD sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X67 a_13970_2496# a_13760_1103# a_14053_2496# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
R1 PAD_A_NOESD_H PAD sky130_fd_pr__res_generic_m4 w=12.4 l=0.035
X68 a_7539_11435# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/NG_PAD_VPMP_H VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.185 ps=1.93 w=0.7 l=0.6
X69 VSSA a_387_12076# a_334_12102# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.199 ps=2.03 w=0.75 l=0.5
X70 VSWITCH a_1225_12852# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/NG_PAD_VPMP_H VSWITCH sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X71 VSWITCH a_1024_12357# a_2162_14426# VSWITCH sky130_fd_pr__pfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.185 ps=1.93 w=0.7 l=0.6
X72 VSSIO_Q a_387_12076# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_4/ROUT VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X73 VCCD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/PG_PAD_VDDIOQ_H_N a_8765_11461# VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X74 a_14397_2496# VCCD a_13902_2778# VSSD sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.9
X75 VCCD a_10643_12610# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_9/A VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.155 pd=1.37 as=0.111 ps=1.37 w=0.42 l=0.5
X76 VSSA a_787_17182# a_2080_14827# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.5
X77 a_9350_10698# VCCD a_8871_10272# VSSD sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X78 a_6543_11435# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_2/Y VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X79 a_324_14186# a_377_12820# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X80 a_593_13760# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_9/Y VSSA VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X81 a_2392_13760# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_7/Y VSSA VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X82 VSSA a_377_12820# a_324_14186# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.398 ps=3.53 w=1.5 l=0.5
X83 a_2080_14827# a_1079_9778# a_184_17734# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X84 VSSD a_7173_10183# a_2250_17651# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.6
X85 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/PG_AMX_VDDA_H_N a_184_18182# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.5
X86 VSSA a_195_17182# w_12765_16869# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.118 pd=1.4 as=0.118 ps=1.4 w=0.42 l=0.5
X87 a_1072_12852# a_689_12820# a_1225_12852# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X88 VDDIO_Q a_2250_17651# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_4/ROUT VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=2.1 pd=15.3 as=2.1 ps=15.3 w=15 l=0.5
X89 a_178_9778# a_282_14802# a_643_9778# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X90 VCCD a_6367_11435# a_6314_11461# VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X91 VSSA sky130_fd_io__gpiov2_ctl_0/sky130_fd_io__com_ctl_hldv2_0/HLD_I_H w_9674_16869# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.118 pd=1.4 as=0.118 ps=1.4 w=0.42 l=0.5
X92 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/NG_PAD_VPMP_H a_231_9686# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.5
X93 a_178_9778# a_1079_9778# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X94 VSWITCH a_1077_11842# a_1024_11940# VSWITCH sky130_fd_pr__pfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=1
X95 VCCD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_7/A a_11131_11430# VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.155 pd=1.37 as=0.14 ps=1.28 w=1 l=0.6
X96 a_2159_13760# VCCD a_2392_13760# VSSA sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X97 a_11523_13190# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_8/A VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X98 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/NG_AMX_VPMP_H a_1225_14186# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.6
X99 VSSA a_231_9686# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/NG_PAD_VPMP_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.5
X100 a_421_13760# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_9/A VSSA VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X101 VCCD ANALOG_EN a_13816_1289# VCCD sky130_fd_pr__pfet_01v8_hvt ad=0.345 pd=2.69 as=0.295 ps=2.59 w=1 l=0.25
X102 a_787_17182# a_229_14828# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X103 VSSD a_10643_12610# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.471 pd=3.65 as=76.3 ps=612 w=0.42 l=0.5
X104 VCCD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_3/Y sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_7/A VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X105 a_7659_11461# a_7539_11435# a_6895_11435# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.185 ps=1.93 w=0.7 l=0.6
X106 VSSD a_3642_14801# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/PG_PAD_VDDIOQ_H_N VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.6
X107 a_2250_17651# a_7173_10183# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
R2 PAD_A_NOESD_H PAD sky130_fd_pr__res_generic_m3 w=12.4 l=0.035
X108 VSSA a_195_17182# w_9674_14653# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.118 pd=1.4 as=0.118 ps=1.4 w=0.42 l=0.5
X109 VDDA a_620_18182# a_184_18182# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=1
X110 a_789_12852# VCCD a_421_13378# VSSA sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X111 a_689_12820# a_1024_11940# VSWITCH VSWITCH sky130_fd_pr__pfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X112 a_14397_2496# a_13816_1289# a_13970_2496# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X113 VSSA sky130_fd_io__gpiov2_ctl_0/sky130_fd_io__com_ctl_hldv2_0/HLD_I_H w_12765_14755# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.118 pd=1.4 as=0.118 ps=1.4 w=0.42 l=0.5
X114 VSSD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_1/Y a_10940_10272# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X115 VSSD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_11/Y a_7370_13247# VSSD sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
X116 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_1/B sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_3/Y a_7625_13629# VSSD sky130_fd_pr__nfet_01v8 ad=0.244 pd=1.42 as=0.101 ps=1.08 w=0.84 l=0.15
X117 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/PG_PAD_VDDIOQ_H_N a_178_9778# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X118 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/PG_PAD_VDDIOQ_H_N a_3642_14801# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X119 a_7621_13247# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_11/Y VCCD VCCD sky130_fd_pr__pfet_01v8_hvt ad=0.176 pd=1.54 as=0.189 ps=1.56 w=1.26 l=0.15
X120 a_7625_13629# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_11/Y VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.101 pd=1.08 as=0.118 ps=1.12 w=0.84 l=0.15
X121 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_7/A sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/PG_PAD_VDDIOQ_H_N a_10705_12172# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.5
X122 a_10643_12610# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_9/A VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.471 ps=3.65 w=0.42 l=0.5
X123 a_14053_2496# VCCD a_14092_2778# VSSD sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.9
X124 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_9/A sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_2/A VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X125 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_8/A sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_2/Y VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X126 VSSD a_6367_11435# a_6314_11461# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.185 ps=1.93 w=0.7 l=0.6
X127 a_7621_13247# a_7370_13247# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_1/B VCCD sky130_fd_pr__pfet_01v8_hvt ad=0.334 pd=3.05 as=0.359 ps=3.09 w=1.26 l=0.15
X128 a_1024_12357# a_2162_14426# VSWITCH VSWITCH sky130_fd_pr__pfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X129 a_14053_2496# a_13760_1103# a_13970_2496# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X130 a_12162_13064# a_334_12102# a_12006_13064# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X131 a_324_14186# a_1225_14186# VSWITCH VSWITCH sky130_fd_pr__pfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X132 VDDA a_497_17084# a_478_17182# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.398 ps=3.53 w=1.5 l=0.5
X133 VSSD a_178_9778# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/PG_PAD_VDDIOQ_H_N VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.6
X134 a_2250_17651# a_7173_10183# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X135 a_10705_12172# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/PG_PAD_VDDIOQ_H_N a_10705_12016# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X136 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/NG_AMX_VPMP_H a_1225_12852# VSWITCH VSWITCH sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X137 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_5/ROUT a_387_12076# VSSIO_Q VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X138 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_5/ROUT a_387_12076# VSSIO_Q VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X139 VSSD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_9/Y a_8871_10272# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X140 a_13970_2496# a_13816_1289# a_14397_2496# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X141 a_10705_11704# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_3/Y VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.471 ps=3.65 w=5 l=0.5
X142 VSSD a_11131_11430# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.471 pd=3.65 as=0 ps=0 w=0.42 l=0.5
X143 VCCD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/PG_PAD_VDDIOQ_H_N a_8300_11461# VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X144 VSSA ENABLE_VSWITCH_H a_342_11805# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.185 ps=1.93 w=0.7 l=0.6
X145 a_421_13378# VCCD a_789_12852# VSSA sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X146 a_14397_2496# a_13816_1289# a_13970_2496# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X147 VSSD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_5/A a_12443_12112# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.471 pd=3.65 as=0.111 ps=1.37 w=0.42 l=0.5
X148 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_5/A sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/PG_PAD_VDDIOQ_H_N a_12897_12172# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.5
X149 VCCD a_6895_11435# a_7015_11461# VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X150 a_8699_10272# VCCD a_9067_10698# VSSD sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X151 a_447_9352# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_8/Y VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X152 a_620_17850# a_184_17734# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=1
X153 VSSD a_7173_10183# a_2250_17651# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.6
X154 a_9877_11799# a_8765_11461# a_8067_11435# VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X155 VSSD a_7173_10183# a_2250_17651# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.6
X156 a_2250_17651# a_7173_10183# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X157 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_4/ROUT a_2250_17651# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=4.2 pd=30.6 as=2.1 ps=15.3 w=15 l=0.5
X158 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/NG_PAD_VPMP_H a_1225_12852# VSWITCH VSWITCH sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X159 VSSD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_9/A a_8699_10272# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X160 VSSD sky130_fd_io__gpiov2_ctl_0/HLD_I_H_N a_13970_2496# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.5
X161 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_4/ROUT a_387_12076# VSSIO_Q VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X162 a_497_17084# a_195_17182# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.5
X163 VSSIO_Q a_387_12076# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_4/ROUT VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X164 a_2080_14827# a_178_9778# a_620_17850# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X165 a_2080_14827# a_1079_9778# a_184_17734# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X166 a_9406_11799# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/NG_PAD_VPMP_H VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X167 a_7173_10183# a_231_9686# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X168 VSSA sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_8/Y a_593_13378# VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X169 a_12897_12172# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/PG_PAD_VDDIOQ_H_N a_12897_12016# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X170 a_620_17850# a_178_9778# a_2080_14827# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X171 a_1072_14186# VCCD a_593_13760# VSSA sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X172 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_5/A a_12443_12112# VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.155 ps=1.37 w=0.42 l=0.5
X173 VDDIO_Q a_3642_14801# a_4110_14801# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.185 ps=1.93 w=0.7 l=0.6
X174 a_12897_11704# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_1/Y VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.471 ps=3.65 w=5 l=0.5
X175 VCCD a_8067_11435# a_6543_11435# VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X176 a_13970_2496# a_13816_1289# a_14397_2496# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X177 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_5/ROUT a_2250_17651# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=2.1 pd=15.3 as=2.1 ps=15.3 w=15 l=0.5
X178 a_447_9352# VCCD a_926_9778# VSSD sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X179 a_497_17084# a_231_9686# a_382_14828# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.5
X180 VDDIO_Q a_2250_17651# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_5/ROUT VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=2.1 pd=15.3 as=2.1 ps=15.3 w=15 l=0.5
X181 VSSD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/PG_PAD_VDDIOQ_H_N a_8473_11461# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X182 VSSD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_8/Y a_447_9352# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X183 VCCD a_6543_11435# a_6367_11435# VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X184 w_9674_16869# a_195_17182# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.118 pd=1.4 as=0.118 ps=1.4 w=0.42 l=0.5
X185 VSSA sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_8/A a_421_13378# VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X186 a_3642_14801# a_282_14802# a_9067_10698# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X187 a_14053_2496# a_13760_1103# a_13970_2496# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X188 VSSA a_1225_12852# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/NG_AMX_VPMP_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.6
X189 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_8/A a_11523_13190# VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.155 ps=1.37 w=0.42 l=0.5
X190 VCCD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_11/Y a_7453_13247# VCCD sky130_fd_pr__pfet_01v8_hvt ad=0.189 pd=1.56 as=0.151 ps=1.5 w=1.26 l=0.15
X191 VSSA sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_0/Y a_2749_13760# VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X192 a_643_9778# a_282_14802# a_178_9778# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X193 a_275_9352# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_8/A VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X194 a_7453_13247# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_3/Y a_7370_13247# VCCD sky130_fd_pr__pfet_01v8_hvt ad=0.151 pd=1.5 as=0.334 ps=3.05 w=1.26 l=0.15
X195 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/NG_PAD_VPMP_H a_1225_14186# VSWITCH VSWITCH sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X196 a_13902_2778# VCCD a_14397_2496# VSSD sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.9
X197 a_195_17182# ENABLE_VDDA_H VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.398 ps=3.53 w=1.5 l=0.5
X198 a_6895_11435# a_7539_11435# VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X199 a_10643_12610# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_9/A VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.155 ps=1.37 w=1 l=0.6
X200 VCCD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/NG_PAD_VPMP_H a_9877_11799# VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X201 VSSA a_1225_14186# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/NG_PAD_VPMP_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.6
X202 a_7173_10183# a_282_14802# a_11173_10272# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X203 w_12765_14755# a_195_17182# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.118 pd=1.4 as=0.118 ps=1.4 w=0.42 l=0.5
X204 a_324_12852# a_689_12820# a_789_12852# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X205 VSSD a_13816_1289# a_13760_1103# VSSD sky130_fd_pr__nfet_01v8 ad=0.263 pd=2.19 as=0.211 ps=2.05 w=0.74 l=0.15
X206 a_787_17182# a_229_14828# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.5
X207 a_184_17734# a_1079_9778# a_2080_14827# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X208 a_6543_11435# a_8067_11435# a_8011_11461# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X209 a_387_12076# a_1024_12357# VSWITCH VSWITCH sky130_fd_pr__pfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.199 ps=2.03 w=0.75 l=2
X210 a_11173_10272# a_282_14802# a_7173_10183# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.398 ps=3.53 w=1.5 l=0.5
X211 a_10406_10767# a_282_14802# a_10350_10272# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.398 ps=3.53 w=1.5 l=0.5
X212 a_789_12852# a_689_12820# a_324_12852# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X213 VSSIO_Q a_387_12076# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_5/ROUT VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X214 VSSA a_497_17084# a_478_17182# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.5
X215 a_926_9778# VCCD a_447_9352# VSSD sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X216 a_7539_11435# a_8300_11461# a_9406_11799# VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X217 a_13970_2496# a_13760_1103# a_14053_2496# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X218 a_11850_13064# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_2/Y VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.471 ps=3.65 w=5 l=0.5
X219 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_5/ROUT a_387_12076# VSSIO_Q VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X220 a_1225_12852# a_689_12820# a_1072_12852# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.398 ps=3.53 w=1.5 l=0.5
X221 VSSD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_8/A a_275_9352# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X222 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_8/A a_2250_17651# a_12162_13064# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.5
X223 VSWITCH ENABLE_VSWITCH_H a_342_11805# VSWITCH sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X224 VSSD a_6543_11435# a_6367_11435# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X225 VCCD a_6367_11435# a_6314_11461# VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X226 VSSD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_5/Y a_10583_10272# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X227 VSWITCH a_324_14186# a_1225_14186# VSWITCH sky130_fd_pr__pfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.185 ps=1.93 w=0.7 l=0.6
X228 VDDA a_620_17850# a_184_17734# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=1
X229 a_9350_10698# a_282_14802# a_4110_14801# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X230 a_1077_11842# a_342_11805# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.5
X231 a_324_12852# a_1225_12852# VSWITCH VSWITCH sky130_fd_pr__pfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X232 VDDIO_Q a_13902_2778# a_231_9686# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.398 ps=3.53 w=1.5 l=0.5
X233 w_12765_14755# a_6367_11435# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_7/ROUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.84 pd=6.56 as=0.84 ps=6.56 w=3 l=0.5
X234 a_9067_10698# a_282_14802# a_3642_14801# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X235 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/NG_AMX_VPMP_H a_1225_14186# VSWITCH VSWITCH sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X236 a_10940_10272# VCCD a_11173_10272# VSSD sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X237 VSSIO_Q a_387_12076# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_5/ROUT VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X238 a_8300_11461# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/PG_AMX_VDDA_H_N VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X239 a_184_17734# a_478_17182# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.5
X240 VSSA a_1225_14186# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/NG_AMX_VPMP_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.6
X241 a_497_17084# a_229_14828# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=1
X242 VSSA a_184_17734# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/PG_AMX_VDDA_H_N VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.5
X243 a_2982_13760# VCCD a_2749_13760# VSSA sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X244 a_789_14186# VCCD a_421_13760# VSSA sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X245 a_7015_11461# a_6895_11435# VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X246 VSWITCH a_1077_11842# a_377_12820# VSWITCH sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.398 ps=3.53 w=1.5 l=0.5
X247 VSSD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/NG_PAD_VPMP_H a_8067_11435# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X248 a_8765_11461# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/PG_AMX_VDDA_H_N VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X249 a_1077_11842# a_231_9686# a_3218_11709# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.5
X250 a_2250_17651# a_7173_10183# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.6
X251 VCCD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_14/Y a_6895_11435# VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X252 a_643_9778# VCCD a_275_9352# VSSD sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X253 VDDIO_Q a_7173_10183# a_2250_17651# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X254 a_324_12852# a_377_12820# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X255 a_14092_2778# VCCD a_14053_2496# VSSD sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.9
X256 VSSD a_8300_11461# a_7539_11435# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.196 pd=1.96 as=0.098 ps=0.98 w=0.7 l=0.6
X257 VSSA a_377_12820# a_324_12852# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.398 ps=3.53 w=1.5 l=0.5
X258 a_184_18182# a_4110_14801# a_3462_14827# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.5
X259 VCCD a_13816_1289# a_13760_1103# VCCD sky130_fd_pr__pfet_01v8_hvt ad=0.345 pd=2.69 as=0.295 ps=2.59 w=1 l=0.25
X260 a_11080_13064# a_6314_11461# a_10924_13064# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X261 a_2162_14426# a_377_12820# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X262 a_10350_10272# a_282_14802# a_10406_10767# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X263 a_13970_2496# sky130_fd_io__gpiov2_ctl_0/HLD_I_H_N VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.5
X264 VCCD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_9/A a_10643_12610# VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X265 VSSA ENABLE_VDDA_H a_382_14828# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.5
X266 a_3462_14827# a_4110_14801# a_184_18182# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X267 a_3642_14801# a_4110_14801# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X268 a_7370_13247# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_3/Y VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.223 ps=2.21 w=0.84 l=0.15
X269 a_4110_14801# a_282_14802# a_9350_10698# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.398 ps=3.53 w=1.5 l=0.5
X270 a_12443_12112# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_5/A VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X271 a_3642_14801# a_231_9686# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X272 VDDIO_Q a_3642_14801# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/PG_PAD_VDDIOQ_H_N VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X273 a_275_9352# VCCD a_643_9778# VSSD sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X274 a_8473_11461# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/PG_AMX_VDDA_H_N a_8300_11461# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.185 ps=1.93 w=0.7 l=0.6
X275 VDDIO_Q a_178_9778# a_1079_9778# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.185 ps=1.93 w=0.7 l=0.6
X276 VSSD a_231_9686# a_3642_14801# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.398 ps=3.53 w=1.5 l=0.5
X277 a_6367_11435# a_6543_11435# VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X278 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_5/A sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_1/Y VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X279 VCCD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_2/Y sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_8/A VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X280 a_10583_10272# VCCD a_10350_10272# VSSD sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X281 VCCD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/PG_PAD_VDDIOQ_H_N a_8300_11461# VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X282 VSSA a_1024_11940# a_689_12820# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.5
X283 a_8938_11461# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/PG_AMX_VDDA_H_N a_8765_11461# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.185 ps=1.93 w=0.7 l=0.6
X284 a_7015_11461# a_6895_11435# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X285 a_421_13760# VCCD a_789_14186# VSSA sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X286 a_1072_14186# a_689_12820# a_1225_14186# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X287 a_3218_11709# a_231_9686# a_1077_11842# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X288 VSSD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_14/Y a_7659_11461# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X289 a_178_9778# a_231_9686# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X290 w_12765_16869# a_7015_11461# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_9/ROUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.84 pd=6.56 as=0.84 ps=6.56 w=3 l=0.5
X291 a_8871_10272# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_9/Y VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X292 VSSD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_7/A a_11131_11430# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.471 pd=3.65 as=0.111 ps=1.37 w=0.42 l=0.5
X293 a_497_17084# a_231_9686# a_382_14828# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X294 VSSD a_7370_13247# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_1/B VSSD sky130_fd_pr__nfet_01v8 ad=0.479 pd=2.82 as=0.244 ps=1.42 w=0.84 l=0.15
X295 a_7367_11461# a_7015_11461# VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X296 VSSD a_231_9686# a_7173_10183# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X297 a_4259_12681# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/NG_PAD_VPMP_H VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.199 ps=2.03 w=0.75 l=0.5
X298 a_184_18182# a_4110_14801# a_3462_14827# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X299 a_382_14828# a_282_14802# a_229_14828# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X300 VSSD a_12443_12112# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.471 pd=3.65 as=0 ps=0 w=0.42 l=0.5
X301 a_593_13378# VCCD a_1072_12852# VSSA sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X302 VSSA sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_9/Y a_593_13760# VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X303 VSSA sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_7/Y a_2392_13760# VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X304 VSSA a_1225_12852# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/NG_PAD_VPMP_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.6
X305 a_2162_14426# a_689_12820# a_2982_13760# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X306 a_8871_10272# VCCD a_9350_10698# VSSD sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X307 a_926_9778# a_282_14802# a_1079_9778# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X308 VDDIO_Q a_178_9778# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/PG_PAD_VDDIOQ_H_N VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X309 VCCD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/PG_PAD_VDDIOQ_H_N a_8765_11461# VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X310 VSSD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_2/A a_11080_13064# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.471 pd=3.65 as=0.7 ps=5.28 w=5 l=0.5
X311 a_12006_13064# a_7367_11461# a_11850_13064# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X312 a_1024_12357# a_689_12820# a_2159_13760# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.398 ps=3.53 w=1.5 l=0.5
X313 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_5/ROUT a_387_12076# VSSIO_Q VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X314 VSSD a_11523_13190# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.111 pd=1.37 as=0 ps=0 w=0.42 l=0.5
X315 a_10705_12016# a_643_12102# a_10705_11860# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X316 a_6543_11435# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_2/Y VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X317 a_3462_14827# a_787_17182# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.5
X318 a_2250_17651# a_7173_10183# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.6
X319 a_2749_13760# VCCD a_2982_13760# VSSA sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X320 VCCD a_8067_11435# a_6543_11435# VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X321 VCCD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_2/A sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_9/A VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X322 a_342_11805# ENABLE_VSWITCH_H VSWITCH VSWITCH sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X323 a_6367_11435# a_6543_11435# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X324 a_387_12076# a_231_9686# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.5
X325 a_13902_2778# a_14092_2778# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.199 ps=2.03 w=0.75 l=0.5
X326 a_593_13378# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_8/Y VSSA VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X327 VSSA sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_9/A a_421_13760# VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X328 VCCD a_6543_11435# a_6367_11435# VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X329 VSWITCH a_324_12852# a_1225_12852# VSWITCH sky130_fd_pr__pfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.185 ps=1.93 w=0.7 l=0.6
X330 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/PG_PAD_VDDIOQ_H_N a_178_9778# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.6
X331 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/PG_PAD_VDDIOQ_H_N a_3642_14801# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.6
X332 a_14397_2496# VCCD a_13902_2778# VSSD sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X333 VDDIO_Q a_7173_10183# a_2250_17651# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X334 VDDIO_Q a_7173_10183# a_2250_17651# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X335 a_13902_2778# sky130_fd_io__gpiov2_ctl_0/sky130_fd_io__com_ctl_hldv2_0/HLD_I_H VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.5
X336 VSWITCH a_1225_12852# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/NG_AMX_VPMP_H VSWITCH sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X337 a_10705_11860# a_4259_12681# a_10705_11704# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X338 a_1077_11842# a_231_9686# a_3218_11709# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X339 a_387_12076# a_1024_12357# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.398 ps=3.53 w=1.5 l=0.5
X340 VSSD a_14092_2778# a_282_14802# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.5
X341 VCCD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_8/A a_11523_13190# VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.155 pd=1.37 as=0.14 ps=1.28 w=1 l=0.6
X342 VSSD sky130_fd_io__gpiov2_ctl_0/HLD_I_H_N a_13970_2496# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.5
X343 VSSD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_8/A a_11523_13190# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.471 pd=3.65 as=0.111 ps=1.37 w=0.42 l=0.5
X344 a_7367_11461# a_7015_11461# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X345 a_421_13378# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_8/A VSSA VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X346 a_13970_2496# sky130_fd_io__gpiov2_ctl_0/HLD_I_H_N VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.5
X347 a_11131_11430# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_7/A VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X348 a_12897_12016# a_643_12102# a_12897_11860# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X349 a_195_17182# ENABLE_VDDA_H VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.5
X350 a_2250_17651# a_7173_10183# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.6
X351 VCCD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/NG_PAD_VPMP_H a_9877_11799# VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X352 VCCD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_3/Y a_7621_13247# VCCD sky130_fd_pr__pfet_01v8_hvt ad=0.479 pd=3.44 as=0.176 ps=1.54 w=1.26 l=0.15
X353 a_382_14828# a_282_14802# a_229_14828# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X354 VSSD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/PG_PAD_VDDIOQ_H_N a_8938_11461# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X355 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_8/ROUT a_7015_11461# w_9674_16869# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.84 pd=6.56 as=0.84 ps=6.56 w=3 l=0.5
X356 VSWITCH a_1225_14186# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/NG_PAD_VPMP_H VSWITCH sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X357 a_3462_14827# a_3642_14801# a_620_18182# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X358 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_7/A sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_3/Y VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X359 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_4/ROUT a_387_12076# VSSIO_Q VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X360 a_8011_11461# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_2/Y VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X361 VDDIO_Q a_10406_10767# a_7173_10183# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.185 ps=1.93 w=0.7 l=0.6
X362 a_620_18182# a_3642_14801# a_3462_14827# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X363 VSSIO_Q a_387_12076# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_4/ROUT VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X364 a_7539_11435# a_8300_11461# a_9406_11799# VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X365 a_282_14802# a_14092_2778# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X366 a_2392_13760# VCCD a_2159_13760# VSSA sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X367 a_12897_11860# a_4259_12681# a_12897_11704# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X368 a_10940_10272# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_1/Y VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X369 VSSA a_1077_11842# a_377_12820# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.5
X370 a_2250_17651# a_7173_10183# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.6
X371 a_4259_12681# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/NG_PAD_VPMP_H VSWITCH VSWITCH sky130_fd_pr__pfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.398 ps=3.53 w=1.5 l=0.5
X372 VDDA a_184_17734# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/PG_AMX_VDDA_H_N VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.5
X373 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_4/ROUT a_2250_17651# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=2.1 pd=15.3 as=2.1 ps=15.3 w=15 l=0.5
X374 a_3218_11709# a_282_14802# a_1024_11940# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X375 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/PG_AMX_VDDA_H_N a_184_17734# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.5
X376 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_4/ROUT a_387_12076# VSSIO_Q VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.4 ps=10.6 w=5 l=0.5
X377 VDDIO_Q a_2250_17651# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_5/ROUT VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=2.1 pd=15.3 as=2.1 ps=15.3 w=15 l=0.5
X378 a_231_9686# a_13902_2778# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.5
X379 a_1024_11940# a_282_14802# a_3218_11709# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X380 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/NG_AMX_VPMP_H a_1225_12852# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.6
X381 a_8300_11461# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/PG_AMX_VDDA_H_N VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X382 a_10583_10272# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_5/Y VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
.ends

.subckt sky130_ef_io__gpiov2_pad DM[0] IB_MODE_SEL ENABLE_H ENABLE_INP_H SLOW VTRIP_SEL
+ ENABLE_VDDIO ENABLE_VDDA_H PAD_A_NOESD_H ANALOG_POL HLD_H_N w_9674_16462# DM[1]
+ w_12765_14348# DM[2] w_9674_14246# PAD_A_ESD_1_H ENABLE_VSWITCH_H TIE_HI_ESD TIE_LO_ESD
+ OE_N w_12765_16462# AMUXBUS_B VSWITCH ANALOG_SEL IN_H VDDIO INP_DIS OUT HLD_OVR
+ VCCD PAD AMUXBUS_A VCCHIB PAD_A_ESD_0_H ANALOG_EN VSSIO VDDA VDDIO_Q VSSIO_Q IN
+ VSSD VSSA
Xsky130_fd_io__top_gpiov2_0 VSSIO_Q PAD_A_NOESD_H ANALOG_POL ENABLE_VDDIO IN_H IN
+ DM[0] DM[1] DM[2] HLD_OVR INP_DIS ENABLE_VDDA_H VTRIP_SEL OE_N OUT SLOW TIE_LO_ESD
+ PAD_A_ESD_0_H ANALOG_SEL ENABLE_INP_H PAD_A_ESD_1_H TIE_HI_ESD ENABLE_H IB_MODE_SEL
+ ENABLE_VSWITCH_H ANALOG_EN sky130_fd_io__top_gpiov2_0/sky130_fd_io__overlay_gpiov2_m4_0/sky130_fd_io__top_gpio_pad_0/b_1500_19531#
+ w_9674_16462# sky130_fd_io__top_gpiov2_0/sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/PG_AMX_VDDA_H_N
+ w_12765_16462# w_12765_14348# w_9674_14246# HLD_H_N VDDIO_Q VSWITCH VSSA VCCHIB
+ VDDIO PAD VDDA AMUXBUS_B VCCD AMUXBUS_A VSSIO VSSD sky130_fd_io__top_gpiov2
.ends

.subckt sky130_ef_io__gpiov2_pad_wrapped IN_H PAD_A_NOESD_H PAD_A_ESD_0_H PAD_A_ESD_1_H
+ DM[2] DM[1] DM[0] IN INP_DIS IB_MODE_SEL ENABLE_H ENABLE_VDDA_H ENABLE_INP_H OE_N
+ TIE_HI_ESD TIE_LO_ESD SLOW VTRIP_SEL HLD_OVR ANALOG_EN ANALOG_SEL ENABLE_VDDIO ENABLE_VSWITCH_H
+ ANALOG_POL OUT VDDIO_Q w_9674_19062# HLD_H_N VSSIO_Q w_12765_19062# VCCD AMUXBUS_B
+ AMUXBUS_A VSSIO VSWITCH VDDA w_12765_16948# VDDIO VSSA w_9674_16846# VSSD PAD VCCHIB
Xgpio DM[0] IB_MODE_SEL ENABLE_H ENABLE_INP_H SLOW VTRIP_SEL ENABLE_VDDIO ENABLE_VDDA_H
+ PAD_A_NOESD_H ANALOG_POL HLD_H_N w_9674_19062# DM[1] w_12765_16948# DM[2] w_9674_16846#
+ PAD_A_ESD_1_H ENABLE_VSWITCH_H TIE_HI_ESD TIE_LO_ESD OE_N w_12765_19062# AMUXBUS_B
+ VSWITCH ANALOG_SEL IN_H VDDIO INP_DIS OUT HLD_OVR VCCD PAD AMUXBUS_A VCCHIB PAD_A_ESD_0_H
+ ANALOG_EN VSSIO VDDA VDDIO_Q VSSIO_Q IN VSSD VSSA sky130_ef_io__gpiov2_pad
.ends

.subckt sky130_fd_sc_hd__buf_16 A VGND VNB VPB VPWR X
X0 VGND A a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 a_109_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VPWR A a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 a_109_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X17 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 VPWR A a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VGND A a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X21 VGND A a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X22 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X23 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X25 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X26 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X27 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X30 a_109_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X31 a_109_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X32 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X33 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X34 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X35 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X36 VPWR A a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X37 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X38 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X39 a_109_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X40 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X41 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X42 a_109_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X43 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
R0 VPWR HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
R1 LO VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
.ends

.subckt constant_block vccd zero one vssd
Xconst_zero_buf const_source/LO vssd vssd vccd vccd zero sky130_fd_sc_hd__buf_16
Xconst_source vssd vssd vccd vccd const_source/HI const_source/LO sky130_fd_sc_hd__conb_1
Xconst_one_buf const_source/HI vssd vssd vccd vccd one sky130_fd_sc_hd__buf_16
.ends

.subckt sky130_fd_io__pad_esd m4_960_20017# m5_1354_20500#
R0 m4_960_20017# m5_1354_20500# sky130_fd_pr__res_generic_m5 w=253 l=0.1
.ends

.subckt sky130_fd_io__com_busses_esd sky130_fd_io__com_bus_hookup_0/VCCHIB sky130_fd_io__pad_esd_0/m5_1354_20500#
+ sky130_fd_io__com_bus_hookup_0/VSSD sky130_fd_io__pad_esd_0/m4_960_20017# sky130_fd_io__com_bus_hookup_0/AMUXBUS_A
+ sky130_fd_io__com_bus_hookup_0/VCCD sky130_fd_io__com_bus_hookup_0/AMUXBUS_B sky130_fd_io__com_bus_hookup_0/VDDIO
+ sky130_fd_io__com_bus_hookup_0/VSSIO sky130_fd_io__com_bus_hookup_0/VSWITCH sky130_fd_io__com_bus_hookup_0/VSSA
+ sky130_fd_io__com_bus_hookup_0/VDDA sky130_fd_io__com_bus_hookup_0/VSSIO_Q sky130_fd_io__com_bus_hookup_0/VDDIO_Q
Xsky130_fd_io__pad_esd_0 sky130_fd_io__pad_esd_0/m4_960_20017# sky130_fd_io__pad_esd_0/m5_1354_20500#
+ sky130_fd_io__pad_esd
.ends

.subckt sky130_fd_io__top_power_lvc_wpad VSSIO_Q VCCHIB VDDA VDDIO_Q P_PAD SRC_BDY_LVC1
+ SRC_BDY_LVC2 BDY2_B2B DRN_LVC2 DRN_LVC1 P_CORE PADISOR PADISOL OGC_LVC AMUXBUS_B
+ VSSIO VDDIO VSSD VSWITCH VCCD AMUXBUS_A VSSA
Xsky130_fd_io__com_busses_esd_0 VCCHIB P_PAD VSSD P_CORE AMUXBUS_A VCCD AMUXBUS_B
+ VDDIO VSSIO VSWITCH VSSA VDDA VSSIO_Q VDDIO_Q sky130_fd_io__com_busses_esd
X0 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X1 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X2 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X3 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.7 pd=5.28 as=687 ps=3.1k w=5 l=8
X4 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X5 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X6 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X7 DRN_LVC1 a_414_306# a_450_404# DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X8 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X9 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X10 a_2872_5340# a_2595_15129# DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X11 SRC_BDY_LVC1 a_414_306# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=1.28k ps=3.48k w=7 l=8
X12 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=5.62 pd=12.2 as=2.92 ps=6.17 w=5 l=0.18
X13 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X14 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X15 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X16 SRC_BDY_LVC2 a_2595_15129# a_2872_5340# SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.4 pd=7.68 as=4.76 ps=15.4 w=7 l=0.18
X17 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X18 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X19 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X20 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.92 pd=6.17 as=5.62 ps=12.2 w=5 l=0.18
X21 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X22 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
R0 a_414_306# DRN_LVC1 sky130_fd_pr__res_generic_po w=0.33 l=1.95k
X23 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X24 a_450_404# a_414_306# DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X25 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X26 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X27 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X28 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X29 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.92 pd=6.17 as=5.62 ps=12.2 w=5 l=0.18
X30 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X31 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X32 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X33 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X34 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X35 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X36 DRN_LVC1 a_414_306# a_450_404# DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X37 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X38 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X39 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.4 pd=7.68 as=0 ps=0 w=7 l=8
X40 DRN_LVC1 a_414_306# a_450_404# DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
R1 a_2183_16816# a_2595_15129# sky130_fd_pr__res_generic_po w=0.33 l=200
X41 SRC_BDY_LVC1 a_414_306# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X42 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X43 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X44 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X45 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=5.62 pd=12.2 as=2.92 ps=6.17 w=5 l=0.18
X46 a_450_404# a_414_306# DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=1.96 ps=14.6 w=7 l=0.18
X47 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X48 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X49 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X50 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.92 pd=6.17 as=5.62 ps=12.2 w=5 l=0.18
X51 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X52 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X53 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
R2 a_1871_4484# a_13955_3836# sky130_fd_pr__res_generic_po w=0.33 l=300
X54 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X55 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X56 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X57 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X58 a_450_404# a_414_306# DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X59 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X60 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X61 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X62 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X63 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X64 DRN_LVC2 a_2595_15129# a_2872_5340# DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X65 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X66 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X67 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X68 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X69 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X70 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X71 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X72 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X73 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X74 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=5.62 pd=12.2 as=2.92 ps=6.17 w=5 l=0.18
X75 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X76 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X77 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X78 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X79 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
D0 SRC_BDY_LVC1 BDY2_B2B sky130_fd_pr__diode_pd2nw_05v5 pj=3.3e+07 area=2.25e+13
X80 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X81 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X82 DRN_LVC2 a_2595_15129# a_2872_5340# DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X83 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X84 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X85 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X86 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.7 pd=5.28 as=0 ps=0 w=5 l=8
X87 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
D1 BDY2_B2B SRC_BDY_LVC1 sky130_fd_pr__diode_pd2nw_05v5 pj=3.3e+07 area=2.25e+13
X88 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X89 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X90 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X91 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X92 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X93 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X94 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X95 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X96 SRC_BDY_LVC1 a_414_306# a_450_404# SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.4 pd=7.68 as=4.76 ps=15.4 w=7 l=0.18
X97 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X98 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X99 SRC_BDY_LVC1 a_414_306# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.4 pd=7.68 as=0 ps=0 w=7 l=8
X100 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X101 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.92 pd=6.17 as=5.62 ps=12.2 w=5 l=0.18
X102 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X103 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X104 DRN_LVC2 a_2595_15129# a_2872_5340# DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X105 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X106 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X107 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X108 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X109 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X110 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X111 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X112 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X113 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X114 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X115 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X116 a_2872_5340# a_2595_15129# DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X117 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X118 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X119 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X120 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X121 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X122 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X123 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X124 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X125 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X126 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X127 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X128 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X129 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.92 pd=6.17 as=5.62 ps=12.2 w=5 l=0.18
X130 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X131 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X132 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X133 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X134 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X135 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X136 SRC_BDY_LVC1 a_414_306# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.4 pd=7.68 as=0 ps=0 w=7 l=8
X137 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X138 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X139 a_2872_5340# a_2595_15129# DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=1.96 ps=14.6 w=7 l=0.18
X140 SRC_BDY_LVC1 a_414_306# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X141 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X142 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X143 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X144 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X145 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X146 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=5.62 pd=12.2 as=2.92 ps=6.17 w=5 l=0.18
X147 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X148 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X149 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X150 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X151 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X152 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X153 SRC_BDY_LVC1 a_414_306# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X154 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X155 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X156 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X157 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X158 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
D2 BDY2_B2B SRC_BDY_LVC1 sky130_fd_pr__diode_pd2nw_05v5 pj=3.3e+07 area=2.25e+13
X159 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X160 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X161 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X162 DRN_LVC1 a_414_306# a_450_404# DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X163 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X164 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X165 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X166 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X167 DRN_LVC2 a_2595_15129# a_2872_5340# DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X168 SRC_BDY_LVC1 a_414_306# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X169 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X170 a_450_404# a_414_306# DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X171 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X172 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X173 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X174 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X175 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X176 DRN_LVC1 a_414_306# a_450_404# DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X177 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X178 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X179 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X180 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X181 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X182 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X183 SRC_BDY_LVC1 a_414_306# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X184 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X185 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X186 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X187 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X188 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X189 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X190 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X191 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X192 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X193 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X194 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X195 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X196 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
D3 BDY2_B2B SRC_BDY_LVC1 sky130_fd_pr__diode_pd2nw_05v5 pj=3.3e+07 area=2.25e+13
X197 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X198 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X199 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X200 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X201 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X202 DRN_LVC1 a_414_306# a_450_404# DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X203 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X204 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X205 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.7 pd=5.28 as=0 ps=0 w=5 l=8
X206 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X207 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X208 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.92 pd=6.17 as=5.62 ps=12.2 w=5 l=0.18
X209 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X210 DRN_LVC1 a_414_306# a_450_404# DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=1.96 pd=14.6 as=0.98 ps=7.28 w=7 l=0.18
X211 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
R3 DRN_LVC2 a_13955_3836# sky130_fd_pr__res_generic_po w=0.33 l=900
X212 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X213 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X214 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
R4 a_1871_4484# a_2183_16816# sky130_fd_pr__res_generic_po w=0.33 l=720
X215 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X216 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X217 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X218 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X219 SRC_BDY_LVC1 a_414_306# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X220 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X221 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X222 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X223 a_2872_5340# a_2595_15129# DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X224 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X225 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X226 a_2872_5340# a_2595_15129# DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X227 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X228 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X229 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X230 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X231 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X232 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X233 a_450_404# a_414_306# DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X234 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X235 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X236 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.92 pd=6.17 as=5.62 ps=12.2 w=5 l=0.18
X237 a_450_404# a_414_306# DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X238 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X239 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X240 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X241 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X242 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X243 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X244 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X245 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X246 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X247 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X248 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X249 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X250 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X251 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X252 DRN_LVC2 a_2595_15129# a_2872_5340# DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=1.96 pd=14.6 as=0.98 ps=7.28 w=7 l=0.18
X253 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X254 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X255 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X256 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X257 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=5.62 pd=12.2 as=2.92 ps=6.17 w=5 l=0.18
X258 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X259 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X260 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X261 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X262 a_2872_5340# a_2595_15129# DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X263 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X264 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
D4 SRC_BDY_LVC1 BDY2_B2B sky130_fd_pr__diode_pd2nw_05v5 pj=3.3e+07 area=2.25e+13
X265 SRC_BDY_LVC2 a_2595_15129# a_2872_5340# SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.4 pd=7.68 as=4.76 ps=15.4 w=7 l=0.18
X266 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X267 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X268 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X269 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X270 SRC_BDY_LVC1 a_414_306# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X271 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X272 DRN_LVC2 a_2595_15129# a_2872_5340# DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X273 a_450_404# a_414_306# DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X274 DRN_LVC2 a_2595_15129# a_2872_5340# DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X275 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X276 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.4 pd=7.68 as=0 ps=0 w=7 l=8
X277 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=5.62 pd=12.2 as=2.92 ps=6.17 w=5 l=0.18
X278 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X279 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X280 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X281 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X282 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X283 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X284 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X285 DRN_LVC2 a_2595_15129# a_2872_5340# DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X286 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X287 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X288 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X289 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X290 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X291 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X292 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X293 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X294 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X295 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X296 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X297 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X298 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X299 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X300 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X301 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X302 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X303 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X304 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X305 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
D5 SRC_BDY_LVC1 BDY2_B2B sky130_fd_pr__diode_pd2nw_05v5 pj=3.3e+07 area=2.25e+13
X306 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.7 pd=5.28 as=0 ps=0 w=5 l=8
X307 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X308 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=5.62 pd=12.2 as=2.92 ps=6.17 w=5 l=0.18
X309 DRN_LVC1 a_414_306# a_450_404# DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=1.96 pd=14.6 as=0.98 ps=7.28 w=7 l=0.18
X310 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X311 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X312 SRC_BDY_LVC1 a_414_306# a_450_404# SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.4 pd=7.68 as=4.76 ps=15.4 w=7 l=0.18
X313 a_2872_5340# a_2595_15129# DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=1.96 ps=14.6 w=7 l=0.18
X314 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X315 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X316 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X317 a_450_404# a_414_306# DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X318 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X319 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.92 pd=6.17 as=5.62 ps=12.2 w=5 l=0.18
X320 DRN_LVC2 a_2595_15129# a_2872_5340# DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=1.96 pd=14.6 as=0.98 ps=7.28 w=7 l=0.18
X321 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X322 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X323 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X324 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X325 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X326 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X327 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X328 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X329 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X330 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X331 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X332 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X333 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X334 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X335 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=5.62 pd=12.2 as=2.92 ps=6.17 w=5 l=0.18
X336 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X337 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X338 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X339 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
D6 SRC_BDY_LVC1 BDY2_B2B sky130_fd_pr__diode_pd2nw_05v5 pj=3.3e+07 area=2.25e+13
X340 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X341 SRC_BDY_LVC1 a_414_306# a_450_404# SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.4 pd=7.68 as=4.76 ps=15.4 w=7 l=0.18
X342 SRC_BDY_LVC1 a_414_306# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.4 pd=7.68 as=0 ps=0 w=7 l=8
X343 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X344 DRN_LVC1 a_414_306# a_450_404# DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X345 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X346 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X347 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X348 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X349 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X350 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
R5 P_CORE PADISOL sky130_fd_pr__res_generic_m3 w=12.2 l=10m
X351 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X352 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X353 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X354 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X355 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X356 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X357 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X358 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X359 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X360 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X361 a_450_404# a_414_306# DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=1.96 ps=14.6 w=7 l=0.18
X362 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X363 SRC_BDY_LVC1 a_414_306# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X364 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X365 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X366 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X367 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X368 SRC_BDY_LVC1 a_414_306# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X369 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X370 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X371 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X372 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=5.62 pd=12.2 as=2.92 ps=6.17 w=5 l=0.18
X373 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X374 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X375 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X376 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X377 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.7 pd=5.28 as=0 ps=0 w=5 l=8
X378 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X379 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X380 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X381 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X382 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X383 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X384 SRC_BDY_LVC1 a_414_306# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X385 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X386 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X387 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X388 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X389 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X390 a_2872_5340# a_2595_15129# DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X391 a_2872_5340# a_2595_15129# DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X392 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X393 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X394 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X395 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=5.62 pd=12.2 as=2.92 ps=6.17 w=5 l=0.18
X396 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
D7 BDY2_B2B SRC_BDY_LVC1 sky130_fd_pr__diode_pd2nw_05v5 pj=3.3e+07 area=2.25e+13
X397 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X398 a_450_404# a_414_306# DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X399 a_2872_5340# a_2595_15129# DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X400 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X401 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X402 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X403 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X404 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X405 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X406 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X407 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X408 SRC_BDY_LVC1 a_414_306# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X409 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X410 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X411 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X412 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X413 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.7 pd=5.28 as=0 ps=0 w=5 l=8
X414 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X415 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X416 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X417 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X418 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X419 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X420 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X421 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X422 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X423 DRN_LVC1 a_414_306# a_450_404# DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X424 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X425 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X426 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X427 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X428 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X429 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X430 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X431 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=1.33 pd=10.5 as=0 ps=0 w=5 l=4
X432 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X433 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X434 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X435 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.92 pd=6.17 as=5.62 ps=12.2 w=5 l=0.18
X436 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X437 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X438 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
R6 P_CORE PADISOR sky130_fd_pr__res_generic_m3 w=12.2 l=10m
X439 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X440 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X441 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X442 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.92 pd=6.17 as=5.62 ps=12.2 w=5 l=0.18
X443 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X444 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X445 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X446 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X447 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X448 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X449 DRN_LVC2 a_2595_15129# a_2872_5340# DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X450 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X451 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X452 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
.ends

.subckt sky130_ef_io__vccd_lvc_clamped_pad VDDA VCCHIB AMUXBUS_B AMUXBUS_A VCCD_PAD
+ VCCD VDDIO VSSD VSSIO VDDIO_Q VSWITCH VSSA VSSIO_Q
Xsky130_fd_io__top_power_lvc_wpad_0 VSSIO_Q VCCHIB VDDA VDDIO_Q VCCD_PAD VSSIO VSSD
+ VSSA VCCD VCCD VCCD sky130_fd_io__top_power_lvc_wpad_0/PADISOR sky130_fd_io__top_power_lvc_wpad_0/PADISOL
+ VSSA AMUXBUS_B VSSIO VDDIO VSSD VSWITCH VCCD AMUXBUS_A VSSA sky130_fd_io__top_power_lvc_wpad
.ends

.subckt sky130_fd_pr__cap_mim_m3_2_W5U4AW c2_n3079_n3000# m4_n3179_n3100#
X0 c2_n3079_n3000# m4_n3179_n3100# sky130_fd_pr__cap_mim_m3_2 l=30 w=30
.ends

.subckt sky130_fd_sc_hvl__buf_8 A VGND VNB VPB VPWR X
X0 X a_45_443# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X1 VGND a_45_443# X VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X2 X a_45_443# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X3 a_45_443# A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.203 ps=1.29 w=0.75 l=0.5
X4 X a_45_443# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X5 VPWR a_45_443# X VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X6 VGND A a_45_443# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.203 pd=1.29 as=0.214 ps=2.07 w=0.75 l=0.5
X7 X a_45_443# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X8 VPWR A a_45_443# VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X9 VPWR A a_45_443# VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=2.06 as=0.428 ps=3.57 w=1.5 l=0.5
X10 VPWR a_45_443# X VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X11 X a_45_443# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X12 VGND a_45_443# X VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X13 VPWR a_45_443# X VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X14 X a_45_443# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X15 VGND A a_45_443# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X16 VGND a_45_443# X VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.214 pd=2.07 as=0.105 ps=1.03 w=0.75 l=0.5
X17 X a_45_443# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X18 VGND a_45_443# X VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X19 X a_45_443# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X20 VPWR a_45_443# X VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X21 a_45_443# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.42 ps=2.06 w=1.5 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_ZEUEFZ a_n683_n200# a_n189_n297# a_29_n297# a_189_n200#
+ a_n901_n200# a_247_n297# a_n407_n297# a_465_n297# a_407_n200# a_n625_n297# a_683_n297#
+ a_625_n200# a_n843_n297# w_n1101_n497# a_843_n200# a_n29_n200# a_n247_n200# a_n465_n200#
X0 a_n247_n200# a_n407_n297# a_n465_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X1 a_843_n200# a_683_n297# a_625_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.8
X2 a_407_n200# a_247_n297# a_189_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X3 a_189_n200# a_29_n297# a_n29_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X4 a_n465_n200# a_n625_n297# a_n683_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X5 a_625_n200# a_465_n297# a_407_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X6 a_n29_n200# a_n189_n297# a_n247_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X7 a_n683_n200# a_n843_n297# a_n901_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.8
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_TGFUGS a_n792_n200# a_298_n200# a_516_n200# a_734_n200#
+ a_n926_n422# a_138_n288# a_n298_n288# a_80_n200# a_356_n288# a_n516_n288# a_574_n288#
+ a_n734_n288# a_n138_n200# a_n356_n200# a_n574_n200# a_n80_n288#
X0 a_80_n200# a_n80_n288# a_n138_n200# a_n926_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X1 a_n574_n200# a_n734_n288# a_n792_n200# a_n926_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.8
X2 a_734_n200# a_574_n288# a_516_n200# a_n926_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.8
X3 a_298_n200# a_138_n288# a_80_n200# a_n926_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X4 a_n138_n200# a_n298_n288# a_n356_n200# a_n926_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X5 a_n356_n200# a_n516_n288# a_n574_n200# a_n926_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X6 a_516_n200# a_356_n288# a_298_n200# a_n926_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p69_S5N9F3 a_n1806_2500# a_n4122_n2932# a_n5280_2500#
+ a_2054_n2932# a_896_n2932# a_4756_2500# a_3598_n2932# a_3212_2500# a_n3736_n2932#
+ a_1668_n2932# a_n1806_n2932# a_5142_n2932# a_896_2500# a_510_n2932# a_n3350_2500#
+ a_n4508_2500# a_3212_n2932# a_n4894_2500# a_n5410_n3062# a_1282_2500# a_4756_n2932#
+ a_2826_2500# a_2826_n2932# a_n2192_n2932# a_n1034_2500# a_n2578_2500# a_n1420_2500#
+ a_n2964_2500# a_n648_n2932# a_n648_2500# a_n5280_n2932# a_n3350_n2932# a_4370_2500#
+ a_1282_n2932# a_124_n2932# a_n1420_n2932# a_n4894_n2932# a_124_2500# a_n2964_n2932#
+ a_n4122_2500# a_2054_2500# a_510_2500# a_n4508_n2932# a_4370_n2932# a_3598_2500#
+ a_3984_2500# a_2440_n2932# a_2440_2500# a_3984_n2932# a_n2192_2500# a_n3736_2500#
+ a_1668_2500# a_n262_n2932# a_n262_2500# a_n1034_n2932# a_5142_2500# a_n2578_n2932#
X0 a_n2578_2500# a_n2578_n2932# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25
X1 a_n1420_2500# a_n1420_n2932# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25
X2 a_n1806_2500# a_n1806_n2932# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25
X3 a_3212_2500# a_3212_n2932# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25
X4 a_3598_2500# a_3598_n2932# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25
X5 a_n2964_2500# a_n2964_n2932# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25
X6 a_2826_2500# a_2826_n2932# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25
X7 a_4370_2500# a_4370_n2932# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25
X8 a_3984_2500# a_3984_n2932# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25
X9 a_n262_2500# a_n262_n2932# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25
X10 a_n3350_2500# a_n3350_n2932# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25
X11 a_n4122_2500# a_n4122_n2932# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25
X12 a_n3736_2500# a_n3736_n2932# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25
X13 a_5142_2500# a_5142_n2932# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25
X14 a_n4894_2500# a_n4894_n2932# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25
X15 a_1282_2500# a_1282_n2932# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25
X16 a_4756_2500# a_4756_n2932# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25
X17 a_124_2500# a_124_n2932# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25
X18 a_510_2500# a_510_n2932# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25
X19 a_896_2500# a_896_n2932# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25
X20 a_n648_2500# a_n648_n2932# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25
X21 a_n5280_2500# a_n5280_n2932# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25
X22 a_n4508_2500# a_n4508_n2932# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25
X23 a_n1034_2500# a_n1034_n2932# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25
X24 a_n2192_2500# a_n2192_n2932# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25
X25 a_2054_2500# a_2054_n2932# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25
X26 a_1668_2500# a_1668_n2932# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25
X27 a_2440_2500# a_2440_n2932# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_3YBPVB a_n80_n297# a_80_n200# w_n338_n497# a_n138_n200#
X0 a_80_n200# a_n80_n297# a_n138_n200# w_n338_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.8
.ends

.subckt sky130_fd_sc_hvl__schmittbuf_1 A VGND VNB VPB VPWR X
X0 X a_117_181# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.316 ps=1.45 w=0.75 l=0.5
X1 a_217_207# a_117_181# a_64_207# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.111 ps=1.37 w=0.42 l=0.5
X2 VPWR A a_231_463# VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.341 pd=1.73 as=0.105 ps=1.03 w=0.75 l=0.5
X3 VGND A a_217_207# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.316 pd=1.45 as=0.0588 ps=0.7 w=0.42 l=0.5
X4 a_78_463# VGND VNB sky130_fd_pr__res_generic_nd__hv w=0.29 l=1.36
X5 a_64_207# VPWR VPB sky130_fd_pr__res_generic_pd__hv w=0.29 l=3.11
X6 X a_117_181# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.341 ps=1.73 w=1.5 l=0.5
X7 a_231_463# A a_117_181# VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.199 ps=2.03 w=0.75 l=0.5
X8 a_231_463# a_117_181# a_78_463# VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.199 ps=2.03 w=0.75 l=0.5
X9 a_217_207# A a_117_181# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_PKVMTM a_80_n200# a_n272_n422# a_n138_n200# a_n80_n288#
X0 a_80_n200# a_n80_n288# a_n138_n200# a_n272_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.8
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_YUHPXE a_n80_n297# a_80_n200# w_n338_n497# a_n138_n200#
X0 a_80_n200# a_n80_n297# a_n138_n200# w_n338_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.8
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_ZK8HQC a_80_n200# a_n272_n422# a_n138_n200# a_n80_n288#
X0 a_80_n200# a_n80_n288# a_n138_n200# a_n272_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.8
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_WRT4AW c1_n3036_n3000# m3_n3136_n3100#
X0 c1_n3036_n3000# m3_n3136_n3100# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_YEUEBV a_n792_n200# a_138_n297# a_n298_n297#
+ a_298_n200# a_356_n297# a_n516_n297# a_574_n297# a_516_n200# a_n734_n297# a_734_n200#
+ a_n80_n297# a_80_n200# a_n138_n200# a_n356_n200# a_n574_n200# w_n992_n497#
X0 a_80_n200# a_n80_n297# a_n138_n200# w_n992_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X1 a_n574_n200# a_n734_n297# a_n792_n200# w_n992_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.8
X2 a_734_n200# a_574_n297# a_516_n200# w_n992_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.8
X3 a_298_n200# a_138_n297# a_80_n200# w_n992_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X4 a_n138_n200# a_n298_n297# a_n356_n200# w_n992_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X5 a_n356_n200# a_n516_n297# a_n574_n200# w_n992_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X6 a_516_n200# a_356_n297# a_298_n200# w_n992_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_YUHPBG a_n80_n297# a_80_n200# w_n338_n497# a_n138_n200#
X0 a_80_n200# a_n80_n297# a_n138_n200# w_n338_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.8
.ends

.subckt sky130_fd_sc_hvl__inv_8 A VGND VNB VPB VPWR Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X2 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.157 pd=1.17 as=0.105 ps=1.03 w=0.75 l=0.5
X3 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X4 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.206 pd=2.05 as=0.105 ps=1.03 w=0.75 l=0.5
X5 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X6 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X7 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X8 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X9 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.157 ps=1.17 w=0.75 l=0.5
X10 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X11 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.398 ps=3.53 w=1.5 l=0.5
X12 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X13 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X14 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X15 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.199 ps=2.03 w=0.75 l=0.5
.ends

.subckt simple_por vdd3v3 vdd1v8 porb_h por_l porb_l vss1v8 vss3v3
Xsky130_fd_pr__cap_mim_m3_2_W5U4AW_0 vss3v3 sky130_fd_sc_hvl__schmittbuf_1_0/A sky130_fd_pr__cap_mim_m3_2_W5U4AW
Xsky130_fd_sc_hvl__buf_8_1 sky130_fd_sc_hvl__inv_8_0/A vss1v8 vss1v8 vdd1v8 vdd1v8
+ porb_l sky130_fd_sc_hvl__buf_8
Xsky130_fd_pr__pfet_g5v0d10v5_ZEUEFZ_0 m1_502_7653# m1_502_7653# m1_502_7653# m1_502_7653#
+ vdd3v3 m1_502_7653# m1_502_7653# m1_502_7653# vdd3v3 m1_502_7653# m1_502_7653# m1_502_7653#
+ m1_502_7653# vdd3v3 vdd3v3 vdd3v3 m1_502_7653# vdd3v3 sky130_fd_pr__pfet_g5v0d10v5_ZEUEFZ
Xsky130_fd_pr__nfet_g5v0d10v5_TGFUGS_0 m1_721_6815# vss3v3 m1_721_6815# vss3v3 vss3v3
+ m1_721_6815# m1_721_6815# m1_721_6815# m1_721_6815# m1_721_6815# m1_721_6815# m1_721_6815#
+ vss3v3 m1_721_6815# vss3v3 m1_721_6815# sky130_fd_pr__nfet_g5v0d10v5_TGFUGS
Xsky130_fd_pr__res_xhigh_po_0p69_S5N9F3_0 li_3322_5813# li_1391_165# vss3v3 li_7567_165#
+ li_6023_165# vdd3v3 li_9111_165# li_8726_5813# li_1391_165# li_6795_165# li_3707_165#
+ vss3v3 li_6410_5813# li_6023_165# li_1778_5813# li_1006_5813# li_8339_165# vss3v3
+ vss3v3 li_6410_5813# li_9883_165# li_7954_5813# li_8339_165# li_2935_165# li_4094_5813#
+ li_2550_5813# li_4094_5813# li_2550_5813# li_4479_165# li_4866_5813# vss3v3 li_2163_165#
+ li_9498_5813# li_6795_165# li_5251_165# li_3707_165# li_619_165# li_5638_5813# li_2163_165#
+ li_1006_5813# li_7182_5813# li_5638_5813# li_619_165# li_9883_165# li_8726_5813#
+ li_9498_5813# li_7567_165# li_7954_5813# li_9111_165# li_3322_5813# li_1778_5813#
+ li_7182_5813# li_5251_165# li_4866_5813# li_4479_165# vss3v3 li_2935_165# sky130_fd_pr__res_xhigh_po_0p69_S5N9F3
Xsky130_fd_pr__pfet_g5v0d10v5_3YBPVB_0 m1_185_6573# m1_721_6815# vdd3v3 m1_2993_7658#
+ sky130_fd_pr__pfet_g5v0d10v5_3YBPVB
Xsky130_fd_pr__pfet_g5v0d10v5_3YBPVB_1 m1_2756_6573# m1_4283_8081# vdd3v3 m1_2756_6573#
+ sky130_fd_pr__pfet_g5v0d10v5_3YBPVB
Xsky130_fd_sc_hvl__schmittbuf_1_0 sky130_fd_sc_hvl__schmittbuf_1_0/A vss3v3 vss3v3
+ vdd3v3 vdd3v3 sky130_fd_sc_hvl__inv_8_0/A sky130_fd_sc_hvl__schmittbuf_1
Xsky130_fd_pr__pfet_g5v0d10v5_3YBPVB_2 m1_2756_6573# sky130_fd_sc_hvl__schmittbuf_1_0/A
+ vdd3v3 m1_6249_7690# sky130_fd_pr__pfet_g5v0d10v5_3YBPVB
Xsky130_fd_pr__pfet_g5v0d10v5_3YBPVB_3 m1_185_6573# m1_502_7653# vdd3v3 m1_185_6573#
+ sky130_fd_pr__pfet_g5v0d10v5_3YBPVB
Xsky130_fd_pr__nfet_g5v0d10v5_PKVMTM_0 m1_2756_6573# vss3v3 vss3v3 m1_721_6815# sky130_fd_pr__nfet_g5v0d10v5_PKVMTM
Xsky130_fd_pr__pfet_g5v0d10v5_YUHPXE_0 m1_4283_8081# m1_6249_7690# vdd3v3 vdd3v3 sky130_fd_pr__pfet_g5v0d10v5_YUHPXE
Xsky130_fd_pr__nfet_g5v0d10v5_ZK8HQC_1 m1_185_6573# vss3v3 vss3v3 li_2550_5813# sky130_fd_pr__nfet_g5v0d10v5_ZK8HQC
Xsky130_fd_pr__cap_mim_m3_1_WRT4AW_0 sky130_fd_sc_hvl__schmittbuf_1_0/A vss3v3 sky130_fd_pr__cap_mim_m3_1_WRT4AW
Xsky130_fd_pr__pfet_g5v0d10v5_YEUEBV_0 vdd3v3 m1_4283_8081# m1_4283_8081# m1_4283_8081#
+ m1_4283_8081# m1_4283_8081# m1_4283_8081# vdd3v3 m1_4283_8081# m1_4283_8081# m1_4283_8081#
+ vdd3v3 m1_4283_8081# vdd3v3 m1_4283_8081# vdd3v3 sky130_fd_pr__pfet_g5v0d10v5_YEUEBV
Xsky130_fd_pr__pfet_g5v0d10v5_YUHPBG_0 m1_502_7653# m1_2993_7658# vdd3v3 vdd3v3 sky130_fd_pr__pfet_g5v0d10v5_YUHPBG
Xsky130_fd_sc_hvl__buf_8_0 sky130_fd_sc_hvl__inv_8_0/A vss3v3 vss3v3 vdd3v3 vdd3v3
+ porb_h sky130_fd_sc_hvl__buf_8
Xsky130_fd_sc_hvl__inv_8_0 sky130_fd_sc_hvl__inv_8_0/A vss1v8 vss1v8 vdd1v8 vdd1v8
+ por_l sky130_fd_sc_hvl__inv_8
.ends

.subckt sky130_fd_io__sio_clamp_pcap_4x5 a_36_36# a_229_118#
X0 a_36_36# a_229_118# a_36_36# a_36_36# sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=10.5 as=2.65 ps=21.1 w=5 l=4
.ends

.subckt sky130_fd_io__esd_rcclamp_nfetcap a_179_100# a_n14_18#
X0 a_n14_18# a_179_100# a_n14_18# a_n14_18# sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=10.5 as=2.65 ps=21.1 w=5 l=8
.ends

.subckt sky130_fd_io__hvc_clampv2 m2_5179_0# w_1040_5785# sky130_fd_io__com_busses_esd_0/sky130_fd_io__pad_esd_0/m5_1354_20500#
+ m3_10082_12712# m3_103_12712# sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDIO_Q
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/AMUXBUS_B sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSIO_Q
+ w_2676_441# sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDIO
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VCCHIB sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSIO
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDA sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSD
+ m3_99_0# sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSWITCH sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VCCD
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/AMUXBUS_A sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSA
Xsky130_fd_io__sio_clamp_pcap_4x5_0[0] w_2676_441# a_1268_5934# sky130_fd_io__sio_clamp_pcap_4x5
Xsky130_fd_io__sio_clamp_pcap_4x5_0[1] w_2676_441# a_1268_5934# sky130_fd_io__sio_clamp_pcap_4x5
Xsky130_fd_io__sio_clamp_pcap_4x5_0[2] w_2676_441# a_1268_5934# sky130_fd_io__sio_clamp_pcap_4x5
Xsky130_fd_io__com_busses_esd_0 sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VCCHIB
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__pad_esd_0/m5_1354_20500# sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSD
+ m3_99_0# sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/AMUXBUS_A
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VCCD sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/AMUXBUS_B
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDIO sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSIO
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSWITCH sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSA
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDA sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSIO_Q
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDIO_Q sky130_fd_io__com_busses_esd
Xsky130_fd_io__sio_clamp_pcap_4x5_1 w_2676_441# a_1268_5934# sky130_fd_io__sio_clamp_pcap_4x5
Xsky130_fd_io__esd_rcclamp_nfetcap_0[0|0] a_1268_5934# w_2676_441# sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[1|0] a_1268_5934# w_2676_441# sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[2|0] a_1268_5934# w_2676_441# sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[0|1] a_1268_5934# w_2676_441# sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[1|1] a_1268_5934# w_2676_441# sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[2|1] a_1268_5934# w_2676_441# sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[0|2] a_1268_5934# w_2676_441# sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[1|2] a_1268_5934# w_2676_441# sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[2|2] a_1268_5934# w_2676_441# sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[0|3] a_1268_5934# w_2676_441# sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[1|3] a_1268_5934# w_2676_441# sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[2|3] a_1268_5934# w_2676_441# sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[0|4] a_1268_5934# w_2676_441# sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[1|4] a_1268_5934# w_2676_441# sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[2|4] a_1268_5934# w_2676_441# sky130_fd_io__esd_rcclamp_nfetcap
X0 a_1368_5960# a_1268_5934# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=1.86 pd=14.5 as=0.98 ps=7.28 w=7 l=0.5
X1 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X2 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X3 w_2676_441# a_1268_5934# a_1368_5960# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X4 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X5 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.4 as=7.55 ps=11.5 w=10 l=0.5
X6 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X7 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X8 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X9 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.4 as=7.55 ps=11.5 w=10 l=0.5
X10 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.86 ps=14.5 w=7 l=0.5
X11 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X12 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X13 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X14 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X15 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X16 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X17 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X18 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X19 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X20 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X21 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X22 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X23 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X24 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.5 as=6.95 ps=21.4 w=10 l=0.5
X25 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X26 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X27 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X28 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.5 as=6.95 ps=21.4 w=10 l=0.5
X29 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X30 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X31 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.4 as=7.55 ps=11.5 w=10 l=0.5
X32 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X33 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X34 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X35 a_1368_5960# a_1268_5934# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X36 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X37 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.4 as=7.55 ps=11.5 w=10 l=0.5
X38 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.5 as=6.95 ps=21.4 w=10 l=0.5
X39 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X40 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X41 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X42 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X43 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X44 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X45 a_1368_5960# a_1268_5934# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X46 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X47 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X48 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X49 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X50 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X51 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X52 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X53 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X54 w_2676_441# a_1268_5934# a_1368_5960# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X55 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X56 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X57 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.5 as=6.95 ps=21.4 w=10 l=0.5
X58 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X59 a_1368_5960# a_1268_5934# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X60 w_2676_441# a_1268_5934# a_1368_5960# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X61 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X62 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X63 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X64 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X65 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X66 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X67 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.4 as=7.55 ps=11.5 w=10 l=0.5
X68 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X69 w_2676_441# a_1268_5934# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=10.5 as=74.2 ps=498 w=5 l=4
X70 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.5 as=6.95 ps=21.4 w=10 l=0.5
X71 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X72 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X73 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X74 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X75 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X76 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X77 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.4 as=7.55 ps=11.5 w=10 l=0.5
X78 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X79 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X80 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X81 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
R0 a_1268_5934# a_1672_8570# sky130_fd_pr__res_generic_po w=0.33 l=470
X82 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X83 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X84 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X85 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X86 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X87 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X88 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X89 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X90 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X91 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X92 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.4 as=7.55 ps=11.5 w=10 l=0.5
X93 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X94 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X95 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X96 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X97 w_2676_441# a_1268_5934# a_1368_5960# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X98 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X99 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X100 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X101 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X102 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X103 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X104 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X105 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.5 as=6.95 ps=21.4 w=10 l=0.5
X106 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X107 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X108 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X109 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X110 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X111 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X112 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X113 w_2676_441# a_1268_5934# a_1368_5960# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X114 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X115 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X116 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X117 a_1368_5960# a_1268_5934# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X118 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X119 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.5 as=6.95 ps=21.4 w=10 l=0.5
X120 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X121 w_2676_441# a_1268_5934# a_1368_5960# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X122 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X123 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X124 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X125 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X126 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X127 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.4 as=7.55 ps=11.5 w=10 l=0.5
R1 m3_99_0# m3_103_12712# sky130_fd_pr__res_generic_m3 w=12.1 l=10m
X128 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.4 as=7.55 ps=11.5 w=10 l=0.5
X129 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X130 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X131 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X132 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
R2 w_1040_5785# a_214_8570# sky130_fd_pr__res_generic_po w=0.33 l=700
X133 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X134 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X135 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X136 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X137 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X138 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X139 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X140 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X141 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X142 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X143 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X144 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X145 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X146 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X147 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.5 as=6.95 ps=21.4 w=10 l=0.5
X148 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X149 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X150 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X151 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=1.86 pd=14.5 as=0.98 ps=7.28 w=7 l=0.5
R3 a_1672_8570# a_214_8570# sky130_fd_pr__res_generic_po w=0.33 l=1.55k
X152 a_1368_5960# a_1268_5934# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X153 w_2676_441# a_1268_5934# a_1368_5960# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X154 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X155 a_1368_5960# a_1268_5934# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.86 ps=14.5 w=7 l=0.5
X156 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X157 a_1368_5960# a_1268_5934# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X158 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X159 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X160 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X161 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X162 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X163 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X164 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X165 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X166 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X167 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X168 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X169 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X170 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
R4 m3_99_0# m3_10082_12712# sky130_fd_pr__res_generic_m3 w=12.1 l=10m
X171 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X172 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.5 as=6.95 ps=21.4 w=10 l=0.5
X173 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X174 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X175 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X176 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X177 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X178 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.4 as=7.55 ps=11.5 w=10 l=0.5
X179 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X180 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X181 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X182 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X183 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X184 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X185 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X186 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X187 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.5 as=6.95 ps=21.4 w=10 l=0.5
X188 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X189 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X190 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X191 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X192 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X193 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X194 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X195 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X196 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.4 as=7.55 ps=11.5 w=10 l=0.5
X197 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X198 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X199 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X200 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X201 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X202 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X203 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X204 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X205 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.5 as=6.95 ps=21.4 w=10 l=0.5
X206 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X207 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
.ends

.subckt sky130_fd_io__top_power_hvc_wpadv2 PADISOR PADISOL SRC_BDY_HVC OGC_HVC AMUXBUS_B
+ VSSIO_Q P_PAD sky130_fd_io__hvc_clampv2_0/m3_103_12712# VDDIO_Q P_CORE sky130_fd_io__hvc_clampv2_0/m3_10082_12712#
+ DRN_HVC VCCHIB VDDIO VDDA VCCD VSWITCH VSSA VSSIO VSSD AMUXBUS_A
Xsky130_fd_io__hvc_clampv2_0 OGC_HVC DRN_HVC P_PAD sky130_fd_io__hvc_clampv2_0/m3_10082_12712#
+ sky130_fd_io__hvc_clampv2_0/m3_103_12712# VDDIO_Q AMUXBUS_B VSSIO_Q SRC_BDY_HVC
+ VDDIO VCCHIB VSSIO VDDA VSSD P_CORE VSWITCH VCCD AMUXBUS_A VSSA sky130_fd_io__hvc_clampv2
.ends

.subckt sky130_ef_io__vddio_hvc_clamped_pad VDDA VSSIO_Q VDDIO VDDIO_Q VSSD VDDIO_PAD
+ VSSA AMUXBUS_B AMUXBUS_A VSWITCH VCCHIB VSSIO VCCD
Xsky130_fd_io__top_power_hvc_wpadv2_2 VDDIO_Q VDDIO_Q VSSIO VDDIO AMUXBUS_B VSSIO_Q
+ VDDIO_PAD VDDIO_Q VDDIO_Q VDDIO VDDIO_Q VDDIO VCCHIB VDDIO VDDA VCCD VSWITCH VSSA
+ VSSIO VSSD AMUXBUS_A sky130_fd_io__top_power_hvc_wpadv2
.ends

.subckt sky130_fd_io__top_ground_hvc_wpad VCCHIB VDDA VDDIO_Q VSSIO_Q G_PAD PADISOR
+ PADISOL DRN_HVC SRC_BDY_HVC OGC_HVC G_CORE AMUXBUS_B VDDIO VSSIO VSSD VSWITCH VCCD
+ AMUXBUS_A VSSA
Xsky130_fd_io__sio_clamp_pcap_4x5_0 SRC_BDY_HVC a_1268_5934# sky130_fd_io__sio_clamp_pcap_4x5
Xsky130_fd_io__com_busses_esd_0 VCCHIB G_PAD VSSD G_CORE AMUXBUS_A VCCD AMUXBUS_B
+ VDDIO VSSIO VSWITCH VSSA VDDA VSSIO_Q VDDIO_Q sky130_fd_io__com_busses_esd
Xsky130_fd_io__sio_clamp_pcap_4x5_1[0] SRC_BDY_HVC a_1268_5934# sky130_fd_io__sio_clamp_pcap_4x5
Xsky130_fd_io__sio_clamp_pcap_4x5_1[1] SRC_BDY_HVC a_1268_5934# sky130_fd_io__sio_clamp_pcap_4x5
Xsky130_fd_io__sio_clamp_pcap_4x5_1[2] SRC_BDY_HVC a_1268_5934# sky130_fd_io__sio_clamp_pcap_4x5
Xsky130_fd_io__esd_rcclamp_nfetcap_0[0|0] a_1268_5934# SRC_BDY_HVC sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[1|0] a_1268_5934# SRC_BDY_HVC sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[2|0] a_1268_5934# SRC_BDY_HVC sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[0|1] a_1268_5934# SRC_BDY_HVC sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[1|1] a_1268_5934# SRC_BDY_HVC sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[2|1] a_1268_5934# SRC_BDY_HVC sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[0|2] a_1268_5934# SRC_BDY_HVC sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[1|2] a_1268_5934# SRC_BDY_HVC sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[2|2] a_1268_5934# SRC_BDY_HVC sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[0|3] a_1268_5934# SRC_BDY_HVC sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[1|3] a_1268_5934# SRC_BDY_HVC sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[2|3] a_1268_5934# SRC_BDY_HVC sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[0|4] a_1268_5934# SRC_BDY_HVC sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[1|4] a_1268_5934# SRC_BDY_HVC sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[2|4] a_1268_5934# SRC_BDY_HVC sky130_fd_io__esd_rcclamp_nfetcap
X0 a_1368_5960# a_1268_5934# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=1.86 pd=14.5 as=0.98 ps=7.28 w=7 l=0.5
X1 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X2 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X3 SRC_BDY_HVC a_1268_5934# a_1368_5960# SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X4 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X5 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.4 as=7.55 ps=11.5 w=10 l=0.5
X6 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X7 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X8 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X9 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.4 as=7.55 ps=11.5 w=10 l=0.5
X10 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.86 ps=14.5 w=7 l=0.5
X11 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X12 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X13 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X14 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X15 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X16 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X17 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X18 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X19 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X20 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X21 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X22 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X23 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X24 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.5 as=6.95 ps=21.4 w=10 l=0.5
X25 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X26 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X27 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X28 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.5 as=6.95 ps=21.4 w=10 l=0.5
X29 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X30 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X31 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.4 as=7.55 ps=11.5 w=10 l=0.5
X32 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X33 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X34 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X35 a_1368_5960# a_1268_5934# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X36 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X37 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.4 as=7.55 ps=11.5 w=10 l=0.5
X38 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.5 as=6.95 ps=21.4 w=10 l=0.5
X39 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X40 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X41 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X42 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X43 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X44 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X45 a_1368_5960# a_1268_5934# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X46 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X47 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X48 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X49 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X50 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X51 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X52 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X53 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
R0 G_CORE PADISOL sky130_fd_pr__res_generic_m3 w=11.8 l=10m
X54 SRC_BDY_HVC a_1268_5934# a_1368_5960# SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X55 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X56 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X57 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.5 as=6.95 ps=21.4 w=10 l=0.5
X58 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X59 a_1368_5960# a_1268_5934# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X60 SRC_BDY_HVC a_1268_5934# a_1368_5960# SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X61 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X62 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X63 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X64 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X65 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X66 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X67 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.4 as=7.55 ps=11.5 w=10 l=0.5
X68 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X69 SRC_BDY_HVC a_1268_5934# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=10.5 as=55.8 ps=443 w=5 l=4
X70 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.5 as=6.95 ps=21.4 w=10 l=0.5
X71 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X72 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X73 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X74 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X75 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X76 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X77 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.4 as=7.55 ps=11.5 w=10 l=0.5
X78 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X79 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X80 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X81 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X82 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X83 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X84 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X85 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X86 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X87 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X88 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X89 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X90 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X91 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X92 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.4 as=7.55 ps=11.5 w=10 l=0.5
X93 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X94 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X95 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X96 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X97 SRC_BDY_HVC a_1268_5934# a_1368_5960# SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X98 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X99 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
R1 G_CORE PADISOR sky130_fd_pr__res_generic_m3 w=11.8 l=10m
X100 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X101 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X102 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X103 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X104 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X105 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.5 as=6.95 ps=21.4 w=10 l=0.5
X106 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X107 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X108 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X109 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X110 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X111 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X112 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X113 SRC_BDY_HVC a_1268_5934# a_1368_5960# SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X114 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X115 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X116 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X117 a_1368_5960# a_1268_5934# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X118 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X119 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.5 as=6.95 ps=21.4 w=10 l=0.5
X120 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X121 SRC_BDY_HVC a_1268_5934# a_1368_5960# SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X122 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X123 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X124 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X125 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X126 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X127 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.4 as=7.55 ps=11.5 w=10 l=0.5
X128 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.4 as=7.55 ps=11.5 w=10 l=0.5
X129 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X130 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X131 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X132 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
R2 DRN_HVC a_214_8638# sky130_fd_pr__res_generic_po w=0.33 l=700
X133 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X134 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X135 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X136 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X137 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X138 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X139 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X140 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X141 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X142 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X143 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X144 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X145 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X146 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X147 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.5 as=6.95 ps=21.4 w=10 l=0.5
X148 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X149 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X150 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X151 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=1.86 pd=14.5 as=0.98 ps=7.28 w=7 l=0.5
R3 a_1672_8638# a_214_8638# sky130_fd_pr__res_generic_po w=0.33 l=1.55k
X152 a_1368_5960# a_1268_5934# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X153 SRC_BDY_HVC a_1268_5934# a_1368_5960# SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X154 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X155 a_1368_5960# a_1268_5934# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.86 ps=14.5 w=7 l=0.5
X156 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X157 a_1368_5960# a_1268_5934# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X158 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
R4 a_1268_5934# a_1672_8638# sky130_fd_pr__res_generic_po w=0.33 l=470
X159 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X160 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X161 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X162 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X163 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X164 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X165 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X166 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X167 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X168 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X169 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X170 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X171 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X172 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.5 as=6.95 ps=21.4 w=10 l=0.5
X173 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X174 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X175 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X176 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X177 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X178 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.4 as=7.55 ps=11.5 w=10 l=0.5
X179 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X180 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X181 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X182 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X183 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X184 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X185 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X186 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X187 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.5 as=6.95 ps=21.4 w=10 l=0.5
X188 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X189 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X190 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X191 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X192 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X193 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X194 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X195 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X196 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.4 as=7.55 ps=11.5 w=10 l=0.5
X197 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X198 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X199 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X200 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X201 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X202 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X203 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X204 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X205 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.5 as=6.95 ps=21.4 w=10 l=0.5
X206 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X207 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
.ends

.subckt sky130_ef_io__vssio_hvc_clamped_pad VDDA VSSD VSSA AMUXBUS_B AMUXBUS_A VSSIO_PAD
+ VDDIO_Q VDDIO VSSIO VSSIO_Q VSWITCH VCCHIB VCCD
Xsky130_fd_io__top_ground_hvc_wpad_2 VCCHIB VDDA VDDIO_Q VSSIO_Q VSSIO_PAD VSSIO_Q
+ VSSIO_Q VDDIO VSSIO VDDIO VSSIO AMUXBUS_B VDDIO VSSIO VSSD VSWITCH VCCD AMUXBUS_A
+ VSSA sky130_fd_io__top_ground_hvc_wpad
.ends

.subckt sky130_ef_io__vdda_hvc_clamped_pad VDDIO_Q VSSIO_Q VSSIO VDDA_PAD AMUXBUS_B
+ AMUXBUS_A VDDA VCCHIB VSSD VSSA VSWITCH VCCD VDDIO
Xsky130_fd_io__top_power_hvc_wpadv2_1 sky130_fd_io__top_power_hvc_wpadv2_1/PADISOR
+ sky130_fd_io__top_power_hvc_wpadv2_1/PADISOL VSSA VDDIO AMUXBUS_B VSSIO_Q VDDA_PAD
+ sky130_fd_io__top_power_hvc_wpadv2_1/sky130_fd_io__hvc_clampv2_0/m3_103_12712# VDDIO_Q
+ VDDA sky130_fd_io__top_power_hvc_wpadv2_1/sky130_fd_io__hvc_clampv2_0/m3_10082_12712#
+ VDDA VCCHIB VDDIO VDDA VCCD VSWITCH VSSA VSSIO VSSD AMUXBUS_A sky130_fd_io__top_power_hvc_wpadv2
.ends

.subckt sky130_fd_io__top_ground_lvc_wpad PADISOR PADISOL VSSIO_Q VCCHIB VDDA VDDIO_Q
+ G_PAD SRC_BDY_LVC1 SRC_BDY_LVC2 BDY2_B2B DRN_LVC2 DRN_LVC1 G_CORE OGC_LVC AMUXBUS_B
+ VSSIO VDDIO VSSD VSWITCH VCCD AMUXBUS_A VSSA
Xsky130_fd_io__com_busses_esd_0 VCCHIB G_PAD VSSD G_CORE AMUXBUS_A VCCD AMUXBUS_B
+ VDDIO VSSIO VSWITCH VSSA VDDA VSSIO_Q VDDIO_Q sky130_fd_io__com_busses_esd
X0 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X1 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X2 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X3 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.7 pd=5.28 as=687 ps=3.1k w=5 l=8
X4 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X5 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X6 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X7 DRN_LVC1 a_414_306# a_450_404# DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X8 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X9 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X10 a_2872_5340# a_2595_15129# DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X11 SRC_BDY_LVC1 a_414_306# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=1.28k ps=3.48k w=7 l=8
X12 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=5.62 pd=12.2 as=2.92 ps=6.17 w=5 l=0.18
X13 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X14 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X15 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X16 SRC_BDY_LVC2 a_2595_15129# a_2872_5340# SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.4 pd=7.68 as=4.76 ps=15.4 w=7 l=0.18
X17 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X18 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X19 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X20 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.92 pd=6.17 as=5.62 ps=12.2 w=5 l=0.18
X21 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X22 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
R0 a_414_306# DRN_LVC1 sky130_fd_pr__res_generic_po w=0.33 l=1.95k
X23 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X24 a_450_404# a_414_306# DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X25 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X26 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X27 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X28 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X29 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.92 pd=6.17 as=5.62 ps=12.2 w=5 l=0.18
X30 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X31 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X32 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X33 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X34 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X35 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X36 DRN_LVC1 a_414_306# a_450_404# DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X37 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X38 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X39 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.4 pd=7.68 as=0 ps=0 w=7 l=8
X40 DRN_LVC1 a_414_306# a_450_404# DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
R1 a_2183_16816# a_2595_15129# sky130_fd_pr__res_generic_po w=0.33 l=200
X41 SRC_BDY_LVC1 a_414_306# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X42 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X43 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X44 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X45 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=5.62 pd=12.2 as=2.92 ps=6.17 w=5 l=0.18
X46 a_450_404# a_414_306# DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=1.96 ps=14.6 w=7 l=0.18
X47 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X48 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X49 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X50 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.92 pd=6.17 as=5.62 ps=12.2 w=5 l=0.18
X51 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X52 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X53 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
R2 a_1871_4484# a_13955_3836# sky130_fd_pr__res_generic_po w=0.33 l=300
X54 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X55 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X56 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X57 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X58 a_450_404# a_414_306# DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X59 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X60 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X61 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X62 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X63 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X64 DRN_LVC2 a_2595_15129# a_2872_5340# DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X65 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X66 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X67 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X68 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X69 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X70 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X71 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X72 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X73 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X74 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=5.62 pd=12.2 as=2.92 ps=6.17 w=5 l=0.18
X75 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X76 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X77 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X78 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X79 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
D0 SRC_BDY_LVC1 BDY2_B2B sky130_fd_pr__diode_pd2nw_05v5 pj=3.3e+07 area=2.25e+13
X80 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X81 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X82 DRN_LVC2 a_2595_15129# a_2872_5340# DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X83 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X84 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X85 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X86 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.7 pd=5.28 as=0 ps=0 w=5 l=8
X87 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
D1 BDY2_B2B SRC_BDY_LVC1 sky130_fd_pr__diode_pd2nw_05v5 pj=3.3e+07 area=2.25e+13
X88 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X89 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X90 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X91 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X92 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X93 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X94 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X95 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X96 SRC_BDY_LVC1 a_414_306# a_450_404# SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.4 pd=7.68 as=4.76 ps=15.4 w=7 l=0.18
X97 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X98 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X99 SRC_BDY_LVC1 a_414_306# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.4 pd=7.68 as=0 ps=0 w=7 l=8
X100 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X101 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.92 pd=6.17 as=5.62 ps=12.2 w=5 l=0.18
X102 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X103 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X104 DRN_LVC2 a_2595_15129# a_2872_5340# DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X105 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X106 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X107 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X108 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X109 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X110 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X111 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X112 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X113 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X114 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X115 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X116 a_2872_5340# a_2595_15129# DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X117 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X118 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X119 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X120 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X121 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X122 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X123 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X124 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X125 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X126 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X127 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X128 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X129 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.92 pd=6.17 as=5.62 ps=12.2 w=5 l=0.18
X130 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X131 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X132 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X133 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X134 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X135 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X136 SRC_BDY_LVC1 a_414_306# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.4 pd=7.68 as=0 ps=0 w=7 l=8
X137 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X138 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X139 a_2872_5340# a_2595_15129# DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=1.96 ps=14.6 w=7 l=0.18
X140 SRC_BDY_LVC1 a_414_306# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X141 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X142 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X143 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X144 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X145 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X146 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=5.62 pd=12.2 as=2.92 ps=6.17 w=5 l=0.18
X147 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X148 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X149 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X150 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X151 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X152 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X153 SRC_BDY_LVC1 a_414_306# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X154 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X155 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X156 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X157 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X158 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
D2 BDY2_B2B SRC_BDY_LVC1 sky130_fd_pr__diode_pd2nw_05v5 pj=3.3e+07 area=2.25e+13
X159 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X160 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X161 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X162 DRN_LVC1 a_414_306# a_450_404# DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X163 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X164 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X165 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X166 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X167 DRN_LVC2 a_2595_15129# a_2872_5340# DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X168 SRC_BDY_LVC1 a_414_306# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X169 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X170 a_450_404# a_414_306# DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X171 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X172 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X173 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X174 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X175 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X176 DRN_LVC1 a_414_306# a_450_404# DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X177 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X178 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X179 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X180 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X181 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X182 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X183 SRC_BDY_LVC1 a_414_306# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X184 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
R3 G_CORE PADISOR sky130_fd_pr__res_generic_m3 w=11.8 l=10m
X185 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X186 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X187 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X188 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X189 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X190 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X191 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X192 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X193 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X194 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X195 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X196 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
D3 BDY2_B2B SRC_BDY_LVC1 sky130_fd_pr__diode_pd2nw_05v5 pj=3.3e+07 area=2.25e+13
X197 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X198 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X199 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X200 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X201 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X202 DRN_LVC1 a_414_306# a_450_404# DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X203 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X204 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X205 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.7 pd=5.28 as=0 ps=0 w=5 l=8
R4 G_CORE PADISOL sky130_fd_pr__res_generic_m3 w=11.8 l=10m
X206 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X207 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X208 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.92 pd=6.17 as=5.62 ps=12.2 w=5 l=0.18
X209 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X210 DRN_LVC1 a_414_306# a_450_404# DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=1.96 pd=14.6 as=0.98 ps=7.28 w=7 l=0.18
X211 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
R5 DRN_LVC2 a_13955_3836# sky130_fd_pr__res_generic_po w=0.33 l=900
X212 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X213 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X214 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
R6 a_1871_4484# a_2183_16816# sky130_fd_pr__res_generic_po w=0.33 l=720
X215 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X216 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X217 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X218 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X219 SRC_BDY_LVC1 a_414_306# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X220 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X221 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X222 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X223 a_2872_5340# a_2595_15129# DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X224 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X225 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X226 a_2872_5340# a_2595_15129# DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X227 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X228 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X229 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X230 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X231 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X232 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X233 a_450_404# a_414_306# DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X234 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X235 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X236 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.92 pd=6.17 as=5.62 ps=12.2 w=5 l=0.18
X237 a_450_404# a_414_306# DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X238 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X239 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X240 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X241 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X242 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X243 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X244 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X245 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X246 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X247 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X248 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X249 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X250 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X251 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X252 DRN_LVC2 a_2595_15129# a_2872_5340# DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=1.96 pd=14.6 as=0.98 ps=7.28 w=7 l=0.18
X253 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X254 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X255 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X256 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X257 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=5.62 pd=12.2 as=2.92 ps=6.17 w=5 l=0.18
X258 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X259 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X260 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X261 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X262 a_2872_5340# a_2595_15129# DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X263 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X264 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
D4 SRC_BDY_LVC1 BDY2_B2B sky130_fd_pr__diode_pd2nw_05v5 pj=3.3e+07 area=2.25e+13
X265 SRC_BDY_LVC2 a_2595_15129# a_2872_5340# SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.4 pd=7.68 as=4.76 ps=15.4 w=7 l=0.18
X266 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X267 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X268 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X269 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X270 SRC_BDY_LVC1 a_414_306# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X271 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X272 DRN_LVC2 a_2595_15129# a_2872_5340# DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X273 a_450_404# a_414_306# DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X274 DRN_LVC2 a_2595_15129# a_2872_5340# DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X275 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X276 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.4 pd=7.68 as=0 ps=0 w=7 l=8
X277 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=5.62 pd=12.2 as=2.92 ps=6.17 w=5 l=0.18
X278 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X279 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X280 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X281 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X282 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X283 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X284 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X285 DRN_LVC2 a_2595_15129# a_2872_5340# DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X286 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X287 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X288 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X289 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X290 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X291 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X292 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X293 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X294 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X295 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X296 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X297 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X298 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X299 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X300 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X301 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X302 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X303 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X304 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X305 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
D5 SRC_BDY_LVC1 BDY2_B2B sky130_fd_pr__diode_pd2nw_05v5 pj=3.3e+07 area=2.25e+13
X306 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.7 pd=5.28 as=0 ps=0 w=5 l=8
X307 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X308 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=5.62 pd=12.2 as=2.92 ps=6.17 w=5 l=0.18
X309 DRN_LVC1 a_414_306# a_450_404# DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=1.96 pd=14.6 as=0.98 ps=7.28 w=7 l=0.18
X310 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X311 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X312 SRC_BDY_LVC1 a_414_306# a_450_404# SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.4 pd=7.68 as=4.76 ps=15.4 w=7 l=0.18
X313 a_2872_5340# a_2595_15129# DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=1.96 ps=14.6 w=7 l=0.18
X314 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X315 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X316 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X317 a_450_404# a_414_306# DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X318 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X319 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.92 pd=6.17 as=5.62 ps=12.2 w=5 l=0.18
X320 DRN_LVC2 a_2595_15129# a_2872_5340# DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=1.96 pd=14.6 as=0.98 ps=7.28 w=7 l=0.18
X321 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X322 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X323 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X324 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X325 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X326 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X327 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X328 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X329 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X330 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X331 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X332 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X333 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X334 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X335 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=5.62 pd=12.2 as=2.92 ps=6.17 w=5 l=0.18
X336 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X337 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X338 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X339 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
D6 SRC_BDY_LVC1 BDY2_B2B sky130_fd_pr__diode_pd2nw_05v5 pj=3.3e+07 area=2.25e+13
X340 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X341 SRC_BDY_LVC1 a_414_306# a_450_404# SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.4 pd=7.68 as=4.76 ps=15.4 w=7 l=0.18
X342 SRC_BDY_LVC1 a_414_306# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.4 pd=7.68 as=0 ps=0 w=7 l=8
X343 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X344 DRN_LVC1 a_414_306# a_450_404# DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X345 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X346 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X347 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X348 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X349 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X350 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X351 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X352 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X353 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X354 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X355 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X356 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X357 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X358 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X359 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X360 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X361 a_450_404# a_414_306# DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=1.96 ps=14.6 w=7 l=0.18
X362 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X363 SRC_BDY_LVC1 a_414_306# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X364 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X365 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X366 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X367 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X368 SRC_BDY_LVC1 a_414_306# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X369 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X370 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X371 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X372 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=5.62 pd=12.2 as=2.92 ps=6.17 w=5 l=0.18
X373 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X374 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X375 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X376 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X377 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.7 pd=5.28 as=0 ps=0 w=5 l=8
X378 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X379 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X380 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X381 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X382 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X383 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X384 SRC_BDY_LVC1 a_414_306# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X385 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X386 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X387 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X388 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X389 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X390 a_2872_5340# a_2595_15129# DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X391 a_2872_5340# a_2595_15129# DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X392 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X393 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X394 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X395 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=5.62 pd=12.2 as=2.92 ps=6.17 w=5 l=0.18
X396 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
D7 BDY2_B2B SRC_BDY_LVC1 sky130_fd_pr__diode_pd2nw_05v5 pj=3.3e+07 area=2.25e+13
X397 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X398 a_450_404# a_414_306# DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X399 a_2872_5340# a_2595_15129# DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X400 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X401 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X402 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X403 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X404 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X405 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X406 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X407 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X408 SRC_BDY_LVC1 a_414_306# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X409 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X410 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X411 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X412 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X413 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.7 pd=5.28 as=0 ps=0 w=5 l=8
X414 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X415 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X416 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X417 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X418 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X419 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X420 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X421 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X422 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X423 DRN_LVC1 a_414_306# a_450_404# DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X424 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X425 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X426 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X427 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X428 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X429 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X430 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X431 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=1.33 pd=10.5 as=0 ps=0 w=5 l=4
X432 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X433 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X434 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X435 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.92 pd=6.17 as=5.62 ps=12.2 w=5 l=0.18
X436 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X437 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X438 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X439 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X440 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X441 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X442 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.92 pd=6.17 as=5.62 ps=12.2 w=5 l=0.18
X443 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X444 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X445 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X446 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X447 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X448 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X449 DRN_LVC2 a_2595_15129# a_2872_5340# DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X450 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X451 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X452 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
.ends

.subckt sky130_ef_io__vssd_lvc_clamped3_pad VDDA VSSIO_Q VSSD1 VCCD VSSD AMUXBUS_B
+ AMUXBUS_A VSSA VSSD_PAD VSWITCH VCCHIB VDDIO VDDIO_Q VSSIO VCCD1
Xsky130_fd_io__top_ground_lvc_wpad_1 sky130_fd_io__top_ground_lvc_wpad_1/PADISOR sky130_fd_io__top_ground_lvc_wpad_1/PADISOL
+ VSSIO_Q VCCHIB VDDA VDDIO_Q VSSD_PAD VSSD1 VSSD1 VSSIO VCCD1 VCCD1 VSSD1 VSSIO AMUXBUS_B
+ VSSIO VDDIO VSSD VSWITCH VCCD AMUXBUS_A VSSA sky130_fd_io__top_ground_lvc_wpad
.ends

.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=2.89
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=2.89
.ends

.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=0.59
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=0.59
.ends

.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=4.73
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=4.73
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=1.05
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=1.05
.ends

.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=1.97
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=1.97
.ends

.subckt user_id_programming mask_rev[0] mask_rev[10] mask_rev[11] mask_rev[12] mask_rev[14]
+ mask_rev[15] mask_rev[16] mask_rev[17] mask_rev[18] mask_rev[19] mask_rev[1] mask_rev[20]
+ mask_rev[21] mask_rev[22] mask_rev[23] mask_rev[24] mask_rev[25] mask_rev[26] mask_rev[27]
+ mask_rev[29] mask_rev[2] mask_rev[30] mask_rev[31] mask_rev[3] mask_rev[4] mask_rev[5]
+ mask_rev[6] mask_rev[7] mask_rev[8] mask_rev[9] mask_rev[28] mask_rev[13] VPWR VGND
Xmask_rev_value\[1\] VGND VGND VPWR VPWR mask_rev_value\[1\]/HI mask_rev[1] sky130_fd_sc_hd__conb_1
XFILLER_6_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmask_rev_value\[30\] VGND VGND VPWR VPWR mask_rev_value\[30\]/HI mask_rev[30] sky130_fd_sc_hd__conb_1
XFILLER_0_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmask_rev_value\[23\] VGND VGND VPWR VPWR mask_rev_value\[23\]/HI mask_rev[23] sky130_fd_sc_hd__conb_1
XFILLER_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmask_rev_value\[16\] VGND VGND VPWR VPWR mask_rev_value\[16\]/HI mask_rev[16] sky130_fd_sc_hd__conb_1
XFILLER_0_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmask_rev_value\[21\] VGND VGND VPWR VPWR mask_rev_value\[21\]/HI mask_rev[21] sky130_fd_sc_hd__conb_1
XFILLER_3_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmask_rev_value\[14\] VGND VGND VPWR VPWR mask_rev_value\[14\]/HI mask_rev[14] sky130_fd_sc_hd__conb_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmask_rev_value\[8\] VGND VGND VPWR VPWR mask_rev_value\[8\]/HI mask_rev[8] sky130_fd_sc_hd__conb_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmask_rev_value\[12\] VGND VGND VPWR VPWR mask_rev_value\[12\]/HI mask_rev[12] sky130_fd_sc_hd__conb_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmask_rev_value\[6\] VGND VGND VPWR VPWR mask_rev_value\[6\]/HI mask_rev[6] sky130_fd_sc_hd__conb_1
XFILLER_1_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmask_rev_value\[28\] VGND VGND VPWR VPWR mask_rev_value\[28\]/HI mask_rev[28] sky130_fd_sc_hd__conb_1
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmask_rev_value\[10\] VGND VGND VPWR VPWR mask_rev_value\[10\]/HI mask_rev[10] sky130_fd_sc_hd__conb_1
XFILLER_1_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmask_rev_value\[4\] VGND VGND VPWR VPWR mask_rev_value\[4\]/HI mask_rev[4] sky130_fd_sc_hd__conb_1
XFILLER_7_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmask_rev_value\[26\] VGND VGND VPWR VPWR mask_rev_value\[26\]/HI mask_rev[26] sky130_fd_sc_hd__conb_1
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmask_rev_value\[19\] VGND VGND VPWR VPWR mask_rev_value\[19\]/HI mask_rev[19] sky130_fd_sc_hd__conb_1
Xmask_rev_value\[2\] VGND VGND VPWR VPWR mask_rev_value\[2\]/HI mask_rev[2] sky130_fd_sc_hd__conb_1
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmask_rev_value\[31\] VGND VGND VPWR VPWR mask_rev_value\[31\]/HI mask_rev[31] sky130_fd_sc_hd__conb_1
Xmask_rev_value\[24\] VGND VGND VPWR VPWR mask_rev_value\[24\]/HI mask_rev[24] sky130_fd_sc_hd__conb_1
Xmask_rev_value\[17\] VGND VGND VPWR VPWR mask_rev_value\[17\]/HI mask_rev[17] sky130_fd_sc_hd__conb_1
XFILLER_5_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmask_rev_value\[0\] VGND VGND VPWR VPWR mask_rev_value\[0\]/HI mask_rev[11] sky130_fd_sc_hd__conb_1
XFILLER_5_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmask_rev_value\[22\] VGND VGND VPWR VPWR mask_rev_value\[22\]/HI mask_rev[22] sky130_fd_sc_hd__conb_1
XFILLER_2_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmask_rev_value\[15\] VGND VGND VPWR VPWR mask_rev_value\[15\]/HI mask_rev[15] sky130_fd_sc_hd__conb_1
XFILLER_2_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmask_rev_value\[9\] VGND VGND VPWR VPWR mask_rev_value\[9\]/HI mask_rev[9] sky130_fd_sc_hd__conb_1
XFILLER_8_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmask_rev_value\[20\] VGND VGND VPWR VPWR mask_rev_value\[20\]/HI mask_rev[20] sky130_fd_sc_hd__conb_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmask_rev_value\[13\] VGND VGND VPWR VPWR mask_rev_value\[13\]/HI mask_rev[13] sky130_fd_sc_hd__conb_1
Xmask_rev_value\[7\] VGND VGND VPWR VPWR mask_rev_value\[7\]/HI mask_rev[7] sky130_fd_sc_hd__conb_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmask_rev_value\[29\] VGND VGND VPWR VPWR mask_rev_value\[29\]/HI mask_rev[29] sky130_fd_sc_hd__conb_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmask_rev_value\[11\] VGND VGND VPWR VPWR mask_rev_value\[11\]/HI mask_rev[0] sky130_fd_sc_hd__conb_1
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmask_rev_value\[5\] VGND VGND VPWR VPWR mask_rev_value\[5\]/HI mask_rev[5] sky130_fd_sc_hd__conb_1
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmask_rev_value\[27\] VGND VGND VPWR VPWR mask_rev_value\[27\]/HI mask_rev[27] sky130_fd_sc_hd__conb_1
XFILLER_6_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmask_rev_value\[3\] VGND VGND VPWR VPWR mask_rev_value\[3\]/HI mask_rev[3] sky130_fd_sc_hd__conb_1
XFILLER_6_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmask_rev_value\[25\] VGND VGND VPWR VPWR mask_rev_value\[25\]/HI mask_rev[25] sky130_fd_sc_hd__conb_1
Xmask_rev_value\[18\] VGND VGND VPWR VPWR mask_rev_value\[18\]/HI mask_rev[18] sky130_fd_sc_hd__conb_1
.ends

.subckt sky130_ef_io__vssd_lvc_clamped_pad VDDA VSSD_PAD VCCD VSWITCH VDDIO VDDIO_Q
+ AMUXBUS_B AMUXBUS_A VSSD VSSIO VSSIO_Q VCCHIB VSSA
Xsky130_fd_io__top_ground_lvc_wpad_1 sky130_fd_io__top_ground_lvc_wpad_1/PADISOR sky130_fd_io__top_ground_lvc_wpad_1/PADISOL
+ VSSIO_Q VCCHIB VDDA VDDIO_Q VSSD_PAD VSSIO VSSD VSSA VCCD VCCD VSSD VSSA AMUXBUS_B
+ VSSIO VDDIO VSSD VSWITCH VCCD AMUXBUS_A VSSA sky130_fd_io__top_ground_lvc_wpad
.ends

.subckt sky130_ef_io__vccd_lvc_clamped3_pad VDDA VCCHIB VSSD1 VDDIO VSWITCH AMUXBUS_B
+ VSSIO AMUXBUS_A VCCD VCCD_PAD VCCD1 VSSD VDDIO_Q VSSA VSSIO_Q
Xsky130_fd_io__top_power_lvc_wpad_0 VSSIO_Q VCCHIB VDDA VDDIO_Q VCCD_PAD VSSD1 VSSD1
+ VSSIO VCCD1 VCCD1 VCCD1 sky130_fd_io__top_power_lvc_wpad_0/PADISOR sky130_fd_io__top_power_lvc_wpad_0/PADISOL
+ VSSIO AMUXBUS_B VSSIO VDDIO VSSD VSWITCH VCCD AMUXBUS_A VSSA sky130_fd_io__top_power_lvc_wpad
.ends

.subckt sky130_fd_sc_hvl__decap_4 VGND VNB VPB VPWR
X0 VGND VPWR VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.412 ps=4.1 w=0.75 l=1
X1 VPWR VGND VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.55 ps=5.1 w=1 l=1
.ends

.subckt sky130_fd_sc_hvl__decap_8 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.275 pd=2.55 as=0.84 ps=7.68 w=1 l=1
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.623 ps=6.16 w=0.75 l=1
X2 VPWR VGND VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0 ps=0 w=1 l=1
X3 VGND VPWR VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0 ps=0 w=0.75 l=1
.ends

.subckt sky130_fd_sc_hvl__diode_2 DIODE VGND VNB VPB VPWR
D0 VNB DIODE sky130_fd_pr__diode_pw2nd_11v0 pj=3.16e+06 area=6.072e+11
.ends

.subckt sky130_fd_sc_hvl__lsbufhv2lv_1 A LVPWR VGND VNB VPB VPWR X
X0 a_30_1337# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.12 ps=1.41 w=0.42 l=0.5
X1 VGND a_30_1337# a_30_207# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.179 pd=1.26 as=0.12 ps=1.41 w=0.42 l=0.5
X2 VGND a_30_207# a_389_141# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.105 ps=1.03 w=0.75 l=0.5
X3 VGND a_30_207# a_389_141# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.199 ps=2.03 w=0.75 l=0.5
X4 a_389_1337# a_30_1337# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.105 ps=1.03 w=0.75 l=0.5
X5 VGND a_30_207# a_389_141# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.199 ps=2.03 w=0.75 l=0.5
X6 VGND A a_30_1337# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.179 pd=1.26 as=0.12 ps=1.41 w=0.42 l=0.5
X7 VGND a_30_1337# a_389_1337# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.199 ps=2.03 w=0.75 l=0.5
X8 a_389_141# a_30_207# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.179 ps=1.26 w=0.75 l=0.5
X9 VGND a_30_1337# a_389_1337# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X10 LVPWR a_389_141# X LVPWR sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.4 as=0.297 ps=2.77 w=1.12 l=0.15
X11 VGND a_389_141# X VNB sky130_fd_pr__nfet_01v8 ad=0.196 pd=2.01 as=0.196 ps=2.01 w=0.74 l=0.15
X12 a_389_1337# a_30_1337# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.179 ps=1.26 w=0.75 l=0.5
X13 LVPWR a_389_1337# a_389_141# LVPWR sky130_fd_pr__pfet_01v8_hvt ad=0.297 pd=2.77 as=0.297 ps=2.77 w=1.12 l=0.15
X14 a_30_207# a_30_1337# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.12 ps=1.41 w=0.42 l=0.5
X15 a_389_1337# a_389_141# LVPWR LVPWR sky130_fd_pr__pfet_01v8_hvt ad=0.297 pd=2.77 as=0.157 ps=1.4 w=1.12 l=0.15
.ends

.subckt xres_buf A X LVPWR LVGND VPWR VGND
XFILLER_0_24 VGND VGND VPWR VPWR sky130_fd_sc_hvl__decap_4
XFILLER_1_0 VGND VGND VPWR VPWR sky130_fd_sc_hvl__decap_8
XFILLER_0_16 VGND VGND VPWR VPWR sky130_fd_sc_hvl__decap_8
XFILLER_1_8 VGND VGND VPWR VPWR sky130_fd_sc_hvl__decap_4
XANTENNA_lvlshiftdown_A A VGND VGND VPWR VPWR sky130_fd_sc_hvl__diode_2
XFILLER_2_0 VGND VGND VPWR VPWR sky130_fd_sc_hvl__decap_8
XFILLER_0_0 VGND VGND VPWR VPWR sky130_fd_sc_hvl__decap_8
XFILLER_0_8 VGND VGND VPWR VPWR sky130_fd_sc_hvl__decap_8
Xlvlshiftdown A LVPWR VGND VGND VPWR VPWR X sky130_fd_sc_hvl__lsbufhv2lv_1
.ends

.subckt sky130_ef_io__vssa_hvc_clamped_pad VSSD VSSA VDDIO VSSA_PAD VCCHIB VSWITCH
+ VSSIO VDDIO_Q VDDA VSSIO_Q VCCD AMUXBUS_B AMUXBUS_A
Xsky130_fd_io__top_ground_hvc_wpad_0 VCCHIB VDDA VDDIO_Q VSSIO_Q VSSA_PAD sky130_fd_io__top_ground_hvc_wpad_0/PADISOR
+ sky130_fd_io__top_ground_hvc_wpad_0/PADISOL VDDA VSSA VDDIO VSSA AMUXBUS_B VDDIO
+ VSSIO VSSD VSWITCH VCCD AMUXBUS_A VSSA sky130_fd_io__top_ground_hvc_wpad
.ends

.subckt sky130_fd_io__com_res_weak_v2 a_n281_1306# a_534_6146#
R0 a_n13_3671# m1_3_3617# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R1 a_n283_3382# a_n283_2797# sky130_fd_pr__res_generic_po w=0.8 l=1.5
R2 m1_n268_3094# a_n283_2797# sky130_fd_pr__res_generic_m1 w=0.66 l=10m
R3 m1_n268_1364# a_n281_1306# sky130_fd_pr__res_generic_m1 w=0.66 l=10m
R4 m1_3_3580# a_n13_2329# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R5 a_n13_3671# a_n13_2329# sky130_fd_pr__res_generic_po w=0.8 l=6
R6 a_n283_2797# a_n283_2447# sky130_fd_pr__res_generic_po w=0.8 l=1.5
R7 a_n283_2447# m1_n268_1924# sky130_fd_pr__res_generic_m1 w=0.66 l=10m
R8 a_n283_2797# m1_n268_2513# sky130_fd_pr__res_generic_m1 w=0.66 l=10m
R9 a_n13_2329# a_n283_3382# sky130_fd_pr__res_generic_po w=0.8 l=6
R10 a_n13_2329# m1_2_2233# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R11 m1_n268_1924# a_n281_1656# sky130_fd_pr__res_generic_m1 w=0.66 l=10m
R12 a_n13_6243# a_534_6146# sky130_fd_pr__res_generic_po w=0.8 l=50
R13 a_n13_6243# a_n13_3671# sky130_fd_pr__res_generic_po w=0.8 l=12
R14 m1_n268_2513# a_n283_2447# sky130_fd_pr__res_generic_m1 w=0.66 l=10m
R15 m1_2_2233# a_n283_3382# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R16 a_n283_2447# a_n281_1656# sky130_fd_pr__res_generic_po w=0.8 l=1.5
R17 a_n283_3382# m1_n268_3094# sky130_fd_pr__res_generic_m1 w=0.66 l=10m
R18 a_n281_1656# m1_n268_1364# sky130_fd_pr__res_generic_m1 w=0.66 l=10m
R19 a_n281_1656# a_n281_1306# sky130_fd_pr__res_generic_po w=0.8 l=1.5
.ends

.subckt sky130_fd_io__xres4v2_in_buf VGND IN_H VDDIO VNORMAL VNORMAL_B PAD ENABLE_HV
+ IN_H_N VCCHIB ENABLE_VDDIO_LV a_n445_2580# m2_288_2575# w_4058_2188# a_n32352_n9635#
Xsky130_fd_io__inv_1_0 VGND VCCHIB VCCHIB VGND sky130_fd_io__inv_1_0/Y ENABLE_VDDIO_LV
+ sky130_fd_io__inv_1
X0 a_n445_2580# sky130_fd_io__inv_1_0/Y VCCHIB VCCHIB sky130_fd_pr__pfet_g5v0d10v5 ad=1.4 pd=10.6 as=0.7 ps=5.28 w=5 l=0.5
X1 VDDIO VNORMAL a_157_2580# VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.4 ps=10.6 w=5 l=0.5
X2 a_469_2037# a_n176_869# a_n232_901# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X3 a_n29280_n8739# VNORMAL_B a_n31524_n8739# VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.4 ps=10.6 w=5 l=0.5
X4 a_n11573_n8777# a_111_449# VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.5
X5 VGND a_n176_869# a_2300_3398# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X6 a_1560_2580# ENABLE_HV VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.84 pd=6.56 as=0.795 ps=6.53 w=3 l=0.5
X7 VGND IN_H_N IN_H VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.5
X8 VGND PAD a_n232_901# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X9 a_n232_901# a_n176_869# a_469_2037# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.6 as=0.7 ps=5.28 w=5 l=0.8
X10 a_2165_2545# a_n176_869# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.84 pd=6.56 as=0.795 ps=6.53 w=3 l=0.5
X11 VGND a_2165_2545# a_2356_3115# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.5
X12 VDDIO a_2356_3115# a_2300_3398# VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.118 ps=1.4 w=0.42 l=0.5
X13 IN_H_N a_2300_3398# VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.84 pd=6.56 as=0.795 ps=6.53 w=3 l=0.5
X14 a_5826_2675# ENABLE_HV VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X15 a_n176_869# PAD w_5030_2188# w_5030_2188# sky130_fd_pr__pfet_g5v0d10v5 ad=0.28 pd=2.56 as=0.28 ps=2.56 w=1 l=0.8
X16 a_n16_901# a_n176_869# a_n232_901# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.6 as=1.4 ps=10.6 w=5 l=0.8
X17 a_1560_2580# ENABLE_HV VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=1.4 pd=10.6 as=1.33 ps=10.5 w=5 l=0.5
X18 a_n232_901# PAD VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X19 IN_H IN_H_N VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.84 pd=6.56 as=0.42 ps=3.28 w=3 l=0.5
X20 VDDIO a_5826_2675# a_111_449# VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.6
X21 IN_H_N a_2300_3398# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.84 pd=6.56 as=0.795 ps=6.53 w=3 l=0.5
X22 VGND a_5826_2675# a_111_449# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.185 ps=1.93 w=0.7 l=0.6
X23 a_2356_3115# a_2165_2545# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X24 VDDIO a_111_449# a_n29280_n8739# VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.5
X25 VDDIO VNORMAL_B a_5826_2675# VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X26 a_n176_869# PAD a_n232_901# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.4 ps=10.6 w=5 l=0.8
X27 a_n9813_4210# VNORMAL_B a_n11573_n8777# VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X28 VGND VNORMAL_B a_5852_3096# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X29 a_2300_3398# a_n176_869# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.5
X30 w_4058_2188# a_111_449# a_n445_2580# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.28 pd=2.56 as=0.28 ps=2.56 w=1 l=0.9
X31 VGND VGND VGND VGND sky130_fd_pr__nfet_05v0_nvt ad=2.65 pd=20.5 as=4.71 ps=36.5 w=10 l=0.9
X32 a_2165_2545# a_n176_869# w_4058_2188# w_4058_2188# sky130_fd_pr__pfet_g5v0d10v5 ad=1.4 pd=10.6 as=1.4 ps=10.6 w=5 l=0.5
X33 IN_H IN_H_N VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.28 pd=2.56 as=0.14 ps=1.28 w=1 l=0.5
X34 IN_H IN_H_N VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.5
X35 a_469_2037# a_n176_869# a_n232_901# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X36 a_n29280_n8739# a_n31524_n8739# VGND sky130_fd_pr__res_generic_nd__hv w=0.29 l=1.08k
X37 VDDIO IN_H_N IN_H VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X38 a_n232_901# PAD a_n176_869# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X39 a_n757_2580# a_111_449# w_5030_2188# VGND sky130_fd_pr__nfet_05v0_nvt ad=2.8 pd=20.6 as=2.8 ps=20.6 w=10 l=0.9
X40 a_n16_901# VNORMAL_B VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=1.4 pd=10.6 as=0.7 ps=5.28 w=5 l=0.5
X41 VCCHIB sky130_fd_io__inv_1_0/Y a_n757_2580# VCCHIB sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.4 ps=10.6 w=5 l=0.5
R0 a_n9813_4210# a_n11573_n8777# sky130_fd_pr__res_generic_po w=0.4 l=714
X42 w_5030_2188# w_5030_2188# w_5030_2188# w_5030_2188# sky130_fd_pr__pfet_g5v0d10v5 ad=0.28 pd=2.56 as=0.84 ps=7.68 w=1 l=0.8
X43 a_n232_901# a_n176_869# a_469_2037# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X44 a_5826_2675# ENABLE_HV VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X45 VDDIO a_5826_2675# a_111_449# VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.6
X46 a_n176_869# PAD a_n31524_n8739# VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=1.4 pd=10.6 as=1.4 ps=10.6 w=5 l=0.5
X47 a_2165_2545# a_n176_869# a_n9813_4210# VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=1.4 pd=10.6 as=0.7 ps=5.28 w=5 l=0.5
X48 a_469_2037# PAD a_157_2580# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.28 pd=2.56 as=0.28 ps=2.56 w=1 l=0.9
X49 a_5852_3096# ENABLE_HV a_5826_2675# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.185 ps=1.93 w=0.7 l=0.6
X50 IN_H IN_H_N VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X51 VDDIO VNORMAL_B a_5826_2675# VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X52 a_2356_3115# a_2300_3398# VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.118 pd=1.4 as=0.0588 ps=0.7 w=0.42 l=0.5
.ends

.subckt sky130_fd_io__xres_inv_hysv2 VCC_IO VSSD OUT_H a_122_112# a_322_144# a_322_604#
X0 a_578_144# a_122_112# a_322_604# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.84 pd=6.56 as=0.42 ps=3.28 w=3 l=1
X1 a_322_144# OUT_H VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.118 pd=1.4 as=0.118 ps=1.4 w=0.42 l=1
X2 a_322_144# a_122_112# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=1
X3 a_578_144# a_122_112# a_322_144# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.28 pd=2.56 as=0.14 ps=1.28 w=1 l=1
X4 OUT_H a_578_144# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.84 pd=6.56 as=0.84 ps=6.56 w=3 l=0.5
X5 VCC_IO OUT_H a_322_604# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.118 pd=1.4 as=0.118 ps=1.4 w=0.42 l=1
X6 OUT_H a_578_144# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.28 pd=2.56 as=0.28 ps=2.56 w=1 l=0.5
X7 a_322_604# a_122_112# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.84 ps=6.56 w=3 l=1
.ends

.subckt sky130_fd_io__gpio_buf_localesdv2 VTRIP_SEL_H VGND OUT_H OUT_VT sky130_fd_io__res250only_small_0/PAD
+ VCC_IO
Xsky130_fd_io__signal_5_sym_hv_local_5term_0 VGND VCC_IO OUT_VT VGND VCC_IO VCC_IO
+ sky130_fd_io__signal_5_sym_hv_local_5term
Xsky130_fd_io__signal_5_sym_hv_local_5term_1 VGND VCC_IO VGND VGND OUT_VT VCC_IO sky130_fd_io__signal_5_sym_hv_local_5term
Xsky130_fd_io__signal_5_sym_hv_local_5term_2 VGND VCC_IO OUT_H VGND VCC_IO VCC_IO
+ sky130_fd_io__signal_5_sym_hv_local_5term
Xsky130_fd_io__signal_5_sym_hv_local_5term_3 VGND VCC_IO VGND VGND OUT_H VCC_IO sky130_fd_io__signal_5_sym_hv_local_5term
Xsky130_fd_io__res250only_small_0 sky130_fd_io__res250only_small_0/PAD OUT_H sky130_fd_io__res250only_small
X0 OUT_VT VTRIP_SEL_H OUT_H VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=1
.ends

.subckt sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2 VCC_IO a_10282_1285# a_5322_1285#
+ a_8980_1457# a_7988_1457# a_2036_1457# a_13940_1457# a_12948_1457# a_12266_1285#
+ a_7306_1285# a_5012_1457# a_3900_1285# a_2908_1285# a_5884_1285# a_14178_1285# a_10844_1285#
+ a_1354_1285# a_7868_1285# a_12828_1285# a_8860_1285# a_13820_1285# a_4330_1285#
+ a_3338_1285# a_6996_1457# a_11956_1457# a_1044_1457# a_11274_1285# a_6314_1285#
+ w_469_785# a_9972_1457# a_4020_1457# a_3028_1457# a_8298_1285# a_13258_1285# a_9290_1285#
+ a_1916_1285# a_6004_1457# a_4892_1285# a_6876_1285# a_924_1285# a_11836_1285# a_2346_1285#
+ a_9852_1285# a_10964_1457#
X0 w_469_785# a_5322_1285# a_5012_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X1 a_9972_1457# a_9852_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X2 w_469_785# a_11274_1285# a_10964_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X3 a_10964_1457# a_10844_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X4 a_6996_1457# a_6876_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X5 w_469_785# a_2346_1285# a_2036_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X6 a_2036_1457# a_1916_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X7 w_469_785# a_12266_1285# a_11956_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X8 w_469_785# a_6314_1285# a_6004_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X9 a_11956_1457# a_11836_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X10 w_469_785# a_9290_1285# a_8980_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X11 a_5012_1457# a_4892_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X12 w_469_785# a_10282_1285# a_9972_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X13 w_469_785# a_4330_1285# a_4020_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X14 a_4020_1457# a_3900_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X15 a_8980_1457# a_8860_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X16 w_469_785# a_3338_1285# a_3028_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X17 w_469_785# a_8298_1285# a_7988_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X18 a_1044_1457# a_924_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.42 ps=11.4 w=5 l=0.6
X19 w_469_785# a_7306_1285# a_6996_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X20 a_13940_1457# a_13820_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=2.97 pd=6.19 as=3.78 ps=11.5 w=5 l=0.6
X21 a_3028_1457# a_2908_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X22 a_7988_1457# a_7868_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X23 w_469_785# a_13258_1285# a_12948_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X24 a_12948_1457# a_12828_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X25 w_469_785# a_14178_1285# a_13940_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.42 pd=11.4 as=2.97 ps=6.19 w=5 l=0.6
X26 w_469_785# a_1354_1285# a_1044_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X27 a_6004_1457# a_5884_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X28 w_469_785# a_11274_1285# a_10964_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X29 w_469_785# a_5322_1285# a_5012_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X30 a_9972_1457# a_9852_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X31 a_10964_1457# a_10844_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X32 w_469_785# a_2346_1285# a_2036_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X33 a_6996_1457# a_6876_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X34 w_469_785# a_6314_1285# a_6004_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X35 a_2036_1457# a_1916_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X36 w_469_785# a_12266_1285# a_11956_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X37 a_11956_1457# a_11836_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X38 a_5012_1457# a_4892_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X39 w_469_785# a_4330_1285# a_4020_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X40 w_469_785# a_9290_1285# a_8980_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X41 a_8980_1457# a_8860_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X42 w_469_785# a_10282_1285# a_9972_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X43 a_1044_1457# a_924_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.42 ps=11.4 w=5 l=0.6
X44 a_4020_1457# a_3900_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X45 w_469_785# a_3338_1285# a_3028_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X46 w_469_785# a_8298_1285# a_7988_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X47 a_3028_1457# a_2908_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X48 a_7988_1457# a_7868_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X49 w_469_785# a_13258_1285# a_12948_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X50 w_469_785# a_7306_1285# a_6996_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X51 a_13940_1457# a_13820_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=2.97 pd=6.19 as=3.78 ps=11.5 w=5 l=0.6
X52 a_12948_1457# a_12828_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X53 w_469_785# a_1354_1285# a_1044_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X54 w_469_785# a_14178_1285# a_13940_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.42 pd=11.4 as=2.97 ps=6.19 w=5 l=0.6
X55 a_6004_1457# a_5884_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
.ends

.subckt sky130_fd_io__gpio_pddrvr_strong_xres4v2 PD_H[2] PD_H[3] TIE_LO_ESD VGND_IO
+ sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_11956_1457# sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_6996_1457#
+ sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_1044_1457# sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_9972_1457#
+ sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_3028_1457# sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_4020_1457#
+ sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_6004_1457# sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_10964_1457#
+ w_335_3259# sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_12948_1457# sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_7988_1457#
+ sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_13940_1457# sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_8980_1457#
+ sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_2036_1457# m1_785_3898# sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_5012_1457#
+ VCC_IO
Xsky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0 VCC_IO PD_H[3] m1_9769_3903# sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_8980_1457#
+ sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_7988_1457# sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_2036_1457#
+ sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_13940_1457# sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_12948_1457#
+ m1_2697_3903# m1_7657_3903# sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_5012_1457#
+ m1_11193_3903# m1_11193_3903# m1_8232_3903# m1_785_3898# PD_H[3] m1_12747_3903#
+ PD_H[2] m1_2135_3903# PD_H[2] m1_785_3898# m1_9769_3903# m1_11193_3903# sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_6996_1457#
+ sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_11956_1457# sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_1044_1457#
+ PD_H[3] m1_8232_3903# w_335_3259# sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_9972_1457#
+ sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_4020_1457# sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_3028_1457#
+ PD_H[2] m1_785_3898# PD_H[3] m1_12747_3903# sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_6004_1457#
+ m1_9769_3903# m1_8232_3903# m1_12747_3903# PD_H[3] m1_12747_3903# PD_H[3] sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_10964_1457#
+ sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2
R0 m2_6804_1099# PD_H[2] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R1 m2_12763_1099# PD_H[2] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R2 m1_2135_3903# m2_1848_1400# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R3 m2_13622_1100# TIE_LO_ESD sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R4 m1_12747_3903# m2_12763_1400# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R5 m2_1260_1100# PD_H[2] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R6 m1_7657_3903# m2_6804_1400# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R7 m2_897_1099# PD_H[2] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R8 m1_12747_3903# m2_13622_1100# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R9 m1_2135_3903# m2_1260_1100# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R10 m1_785_3898# m2_897_1400# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R11 m2_12189_1099# TIE_LO_ESD sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R12 m2_9986_1099# PD_H[2] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R13 m2_413_1100# TIE_LO_ESD sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R14 m2_3095_1099# PD_H[3] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R15 m2_9366_1099# TIE_LO_ESD sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R16 m1_11193_3903# m2_12189_1400# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R17 m1_9769_3903# m2_9986_1400# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R18 m1_785_3898# m2_413_1100# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R19 m1_2697_3903# m2_3095_1400# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R20 m1_8232_3903# m2_9366_1400# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R21 m2_11758_1100# PD_H[3] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R22 m1_11193_3903# m2_11758_1100# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R23 m2_8935_1100# PD_H[3] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R24 m2_10846_1099# TIE_LO_ESD sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R25 m2_656_1099# PD_H[3] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R26 m2_11329_1099# PD_H[2] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R27 m2_1565_1099# PD_H[3] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R28 m2_3378_1099# TIE_LO_ESD sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R29 m1_8232_3903# m2_8935_1100# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R30 m1_9769_3903# m2_10846_1400# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R31 m1_11193_3903# m2_11329_1400# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R32 m2_8506_1099# PD_H[2] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R33 m2_10415_1100# PD_H[3] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R34 m1_785_3898# m2_656_1400# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R35 m2_7664_1099# TIE_LO_ESD sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R36 m1_2135_3903# m2_1565_1400# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R37 m1_2697_3903# m2_3378_1400# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R38 m1_8232_3903# m2_8506_1400# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R39 m1_9769_3903# m2_10415_1100# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R40 m1_7657_3903# m2_7664_1400# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R41 m2_7233_1100# PD_H[3] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R42 m2_13193_1099# PD_H[3] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R43 m2_2790_1100# PD_H[2] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R44 m1_7657_3903# m2_7233_1100# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R45 m1_12747_3903# m2_13193_1400# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R46 TIE_LO_ESD VGND_IO sky130_fd_pr__res_generic_po w=0.5 l=10.2
R47 m2_1848_1099# TIE_LO_ESD sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R48 m1_2697_3903# m2_2790_1100# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
.ends

.subckt sky130_fd_io__tk_tie_r_out_esd A B
R0 A B sky130_fd_pr__res_generic_po w=0.5 l=10.2
.ends

.subckt sky130_fd_io__xres2v2_rcfilter_lpfv2 IN VCC_IO a_9105_2295# a_1381_4189# a_7373_4189#
+ a_3949_4189# a_2237_4189# a_525_4189# a_472_471# a_7393_2295# a_472_1087# a_8249_2295#
+ a_5661_4189# a_472_779# a_336_26# a_472_317# a_472_1549# a_6517_4189# a_6537_2295#
+ a_9941_4189# a_472_163# a_3093_4189# a_472_1395# a_4805_4189# a_9961_2295# a_9085_4189#
+ a_472_1857#
X0 a_472_317# a_472_1087# a_472_317# a_336_26# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=25.3 ps=189 w=7 l=4
X1 a_9941_4189# a_9941_4189# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R0 m1_14480_2172# a_11618_2147# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R1 a_11618_3071# m1_14484_3300# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R2 m1_14480_4922# a_7373_4189# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R3 IN m1_14484_4202# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R4 m1_11613_5471# a_7373_4189# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R5 m1_14328_5846# a_5661_4189# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X2 a_3382_6882# a_7373_4189# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
X3 a_7373_4189# a_7373_4189# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R6 a_472_6420# m1_3338_6444# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R7 m1_14480_5846# a_5661_4189# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R8 m1_3363_1728# a_3382_1703# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R9 m1_14480_3096# a_11618_3071# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R10 a_7373_4189# m1_14484_5126# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R11 a_472_317# m1_3338_341# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R12 a_472_7344# m1_3338_7368# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R13 a_472_1395# m1_467_1384# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R14 a_472_779# m1_467_769# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
X4 VCC_IO a_2237_4189# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=25.3 ps=189 w=7 l=4
X5 a_11618_3379# a_11618_3379# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R15 m1_3334_1112# a_472_1087# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R16 a_472_1857# m1_5939_1932# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R17 m1_3363_496# a_3382_471# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X6 a_472_7036# a_3382_7190# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
X7 a_472_317# a_12884_625# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
R18 a_11618_2455# m1_14484_2684# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X8 a_9085_4189# a_9085_4189# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R19 a_472_1395# m1_10927_1419# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X9 a_6517_4189# a_6517_4189# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R20 a_472_6728# m1_3338_6752# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X10 a_472_6728# a_472_6728# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R21 a_7373_4189# m1_14484_5434# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R22 a_472_317# m1_5624_734# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X11 a_472_317# a_7393_2295# a_472_317# a_336_26# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=4
R23 a_472_7652# m1_3338_7676# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X12 a_11618_3687# a_11618_3687# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R24 a_472_317# m1_6480_426# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R25 m1_3363_1112# a_3382_1087# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X13 a_3382_7190# a_9085_4189# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
X14 a_472_317# a_12884_933# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
R26 a_11618_2763# m1_14484_2992# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R27 m1_14299_5846# a_472_1395# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R28 m1_467_432# a_472_317# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R29 a_472_317# m1_4825_1042# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X15 VCC_IO a_7373_4189# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=4
R30 a_472_317# m1_6537_426# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R31 a_472_317# m1_4768_1042# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X16 a_472_6728# a_12884_6728# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
X17 a_472_1549# a_3382_1703# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R32 a_6517_4189# m1_14484_5742# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X18 a_472_6112# a_472_6112# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
X19 a_7373_4189# a_7373_4189# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
X20 a_472_317# a_8249_2295# a_472_317# a_336_26# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=4
R33 a_472_7036# m1_3338_7060# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X21 a_472_7036# a_472_7036# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R34 a_472_471# m1_467_461# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R35 a_472_7344# m1_3338_7419# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X22 a_472_1087# a_3382_1087# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R36 m1_2201_1652# a_472_1549# sky130_fd_pr__res_generic_m1 w=0.29 l=10m
R37 a_472_317# m1_3338_700# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X23 VCC_IO a_7373_4189# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=4
X24 a_3382_1703# a_11618_2147# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
R38 m1_10929_804# a_472_779# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X25 a_472_6420# a_472_6420# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
X26 a_472_6112# a_12884_6112# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
X27 a_472_779# a_3382_779# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R39 a_7373_4189# m1_11741_5169# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R40 a_472_6728# m1_3338_6803# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X28 a_472_7344# a_472_7344# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
X29 a_472_7036# a_12884_7036# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
R41 a_472_7652# m1_3338_7727# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X30 a_472_1395# a_3382_1395# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R42 a_472_317# m1_2201_1681# sky130_fd_pr__res_generic_m1 w=0.29 l=10m
X31 a_472_317# a_472_779# a_472_317# a_336_26# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=4
X32 a_3382_1087# a_11618_2763# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
R43 m1_10929_188# a_472_163# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X33 a_11618_2147# a_12884_1857# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R44 a_472_1549# m1_466_1664# sky130_fd_pr__res_generic_m1 w=0.29 l=0.31
X34 a_472_317# a_472_1857# a_472_317# a_336_26# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=4
X35 a_472_317# a_472_471# a_472_317# a_336_26# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=4
R45 a_472_6112# m1_3338_6187# sky130_fd_pr__res_generic_m1 w=0.29 l=0.31
R46 m1_3334_6907# a_472_6728# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X36 a_472_6420# a_12884_6420# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
X37 a_472_7652# a_472_7652# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
X38 a_472_7344# a_12884_7344# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
X39 a_472_163# a_3382_163# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
X40 VCC_IO a_3949_4189# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=4
X41 VCC_IO a_5661_4189# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=4
X42 a_3382_1395# a_11618_2455# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
R47 m1_10929_496# a_472_471# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X43 a_11618_2455# a_12884_1549# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R48 a_472_7036# m1_3338_7111# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X44 a_11618_3379# a_12884_625# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R49 a_472_6420# m1_3338_6495# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R50 a_472_317# m1_3338_392# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X45 a_7373_4189# a_12884_6728# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
X46 a_472_317# a_6537_2295# a_472_317# a_336_26# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=4
R51 m1_3363_6907# a_3382_6882# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X47 a_472_7652# a_12884_7652# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
X48 a_9085_4189# a_12884_7344# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R52 a_11618_2147# m1_14484_2325# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X49 a_472_471# a_3382_471# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R53 m1_10958_804# a_472_1395# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R54 a_11618_3071# m1_14484_3249# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R55 m1_3334_7215# a_472_7036# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R56 a_472_317# m1_3338_1265# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X50 a_11618_2763# a_12884_1241# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R57 a_472_1395# m1_10927_1470# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X51 VCC_IO a_6517_4189# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=4
R58 m1_3334_6599# a_472_6420# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X52 a_11618_3687# a_12884_317# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R59 a_472_317# m1_3113_1350# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R60 a_9941_4189# m1_14484_4459# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X53 a_3382_779# a_11618_3071# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
X54 a_6517_4189# a_12884_6420# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R61 a_472_317# m1_3056_1350# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R62 m1_10958_188# a_472_1395# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X55 a_7373_4189# a_12884_7036# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
X56 a_472_317# a_9105_2295# a_472_317# a_336_26# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=4
R63 a_11618_2455# m1_14484_2633# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X57 a_472_317# a_472_1549# a_472_317# a_336_26# sky130_fd_pr__nfet_g5v0d10v5 ad=1.86 pd=14.5 as=0 ps=0 w=7 l=4
R64 a_11618_3379# m1_14484_3557# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X58 a_472_317# a_472_1395# a_472_317# a_336_26# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=4
R65 a_472_1549# m1_3338_1573# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X59 a_472_1549# a_472_1549# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R66 m1_3334_7523# a_472_7344# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R67 a_5661_4189# m1_11613_5808# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R68 m1_3363_7215# a_3382_7190# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R69 m1_14509_2480# a_12884_1549# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R70 m1_3363_6599# a_3382_6574# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R71 m1_10929_1728# a_472_1549# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R72 a_9085_4189# m1_14484_4767# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X60 VCC_IO a_3093_4189# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=4
R73 m1_14509_4306# a_12884_7652# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R74 m1_3334_804# a_472_779# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R75 a_472_317# m1_3338_1008# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X61 VCC_IO a_525_4189# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=1.86 pd=14.5 as=0 ps=0 w=7 l=4
X62 a_5661_4189# a_12884_6112# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
X63 a_11618_3071# a_12884_933# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R76 m1_10958_496# a_472_1395# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R77 a_11618_2763# m1_14484_2941# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R78 m1_11613_4547# a_9941_4189# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R79 m1_14509_5230# a_12884_6728# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X64 a_472_7652# a_3382_7806# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R80 m1_1345_1960# a_472_1857# sky130_fd_pr__res_generic_m1 w=0.29 l=10m
X65 a_3382_163# a_11618_3687# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
X66 a_472_317# a_472_317# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R81 a_472_1857# m1_3338_1881# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R82 a_11618_3687# m1_14484_3865# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X67 a_472_1857# a_472_1857# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
X68 a_472_1549# a_12884_1549# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
R83 m1_3334_7831# a_472_7652# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R84 m1_14509_3404# a_12884_625# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X69 a_9941_4189# a_12884_7652# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
X70 a_11618_2455# a_11618_2455# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R85 m1_3363_7523# a_3382_7498# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R86 m1_3334_188# a_472_163# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R87 m1_14509_2788# a_12884_1241# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X71 a_472_6112# a_3382_6266# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R88 a_472_1549# m1_595_1664# sky130_fd_pr__res_generic_m1 w=0.29 l=0.31
X72 a_472_317# a_472_163# a_472_317# a_336_26# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=4
R89 m1_14509_4614# a_12884_7344# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R90 m1_3334_6291# a_472_6112# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R91 a_472_317# m1_3338_1316# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R92 m1_10958_1728# a_472_1395# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R93 a_9085_4189# m1_11613_4576# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R94 a_472_317# m1_1345_1989# sky130_fd_pr__res_generic_m1 w=0.29 l=10m
R95 m1_10929_1112# a_472_1087# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R96 IN m1_14484_4151# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R97 m1_11613_4855# a_9085_4189# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R98 m1_14509_5538# a_12884_6420# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X73 a_3382_7806# IN a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
X74 a_3382_471# a_11618_3379# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
R99 m1_14480_2480# a_11618_2455# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R100 a_9941_4189# m1_14484_4510# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R101 a_7373_4189# m1_14484_5075# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R102 m1_11613_5779# a_6517_4189# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
X75 a_472_317# a_472_317# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
X76 a_472_1857# a_12884_1857# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
R103 m1_14509_3712# a_12884_317# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R104 a_472_317# m1_3338_649# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X77 VCC_IO a_4805_4189# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=4
X78 a_11618_2763# a_11618_2763# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R105 m1_3363_7831# a_3382_7806# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R106 m1_14480_4306# a_9941_4189# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R107 a_472_1857# m1_5939_1881# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R108 m1_3334_496# a_472_471# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X79 a_472_6420# a_3382_6574# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
X80 a_3382_6266# a_6517_4189# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
X81 a_472_317# a_472_317# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R109 m1_3334_1420# a_472_1395# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R110 m1_14480_5230# a_7373_4189# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R111 a_11618_3379# m1_14484_3608# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R112 a_6517_4189# m1_11613_5500# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
X82 a_472_7344# a_3382_7498# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R113 a_472_1549# m1_3338_1624# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R114 m1_14509_2172# a_12884_1857# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R115 m1_14509_4922# a_12884_7036# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R116 m1_467_1047# a_472_317# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R117 a_7373_4189# m1_11613_4884# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R118 a_472_317# m1_5681_734# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R119 m1_3363_6291# a_3382_6266# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R120 m1_14480_3404# a_11618_3379# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R121 m1_14509_5846# a_12884_6112# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R122 m1_14509_3096# a_12884_933# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R123 m1_10958_1112# a_472_1395# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R124 m1_14480_2788# a_11618_2763# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R125 a_9085_4189# m1_14484_4818# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X83 a_472_317# a_9961_2295# a_472_317# a_336_26# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=4
X84 a_472_317# a_472_317# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R126 a_7373_4189# m1_14484_5383# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R127 a_472_317# m1_3338_957# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X85 IN IN a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R128 m1_14480_4614# a_9085_4189# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R129 m1_3363_804# a_3382_779# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X86 VCC_IO a_9085_4189# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=4
X87 a_472_6728# a_3382_6882# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
X88 a_3382_6574# a_7373_4189# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
R130 m1_3334_1728# a_472_1549# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X89 a_472_317# a_12884_1241# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
R131 a_472_6112# m1_3338_6136# sky130_fd_pr__res_generic_m1 w=0.29 l=0.31
R132 m1_14480_5538# a_6517_4189# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X90 VCC_IO a_1381_4189# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=4
X91 a_11618_2147# a_11618_2147# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R133 a_472_1857# m1_3338_1932# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R134 m1_3363_1420# a_3382_1395# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R135 a_472_1087# m1_467_1076# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R136 a_11618_3687# m1_14484_3916# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X92 a_3382_7498# a_9941_4189# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
X93 VCC_IO a_9941_4189# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=4
R137 m1_467_1355# a_472_317# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R138 a_7373_4189# m1_11612_5169# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X94 a_11618_3071# a_11618_3071# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R139 m1_14480_3712# a_11618_3687# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R140 m1_467_740# a_472_317# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R141 m1_3363_188# a_3382_163# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X95 a_472_317# a_12884_317# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
R142 a_11618_2147# m1_14484_2376# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R143 a_6517_4189# m1_14484_5691# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
.ends

.subckt sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2 w_415_600# a_4969_1552# a_2303_1380#
+ a_5961_1552# a_13777_1380# a_8817_1380# a_4287_1380# a_10921_1552# a_7945_1552#
+ a_12905_1552# a_7263_1380# a_12223_1380# a_9929_1552# a_9247_1380# a_2865_1380#
+ a_1993_1552# a_5841_1380# a_4849_1380# a_10801_1380# a_14135_1380# a_1311_1380#
+ a_3977_1552# a_12785_1380# a_7825_1380# a_3295_1380# a_6953_1552# a_9809_1380# a_11913_1552#
+ a_1001_1552# a_6271_1380# a_5279_1380# a_11231_1380# a_10239_1380# a_13897_1552#
+ a_8937_1552# a_8255_1380# a_1873_1380# a_13215_1380# a_3857_1380# a_2985_1552# a_11793_1380#
+ a_881_1380# a_6833_1380#
X0 a_13897_1552# a_13777_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.97 pd=6.19 as=3.78 ps=11.5 w=5 l=0.6
X1 a_4969_1552# a_4849_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X2 a_8937_1552# a_8817_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X3 w_415_600# a_10239_1380# a_9929_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X4 a_1993_1552# a_1873_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X5 w_415_600# a_3295_1380# a_2985_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X6 w_415_600# a_14135_1380# a_13897_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=4.3 pd=11.7 as=2.97 ps=6.19 w=5 l=0.6
X7 a_5961_1552# a_5841_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X8 w_415_600# a_2303_1380# a_1993_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X9 w_415_600# a_7263_1380# a_6953_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X10 a_4969_1552# a_4849_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X11 w_415_600# a_11231_1380# a_10921_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X12 a_12905_1552# a_12785_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X13 w_415_600# a_10239_1380# a_9929_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X14 a_8937_1552# a_8817_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X15 w_415_600# a_3295_1380# a_2985_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X16 w_415_600# a_2303_1380# a_1993_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X17 w_415_600# a_7263_1380# a_6953_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X18 a_12905_1552# a_12785_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X19 a_3977_1552# a_3857_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X20 a_7945_1552# a_7825_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X21 w_415_600# a_13215_1380# a_12905_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X22 w_415_600# a_1311_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X23 w_415_600# a_6271_1380# a_5961_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X24 a_3977_1552# a_3857_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X25 w_415_600# a_5279_1380# a_4969_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X26 a_11913_1552# a_11793_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X27 a_7945_1552# a_7825_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X28 w_415_600# a_9247_1380# a_8937_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X29 a_10921_1552# a_10801_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X30 w_415_600# a_13215_1380# a_12905_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X31 w_415_600# a_1311_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X32 w_415_600# a_6271_1380# a_5961_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X33 a_1001_1552# a_881_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=4.32 ps=11.7 w=5 l=0.6
X34 a_2985_1552# a_2865_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X35 w_415_600# a_5279_1380# a_4969_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X36 a_11913_1552# a_11793_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X37 a_10921_1552# a_10801_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X38 a_6953_1552# a_6833_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X39 w_415_600# a_9247_1380# a_8937_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X40 w_415_600# a_12223_1380# a_11913_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X41 a_1001_1552# a_881_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=4.32 ps=11.7 w=5 l=0.6
X42 a_9929_1552# a_9809_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X43 a_2985_1552# a_2865_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X44 w_415_600# a_4287_1380# a_3977_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X45 a_6953_1552# a_6833_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X46 w_415_600# a_8255_1380# a_7945_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X47 w_415_600# a_12223_1380# a_11913_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X48 a_13897_1552# a_13777_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.97 pd=6.19 as=3.78 ps=11.5 w=5 l=0.6
X49 a_9929_1552# a_9809_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X50 a_1993_1552# a_1873_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X51 w_415_600# a_4287_1380# a_3977_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X52 w_415_600# a_14135_1380# a_13897_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=4.3 pd=11.7 as=2.97 ps=6.19 w=5 l=0.6
X53 w_415_600# a_8255_1380# a_7945_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X54 a_5961_1552# a_5841_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X55 w_415_600# a_11231_1380# a_10921_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
.ends

.subckt sky130_fd_io__gpio_pudrvr_strong_axres4v2 PU_H_N[3] PU_H_N[2] sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_11913_1552#
+ sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_8937_1552# sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_13897_1552#
+ TIE_HI_ESD sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_2985_1552# sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_4969_1552#
+ sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_5961_1552# sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_10921_1552#
+ sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_7945_1552# sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_12905_1552#
+ VNB sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_9929_1552# li_11868_461#
+ sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_1993_1552# sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_3977_1552#
+ sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/w_415_600# sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_6953_1552#
+ a_14575_48# sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_1001_1552#
Xsky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0 sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/w_415_600#
+ sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_4969_1552# PU_H_N[2] sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_5961_1552#
+ m1_14229_1478# m1_8837_1478# PU_H_N[3] sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_10921_1552#
+ sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_7945_1552# sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_12905_1552#
+ PU_H_N[3] m1_11745_1478# sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_9929_1552#
+ m1_8837_1478# PU_H_N[2] sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_1993_1552#
+ PU_H_N[3] PU_H_N[3] m1_10391_1478# m1_14229_1478# PU_H_N[2] sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_3977_1552#
+ PU_H_N[2] PU_H_N[3] PU_H_N[2] sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_6953_1552#
+ m1_10391_1478# sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_11913_1552# sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_1001_1552#
+ PU_H_N[3] PU_H_N[3] m1_11745_1478# m1_10391_1478# sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_13897_1552#
+ sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_8937_1552# m1_8837_1478# PU_H_N[2]
+ m1_13667_1478# PU_H_N[3] sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_2985_1552#
+ m1_11745_1478# PU_H_N[2] PU_H_N[3] sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2
R0 m1_14229_1478# m2_14532_958# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R1 m1_13667_1478# m2_13593_958# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R2 TIE_HI_ESD a_14575_48# sky130_fd_pr__res_generic_po w=0.5 l=10.2
R3 m2_9839_n208# PU_H_N[2] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R4 m1_10391_1478# m2_10945_92# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R5 m2_11422_n209# PU_H_N[2] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R6 m1_13667_1478# m2_14075_958# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R7 m1_11745_1478# m2_12267_n279# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R8 m1_11745_1478# m2_12510_21# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R9 m1_8837_1478# m2_9605_92# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R10 m2_10945_n209# TIE_HI_ESD sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R11 m1_8837_1478# m2_9363_92# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R12 m1_10391_1478# m2_11422_92# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R13 m2_9605_n209# PU_H_N[3] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R14 m2_12510_n280# PU_H_N[3] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R15 m2_14769_657# PU_H_N[2] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R16 m2_11186_n208# PU_H_N[3] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R17 m2_13837_658# PU_H_N[3] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R18 m2_14286_658# TIE_HI_ESD sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R19 m2_14532_657# PU_H_N[3] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R20 m1_10391_1478# m2_11186_n208# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R21 m2_13593_657# TIE_HI_ESD sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R22 m2_12751_n280# PU_H_N[2] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R23 m1_13667_1478# m2_13837_658# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R24 m1_14229_1478# m2_14769_958# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R25 m1_11745_1478# m2_12751_21# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R26 m2_9363_n209# TIE_HI_ESD sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R27 m2_12267_n279# TIE_HI_ESD sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R28 m1_8837_1478# m2_9839_n208# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R29 m1_14229_1478# m2_14286_658# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R30 m2_14075_657# PU_H_N[2] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
.ends

.subckt sky130_fd_io__top_xres4v2 XRES_H_N FILT_IN_H ENABLE_VDDIO TIE_WEAK_HI_H ENABLE_H
+ PULLUP_H EN_VDDIO_SIG_H TIE_LO_ESD TIE_HI_ESD DISABLE_PULLUP_H INP_SEL_H VSSA VSSD
+ AMUXBUS_B AMUXBUS_A VDDIO_Q VDDIO VSWITCH VDDA VCCD VCCHIB VSSIO_Q VSSIO PAD PAD_A_ESD_H
Xsky130_fd_io__com_res_weak_v2_0 PULLUP_H a_5670_7125# sky130_fd_io__com_res_weak_v2
Xsky130_fd_io__com_res_weak_0 VDDIO sky130_fd_io__com_res_weak_0/RB li_7794_26629#
+ li_9658_25954# li_12154_26629# li_8568_25954# li_11000_25954# sky130_fd_io__com_res_weak
Xsky130_fd_io__xres4v2_in_buf_0 VSSD sky130_fd_io__xres4v2_in_buf_0/IN_H VDDIO_Q EN_VDDIO_SIG_H
+ sky130_fd_io__xres4v2_in_buf_0/VNORMAL_B sky130_fd_io__xres4v2_in_buf_0/PAD ENABLE_H
+ sky130_fd_io__xres4v2_in_buf_0/IN_H_N VCCHIB ENABLE_VDDIO m1_3250_3609# EN_VDDIO_SIG_H
+ m1_1351_2970# VSSD sky130_fd_io__xres4v2_in_buf
Xsky130_fd_io__xres_inv_hysv2_0 VDDIO_Q VSSD sky130_fd_io__xres_inv_hysv2_0/OUT_H
+ m1_6377_8979# li_6043_2944# li_5552_2976# sky130_fd_io__xres_inv_hysv2
Xsky130_fd_io__gpio_buf_localesdv2_0 VSSD VSSD sky130_fd_io__xres4v2_in_buf_0/PAD
+ sky130_fd_io__gpio_buf_localesdv2_0/OUT_VT PAD VDDIO sky130_fd_io__gpio_buf_localesdv2
Xsky130_fd_io__gpio_pddrvr_strong_xres4v2_0 sky130_fd_io__gpio_pddrvr_strong_xres4v2_0/PD_H[3]
+ sky130_fd_io__gpio_pddrvr_strong_xres4v2_0/PD_H[3] sky130_fd_io__gpio_pddrvr_strong_xres4v2_0/PD_H[3]
+ VSSIO PAD PAD PAD PAD PAD PAD PAD PAD VSSIO PAD PAD PAD PAD PAD m1_915_33059# PAD
+ VDDIO sky130_fd_io__gpio_pddrvr_strong_xres4v2
Xsky130_fd_io__tk_tie_r_out_esd_0 VDDIO TIE_HI_ESD sky130_fd_io__tk_tie_r_out_esd
Xsky130_fd_io__tk_tie_r_out_esd_1 VSSIO TIE_LO_ESD sky130_fd_io__tk_tie_r_out_esd
Xsky130_fd_io__res250only_small_0 TIE_WEAK_HI_H sky130_fd_io__com_res_weak_0/RB sky130_fd_io__res250only_small
Xsky130_fd_io__res250only_small_1 PAD PAD_A_ESD_H sky130_fd_io__res250only_small
Xsky130_fd_io__xres2v2_rcfilter_lpfv2_0 sky130_fd_io__xres2v2_rcfilter_lpfv2_0/IN
+ VDDIO_Q m1_10468_10072# m1_6377_8979# m1_10468_9216# m1_10468_4936# m1_10468_3224#
+ m1_10468_1512# m1_10468_4936# m1_10468_9216# m1_10468_3224# m1_10468_9216# m1_10468_6648#
+ m1_10468_4080# VSSD VSSD m1_10468_1512# m1_10468_7504# m1_10468_7504# m1_10468_10928#
+ m1_10468_5792# m1_10468_4080# m1_6377_8979# m1_10468_5792# m1_10468_10928# m1_10468_10072#
+ m1_10468_6648# sky130_fd_io__xres2v2_rcfilter_lpfv2
Xsky130_fd_io__gpio_pudrvr_strong_axres4v2_0 sky130_fd_io__gpio_pudrvr_strong_axres4v2_0/PU_H_N[3]
+ sky130_fd_io__gpio_pudrvr_strong_axres4v2_0/PU_H_N[3] PAD PAD PAD sky130_fd_io__gpio_pudrvr_strong_axres4v2_0/PU_H_N[3]
+ PAD PAD PAD PAD PAD PAD VSSD PAD VSSD PAD PAD VDDIO PAD VDDIO PAD sky130_fd_io__gpio_pudrvr_strong_axres4v2
X0 a_5670_7125# a_5551_5929# VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.5
X1 XRES_H_N a_5556_4246# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X2 VDDIO_Q a_5556_4246# XRES_H_N VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X3 FILT_IN_H a_3226_2008# sky130_fd_io__xres2v2_rcfilter_lpfv2_0/IN VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.84 pd=6.56 as=0.84 ps=6.56 w=3 l=0.5
X4 VDDIO_Q EN_VDDIO_SIG_H sky130_fd_io__xres4v2_in_buf_0/VNORMAL_B VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X5 VSSD DISABLE_PULLUP_H a_5525_5809# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X6 VSSD a_5525_5809# a_5551_5929# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X7 VSSD INP_SEL_H a_3226_2008# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X8 VDDIO_Q a_5556_4246# XRES_H_N VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X9 a_5525_5809# DISABLE_PULLUP_H VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X10 a_5525_5809# DISABLE_PULLUP_H VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X11 a_3226_2008# INP_SEL_H VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X12 VSSD a_5556_4246# XRES_H_N VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X13 a_5551_5929# a_5525_5809# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.185 ps=1.93 w=0.7 l=0.6
X14 a_5556_4246# sky130_fd_io__xres_inv_hysv2_0/OUT_H VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X15 XRES_H_N a_5556_4246# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X16 VDDIO_Q a_5556_4246# XRES_H_N VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X17 VDDIO_Q a_5556_4246# XRES_H_N VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X18 VDDIO a_5551_5929# a_5670_7125# VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.5
X19 XRES_H_N a_5556_4246# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X20 VSSD a_5556_4246# XRES_H_N VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X21 VDDIO_Q a_5556_4246# XRES_H_N VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X22 sky130_fd_io__xres2v2_rcfilter_lpfv2_0/IN a_3226_2008# sky130_fd_io__xres4v2_in_buf_0/IN_H VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.84 pd=6.56 as=0.84 ps=6.56 w=3 l=0.5
X23 XRES_H_N a_5556_4246# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X24 VDDIO_Q EN_VDDIO_SIG_H sky130_fd_io__xres4v2_in_buf_0/VNORMAL_B VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X25 sky130_fd_io__xres4v2_in_buf_0/VNORMAL_B EN_VDDIO_SIG_H VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X26 XRES_H_N a_5556_4246# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X27 VDDIO a_5525_5809# a_5551_5929# VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X28 VDDIO a_5525_5809# a_5551_5929# VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X29 VDDIO a_5551_5929# a_5670_7125# VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X30 a_5670_7125# a_5551_5929# VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X31 VDDIO DISABLE_PULLUP_H a_5525_5809# VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X32 VDDIO DISABLE_PULLUP_H a_5525_5809# VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X33 a_5556_4246# sky130_fd_io__xres_inv_hysv2_0/OUT_H VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X34 a_3226_2008# INP_SEL_H VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X35 VDDIO_Q INP_SEL_H a_3226_2008# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X36 XRES_H_N a_5556_4246# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X37 a_5551_5929# a_5525_5809# VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X38 a_5551_5929# a_5525_5809# VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X39 VDDIO_Q a_5556_4246# XRES_H_N VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X40 XRES_H_N a_5556_4246# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X41 VSSD a_5556_4246# XRES_H_N VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X42 FILT_IN_H INP_SEL_H sky130_fd_io__xres2v2_rcfilter_lpfv2_0/IN VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.84 pd=6.56 as=0.84 ps=6.56 w=3 l=0.5
X43 VSSD EN_VDDIO_SIG_H sky130_fd_io__xres4v2_in_buf_0/VNORMAL_B VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X44 sky130_fd_io__xres4v2_in_buf_0/VNORMAL_B EN_VDDIO_SIG_H VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X45 XRES_H_N a_5556_4246# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X46 a_3226_2008# INP_SEL_H VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.185 ps=1.93 w=0.7 l=0.6
X47 a_5525_5809# DISABLE_PULLUP_H VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X48 sky130_fd_io__xres2v2_rcfilter_lpfv2_0/IN INP_SEL_H sky130_fd_io__xres4v2_in_buf_0/IN_H VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.84 pd=6.56 as=0.84 ps=6.56 w=3 l=0.5
X49 VDDIO_Q a_5556_4246# XRES_H_N VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X50 VDDIO_Q INP_SEL_H a_3226_2008# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X51 VSSD a_5556_4246# XRES_H_N VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X52 XRES_H_N a_5556_4246# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X53 a_5556_4246# sky130_fd_io__xres_inv_hysv2_0/OUT_H VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X54 XRES_H_N a_5556_4246# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.185 ps=1.93 w=0.7 l=0.6
X55 XRES_H_N a_5556_4246# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X56 VDDIO_Q a_5556_4246# XRES_H_N VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X57 sky130_fd_io__xres4v2_in_buf_0/VNORMAL_B EN_VDDIO_SIG_H VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X58 XRES_H_N a_5556_4246# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
.ends

.subckt chip_io_openframe vddio_pad vssio_pad vdda1_pad2 vccd2_pad vddio vccd vdda
+ vdda1 vdda2 vccd1 vccd2 porb_l por_l resetb_h resetb_l mask_rev[31] mask_rev[30]
+ mask_rev[29] mask_rev[28] mask_rev[27] mask_rev[26] mask_rev[25] mask_rev[24] mask_rev[23]
+ mask_rev[22] mask_rev[21] mask_rev[20] mask_rev[19] mask_rev[18] mask_rev[17] mask_rev[16]
+ mask_rev[15] mask_rev[14] mask_rev[13] mask_rev[12] mask_rev[11] mask_rev[10] mask_rev[9]
+ mask_rev[8] mask_rev[7] mask_rev[6] mask_rev[5] mask_rev[4] mask_rev[3] mask_rev[2]
+ mask_rev[1] mask_rev[0] gpio[36] gpio_out[41] gpio_out[39] gpio_out[38] gpio_out[37]
+ gpio_out[36] gpio_out[35] gpio_out[33] gpio_out[32] gpio_out[30] gpio_out[26] gpio_out[23]
+ gpio_out[18] gpio_out[17] gpio_out[16] gpio_out[15] gpio_out[13] gpio_out[12] gpio_oeb[43]
+ gpio_oeb[42] gpio_oeb[41] gpio_oeb[37] gpio_oeb[34] gpio_oeb[29] gpio_oeb[28] gpio_oeb[27]
+ gpio_oeb[26] gpio_oeb[25] gpio_oeb[24] gpio_oeb[23] gpio_oeb[22] gpio_oeb[21] gpio_oeb[20]
+ gpio_oeb[18] gpio_oeb[17] gpio_oeb[16] gpio_oeb[15] gpio_oeb[14] gpio_oeb[13] gpio_oeb[6]
+ gpio_oeb[3] gpio_oeb[0] gpio_inp_dis[39] gpio_inp_dis[37] gpio_inp_dis[36] gpio_inp_dis[33]
+ gpio_inp_dis[32] gpio_inp_dis[22] gpio_inp_dis[21] gpio_inp_dis[20] gpio_inp_dis[18]
+ gpio_inp_dis[15] gpio_inp_dis[14] gpio_inp_dis[12] gpio_inp_dis[11] gpio_inp_dis[8]
+ gpio_inp_dis[4] gpio_ib_mode_sel[43] gpio_ib_mode_sel[42] gpio_ib_mode_sel[40] gpio_ib_mode_sel[39]
+ gpio_ib_mode_sel[38] gpio_ib_mode_sel[37] gpio_ib_mode_sel[36] gpio_ib_mode_sel[35]
+ gpio_ib_mode_sel[34] gpio_ib_mode_sel[33] gpio_ib_mode_sel[32] gpio_ib_mode_sel[31]
+ gpio_ib_mode_sel[30] gpio_ib_mode_sel[26] gpio_ib_mode_sel[25] gpio_ib_mode_sel[24]
+ gpio_ib_mode_sel[23] gpio_ib_mode_sel[22] gpio_ib_mode_sel[21] gpio_ib_mode_sel[20]
+ gpio_ib_mode_sel[18] gpio_ib_mode_sel[15] gpio_ib_mode_sel[14] gpio_ib_mode_sel[10]
+ gpio_ib_mode_sel[8] gpio_ib_mode_sel[7] gpio_ib_mode_sel[6] gpio_ib_mode_sel[5]
+ gpio_ib_mode_sel[4] gpio_vtrip_sel[42] gpio_vtrip_sel[41] gpio_vtrip_sel[40] gpio_vtrip_sel[37]
+ gpio_vtrip_sel[36] gpio_vtrip_sel[34] gpio_vtrip_sel[33] gpio_vtrip_sel[32] gpio_vtrip_sel[30]
+ gpio_vtrip_sel[29] gpio_vtrip_sel[19] gpio_vtrip_sel[18] gpio_vtrip_sel[17] gpio_vtrip_sel[16]
+ gpio_vtrip_sel[15] gpio_vtrip_sel[14] gpio_vtrip_sel[13] gpio_vtrip_sel[12] gpio_vtrip_sel[5]
+ gpio_vtrip_sel[4] gpio_vtrip_sel[3] gpio_vtrip_sel[2] gpio_vtrip_sel[1] gpio_vtrip_sel[0]
+ gpio_slow_sel[34] gpio_slow_sel[33] gpio_slow_sel[32] gpio_slow_sel[31] gpio_slow_sel[30]
+ gpio_slow_sel[29] gpio_slow_sel[24] gpio_slow_sel[23] gpio_slow_sel[22] gpio_slow_sel[21]
+ gpio_slow_sel[20] gpio_slow_sel[17] gpio_slow_sel[16] gpio_slow_sel[15] gpio_slow_sel[14]
+ gpio_slow_sel[13] gpio_slow_sel[12] gpio_slow_sel[11] gpio_slow_sel[10] gpio_slow_sel[9]
+ gpio_slow_sel[8] gpio_slow_sel[5] gpio_holdover[43] gpio_holdover[42] gpio_holdover[32]
+ gpio_holdover[31] gpio_holdover[29] gpio_holdover[28] gpio_holdover[27] gpio_holdover[24]
+ gpio_holdover[21] gpio_holdover[20] gpio_holdover[15] gpio_holdover[14] gpio_holdover[13]
+ gpio_holdover[12] gpio_holdover[11] gpio_holdover[10] gpio_holdover[9] gpio_holdover[8]
+ gpio_holdover[7] gpio_holdover[6] gpio_holdover[4] gpio_holdover[3] gpio_holdover[2]
+ gpio_holdover[0] gpio_analog_en[38] gpio_analog_en[37] gpio_analog_en[36] gpio_analog_en[35]
+ gpio_analog_en[34] gpio_analog_en[33] gpio_analog_en[31] gpio_analog_en[30] gpio_analog_en[26]
+ gpio_analog_en[25] gpio_analog_en[19] gpio_analog_en[17] gpio_analog_en[16] gpio_analog_en[15]
+ gpio_analog_en[14] gpio_analog_en[13] gpio_analog_en[12] gpio_analog_en[11] gpio_analog_en[10]
+ gpio_analog_en[7] gpio_analog_en[6] gpio_analog_en[5] gpio_analog_en[3] gpio_analog_en[2]
+ gpio_analog_en[1] gpio_analog_sel[36] gpio_analog_sel[35] gpio_analog_sel[34] gpio_analog_sel[33]
+ gpio_analog_sel[32] gpio_analog_sel[31] gpio_analog_sel[30] gpio_analog_sel[19]
+ gpio_analog_sel[18] gpio_analog_sel[17] gpio_analog_sel[16] gpio_analog_sel[8] gpio_analog_sel[7]
+ gpio_analog_sel[6] gpio_analog_pol[39] gpio_analog_pol[38] gpio_analog_pol[37] gpio_analog_pol[36]
+ gpio_analog_pol[32] gpio_analog_pol[31] gpio_analog_pol[30] gpio_analog_pol[27]
+ gpio_analog_pol[26] gpio_analog_pol[25] gpio_analog_pol[19] gpio_analog_pol[9] gpio_analog_pol[6]
+ gpio_analog_pol[5] gpio_analog_pol[4] gpio_analog_pol[3] gpio_analog_pol[2] gpio_dm0[43]
+ gpio_dm0[42] gpio_dm0[39] gpio_dm0[30] gpio_dm0[27] gpio_dm0[23] gpio_dm0[22] gpio_dm0[13]
+ gpio_dm0[12] gpio_dm0[10] gpio_dm0[9] gpio_dm0[8] gpio_dm0[7] gpio_dm0[6] gpio_dm0[5]
+ gpio_dm0[4] gpio_dm0[3] gpio_dm1[43] gpio_dm1[42] gpio_dm1[41] gpio_dm1[39] gpio_dm1[38]
+ gpio_dm1[29] gpio_dm1[28] gpio_dm1[27] gpio_dm1[26] gpio_dm1[25] gpio_dm1[24] gpio_dm1[23]
+ gpio_dm1[22] gpio_dm1[21] gpio_dm1[20] gpio_dm1[16] gpio_dm1[15] gpio_dm1[11] gpio_dm1[10]
+ gpio_dm1[2] gpio_dm1[1] gpio_dm1[0] gpio_dm2[39] gpio_dm2[38] gpio_dm2[37] gpio_dm2[36]
+ gpio_dm2[24] gpio_dm2[16] gpio_dm2[15] gpio_dm2[14] gpio_dm2[11] gpio_dm2[10] gpio_dm2[9]
+ gpio_dm2[8] gpio_dm2[7] gpio_dm2[6] gpio_dm2[5] gpio_dm2[4] gpio_dm2[3] gpio_dm2[2]
+ gpio_dm2[1] gpio_dm2[0] gpio_in[42] gpio_in[39] gpio_in[38] gpio_in[37] gpio_in[35]
+ gpio_in[34] gpio_in[32] gpio_in[31] gpio_in[28] gpio_in[25] gpio_in[22] gpio_in[19]
+ gpio_in[18] gpio_in[17] gpio_in[16] gpio_in[14] gpio_in[13] gpio_in[11] gpio_in[10]
+ gpio_in[9] gpio_in[7] gpio_in[4] gpio_in[1] gpio_in_h[40] gpio_in_h[39] gpio_in_h[38]
+ gpio_in_h[37] gpio_in_h[36] gpio_in_h[34] gpio_in_h[33] gpio_in_h[31] gpio_in_h[30]
+ gpio_in_h[20] gpio_in_h[19] gpio_in_h[18] gpio_in_h[17] gpio_in_h[16] gpio_in_h[15]
+ gpio_in_h[14] gpio_in_h[13] gpio_in_h[12] gpio_in_h[11] gpio_in_h[10] gpio_in_h[6]
+ gpio_in_h[3] gpio_in_h[0] gpio_loopback_zero[43] gpio_loopback_zero[42] gpio_loopback_zero[41]
+ gpio_loopback_zero[40] gpio_loopback_zero[39] gpio_loopback_zero[38] gpio_loopback_zero[37]
+ gpio_loopback_zero[36] gpio_loopback_zero[35] gpio_loopback_zero[34] gpio_loopback_zero[33]
+ gpio_loopback_zero[32] gpio_loopback_zero[31] gpio_loopback_zero[30] gpio_loopback_zero[29]
+ gpio_loopback_zero[28] gpio_loopback_zero[27] gpio_loopback_zero[26] gpio_loopback_zero[25]
+ gpio_loopback_zero[24] gpio_loopback_zero[23] gpio_loopback_zero[22] gpio_loopback_zero[21]
+ gpio_loopback_zero[20] gpio_loopback_zero[19] gpio_loopback_zero[18] gpio_loopback_zero[17]
+ gpio_loopback_zero[16] gpio_loopback_zero[15] gpio_loopback_zero[14] gpio_loopback_zero[13]
+ gpio_loopback_zero[12] gpio_loopback_zero[11] gpio_loopback_zero[10] gpio_loopback_zero[9]
+ gpio_loopback_zero[8] gpio_loopback_zero[7] gpio_loopback_zero[6] gpio_loopback_zero[5]
+ gpio_loopback_zero[4] gpio_loopback_zero[3] gpio_loopback_zero[2] gpio_loopback_zero[1]
+ gpio_loopback_zero[0] gpio_loopback_one[43] gpio_loopback_one[42] gpio_loopback_one[41]
+ gpio_loopback_one[38] gpio_loopback_one[36] gpio_loopback_one[35] gpio_loopback_one[31]
+ gpio_loopback_one[30] gpio_loopback_one[29] gpio_loopback_one[28] gpio_loopback_one[27]
+ gpio_loopback_one[26] gpio_loopback_one[25] gpio_loopback_one[24] gpio_loopback_one[22]
+ gpio_loopback_one[21] gpio_loopback_one[14] gpio_loopback_one[11] gpio_loopback_one[8]
+ gpio_loopback_one[3] analog_io[39] analog_io[36] analog_io[35] analog_io[33] analog_io[30]
+ analog_io[28] analog_io[26] analog_io[20] analog_io[19] analog_io[18] analog_io[17]
+ analog_io[15] analog_io[14] analog_io[13] analog_io[10] analog_io[7] analog_io[5]
+ analog_io[2] analog_noesd_io[43] analog_noesd_io[42] analog_noesd_io[41] analog_noesd_io[40]
+ analog_noesd_io[39] analog_noesd_io[38] analog_noesd_io[37] analog_noesd_io[34]
+ analog_noesd_io[28] analog_noesd_io[27] analog_noesd_io[26] analog_noesd_io[25]
+ analog_noesd_io[23] analog_noesd_io[22] analog_noesd_io[21] analog_noesd_io[16]
+ analog_noesd_io[12] analog_noesd_io[6] analog_noesd_io[1] analog_noesd_io[0] w_694469_865869#
+ gpio_analog_pol[20] w_23367_407274# w_694469_100152# w_23367_534874# gpio_out[0]
+ w_137274_1012253# area1_gpio_pad[11]/PAD_A_ESD_1_H sky130_ef_io__gpiov2_pad_wrapped_17/PAD_A_ESD_1_H
+ sky130_ef_io__gpiov2_pad_wrapped_2/PAD_A_ESD_1_H w_188674_1014469# w_404752_21253#
+ w_459552_23367# gpio_vtrip_sel[39] gpio_analog_pol[21] area1_gpio_pad[5]/PAD_A_ESD_1_H
+ w_485565_1014469# w_291674_1014469# w_638765_1014469# w_23367_280765# gpio_inp_dis[0]
+ analog_noesd_io[29] gpio_analog_pol[22] gpio_dm0[16] w_692253_776670# w_23367_710765#
+ w_692355_547952# gpio_analog_pol[23] w_23367_537965# area1_gpio_pad[15]/PAD_A_ESD_1_H
+ w_21151_364074# analog_noesd_io[3] w_21253_966965# gpio_out[3] gpio_in_h[41] area1_gpio_pad[9]/PAD_A_ESD_1_H
+ gpio_analog_pol[24] gpio_inp_dis[42] w_459552_21253# w_694469_145352# w_692355_593152#
+ w_485565_1012355# w_694469_951752# w_694469_190352# w_638765_1012355# gpio_vtrip_sel[6]
+ w_349952_23367# gpio_inp_dis[27] w_692355_325552# gpio_in_h[42] gpio_dm1[8] sky130_ef_io__gpiov2_pad_wrapped_5/PAD_A_ESD_1_H
+ w_189869_23367# gpio_slow_sel[36] w_694469_235552# w_21151_794074# w_692355_683352#
+ w_21253_194365# gpio_holdover[37] w_694469_280552# w_85874_1014469# sky130_ef_io__gpiov2_pad_wrapped_5/HLD_H_N
+ gpio_inp_dis[29] gpio_in_h[43] gpio_dm1[7] sky130_ef_io__gpiov2_pad_wrapped_12/PAD_A_ESD_1_H
+ gpio_out[6] w_21253_624365# w_482474_1012253# gpio_ib_mode_sel[27] gpio_holdover[33]
+ w_295152_23367# w_635674_1012253# gpio_dm2[23] w_349952_21253# w_23367_578074# analog_io[43]
+ w_692253_551270# gpio_dm1[6] w_694469_370752# area0_gpio_pad[3]/PAD_A_ESD_1_H w_189869_21253#
+ gpio_holdover[18] gpio_ib_mode_sel[29] gpio_inp_dis[24] area1_gpio_pad[3]/HLD_H_N
+ gpio_vtrip_sel[20] sky130_ef_io__gpiov2_pad_wrapped_12/HLD_H_N analog_io[23] w_21151_277674#
+ area1_gpio_pad[2]/PAD_A_ESD_1_H gpio_dm0[15] gpio_oeb[30] gpio_dm1[5] analog_noesd_io[8]
+ gpio_slow_sel[19] gpio_ib_mode_sel[28] gpio_holdover[39] w_692253_641470# sky130_ef_io__gpiov2_pad_wrapped_8/PAD_A_ESD_1_H
+ w_692253_955070# w_295152_21253# w_294765_1014469# gpio_dm0[38] sky130_ef_io__gpiov2_pad_wrapped_6/HLD_H_N
+ w_21151_707674# gpio_inp_dis[7] w_23367_234474# gpio_dm1[9] w_692355_100152# w_694469_776669#
+ gpio_analog_pol[29] w_393474_1014469# w_21151_963874# gpio_dm1[4] gpio_out[20] sky130_ef_io__gpiov2_pad_wrapped_15/PAD_A_ESD_1_H
+ gpio_inp_dis[3] area1_gpio_pad[12]/PAD_A_ESD_1_H w_692253_596470# gpio_analog_en[9]
+ analog_io[27] sky130_ef_io__gpiov2_pad_wrapped_0/PAD_A_ESD_1_H w_692253_731670#
+ gpio_loopback_one[4] w_21253_280765# area1_gpio_pad[6]/PAD_A_ESD_1_H w_692253_328870#
+ gpio_dm1[3] analog_noesd_io[31] w_23367_410365# gpio_vtrip_sel[21] gpio_oeb[33]
+ w_21253_710765# area1_gpio_pad[0]/HLD_H_N gpio_dm0[2] w_294765_1012355# w_462869_23367#
+ w_23367_237565# w_21253_537965# sky130_ef_io__gpiov2_pad_wrapped_6/TIE_LO_ESD gpio_in[2]
+ w_23367_664474# w_692253_686670# w_21151_191274# w_692253_374070# area1_gpio_pad[5]/TIE_LO_ESD
+ area1_gpio_pad[16]/PAD_A_ESD_1_H analog_noesd_io[5] gpio_in[5] w_692355_145352#
+ w_21151_621274# gpio_dm0[1] analog_noesd_io[13] area1_gpio_pad[9]/HLD_H_N gpio_analog_pol[28]
+ sky130_ef_io__gpiov2_pad_wrapped_13/HLD_H_N w_692355_951752# w_692355_190352# gpio_dm2[22]
+ gpio_analog_sel[20] gpio_analog_en[39] analog_io[4] w_694469_862552# gpio_in[8]
+ w_88965_1014469# gpio_loopback_one[12] area1_gpio_pad[0]/TIE_LO_ESD w_188674_1012253#
+ gpio_analog_sel[21] gpio_dm2[43] gpio_oeb[36] gpio_dm0[0] sky130_ef_io__gpiov2_pad_wrapped_18/PAD_A_ESD_1_H
+ gpio_loopback_one[32] w_291674_1012253# gpio_vtrip_sel[43] gpio_out[42] sky130_ef_io__gpiov2_pad_wrapped_3/PAD_A_ESD_1_H
+ w_462869_21253# w_23367_667565# analog_io[40] gpio_out[2] gpio_inp_dis[43] w_692355_235552#
+ w_694469_551269# gpio_oeb[2] gpio_vtrip_sel[22] w_23367_320874# gpio_loopback_one[37]
+ area1_gpio_pad[8]/TIE_LO_ESD gpio_analog_sel[22] area1_gpio_pad[7]/HLD_H_N w_692355_280552#
+ area0_gpio_pad[0]/PAD_A_ESD_1_H gpio_holdover[36] gpio_dm0[14] analog_noesd_io[17]
+ gpio_inp_dis[9] gpio_in[26] gpio_inp_dis[28] gpio_analog_sel[23] sky130_ef_io__gpiov2_pad_wrapped_10/PAD_A_ESD_1_H
+ gpio_out[29] gpio_out[27] gpio_ib_mode_sel[3] w_88965_1012355# gpio_dm1[14] w_692253_103470#
+ sky130_ef_io__gpiov2_pad_wrapped_13/TIE_LO_ESD w_140365_1014469# sky130_ef_io__gpiov2_pad_wrapped_10/TIE_LO_ESD
+ w_694469_641469# w_694469_955069# area1_gpio_pad[2]/TIE_LO_ESD gpio_analog_sel[24]
+ gpio_slow_sel[35] gpio_slow_sel[25] gpio_analog_en[40] analog_noesd_io[2] w_692355_370752#
+ gpio_ib_mode_sel[2] analog_noesd_io[36] w_23367_323965# gpio_dm2[27] gpio_slow_sel[1]
+ analog_io[11] w_23367_750874# area0_gpio_pad[4]/PAD_A_ESD_1_H sky130_ef_io__gpiov2_pad_wrapped_3/HLD_H_N
+ analog_io[1] gpio_analog_sel[25] gpio_oeb[5] gpio_loopback_one[0] gpio_ib_mode_sel[13]
+ gpio_out[5] gpio_loopback_one[15] w_396565_1014469# gpio_ib_mode_sel[1] gpio_oeb[19]
+ gpio_dm0[21] w_240074_1014469# analog_io[24] w_694469_596469# gpio_slow_sel[26]
+ w_23367_581165# gpio_loopback_one[5] gpio_vtrip_sel[23] gpio_analog_pol[10] gpio_in[23]
+ w_694469_731669# sky130_ef_io__gpiov2_pad_wrapped_7/HLD_H_N gpio_analog_sel[26]
+ gpio_analog_sel[5] area1_gpio_pad[3]/PAD_A_ESD_1_H gpio_inp_dis[40] sky130_ef_io__gpiov2_pad_wrapped_6/PAD_A_ESD_1_H
+ gpio_in_h[2] gpio_ib_mode_sel[0] w_21151_407274# w_186552_23367# w_517669_23367#
+ w_21151_534874# gpio_analog_pol[1] gpio_out[24] w_85874_1012253# gpio_inp_dis[6]
+ analog_noesd_io[19] gpio_analog_pol[40] gpio_in[29] w_694469_328869# w_140365_1012355#
+ gpio_analog_pol[11] gpio_inp_dis[25] gpio_analog_sel[27] gpio_slow_sel[27] sky130_ef_io__gpiov2_pad_wrapped_9/HLD_H_N
+ w_692253_148670# gpio_analog_pol[41] gpio_inp_dis[2] w_23367_753965# gpio_in[43]
+ w_694469_686669# gpio_dm2[21] gpio_analog_pol[12] gpio_holdover[40] sky130_ef_io__gpiov2_pad_wrapped_13/PAD_A_ESD_1_H
+ w_692253_193670# gpio_analog_sel[9] gpio_slow_sel[4] gpio_analog_en[41] area1_gpio_pad[13]/PAD_A_ESD_1_H
+ w_694469_374069# analog_io[9] gpio_oeb[8] w_396565_1012355# gpio_analog_en[20] analog_noesd_io[10]
+ gpio_out[8] gpio_analog_pol[42] gpio_holdover[25] gpio_analog_pol[13] area1_gpio_pad[7]/PAD_A_ESD_1_H
+ gpio_dm2[42] w_21253_410365# w_694469_638152# analog_noesd_io[33] sky130_ef_io__gpiov2_pad_wrapped_15/TIE_LO_ESD
+ gpio_inp_dis[16] gpio_in[20] w_186552_21253# gpio_in_h[5] w_517669_21253# w_21253_237565#
+ gpio_analog_pol[43] w_692253_238870# w_23367_364074# gpio_dm0[37] gpio_analog_pol[14]
+ gpio_vtrip_sel[24] gpio_out[21] sky130_ef_io__gpiov2_pad_wrapped_16/HLD_H_N analog_io[32]
+ w_692253_283870# gpio_loopback_one[18] sky130_ef_io__gpiov2_pad_wrapped_10/HLD_H_N
+ gpio_analog_sel[4] gpio_dm0[26] w_533874_1014469# gpio_loopback_one[33] gpio_vtrip_sel[28]
+ gpio_analog_pol[0] gpio_analog_pol[15] area1_gpio_pad[17]/PAD_A_ESD_1_H analog_noesd_io[7]
+ sky130_ef_io__gpiov2_pad_wrapped_9/PAD_A_ESD_1_H gpio_holdover[16] gpio_out[10]
+ gpio_dm1[37] gpio_slow_sel[28] sky130_ef_io__gpiov2_pad_wrapped_14/HLD_H_N w_694469_728352#
+ gpio_in[40] gpio_slow_sel[7] analog_noesd_io[14] w_692355_862552# gpio_dm0[36] gpio_dm1[13]
+ gpio_oeb[32] gpio_analog_sel[29] w_393474_1012253# gpio_vtrip_sel[8] w_694469_773352#
+ analog_io[6] gpio_inp_dis[35] gpio_analog_pol[16] gpio_loopback_one[10] area0_gpio_pad[0]/HLD_H_N
+ gpio_analog_en[42] gpio_slow_sel[38] w_23367_367165# sky130_ef_io__gpiov2_pad_wrapped_12/TIE_LO_ESD
+ gpio_dm2[26] w_21253_667565# gpio_analog_en[21] gpio_dm1[36] gpio_in_h[29] gpio_dm2[13]
+ sky130_ef_io__gpiov2_pad_wrapped_16/PAD_A_ESD_1_H w_23367_794074# w_694469_103469#
+ gpio_in[0] gpio_analog_pol[17] gpio_inp_dis[31] gpio_in_h[8] sky130_ef_io__gpiov2_pad_wrapped_1/PAD_A_ESD_1_H
+ gpio_in_h[21] gpio_dm0[35] w_137274_1014469# w_353269_23367# gpio_holdover[22] gpio_dm0[20]
+ area1_gpio_pad[10]/HLD_H_N analog_io[41] gpio_ib_mode_sel[17] gpio_holdover[35]
+ gpio_in[3] gpio_analog_pol[18] gpio_inp_dis[13] area0_gpio_pad[1]/PAD_A_ESD_1_H
+ sky130_ef_io__gpiov2_pad_wrapped_17/HLD_H_N analog_noesd_io[30] gpio_slow_sel[39]
+ analog_noesd_io[18] gpio_loopback_one[1] area0_gpio_pad[2]/HLD_H_N gpio_ib_mode_sel[12]
+ gpio_analog_sel[3] gpio_dm1[35] area1_gpio_pad[11]/HLD_H_N w_21151_578074# gpio_dm0[41]
+ area1_gpio_pad[4]/HLD_H_N gpio_in[6] gpio_in_h[22] gpio_dm0[34] analog_io[21] gpio_analog_en[29]
+ vccd_pad gpio_oeb[35] analog_io[29] gpio_loopback_one[6] w_243165_1014469# gpio_dm0[18]
+ gpio_out[43] area0_gpio_pad[3]/HLD_H_N gpio_out[1] area1_gpio_pad[0]/PAD_A_ESD_1_H
+ area1_gpio_pad[8]/HLD_H_N sky130_ef_io__gpiov2_pad_wrapped_0/HLD_H_N gpio_oeb[1]
+ gpio_dm2[35] area0_gpio_pad[0]/TIE_LO_ESD gpio_analog_sel[28] w_23367_797165# gpio_slow_sel[40]
+ analog_noesd_io[4] gpio_dm2[20] gpio_dm1[34] resetb_pad w_21253_323965# gpio_analog_pol[35]
+ gpio_in_h[32] gpio_in[27] gpio_inp_dis[19] gpio_in_h[23] area0_gpio_pad[4]/HLD_H_N
+ gpio_dm0[33] sky130_ef_io__gpiov2_pad_wrapped_8/TIE_LO_ESD gpio_analog_en[43] gpio_dm1[18]
+ w_353269_21253# sky130_ef_io__gpiov2_pad_wrapped_4/HLD_H_N area1_gpio_pad[13]/HLD_H_N
+ area0_gpio_pad[1]/TIE_LO_ESD analog_io[3] analog_io[12] area0_gpio_pad[5]/PAD_A_ESD_1_H
+ w_23367_277674# gpio_analog_en[22] w_694469_148669# gpio_out[28] analog_io[37] gpio_loopback_one[13]
+ gpio_dm2[41] sky130_ef_io__gpiov2_pad_wrapped_3/TIE_LO_ESD gpio_out[9] w_21253_581165#
+ gpio_dm2[34] w_694469_193669# area0_gpio_pad[5]/HLD_H_N vdda1_pad area1_gpio_pad[10]/PAD_A_ESD_1_H
+ gpio_slow_sel[41] area1_gpio_pad[14]/HLD_H_N sky130_ef_io__gpiov2_pad_wrapped_17/TIE_LO_ESD
+ sky130_ef_io__gpiov2_pad_wrapped_8/HLD_H_N analog_io[25] gpio_dm1[33] gpio_loopback_one[9]
+ w_23367_707674# gpio_dm2[18] w_21151_234474# gpio_in_h[24] gpio_dm0[32] gpio_holdover[19]
+ sky130_ef_io__gpiov2_pad_wrapped_4/PAD_A_ESD_1_H area1_gpio_pad[4]/PAD_A_ESD_1_H
+ gpio_vtrip_sel[26] sky130_ef_io__gpiov2_pad_wrapped_18/HLD_H_N vddio_pad2 gpio_inp_dis[5]
+ gpio_dm0[25] w_243165_1012355# vdda_pad w_23367_963874# gpio_analog_sel[2] gpio_out[40]
+ gpio_inp_dis[10] gpio_slow_sel[0] analog_noesd_io[20] area0_gpio_pad[3]/TIE_LO_ESD
+ area1_gpio_pad[9]/TIE_LO_ESD gpio_loopback_one[19] gpio_dm2[33] area1_gpio_pad[12]/TIE_LO_ESD
+ sky130_ef_io__gpiov2_pad_wrapped_0/TIE_LO_ESD gpio[23] gpio_oeb[4] area1_gpio_pad[6]/HLD_H_N
+ gpio_slow_sel[42] w_694469_238869# w_21253_753965# gpio_dm1[32] gpio_loopback_one[39]
+ vssd1 area0_gpio_pad[1]/HLD_H_N gpio_inp_dis[1] gpio_analog_en[27] area1_gpio_pad[10]/TIE_LO_ESD
+ gpio_loopback_one[34] w_694469_283869# gpio_in_h[35] gpio_in_h[25] area1_gpio_pad[16]/HLD_H_N
+ gpio_dm0[31] analog_io[16] gpio_loopback_one[20] vssd2 gpio_dm1[12] w_692253_865870#
+ gpio_inp_dis[41] sky130_ef_io__gpiov2_pad_wrapped_11/PAD_A_ESD_1_H gpio_in[24] gpio_oeb[9]
+ gpio_ib_mode_sel[19] gpio_in[15] area1_gpio_pad[13]/TIE_LO_ESD w_536965_1014469#
+ gpio_holdover[5] area1_gpio_pad[5]/HLD_H_N area1_gpio_pad[14]/PAD_A_ESD_1_H gpio_in_h[1]
+ gpio_analog_pol[34] w_298469_23367# w_191765_1014469# gpio_dm2[32] gpio_inp_dis[26]
+ w_694469_547952# w_482474_1014469# gpio_out[25] area1_gpio_pad[17]/HLD_H_N area0_gpio_pad[2]/TIE_LO_ESD
+ gpio_out[31] w_692355_638152# vssa2_pad gpio_slow_sel[43] analog_noesd_io[11] gpio[8]
+ gpio_analog_sel[38] w_635674_1014469# gpio_dm1[31] gpio_dm2[25] gpio_dm2[12] area1_gpio_pad[14]/TIE_LO_ESD
+ w_21151_664474# area1_gpio_pad[8]/PAD_A_ESD_1_H gpio_analog_en[23] gpio_loopback_one[17]
+ vdda2_pad gpio_holdover[1] area1_gpio_pad[3]/TIE_LO_ESD analog_noesd_io[35] area1_gpio_pad[1]/HLD_H_N
+ gpio[2] gpio_in_h[26] sky130_ef_io__gpiov2_pad_wrapped_16/TIE_LO_ESD area1_gpio_pad[1]/TIE_LO_ESD
+ sky130_ef_io__gpiov2_pad_wrapped_5/TIE_LO_ESD w_23367_191274# w_23367_966965# gpio_slow_sel[37]
+ vssd_pad gpio_holdover[41] analog_noesd_io[24] w_240074_1012253# gpio_dm0[19] gpio[40]
+ w_408069_23367# area1_gpio_pad[18]/HLD_H_N gpio_vtrip_sel[10] sky130_ef_io__gpiov2_pad_wrapped_18/TIE_LO_ESD
+ analog_io[0] gpio_analog_sel[39] gpio_out[14] sky130_ef_io__gpiov2_pad_wrapped_11/HLD_H_N
+ analog_io[34] gpio_analog_sel[10] w_694469_593152# sky130_ef_io__gpiov2_pad_wrapped_11/TIE_LO_ESD
+ gpio_in[30] gpio_slow_sel[3] gpio_dm2[31] gpio[30] w_23367_621274# gpio_slow_sel[2]
+ gpio[35] area1_gpio_pad[4]/TIE_LO_ESD gpio_holdover[26] gpio_vtrip_sel[27] gpio[3]
+ gpio_oeb[7] gpio_dm1[30] gpio[17] area1_gpio_pad[15]/HLD_H_N gpio_out[7] gpio_analog_sel[1]
+ vssd1_pad gpio_dm0[40] analog_io[38] gpio_vtrip_sel[7] gpio_ib_mode_sel[16] gpio_analog_sel[40]
+ gpio[29] gpio_dm1[19] gpio_in_h[27] gpio_dm0[29] w_692355_728352# sky130_ef_io__gpiov2_pad_wrapped_15/HLD_H_N
+ gpio_vtrip_sel[31] gpio_in[33] gpio_loopback_one[40] gpio[27] gpio_inp_dis[17] gpio_analog_sel[11]
+ sky130_ef_io__gpiov2_pad_wrapped_7/PAD_A_ESD_1_H gpio_analog_pol[8] area1_gpio_pad[16]/TIE_LO_ESD
+ area1_gpio_pad[18]/PAD_A_ESD_1_H sky130_ef_io__gpiov2_pad_wrapped_1/TIE_LO_ESD w_514352_23367#
+ sky130_ef_io__gpiov2_pad_wrapped_9/TIE_LO_ESD w_694469_325552# gpio_oeb[10] w_536965_1012355#
+ w_692355_773352# vssio_pad2 gpio_dm0[17] gpio_in[21] gpio[26] gpio_loopback_one[2]
+ w_298469_21253# gpio_inp_dis[34] gpio_in[12] w_191765_1012355# analog_noesd_io[15]
+ gpio_ib_mode_sel[11] gpio_oeb[38] gpio_in_h[4] area1_gpio_pad[15]/TIE_LO_ESD sky130_ef_io__gpiov2_pad_wrapped_4/TIE_LO_ESD
+ analog_io[8] gpio_dm2[30] gpio_in[36] sky130_ef_io__gpiov2_pad_wrapped_2/HLD_H_N
+ gpio_analog_sel[41] gpio_dm1[40] gpio_out[22] gpio_analog_sel[37] gpio_analog_sel[12]
+ gpio[18] area1_gpio_pad[17]/TIE_LO_ESD gpio[14] gpio_dm2[19] gpio[16] vccd1_pad
+ w_694469_683352# gpio_vtrip_sel[35] w_21253_367165# area0_gpio_pad[4]/TIE_LO_ESD
+ gpio_out[34] gpio_loopback_one[7] w_23367_194365# analog_noesd_io[9] gpio[39] w_21151_320874#
+ gpio_inp_dis[38] gpio_analog_pol[33] gpio_analog_en[0] gpio_in_h[9] gpio_dm0[28]
+ gpio_analog_en[18] gpio_loopback_one[23] gpio_inp_dis[30] gpio_dm1[17] vssd2_pad
+ gpio[37] gpio[38] sky130_ef_io__gpiov2_pad_wrapped_14/PAD_A_ESD_1_H gpio_holdover[17]
+ gpio[15] gpio_vtrip_sel[25] gpio_oeb[11] area1_gpio_pad[2]/HLD_H_N gpio[10] w_408069_21253#
+ gpio_analog_sel[42] gpio_analog_sel[13] area1_gpio_pad[18]/TIE_LO_ESD w_23367_624365#
+ gpio_slow_sel[18] gpio_out[11] gpio[6] vssa1_pad gpio_inp_dis[23] gpio_oeb[39] gpio_analog_en[24]
+ gpio_dm2[40] gpio_holdover[34] gpio_in[41] gpio[20] gpio_dm2[29] area1_gpio_pad[6]/TIE_LO_ESD
+ gpio_loopback_one[16] gpio_slow_sel[6] analog_io[42] gpio_out[4] area0_gpio_pad[5]/TIE_LO_ESD
+ gpio_oeb[31] sky130_ef_io__gpiov2_pad_wrapped_7/TIE_LO_ESD gpio_analog_en[4] gpio[0]
+ gpio[1] gpio[7] gpio_ib_mode_sel[41] gpio_vtrip_sel[11] gpio_dm2[17] gpio_analog_en[28]
+ gpio[43] gpio_analog_sel[43] gpio[34] gpio_vtrip_sel[38] vssa gpio_analog_sel[14]
+ gpio[19] analog_noesd_io[32] area0_gpio_pad[2]/PAD_A_ESD_1_H gpio_holdover[38] gpio[41]
+ w_514352_21253# gpio_holdover[30] w_533874_1012253# gpio_oeb[12] gpio[32] gpio_dm0[24]
+ gpio_vtrip_sel[9] gpio_dm0[11] gpio[25] gpio[33] area1_gpio_pad[11]/TIE_LO_ESD gpio_analog_sel[0]
+ gpio_oeb[40] gpio_in_h[28] sky130_ef_io__gpiov2_pad_wrapped_14/TIE_LO_ESD w_404752_23367#
+ analog_io[22] vssa1_pad2 analog_io[31] gpio[22] gpio_holdover[23] gpio_analog_en[8]
+ gpio_dm2[28] gpio_in_h[7] sky130_ef_io__gpiov2_pad_wrapped_1/HLD_H_N gpio_analog_sel[15]
+ gpio[4] vssd porb_h gpio_analog_en[32] gpio_analog_pol[7] gpio[24] vssa_pad sky130_ef_io__gpiov2_pad_wrapped_2/TIE_LO_ESD
+ gpio[11] area1_gpio_pad[7]/TIE_LO_ESD vssio area1_gpio_pad[12]/HLD_H_N gpio[31]
+ gpio[9] gpio[42] w_21253_797165# FILLER_9/VSSIO_Q gpio_out[19] gpio[5] vssa2 w_21151_750874#
+ vssa1 area1_gpio_pad[1]/PAD_A_ESD_1_H gpio[28] gpio[13] gpio[21] gpio_ib_mode_sel[9]
+ gpio[12]
Xarea1_gpio_pad[9] gpio_in_h[9] analog_noesd_io[9] analog_io[9] area1_gpio_pad[9]/PAD_A_ESD_1_H
+ gpio_dm2[9] gpio_dm1[9] gpio_dm0[9] gpio_in[9] gpio_inp_dis[9] gpio_ib_mode_sel[9]
+ porb_h porb_h area1_gpio_pad[9]/TIE_LO_ESD gpio_oeb[9] area1_gpio_pad[9]/HLD_H_N
+ area1_gpio_pad[9]/TIE_LO_ESD gpio_slow_sel[9] gpio_vtrip_sel[9] gpio_holdover[9]
+ gpio_analog_en[9] gpio_analog_sel[9] gpio_loopback_one[9] area1_gpio_pad[9]/TIE_LO_ESD
+ gpio_analog_pol[9] gpio_out[9] FILLER_9/VDDIO_Q w_694469_641469# area1_gpio_pad[9]/HLD_H_N
+ FILLER_9/VSSIO_Q w_694469_638152# vccd FILLER_9/AMUXBUS_B FILLER_9/AMUXBUS_A vssio
+ vddio vdda1 w_692355_638152# vddio vssa1 w_692253_641470# vssd gpio[9] vccd sky130_ef_io__gpiov2_pad_wrapped
Xsky130_ef_io__gpiov2_pad_wrapped_9 gpio_in_h[28] analog_noesd_io[28] analog_io[28]
+ sky130_ef_io__gpiov2_pad_wrapped_9/PAD_A_ESD_1_H gpio_dm2[28] gpio_dm1[28] gpio_dm0[28]
+ gpio_in[28] gpio_inp_dis[28] gpio_ib_mode_sel[28] porb_h porb_h sky130_ef_io__gpiov2_pad_wrapped_9/TIE_LO_ESD
+ gpio_oeb[28] sky130_ef_io__gpiov2_pad_wrapped_9/HLD_H_N sky130_ef_io__gpiov2_pad_wrapped_9/TIE_LO_ESD
+ gpio_slow_sel[28] gpio_vtrip_sel[28] gpio_holdover[28] gpio_analog_en[28] gpio_analog_sel[28]
+ gpio_loopback_one[28] sky130_ef_io__gpiov2_pad_wrapped_9/TIE_LO_ESD gpio_analog_pol[28]
+ gpio_out[28] FILLER_9/VDDIO_Q w_21151_664474# sky130_ef_io__gpiov2_pad_wrapped_9/HLD_H_N
+ FILLER_9/VSSIO_Q w_21253_667565# vccd FILLER_9/AMUXBUS_B FILLER_9/AMUXBUS_A vssio
+ vddio vdda2 w_23367_667565# vddio vssa2 w_23367_664474# vssd gpio[28] vccd sky130_ef_io__gpiov2_pad_wrapped
Xconstant_value_inst[41] vccd gpio_loopback_zero[41] gpio_loopback_one[41] vssd constant_block
Xmgmt_vccd_lvclamp_pad vdda vccd FILLER_9/AMUXBUS_B FILLER_9/AMUXBUS_A vccd_pad vccd
+ vddio vssd vssio FILLER_9/VDDIO_Q vddio vssa FILLER_9/VSSIO_Q sky130_ef_io__vccd_lvc_clamped_pad
Xconstant_value_inst[24] vccd gpio_loopback_zero[24] gpio_loopback_one[24] vssd constant_block
Xarea1_gpio_pad[8] gpio_in_h[27] analog_noesd_io[27] analog_io[27] area1_gpio_pad[8]/PAD_A_ESD_1_H
+ gpio_dm2[27] gpio_dm1[27] gpio_dm0[27] gpio_in[27] gpio_inp_dis[27] gpio_ib_mode_sel[27]
+ porb_h porb_h area1_gpio_pad[8]/TIE_LO_ESD gpio_oeb[27] area1_gpio_pad[8]/HLD_H_N
+ area1_gpio_pad[8]/TIE_LO_ESD gpio_slow_sel[27] gpio_vtrip_sel[27] gpio_holdover[27]
+ gpio_analog_en[27] gpio_analog_sel[27] gpio_loopback_one[27] area1_gpio_pad[8]/TIE_LO_ESD
+ gpio_analog_pol[27] gpio_out[27] FILLER_9/VDDIO_Q w_21151_707674# area1_gpio_pad[8]/HLD_H_N
+ FILLER_9/VSSIO_Q w_21253_710765# vccd FILLER_9/AMUXBUS_B FILLER_9/AMUXBUS_A vssio
+ vddio vdda2 w_23367_710765# vddio vssa2 w_23367_707674# vssd gpio[27] vccd sky130_ef_io__gpiov2_pad_wrapped
Xconstant_value_inst[40] vccd gpio_loopback_zero[40] gpio_loopback_one[40] vssd constant_block
Xconstant_value_inst[23] vccd gpio_loopback_zero[23] gpio_loopback_one[23] vssd constant_block
Xarea1_gpio_pad[7] gpio_in_h[26] analog_noesd_io[26] analog_io[26] area1_gpio_pad[7]/PAD_A_ESD_1_H
+ gpio_dm2[26] gpio_dm1[26] gpio_dm0[26] gpio_in[26] gpio_inp_dis[26] gpio_ib_mode_sel[26]
+ porb_h porb_h area1_gpio_pad[7]/TIE_LO_ESD gpio_oeb[26] area1_gpio_pad[7]/HLD_H_N
+ area1_gpio_pad[7]/TIE_LO_ESD gpio_slow_sel[26] gpio_vtrip_sel[26] gpio_holdover[26]
+ gpio_analog_en[26] gpio_analog_sel[26] gpio_loopback_one[26] area1_gpio_pad[7]/TIE_LO_ESD
+ gpio_analog_pol[26] gpio_out[26] FILLER_9/VDDIO_Q w_21151_750874# area1_gpio_pad[7]/HLD_H_N
+ FILLER_9/VSSIO_Q w_21253_753965# vccd FILLER_9/AMUXBUS_B FILLER_9/AMUXBUS_A vssio
+ vddio vdda2 w_23367_753965# vddio vssa2 w_23367_750874# vssd gpio[26] vccd sky130_ef_io__gpiov2_pad_wrapped
Xconstant_value_inst[22] vccd gpio_loopback_zero[22] gpio_loopback_one[22] vssd constant_block
Xarea1_gpio_pad[6] gpio_in_h[25] analog_noesd_io[25] analog_io[25] area1_gpio_pad[6]/PAD_A_ESD_1_H
+ gpio_dm2[25] gpio_dm1[25] gpio_dm0[25] gpio_in[25] gpio_inp_dis[25] gpio_ib_mode_sel[25]
+ porb_h porb_h area1_gpio_pad[6]/TIE_LO_ESD gpio_oeb[25] area1_gpio_pad[6]/HLD_H_N
+ area1_gpio_pad[6]/TIE_LO_ESD gpio_slow_sel[25] gpio_vtrip_sel[25] gpio_holdover[25]
+ gpio_analog_en[25] gpio_analog_sel[25] gpio_loopback_one[25] area1_gpio_pad[6]/TIE_LO_ESD
+ gpio_analog_pol[25] gpio_out[25] FILLER_9/VDDIO_Q w_21151_794074# area1_gpio_pad[6]/HLD_H_N
+ FILLER_9/VSSIO_Q w_21253_797165# vccd FILLER_9/AMUXBUS_B FILLER_9/AMUXBUS_A vssio
+ vddio vdda2 w_23367_797165# vddio vssa2 w_23367_794074# vssd gpio[25] vccd sky130_ef_io__gpiov2_pad_wrapped
Xconstant_value_inst[21] vccd gpio_loopback_zero[21] gpio_loopback_one[21] vssd constant_block
Xarea1_gpio_pad[5] gpio_in_h[24] analog_noesd_io[24] analog_io[24] area1_gpio_pad[5]/PAD_A_ESD_1_H
+ gpio_dm2[24] gpio_dm1[24] gpio_dm0[24] gpio_in[24] gpio_inp_dis[24] gpio_ib_mode_sel[24]
+ porb_h porb_h area1_gpio_pad[5]/TIE_LO_ESD gpio_oeb[24] area1_gpio_pad[5]/HLD_H_N
+ area1_gpio_pad[5]/TIE_LO_ESD gpio_slow_sel[24] gpio_vtrip_sel[24] gpio_holdover[24]
+ gpio_analog_en[24] gpio_analog_sel[24] gpio_loopback_one[24] area1_gpio_pad[5]/TIE_LO_ESD
+ gpio_analog_pol[24] gpio_out[24] FILLER_9/VDDIO_Q w_21151_963874# area1_gpio_pad[5]/HLD_H_N
+ FILLER_9/VSSIO_Q w_21253_966965# vccd FILLER_9/AMUXBUS_B FILLER_9/AMUXBUS_A vssio
+ vddio vdda2 w_23367_966965# vddio vssa2 w_23367_963874# vssd gpio[24] vccd sky130_ef_io__gpiov2_pad_wrapped
Xconstant_value_inst[20] vccd gpio_loopback_zero[20] gpio_loopback_one[20] vssd constant_block
Xpor vddio vccd porb_h por_l porb_l vssd vssio simple_por
Xarea0_gpio_pad[5] gpio_in_h[43] analog_noesd_io[43] analog_io[43] area0_gpio_pad[5]/PAD_A_ESD_1_H
+ gpio_dm2[43] gpio_dm1[43] gpio_dm0[43] gpio_in[43] gpio_inp_dis[43] gpio_ib_mode_sel[43]
+ porb_h porb_h area0_gpio_pad[5]/TIE_LO_ESD gpio_oeb[43] area0_gpio_pad[5]/HLD_H_N
+ area0_gpio_pad[5]/TIE_LO_ESD gpio_slow_sel[43] gpio_vtrip_sel[43] gpio_holdover[43]
+ gpio_analog_en[43] gpio_analog_sel[43] gpio_loopback_one[43] area0_gpio_pad[5]/TIE_LO_ESD
+ gpio_analog_pol[43] gpio_out[43] FILLER_9/VDDIO_Q w_517669_21253# area0_gpio_pad[5]/HLD_H_N
+ FILLER_9/VSSIO_Q w_514352_21253# vccd FILLER_9/AMUXBUS_B FILLER_9/AMUXBUS_A vssio
+ vddio vdda w_514352_23367# vddio vssa w_517669_23367# vssd gpio[43] vccd sky130_ef_io__gpiov2_pad_wrapped
Xarea1_gpio_pad[4] gpio_in_h[23] analog_noesd_io[23] analog_io[23] area1_gpio_pad[4]/PAD_A_ESD_1_H
+ gpio_dm2[23] gpio_dm1[23] gpio_dm0[23] gpio_in[23] gpio_inp_dis[23] gpio_ib_mode_sel[23]
+ porb_h porb_h area1_gpio_pad[4]/TIE_LO_ESD gpio_oeb[23] area1_gpio_pad[4]/HLD_H_N
+ area1_gpio_pad[4]/TIE_LO_ESD gpio_slow_sel[23] gpio_vtrip_sel[23] gpio_holdover[23]
+ gpio_analog_en[23] gpio_analog_sel[23] gpio_loopback_one[23] area1_gpio_pad[4]/TIE_LO_ESD
+ gpio_analog_pol[23] gpio_out[23] FILLER_9/VDDIO_Q w_85874_1014469# area1_gpio_pad[4]/HLD_H_N
+ FILLER_9/VSSIO_Q w_88965_1014469# vccd FILLER_9/AMUXBUS_B FILLER_9/AMUXBUS_A vssio
+ vddio vdda2 w_88965_1012355# vddio vssa2 w_85874_1012253# vssd gpio[23] vccd sky130_ef_io__gpiov2_pad_wrapped
Xarea1_gpio_pad[18] gpio_in_h[18] analog_noesd_io[18] analog_io[18] area1_gpio_pad[18]/PAD_A_ESD_1_H
+ gpio_dm2[18] gpio_dm1[18] gpio_dm0[18] gpio_in[18] gpio_inp_dis[18] gpio_ib_mode_sel[18]
+ porb_h porb_h area1_gpio_pad[18]/TIE_LO_ESD gpio_oeb[18] area1_gpio_pad[18]/HLD_H_N
+ area1_gpio_pad[18]/TIE_LO_ESD gpio_slow_sel[18] gpio_vtrip_sel[18] gpio_holdover[18]
+ gpio_analog_en[18] gpio_analog_sel[18] gpio_loopback_one[18] area1_gpio_pad[18]/TIE_LO_ESD
+ gpio_analog_pol[18] gpio_out[18] FILLER_9/VDDIO_Q w_393474_1014469# area1_gpio_pad[18]/HLD_H_N
+ FILLER_9/VSSIO_Q w_396565_1014469# vccd FILLER_9/AMUXBUS_B FILLER_9/AMUXBUS_A vssio
+ vddio vdda1 w_396565_1012355# vddio vssa1 w_393474_1012253# vssd gpio[18] vccd sky130_ef_io__gpiov2_pad_wrapped
Xarea0_gpio_pad[4] gpio_in_h[42] analog_noesd_io[42] analog_io[42] area0_gpio_pad[4]/PAD_A_ESD_1_H
+ gpio_dm2[42] gpio_dm1[42] gpio_dm0[42] gpio_in[42] gpio_inp_dis[42] gpio_ib_mode_sel[42]
+ porb_h porb_h area0_gpio_pad[4]/TIE_LO_ESD gpio_oeb[42] area0_gpio_pad[4]/HLD_H_N
+ area0_gpio_pad[4]/TIE_LO_ESD gpio_slow_sel[42] gpio_vtrip_sel[42] gpio_holdover[42]
+ gpio_analog_en[42] gpio_analog_sel[42] gpio_loopback_one[42] area0_gpio_pad[4]/TIE_LO_ESD
+ gpio_analog_pol[42] gpio_out[42] FILLER_9/VDDIO_Q w_462869_21253# area0_gpio_pad[4]/HLD_H_N
+ FILLER_9/VSSIO_Q w_459552_21253# vccd FILLER_9/AMUXBUS_B FILLER_9/AMUXBUS_A vssio
+ vddio vdda w_459552_23367# vddio vssa w_462869_23367# vssd gpio[42] vccd sky130_ef_io__gpiov2_pad_wrapped
Xmgmt_vddio_hvclamp_pad\[0\] vdda FILLER_9/VSSIO_Q vddio FILLER_9/VDDIO_Q vssd vddio_pad
+ vssa FILLER_9/AMUXBUS_B FILLER_9/AMUXBUS_A vddio vccd vssio vccd sky130_ef_io__vddio_hvc_clamped_pad
Xarea1_gpio_pad[3] gpio_in_h[22] analog_noesd_io[22] analog_io[22] area1_gpio_pad[3]/PAD_A_ESD_1_H
+ gpio_dm2[22] gpio_dm1[22] gpio_dm0[22] gpio_in[22] gpio_inp_dis[22] gpio_ib_mode_sel[22]
+ porb_h porb_h area1_gpio_pad[3]/TIE_LO_ESD gpio_oeb[22] area1_gpio_pad[3]/HLD_H_N
+ area1_gpio_pad[3]/TIE_LO_ESD gpio_slow_sel[22] gpio_vtrip_sel[22] gpio_holdover[22]
+ gpio_analog_en[22] gpio_analog_sel[22] gpio_loopback_one[22] area1_gpio_pad[3]/TIE_LO_ESD
+ gpio_analog_pol[22] gpio_out[22] FILLER_9/VDDIO_Q w_137274_1014469# area1_gpio_pad[3]/HLD_H_N
+ FILLER_9/VSSIO_Q w_140365_1014469# vccd FILLER_9/AMUXBUS_B FILLER_9/AMUXBUS_A vssio
+ vddio vdda2 w_140365_1012355# vddio vssa2 w_137274_1012253# vssd gpio[22] vccd sky130_ef_io__gpiov2_pad_wrapped
Xarea1_gpio_pad[17] gpio_in_h[17] analog_noesd_io[17] analog_io[17] area1_gpio_pad[17]/PAD_A_ESD_1_H
+ gpio_dm2[17] gpio_dm1[17] gpio_dm0[17] gpio_in[17] gpio_inp_dis[17] gpio_ib_mode_sel[17]
+ porb_h porb_h area1_gpio_pad[17]/TIE_LO_ESD gpio_oeb[17] area1_gpio_pad[17]/HLD_H_N
+ area1_gpio_pad[17]/TIE_LO_ESD gpio_slow_sel[17] gpio_vtrip_sel[17] gpio_holdover[17]
+ gpio_analog_en[17] gpio_analog_sel[17] gpio_loopback_one[17] area1_gpio_pad[17]/TIE_LO_ESD
+ gpio_analog_pol[17] gpio_out[17] FILLER_9/VDDIO_Q w_482474_1014469# area1_gpio_pad[17]/HLD_H_N
+ FILLER_9/VSSIO_Q w_485565_1014469# vccd FILLER_9/AMUXBUS_B FILLER_9/AMUXBUS_A vssio
+ vddio vdda1 w_485565_1012355# vddio vssa1 w_482474_1012253# vssd gpio[17] vccd sky130_ef_io__gpiov2_pad_wrapped
Xmgmt_vssio_hvclamp_pad\[1\] vdda2 vssd vssa2 FILLER_9/AMUXBUS_B FILLER_9/AMUXBUS_A
+ vssio_pad2 FILLER_9/VDDIO_Q vddio vssio FILLER_9/VSSIO_Q vddio vccd vccd sky130_ef_io__vssio_hvc_clamped_pad
Xarea0_gpio_pad[3] gpio_in_h[41] analog_noesd_io[41] analog_io[41] area0_gpio_pad[3]/PAD_A_ESD_1_H
+ gpio_dm2[41] gpio_dm1[41] gpio_dm0[41] gpio_in[41] gpio_inp_dis[41] gpio_ib_mode_sel[41]
+ porb_h porb_h area0_gpio_pad[3]/TIE_LO_ESD gpio_oeb[41] area0_gpio_pad[3]/HLD_H_N
+ area0_gpio_pad[3]/TIE_LO_ESD gpio_slow_sel[41] gpio_vtrip_sel[41] gpio_holdover[41]
+ gpio_analog_en[41] gpio_analog_sel[41] gpio_loopback_one[41] area0_gpio_pad[3]/TIE_LO_ESD
+ gpio_analog_pol[41] gpio_out[41] FILLER_9/VDDIO_Q w_408069_21253# area0_gpio_pad[3]/HLD_H_N
+ FILLER_9/VSSIO_Q w_404752_21253# vccd FILLER_9/AMUXBUS_B FILLER_9/AMUXBUS_A vssio
+ vddio vdda w_404752_23367# vddio vssa w_408069_23367# vssd gpio[41] vccd sky130_ef_io__gpiov2_pad_wrapped
Xarea1_gpio_pad[2] gpio_in_h[21] analog_noesd_io[21] analog_io[21] area1_gpio_pad[2]/PAD_A_ESD_1_H
+ gpio_dm2[21] gpio_dm1[21] gpio_dm0[21] gpio_in[21] gpio_inp_dis[21] gpio_ib_mode_sel[21]
+ porb_h porb_h area1_gpio_pad[2]/TIE_LO_ESD gpio_oeb[21] area1_gpio_pad[2]/HLD_H_N
+ area1_gpio_pad[2]/TIE_LO_ESD gpio_slow_sel[21] gpio_vtrip_sel[21] gpio_holdover[21]
+ gpio_analog_en[21] gpio_analog_sel[21] gpio_loopback_one[21] area1_gpio_pad[2]/TIE_LO_ESD
+ gpio_analog_pol[21] gpio_out[21] FILLER_9/VDDIO_Q w_188674_1014469# area1_gpio_pad[2]/HLD_H_N
+ FILLER_9/VSSIO_Q w_191765_1014469# vccd FILLER_9/AMUXBUS_B FILLER_9/AMUXBUS_A vssio
+ vddio vdda2 w_191765_1012355# vddio vssa2 w_188674_1012253# vssd gpio[21] vccd sky130_ef_io__gpiov2_pad_wrapped
Xarea1_gpio_pad[16] gpio_in_h[16] analog_noesd_io[16] analog_io[16] area1_gpio_pad[16]/PAD_A_ESD_1_H
+ gpio_dm2[16] gpio_dm1[16] gpio_dm0[16] gpio_in[16] gpio_inp_dis[16] gpio_ib_mode_sel[16]
+ porb_h porb_h area1_gpio_pad[16]/TIE_LO_ESD gpio_oeb[16] area1_gpio_pad[16]/HLD_H_N
+ area1_gpio_pad[16]/TIE_LO_ESD gpio_slow_sel[16] gpio_vtrip_sel[16] gpio_holdover[16]
+ gpio_analog_en[16] gpio_analog_sel[16] gpio_loopback_one[16] area1_gpio_pad[16]/TIE_LO_ESD
+ gpio_analog_pol[16] gpio_out[16] FILLER_9/VDDIO_Q w_533874_1014469# area1_gpio_pad[16]/HLD_H_N
+ FILLER_9/VSSIO_Q w_536965_1014469# vccd FILLER_9/AMUXBUS_B FILLER_9/AMUXBUS_A vssio
+ vddio vdda1 w_536965_1012355# vddio vssa1 w_533874_1012253# vssd gpio[16] vccd sky130_ef_io__gpiov2_pad_wrapped
Xarea0_gpio_pad[2] gpio_in_h[40] analog_noesd_io[40] analog_io[40] area0_gpio_pad[2]/PAD_A_ESD_1_H
+ gpio_dm2[40] gpio_dm1[40] gpio_dm0[40] gpio_in[40] gpio_inp_dis[40] gpio_ib_mode_sel[40]
+ porb_h porb_h area0_gpio_pad[2]/TIE_LO_ESD gpio_oeb[40] area0_gpio_pad[2]/HLD_H_N
+ area0_gpio_pad[2]/TIE_LO_ESD gpio_slow_sel[40] gpio_vtrip_sel[40] gpio_holdover[40]
+ gpio_analog_en[40] gpio_analog_sel[40] gpio_loopback_one[40] area0_gpio_pad[2]/TIE_LO_ESD
+ gpio_analog_pol[40] gpio_out[40] FILLER_9/VDDIO_Q w_353269_21253# area0_gpio_pad[2]/HLD_H_N
+ FILLER_9/VSSIO_Q w_349952_21253# vccd FILLER_9/AMUXBUS_B FILLER_9/AMUXBUS_A vssio
+ vddio vdda w_349952_23367# vddio vssa w_353269_23367# vssd gpio[40] vccd sky130_ef_io__gpiov2_pad_wrapped
Xarea1_gpio_pad[1] gpio_in_h[20] analog_noesd_io[20] analog_io[20] area1_gpio_pad[1]/PAD_A_ESD_1_H
+ gpio_dm2[20] gpio_dm1[20] gpio_dm0[20] gpio_in[20] gpio_inp_dis[20] gpio_ib_mode_sel[20]
+ porb_h porb_h area1_gpio_pad[1]/TIE_LO_ESD gpio_oeb[20] area1_gpio_pad[1]/HLD_H_N
+ area1_gpio_pad[1]/TIE_LO_ESD gpio_slow_sel[20] gpio_vtrip_sel[20] gpio_holdover[20]
+ gpio_analog_en[20] gpio_analog_sel[20] gpio_loopback_one[20] area1_gpio_pad[1]/TIE_LO_ESD
+ gpio_analog_pol[20] gpio_out[20] FILLER_9/VDDIO_Q w_240074_1014469# area1_gpio_pad[1]/HLD_H_N
+ FILLER_9/VSSIO_Q w_243165_1014469# vccd FILLER_9/AMUXBUS_B FILLER_9/AMUXBUS_A vssio
+ vddio vdda2 w_243165_1012355# vddio vssa2 w_240074_1012253# vssd gpio[20] vccd sky130_ef_io__gpiov2_pad_wrapped
Xarea1_gpio_pad[15] gpio_in_h[15] analog_noesd_io[15] analog_io[15] area1_gpio_pad[15]/PAD_A_ESD_1_H
+ gpio_dm2[15] gpio_dm1[15] gpio_dm0[15] gpio_in[15] gpio_inp_dis[15] gpio_ib_mode_sel[15]
+ porb_h porb_h area1_gpio_pad[15]/TIE_LO_ESD gpio_oeb[15] area1_gpio_pad[15]/HLD_H_N
+ area1_gpio_pad[15]/TIE_LO_ESD gpio_slow_sel[15] gpio_vtrip_sel[15] gpio_holdover[15]
+ gpio_analog_en[15] gpio_analog_sel[15] gpio_loopback_one[15] area1_gpio_pad[15]/TIE_LO_ESD
+ gpio_analog_pol[15] gpio_out[15] FILLER_9/VDDIO_Q w_635674_1014469# area1_gpio_pad[15]/HLD_H_N
+ FILLER_9/VSSIO_Q w_638765_1014469# vccd FILLER_9/AMUXBUS_B FILLER_9/AMUXBUS_A vssio
+ vddio vdda1 w_638765_1012355# vddio vssa1 w_635674_1012253# vssd gpio[15] vccd sky130_ef_io__gpiov2_pad_wrapped
Xuser2_vdda_hvclamp_pad FILLER_9/VDDIO_Q FILLER_9/VSSIO_Q vssio vdda2_pad FILLER_9/AMUXBUS_B
+ FILLER_9/AMUXBUS_A vdda2 vccd vssd vssa2 vddio vccd vddio sky130_ef_io__vdda_hvc_clamped_pad
Xarea0_gpio_pad[1] gpio_in_h[39] analog_noesd_io[39] analog_io[39] area0_gpio_pad[1]/PAD_A_ESD_1_H
+ gpio_dm2[39] gpio_dm1[39] gpio_dm0[39] gpio_in[39] gpio_inp_dis[39] gpio_ib_mode_sel[39]
+ porb_h porb_h area0_gpio_pad[1]/TIE_LO_ESD gpio_oeb[39] area0_gpio_pad[1]/HLD_H_N
+ area0_gpio_pad[1]/TIE_LO_ESD gpio_slow_sel[39] gpio_vtrip_sel[39] gpio_holdover[39]
+ gpio_analog_en[39] gpio_analog_sel[39] gpio_loopback_one[39] area0_gpio_pad[1]/TIE_LO_ESD
+ gpio_analog_pol[39] gpio_out[39] FILLER_9/VDDIO_Q w_298469_21253# area0_gpio_pad[1]/HLD_H_N
+ FILLER_9/VSSIO_Q w_295152_21253# vccd FILLER_9/AMUXBUS_B FILLER_9/AMUXBUS_A vssio
+ vddio vdda w_295152_23367# vddio vssa w_298469_23367# vssd gpio[39] vccd sky130_ef_io__gpiov2_pad_wrapped
Xarea1_gpio_pad[0] gpio_in_h[19] analog_noesd_io[19] analog_io[19] area1_gpio_pad[0]/PAD_A_ESD_1_H
+ gpio_dm2[19] gpio_dm1[19] gpio_dm0[19] gpio_in[19] gpio_inp_dis[19] gpio_ib_mode_sel[19]
+ porb_h porb_h area1_gpio_pad[0]/TIE_LO_ESD gpio_oeb[19] area1_gpio_pad[0]/HLD_H_N
+ area1_gpio_pad[0]/TIE_LO_ESD gpio_slow_sel[19] gpio_vtrip_sel[19] gpio_holdover[19]
+ gpio_analog_en[19] gpio_analog_sel[19] gpio_loopback_one[19] area1_gpio_pad[0]/TIE_LO_ESD
+ gpio_analog_pol[19] gpio_out[19] FILLER_9/VDDIO_Q w_291674_1014469# area1_gpio_pad[0]/HLD_H_N
+ FILLER_9/VSSIO_Q w_294765_1014469# vccd FILLER_9/AMUXBUS_B FILLER_9/AMUXBUS_A vssio
+ vddio vdda2 w_294765_1012355# vddio vssa2 w_291674_1012253# vssd gpio[19] vccd sky130_ef_io__gpiov2_pad_wrapped
Xarea1_gpio_pad[14] gpio_in_h[14] analog_noesd_io[14] analog_io[14] area1_gpio_pad[14]/PAD_A_ESD_1_H
+ gpio_dm2[14] gpio_dm1[14] gpio_dm0[14] gpio_in[14] gpio_inp_dis[14] gpio_ib_mode_sel[14]
+ porb_h porb_h area1_gpio_pad[14]/TIE_LO_ESD gpio_oeb[14] area1_gpio_pad[14]/HLD_H_N
+ area1_gpio_pad[14]/TIE_LO_ESD gpio_slow_sel[14] gpio_vtrip_sel[14] gpio_holdover[14]
+ gpio_analog_en[14] gpio_analog_sel[14] gpio_loopback_one[14] area1_gpio_pad[14]/TIE_LO_ESD
+ gpio_analog_pol[14] gpio_out[14] FILLER_9/VDDIO_Q w_694469_955069# area1_gpio_pad[14]/HLD_H_N
+ FILLER_9/VSSIO_Q w_694469_951752# vccd FILLER_9/AMUXBUS_B FILLER_9/AMUXBUS_A vssio
+ vddio vdda1 w_692355_951752# vddio vssa1 w_692253_955070# vssd gpio[14] vccd sky130_ef_io__gpiov2_pad_wrapped
Xarea0_gpio_pad[0] gpio_in_h[38] analog_noesd_io[38] analog_io[38] area0_gpio_pad[0]/PAD_A_ESD_1_H
+ gpio_dm2[38] gpio_dm0[38] gpio_dm1[38] gpio_in[38] gpio_inp_dis[38] gpio_ib_mode_sel[38]
+ porb_h porb_h area0_gpio_pad[0]/TIE_LO_ESD gpio_oeb[38] area0_gpio_pad[0]/HLD_H_N
+ area0_gpio_pad[0]/TIE_LO_ESD gpio_slow_sel[38] gpio_vtrip_sel[38] gpio_holdover[38]
+ gpio_analog_en[38] gpio_analog_sel[38] gpio_loopback_one[38] area0_gpio_pad[0]/TIE_LO_ESD
+ gpio_analog_pol[38] gpio_out[38] FILLER_9/VDDIO_Q w_189869_21253# area0_gpio_pad[0]/HLD_H_N
+ FILLER_9/VSSIO_Q w_186552_21253# vccd FILLER_9/AMUXBUS_B FILLER_9/AMUXBUS_A vssio
+ vddio vdda w_186552_23367# vddio vssa w_189869_23367# vssd gpio[38] vccd sky130_ef_io__gpiov2_pad_wrapped
Xconstant_value_xres_inst vccd constant_value_xres_inst/zero constant_value_xres_inst/one
+ vssd constant_block
Xarea1_gpio_pad[13] gpio_in_h[13] analog_noesd_io[13] analog_io[13] area1_gpio_pad[13]/PAD_A_ESD_1_H
+ gpio_dm2[13] gpio_dm1[13] gpio_dm0[13] gpio_in[13] gpio_inp_dis[13] gpio_ib_mode_sel[13]
+ porb_h porb_h area1_gpio_pad[13]/TIE_LO_ESD gpio_oeb[13] area1_gpio_pad[13]/HLD_H_N
+ area1_gpio_pad[13]/TIE_LO_ESD gpio_slow_sel[13] gpio_vtrip_sel[13] gpio_holdover[13]
+ gpio_analog_en[13] gpio_analog_sel[13] gpio_loopback_one[13] area1_gpio_pad[13]/TIE_LO_ESD
+ gpio_analog_pol[13] gpio_out[13] FILLER_9/VDDIO_Q w_694469_865869# area1_gpio_pad[13]/HLD_H_N
+ FILLER_9/VSSIO_Q w_694469_862552# vccd FILLER_9/AMUXBUS_B FILLER_9/AMUXBUS_A vssio
+ vddio vdda1 w_692355_862552# vddio vssa1 w_692253_865870# vssd gpio[13] vccd sky130_ef_io__gpiov2_pad_wrapped
Xuser1_vssd_lvclamp_pad vdda1 FILLER_9/VSSIO_Q vssd1 vccd vssd FILLER_9/AMUXBUS_B
+ FILLER_9/AMUXBUS_A vssa1 vssd1_pad vddio vccd vddio FILLER_9/VDDIO_Q vssio vccd1
+ sky130_ef_io__vssd_lvc_clamped3_pad
Xarea1_gpio_pad[12] gpio_in_h[12] analog_noesd_io[12] analog_io[12] area1_gpio_pad[12]/PAD_A_ESD_1_H
+ gpio_dm2[12] gpio_dm1[12] gpio_dm0[12] gpio_in[12] gpio_inp_dis[12] gpio_ib_mode_sel[12]
+ porb_h porb_h area1_gpio_pad[12]/TIE_LO_ESD gpio_oeb[12] area1_gpio_pad[12]/HLD_H_N
+ area1_gpio_pad[12]/TIE_LO_ESD gpio_slow_sel[12] gpio_vtrip_sel[12] gpio_holdover[12]
+ gpio_analog_en[12] gpio_analog_sel[12] gpio_loopback_one[12] area1_gpio_pad[12]/TIE_LO_ESD
+ gpio_analog_pol[12] gpio_out[12] FILLER_9/VDDIO_Q w_694469_776669# area1_gpio_pad[12]/HLD_H_N
+ FILLER_9/VSSIO_Q w_694469_773352# vccd FILLER_9/AMUXBUS_B FILLER_9/AMUXBUS_A vssio
+ vddio vdda1 w_692355_773352# vddio vssa1 w_692253_776670# vssd gpio[12] vccd sky130_ef_io__gpiov2_pad_wrapped
Xconstant_value_inst[39] vccd gpio_loopback_zero[39] gpio_loopback_one[39] vssd constant_block
Xuser_id_value mask_rev[0] mask_rev[10] mask_rev[11] mask_rev[12] mask_rev[14] mask_rev[15]
+ mask_rev[16] mask_rev[17] mask_rev[18] mask_rev[19] mask_rev[1] mask_rev[20] mask_rev[21]
+ mask_rev[22] mask_rev[23] mask_rev[24] mask_rev[25] mask_rev[26] mask_rev[27] mask_rev[29]
+ mask_rev[2] mask_rev[30] mask_rev[31] mask_rev[3] mask_rev[4] mask_rev[5] mask_rev[6]
+ mask_rev[7] mask_rev[8] mask_rev[9] mask_rev[28] mask_rev[13] vccd vssd user_id_programming
Xarea1_gpio_pad[11] gpio_in_h[11] analog_noesd_io[11] analog_io[11] area1_gpio_pad[11]/PAD_A_ESD_1_H
+ gpio_dm2[11] gpio_dm1[11] gpio_dm0[11] gpio_in[11] gpio_inp_dis[11] gpio_ib_mode_sel[11]
+ porb_h porb_h area1_gpio_pad[11]/TIE_LO_ESD gpio_oeb[11] area1_gpio_pad[11]/HLD_H_N
+ area1_gpio_pad[11]/TIE_LO_ESD gpio_slow_sel[11] gpio_vtrip_sel[11] gpio_holdover[11]
+ gpio_analog_en[11] gpio_analog_sel[11] gpio_loopback_one[11] area1_gpio_pad[11]/TIE_LO_ESD
+ gpio_analog_pol[11] gpio_out[11] FILLER_9/VDDIO_Q w_694469_731669# area1_gpio_pad[11]/HLD_H_N
+ FILLER_9/VSSIO_Q w_694469_728352# vccd FILLER_9/AMUXBUS_B FILLER_9/AMUXBUS_A vssio
+ vddio vdda1 w_692355_728352# vddio vssa1 w_692253_731670# vssd gpio[11] vccd sky130_ef_io__gpiov2_pad_wrapped
Xuser1_vdda_hvclamp_pad\[0\] FILLER_9/VDDIO_Q FILLER_9/VSSIO_Q vssio vdda1_pad FILLER_9/AMUXBUS_B
+ FILLER_9/AMUXBUS_A vdda1 vccd vssd vssa1 vddio vccd vddio sky130_ef_io__vdda_hvc_clamped_pad
Xmgmt_vssd_lvclamp_pad vdda vssd_pad vccd vddio vddio FILLER_9/VDDIO_Q FILLER_9/AMUXBUS_B
+ FILLER_9/AMUXBUS_A vssd vssio FILLER_9/VSSIO_Q vccd vssa sky130_ef_io__vssd_lvc_clamped_pad
Xconstant_value_inst[38] vccd gpio_loopback_zero[38] gpio_loopback_one[38] vssd constant_block
Xuser2_vccd_lvclamp_pad vdda2 vccd vssd2 vddio vddio FILLER_9/AMUXBUS_B vssio FILLER_9/AMUXBUS_A
+ vccd vccd2_pad vccd2 vssd FILLER_9/VDDIO_Q vssa2 FILLER_9/VSSIO_Q sky130_ef_io__vccd_lvc_clamped3_pad
Xarea1_gpio_pad[10] gpio_in_h[10] analog_noesd_io[10] analog_io[10] area1_gpio_pad[10]/PAD_A_ESD_1_H
+ gpio_dm2[10] gpio_dm1[10] gpio_dm0[10] gpio_in[10] gpio_inp_dis[10] gpio_ib_mode_sel[10]
+ porb_h porb_h area1_gpio_pad[10]/TIE_LO_ESD gpio_oeb[10] area1_gpio_pad[10]/HLD_H_N
+ area1_gpio_pad[10]/TIE_LO_ESD gpio_slow_sel[10] gpio_vtrip_sel[10] gpio_holdover[10]
+ gpio_analog_en[10] gpio_analog_sel[10] gpio_loopback_one[10] area1_gpio_pad[10]/TIE_LO_ESD
+ gpio_analog_pol[10] gpio_out[10] FILLER_9/VDDIO_Q w_694469_686669# area1_gpio_pad[10]/HLD_H_N
+ FILLER_9/VSSIO_Q w_694469_683352# vccd FILLER_9/AMUXBUS_B FILLER_9/AMUXBUS_A vssio
+ vddio vdda1 w_692355_683352# vddio vssa1 w_692253_686670# vssd gpio[10] vccd sky130_ef_io__gpiov2_pad_wrapped
Xxres_buf_0 resetb_h resetb_l vccd vssd vddio vssio xres_buf
Xconstant_value_inst[37] vccd gpio_loopback_zero[37] gpio_loopback_one[37] vssd constant_block
Xmgmt_vssa_hvclamp_pad vssd vssa vddio vssa_pad vccd vddio vssio FILLER_9/VDDIO_Q
+ vdda FILLER_9/VSSIO_Q vccd FILLER_9/AMUXBUS_B FILLER_9/AMUXBUS_A sky130_ef_io__vssa_hvc_clamped_pad
Xuser1_vssa_hvclamp_pad\[1\] vssd vssa1 vddio vssa1_pad2 vccd vddio vssio FILLER_9/VDDIO_Q
+ vdda1 FILLER_9/VSSIO_Q vccd FILLER_9/AMUXBUS_B FILLER_9/AMUXBUS_A sky130_ef_io__vssa_hvc_clamped_pad
Xconstant_value_inst[36] vccd gpio_loopback_zero[36] gpio_loopback_one[36] vssd constant_block
Xconstant_value_inst[19] vccd gpio_loopback_zero[19] gpio_loopback_one[19] vssd constant_block
Xconstant_value_inst[35] vccd gpio_loopback_zero[35] gpio_loopback_one[35] vssd constant_block
Xconstant_value_inst[18] vccd gpio_loopback_zero[18] gpio_loopback_one[18] vssd constant_block
Xconstant_value_inst[34] vccd gpio_loopback_zero[34] gpio_loopback_one[34] vssd constant_block
Xconstant_value_inst[17] vccd gpio_loopback_zero[17] gpio_loopback_one[17] vssd constant_block
Xconstant_value_inst[33] vccd gpio_loopback_zero[33] gpio_loopback_one[33] vssd constant_block
Xconstant_value_inst[16] vccd gpio_loopback_zero[16] gpio_loopback_one[16] vssd constant_block
Xconstant_value_inst[32] vccd gpio_loopback_zero[32] gpio_loopback_one[32] vssd constant_block
Xconstant_value_inst[15] vccd gpio_loopback_zero[15] gpio_loopback_one[15] vssd constant_block
Xconstant_value_inst[31] vccd gpio_loopback_zero[31] gpio_loopback_one[31] vssd constant_block
Xconstant_value_inst[14] vccd gpio_loopback_zero[14] gpio_loopback_one[14] vssd constant_block
Xconstant_value_inst[9] vccd gpio_loopback_zero[9] gpio_loopback_one[9] vssd constant_block
Xconstant_value_inst[30] vccd gpio_loopback_zero[30] gpio_loopback_one[30] vssd constant_block
Xconstant_value_inst[13] vccd gpio_loopback_zero[13] gpio_loopback_one[13] vssd constant_block
Xconstant_value_inst[8] vccd gpio_loopback_zero[8] gpio_loopback_one[8] vssd constant_block
Xconstant_value_inst[12] vccd gpio_loopback_zero[12] gpio_loopback_one[12] vssd constant_block
Xconstant_value_inst[7] vccd gpio_loopback_zero[7] gpio_loopback_one[7] vssd constant_block
Xmgmt_vddio_hvclamp_pad\[1\] vdda2 FILLER_9/VSSIO_Q vddio FILLER_9/VDDIO_Q vssd vddio_pad2
+ vssa2 FILLER_9/AMUXBUS_B FILLER_9/AMUXBUS_A vddio vccd vssio vccd sky130_ef_io__vddio_hvc_clamped_pad
Xconstant_value_inst[11] vccd gpio_loopback_zero[11] gpio_loopback_one[11] vssd constant_block
Xconstant_value_inst[6] vccd gpio_loopback_zero[6] gpio_loopback_one[6] vssd constant_block
Xconstant_value_inst[10] vccd gpio_loopback_zero[10] gpio_loopback_one[10] vssd constant_block
Xconstant_value_inst[5] vccd gpio_loopback_zero[5] gpio_loopback_one[5] vssd constant_block
Xsky130_ef_io__gpiov2_pad_wrapped_10 gpio_in_h[8] analog_noesd_io[8] analog_io[8]
+ sky130_ef_io__gpiov2_pad_wrapped_10/PAD_A_ESD_1_H gpio_dm2[8] gpio_dm1[8] gpio_dm0[8]
+ gpio_in[8] gpio_inp_dis[8] gpio_ib_mode_sel[8] porb_h porb_h sky130_ef_io__gpiov2_pad_wrapped_10/TIE_LO_ESD
+ gpio_oeb[8] sky130_ef_io__gpiov2_pad_wrapped_10/HLD_H_N sky130_ef_io__gpiov2_pad_wrapped_10/TIE_LO_ESD
+ gpio_slow_sel[8] gpio_vtrip_sel[8] gpio_holdover[8] gpio_analog_en[8] gpio_analog_sel[8]
+ gpio_loopback_one[8] sky130_ef_io__gpiov2_pad_wrapped_10/TIE_LO_ESD gpio_analog_pol[8]
+ gpio_out[8] FILLER_9/VDDIO_Q w_694469_596469# sky130_ef_io__gpiov2_pad_wrapped_10/HLD_H_N
+ FILLER_9/VSSIO_Q w_694469_593152# vccd FILLER_9/AMUXBUS_B FILLER_9/AMUXBUS_A vssio
+ vddio vdda1 w_692355_593152# vddio vssa1 w_692253_596470# vssd gpio[8] vccd sky130_ef_io__gpiov2_pad_wrapped
Xconstant_value_inst[4] vccd gpio_loopback_zero[4] gpio_loopback_one[4] vssd constant_block
Xsky130_ef_io__gpiov2_pad_wrapped_11 gpio_in_h[7] analog_noesd_io[7] analog_io[7]
+ sky130_ef_io__gpiov2_pad_wrapped_11/PAD_A_ESD_1_H gpio_dm2[7] gpio_dm1[7] gpio_dm0[7]
+ gpio_in[7] gpio_inp_dis[7] gpio_ib_mode_sel[7] porb_h porb_h sky130_ef_io__gpiov2_pad_wrapped_11/TIE_LO_ESD
+ gpio_oeb[7] sky130_ef_io__gpiov2_pad_wrapped_11/HLD_H_N sky130_ef_io__gpiov2_pad_wrapped_11/TIE_LO_ESD
+ gpio_slow_sel[7] gpio_vtrip_sel[7] gpio_holdover[7] gpio_analog_en[7] gpio_analog_sel[7]
+ gpio_loopback_one[7] sky130_ef_io__gpiov2_pad_wrapped_11/TIE_LO_ESD gpio_analog_pol[7]
+ gpio_out[7] FILLER_9/VDDIO_Q w_694469_551269# sky130_ef_io__gpiov2_pad_wrapped_11/HLD_H_N
+ FILLER_9/VSSIO_Q w_694469_547952# vccd FILLER_9/AMUXBUS_B FILLER_9/AMUXBUS_A vssio
+ vddio vdda1 w_692355_547952# vddio vssa1 w_692253_551270# vssd gpio[7] vccd sky130_ef_io__gpiov2_pad_wrapped
Xuser2_vssd_lvclamp_pad vdda2 FILLER_9/VSSIO_Q vssd2 vccd vssd FILLER_9/AMUXBUS_B
+ FILLER_9/AMUXBUS_A vssa2 vssd2_pad vddio vccd vddio FILLER_9/VDDIO_Q vssio vccd2
+ sky130_ef_io__vssd_lvc_clamped3_pad
Xconstant_value_inst[3] vccd gpio_loopback_zero[3] gpio_loopback_one[3] vssd constant_block
Xmgmt_vssio_hvclamp_pad\[0\] vdda vssd vssa FILLER_9/AMUXBUS_B FILLER_9/AMUXBUS_A
+ vssio_pad FILLER_9/VDDIO_Q vddio vssio FILLER_9/VSSIO_Q vddio vccd vccd sky130_ef_io__vssio_hvc_clamped_pad
Xsky130_ef_io__gpiov2_pad_wrapped_12 gpio_in_h[6] analog_noesd_io[6] analog_io[6]
+ sky130_ef_io__gpiov2_pad_wrapped_12/PAD_A_ESD_1_H gpio_dm2[6] gpio_dm1[6] gpio_dm0[6]
+ gpio_in[6] gpio_inp_dis[6] gpio_ib_mode_sel[6] porb_h porb_h sky130_ef_io__gpiov2_pad_wrapped_12/TIE_LO_ESD
+ gpio_oeb[6] sky130_ef_io__gpiov2_pad_wrapped_12/HLD_H_N sky130_ef_io__gpiov2_pad_wrapped_12/TIE_LO_ESD
+ gpio_slow_sel[6] gpio_vtrip_sel[6] gpio_holdover[6] gpio_analog_en[6] gpio_analog_sel[6]
+ gpio_loopback_one[6] sky130_ef_io__gpiov2_pad_wrapped_12/TIE_LO_ESD gpio_analog_pol[6]
+ gpio_out[6] FILLER_9/VDDIO_Q w_694469_374069# sky130_ef_io__gpiov2_pad_wrapped_12/HLD_H_N
+ FILLER_9/VSSIO_Q w_694469_370752# vccd FILLER_9/AMUXBUS_B FILLER_9/AMUXBUS_A vssio
+ vddio vdda1 w_692355_370752# vddio vssa1 w_692253_374070# vssd gpio[6] vccd sky130_ef_io__gpiov2_pad_wrapped
Xuser2_vssa_hvclamp_pad vssd vssa2 vddio vssa2_pad vccd vddio vssio FILLER_9/VDDIO_Q
+ vdda2 FILLER_9/VSSIO_Q vccd FILLER_9/AMUXBUS_B FILLER_9/AMUXBUS_A sky130_ef_io__vssa_hvc_clamped_pad
Xsky130_ef_io__gpiov2_pad_wrapped_0 gpio_in_h[37] analog_noesd_io[37] analog_io[37]
+ sky130_ef_io__gpiov2_pad_wrapped_0/PAD_A_ESD_1_H gpio_dm2[37] gpio_dm1[37] gpio_dm0[37]
+ gpio_in[37] gpio_inp_dis[37] gpio_ib_mode_sel[37] porb_h porb_h sky130_ef_io__gpiov2_pad_wrapped_0/TIE_LO_ESD
+ gpio_oeb[37] sky130_ef_io__gpiov2_pad_wrapped_0/HLD_H_N sky130_ef_io__gpiov2_pad_wrapped_0/TIE_LO_ESD
+ gpio_slow_sel[37] gpio_vtrip_sel[37] gpio_holdover[37] gpio_analog_en[37] gpio_analog_sel[37]
+ gpio_loopback_one[37] sky130_ef_io__gpiov2_pad_wrapped_0/TIE_LO_ESD gpio_analog_pol[37]
+ gpio_out[37] FILLER_9/VDDIO_Q w_21151_191274# sky130_ef_io__gpiov2_pad_wrapped_0/HLD_H_N
+ FILLER_9/VSSIO_Q w_21253_194365# vccd FILLER_9/AMUXBUS_B FILLER_9/AMUXBUS_A vssio
+ vddio vdda2 w_23367_194365# vddio vssa2 w_23367_191274# vssd gpio[37] vccd sky130_ef_io__gpiov2_pad_wrapped
Xconstant_value_inst[2] vccd gpio_loopback_zero[2] gpio_loopback_one[2] vssd constant_block
Xsky130_ef_io__gpiov2_pad_wrapped_13 gpio_in_h[5] analog_noesd_io[5] analog_io[5]
+ sky130_ef_io__gpiov2_pad_wrapped_13/PAD_A_ESD_1_H gpio_dm2[5] gpio_dm1[5] gpio_dm0[5]
+ gpio_in[5] gpio_inp_dis[5] gpio_ib_mode_sel[5] porb_h porb_h sky130_ef_io__gpiov2_pad_wrapped_13/TIE_LO_ESD
+ gpio_oeb[5] sky130_ef_io__gpiov2_pad_wrapped_13/HLD_H_N sky130_ef_io__gpiov2_pad_wrapped_13/TIE_LO_ESD
+ gpio_slow_sel[5] gpio_vtrip_sel[5] gpio_holdover[5] gpio_analog_en[5] gpio_analog_sel[5]
+ gpio_loopback_one[5] sky130_ef_io__gpiov2_pad_wrapped_13/TIE_LO_ESD gpio_analog_pol[5]
+ gpio_out[5] FILLER_9/VDDIO_Q w_694469_328869# sky130_ef_io__gpiov2_pad_wrapped_13/HLD_H_N
+ FILLER_9/VSSIO_Q w_694469_325552# vccd FILLER_9/AMUXBUS_B FILLER_9/AMUXBUS_A vssio
+ vddio vdda1 w_692355_325552# vddio vssa1 w_692253_328870# vssd gpio[5] vccd sky130_ef_io__gpiov2_pad_wrapped
Xconstant_value_inst[1] vccd gpio_loopback_zero[1] gpio_loopback_one[1] vssd constant_block
Xsky130_ef_io__gpiov2_pad_wrapped_1 gpio_in_h[36] analog_noesd_io[36] analog_io[36]
+ sky130_ef_io__gpiov2_pad_wrapped_1/PAD_A_ESD_1_H gpio_dm2[36] gpio_dm1[36] gpio_dm0[36]
+ gpio_in[36] gpio_inp_dis[36] gpio_ib_mode_sel[36] porb_h porb_h sky130_ef_io__gpiov2_pad_wrapped_1/TIE_LO_ESD
+ gpio_oeb[36] sky130_ef_io__gpiov2_pad_wrapped_1/HLD_H_N sky130_ef_io__gpiov2_pad_wrapped_1/TIE_LO_ESD
+ gpio_slow_sel[36] gpio_vtrip_sel[36] gpio_holdover[36] gpio_analog_en[36] gpio_analog_sel[36]
+ gpio_loopback_one[36] sky130_ef_io__gpiov2_pad_wrapped_1/TIE_LO_ESD gpio_analog_pol[36]
+ gpio_out[36] FILLER_9/VDDIO_Q w_21151_234474# sky130_ef_io__gpiov2_pad_wrapped_1/HLD_H_N
+ FILLER_9/VSSIO_Q w_21253_237565# vccd FILLER_9/AMUXBUS_B FILLER_9/AMUXBUS_A vssio
+ vddio vdda2 w_23367_237565# vddio vssa2 w_23367_234474# vssd gpio[36] vccd sky130_ef_io__gpiov2_pad_wrapped
Xsky130_ef_io__gpiov2_pad_wrapped_14 gpio_in_h[4] analog_noesd_io[4] analog_io[4]
+ sky130_ef_io__gpiov2_pad_wrapped_14/PAD_A_ESD_1_H gpio_dm2[4] gpio_dm1[4] gpio_dm0[4]
+ gpio_in[4] gpio_inp_dis[4] gpio_ib_mode_sel[4] porb_h porb_h sky130_ef_io__gpiov2_pad_wrapped_14/TIE_LO_ESD
+ gpio_oeb[4] sky130_ef_io__gpiov2_pad_wrapped_14/HLD_H_N sky130_ef_io__gpiov2_pad_wrapped_14/TIE_LO_ESD
+ gpio_slow_sel[4] gpio_vtrip_sel[4] gpio_holdover[4] gpio_analog_en[4] gpio_analog_sel[4]
+ gpio_loopback_one[4] sky130_ef_io__gpiov2_pad_wrapped_14/TIE_LO_ESD gpio_analog_pol[4]
+ gpio_out[4] FILLER_9/VDDIO_Q w_694469_283869# sky130_ef_io__gpiov2_pad_wrapped_14/HLD_H_N
+ FILLER_9/VSSIO_Q w_694469_280552# vccd FILLER_9/AMUXBUS_B FILLER_9/AMUXBUS_A vssio
+ vddio vdda1 w_692355_280552# vddio vssa1 w_692253_283870# vssd gpio[4] vccd sky130_ef_io__gpiov2_pad_wrapped
Xuser1_vdda_hvclamp_pad\[1\] FILLER_9/VDDIO_Q FILLER_9/VSSIO_Q vssio vdda1_pad2 FILLER_9/AMUXBUS_B
+ FILLER_9/AMUXBUS_A vdda1 vccd vssd vssa1 vddio vccd vddio sky130_ef_io__vdda_hvc_clamped_pad
Xconstant_value_inst[0] vccd gpio_loopback_zero[0] gpio_loopback_one[0] vssd constant_block
Xsky130_ef_io__gpiov2_pad_wrapped_2 gpio_in_h[35] analog_noesd_io[35] analog_io[35]
+ sky130_ef_io__gpiov2_pad_wrapped_2/PAD_A_ESD_1_H gpio_dm2[35] gpio_dm1[35] gpio_dm0[35]
+ gpio_in[35] gpio_inp_dis[35] gpio_ib_mode_sel[35] porb_h porb_h sky130_ef_io__gpiov2_pad_wrapped_2/TIE_LO_ESD
+ gpio_oeb[35] sky130_ef_io__gpiov2_pad_wrapped_2/HLD_H_N sky130_ef_io__gpiov2_pad_wrapped_2/TIE_LO_ESD
+ gpio_slow_sel[35] gpio_vtrip_sel[35] gpio_holdover[35] gpio_analog_en[35] gpio_analog_sel[35]
+ gpio_loopback_one[35] sky130_ef_io__gpiov2_pad_wrapped_2/TIE_LO_ESD gpio_analog_pol[35]
+ gpio_out[35] FILLER_9/VDDIO_Q w_21151_277674# sky130_ef_io__gpiov2_pad_wrapped_2/HLD_H_N
+ FILLER_9/VSSIO_Q w_21253_280765# vccd FILLER_9/AMUXBUS_B FILLER_9/AMUXBUS_A vssio
+ vddio vdda2 w_23367_280765# vddio vssa2 w_23367_277674# vssd gpio[35] vccd sky130_ef_io__gpiov2_pad_wrapped
Xsky130_ef_io__gpiov2_pad_wrapped_15 gpio_in_h[3] analog_noesd_io[3] analog_io[3]
+ sky130_ef_io__gpiov2_pad_wrapped_15/PAD_A_ESD_1_H gpio_dm2[3] gpio_dm1[3] gpio_dm0[3]
+ gpio_in[3] gpio_inp_dis[3] gpio_ib_mode_sel[3] porb_h porb_h sky130_ef_io__gpiov2_pad_wrapped_15/TIE_LO_ESD
+ gpio_oeb[3] sky130_ef_io__gpiov2_pad_wrapped_15/HLD_H_N sky130_ef_io__gpiov2_pad_wrapped_15/TIE_LO_ESD
+ gpio_slow_sel[3] gpio_vtrip_sel[3] gpio_holdover[3] gpio_analog_en[3] gpio_analog_sel[3]
+ gpio_loopback_one[3] sky130_ef_io__gpiov2_pad_wrapped_15/TIE_LO_ESD gpio_analog_pol[3]
+ gpio_out[3] FILLER_9/VDDIO_Q w_694469_238869# sky130_ef_io__gpiov2_pad_wrapped_15/HLD_H_N
+ FILLER_9/VSSIO_Q w_694469_235552# vccd FILLER_9/AMUXBUS_B FILLER_9/AMUXBUS_A vssio
+ vddio vdda1 w_692355_235552# vddio vssa1 w_692253_238870# vssd gpio[3] vccd sky130_ef_io__gpiov2_pad_wrapped
Xsky130_ef_io__gpiov2_pad_wrapped_3 gpio_in_h[34] analog_noesd_io[34] analog_io[34]
+ sky130_ef_io__gpiov2_pad_wrapped_3/PAD_A_ESD_1_H gpio_dm2[34] gpio_dm1[34] gpio_dm0[34]
+ gpio_in[34] gpio_inp_dis[34] gpio_ib_mode_sel[34] porb_h porb_h sky130_ef_io__gpiov2_pad_wrapped_3/TIE_LO_ESD
+ gpio_oeb[34] sky130_ef_io__gpiov2_pad_wrapped_3/HLD_H_N sky130_ef_io__gpiov2_pad_wrapped_3/TIE_LO_ESD
+ gpio_slow_sel[34] gpio_vtrip_sel[34] gpio_holdover[34] gpio_analog_en[34] gpio_analog_sel[34]
+ gpio_loopback_one[34] sky130_ef_io__gpiov2_pad_wrapped_3/TIE_LO_ESD gpio_analog_pol[34]
+ gpio_out[34] FILLER_9/VDDIO_Q w_21151_320874# sky130_ef_io__gpiov2_pad_wrapped_3/HLD_H_N
+ FILLER_9/VSSIO_Q w_21253_323965# vccd FILLER_9/AMUXBUS_B FILLER_9/AMUXBUS_A vssio
+ vddio vdda2 w_23367_323965# vddio vssa2 w_23367_320874# vssd gpio[34] vccd sky130_ef_io__gpiov2_pad_wrapped
Xsky130_ef_io__gpiov2_pad_wrapped_16 gpio_in_h[2] analog_noesd_io[2] analog_io[2]
+ sky130_ef_io__gpiov2_pad_wrapped_16/PAD_A_ESD_1_H gpio_dm2[2] gpio_dm1[2] gpio_dm0[2]
+ gpio_in[2] gpio_inp_dis[2] gpio_ib_mode_sel[2] porb_h porb_h sky130_ef_io__gpiov2_pad_wrapped_16/TIE_LO_ESD
+ gpio_oeb[2] sky130_ef_io__gpiov2_pad_wrapped_16/HLD_H_N sky130_ef_io__gpiov2_pad_wrapped_16/TIE_LO_ESD
+ gpio_slow_sel[2] gpio_vtrip_sel[2] gpio_holdover[2] gpio_analog_en[2] gpio_analog_sel[2]
+ gpio_loopback_one[2] sky130_ef_io__gpiov2_pad_wrapped_16/TIE_LO_ESD gpio_analog_pol[2]
+ gpio_out[2] FILLER_9/VDDIO_Q w_694469_193669# sky130_ef_io__gpiov2_pad_wrapped_16/HLD_H_N
+ FILLER_9/VSSIO_Q w_694469_190352# vccd FILLER_9/AMUXBUS_B FILLER_9/AMUXBUS_A vssio
+ vddio vdda1 w_692355_190352# vddio vssa1 w_692253_193670# vssd gpio[2] vccd sky130_ef_io__gpiov2_pad_wrapped
Xsky130_ef_io__gpiov2_pad_wrapped_4 gpio_in_h[33] analog_noesd_io[33] analog_io[33]
+ sky130_ef_io__gpiov2_pad_wrapped_4/PAD_A_ESD_1_H gpio_dm2[33] gpio_dm1[33] gpio_dm0[33]
+ gpio_in[33] gpio_inp_dis[33] gpio_ib_mode_sel[33] porb_h porb_h sky130_ef_io__gpiov2_pad_wrapped_4/TIE_LO_ESD
+ gpio_oeb[33] sky130_ef_io__gpiov2_pad_wrapped_4/HLD_H_N sky130_ef_io__gpiov2_pad_wrapped_4/TIE_LO_ESD
+ gpio_slow_sel[33] gpio_vtrip_sel[33] gpio_holdover[33] gpio_analog_en[33] gpio_analog_sel[33]
+ gpio_loopback_one[33] sky130_ef_io__gpiov2_pad_wrapped_4/TIE_LO_ESD gpio_analog_pol[33]
+ gpio_out[33] FILLER_9/VDDIO_Q w_21151_364074# sky130_ef_io__gpiov2_pad_wrapped_4/HLD_H_N
+ FILLER_9/VSSIO_Q w_21253_367165# vccd FILLER_9/AMUXBUS_B FILLER_9/AMUXBUS_A vssio
+ vddio vdda2 w_23367_367165# vddio vssa2 w_23367_364074# vssd gpio[33] vccd sky130_ef_io__gpiov2_pad_wrapped
Xconstant_value_inst[29] vccd gpio_loopback_zero[29] gpio_loopback_one[29] vssd constant_block
Xsky130_ef_io__gpiov2_pad_wrapped_17 gpio_in_h[1] analog_noesd_io[1] analog_io[1]
+ sky130_ef_io__gpiov2_pad_wrapped_17/PAD_A_ESD_1_H gpio_dm2[1] gpio_dm1[1] gpio_dm0[1]
+ gpio_in[1] gpio_inp_dis[1] gpio_ib_mode_sel[1] porb_h porb_h sky130_ef_io__gpiov2_pad_wrapped_17/TIE_LO_ESD
+ gpio_oeb[1] sky130_ef_io__gpiov2_pad_wrapped_17/HLD_H_N sky130_ef_io__gpiov2_pad_wrapped_17/TIE_LO_ESD
+ gpio_slow_sel[1] gpio_vtrip_sel[1] gpio_holdover[1] gpio_analog_en[1] gpio_analog_sel[1]
+ gpio_loopback_one[1] sky130_ef_io__gpiov2_pad_wrapped_17/TIE_LO_ESD gpio_analog_pol[1]
+ gpio_out[1] FILLER_9/VDDIO_Q w_694469_148669# sky130_ef_io__gpiov2_pad_wrapped_17/HLD_H_N
+ FILLER_9/VSSIO_Q w_694469_145352# vccd FILLER_9/AMUXBUS_B FILLER_9/AMUXBUS_A vssio
+ vddio vdda1 w_692355_145352# vddio vssa1 w_692253_148670# vssd gpio[1] vccd sky130_ef_io__gpiov2_pad_wrapped
Xmgmt_vdda_hvclamp_pad FILLER_9/VDDIO_Q FILLER_9/VSSIO_Q vssio vdda_pad FILLER_9/AMUXBUS_B
+ FILLER_9/AMUXBUS_A vdda vccd vssd vssa vddio vccd vddio sky130_ef_io__vdda_hvc_clamped_pad
Xmaster_resetb_pad resetb_h xres_vss_loop constant_value_xres_inst/one xresloop porb_h
+ xres_vss_loop xres_vss_loop xres_vss_loop master_resetb_pad/TIE_HI_ESD xres_vss_loop
+ xres_vss_loop vssa vssd FILLER_9/AMUXBUS_B FILLER_9/AMUXBUS_A FILLER_9/VDDIO_Q vddio
+ vddio vdda vccd vccd FILLER_9/VSSIO_Q vssio resetb_pad xresloop sky130_fd_io__top_xres4v2
Xsky130_ef_io__gpiov2_pad_wrapped_5 gpio_in_h[32] analog_noesd_io[32] analog_io[32]
+ sky130_ef_io__gpiov2_pad_wrapped_5/PAD_A_ESD_1_H gpio_dm2[32] gpio_dm1[32] gpio_dm0[32]
+ gpio_in[32] gpio_inp_dis[32] gpio_ib_mode_sel[32] porb_h porb_h sky130_ef_io__gpiov2_pad_wrapped_5/TIE_LO_ESD
+ gpio_oeb[32] sky130_ef_io__gpiov2_pad_wrapped_5/HLD_H_N sky130_ef_io__gpiov2_pad_wrapped_5/TIE_LO_ESD
+ gpio_slow_sel[32] gpio_vtrip_sel[32] gpio_holdover[32] gpio_analog_en[32] gpio_analog_sel[32]
+ gpio_loopback_one[32] sky130_ef_io__gpiov2_pad_wrapped_5/TIE_LO_ESD gpio_analog_pol[32]
+ gpio_out[32] FILLER_9/VDDIO_Q w_21151_407274# sky130_ef_io__gpiov2_pad_wrapped_5/HLD_H_N
+ FILLER_9/VSSIO_Q w_21253_410365# vccd FILLER_9/AMUXBUS_B FILLER_9/AMUXBUS_A vssio
+ vddio vdda2 w_23367_410365# vddio vssa2 w_23367_407274# vssd gpio[32] vccd sky130_ef_io__gpiov2_pad_wrapped
Xconstant_value_inst[28] vccd gpio_loopback_zero[28] gpio_loopback_one[28] vssd constant_block
Xsky130_ef_io__gpiov2_pad_wrapped_18 gpio_in_h[0] analog_noesd_io[0] analog_io[0]
+ sky130_ef_io__gpiov2_pad_wrapped_18/PAD_A_ESD_1_H gpio_dm2[0] gpio_dm1[0] gpio_dm0[0]
+ gpio_in[0] gpio_inp_dis[0] gpio_ib_mode_sel[0] porb_h porb_h sky130_ef_io__gpiov2_pad_wrapped_18/TIE_LO_ESD
+ gpio_oeb[0] sky130_ef_io__gpiov2_pad_wrapped_18/HLD_H_N sky130_ef_io__gpiov2_pad_wrapped_18/TIE_LO_ESD
+ gpio_slow_sel[0] gpio_vtrip_sel[0] gpio_holdover[0] gpio_analog_en[0] gpio_analog_sel[0]
+ gpio_loopback_one[0] sky130_ef_io__gpiov2_pad_wrapped_18/TIE_LO_ESD gpio_analog_pol[0]
+ gpio_out[0] FILLER_9/VDDIO_Q w_694469_103469# sky130_ef_io__gpiov2_pad_wrapped_18/HLD_H_N
+ FILLER_9/VSSIO_Q w_694469_100152# vccd FILLER_9/AMUXBUS_B FILLER_9/AMUXBUS_A vssio
+ vddio vdda1 w_692355_100152# vddio vssa1 w_692253_103470# vssd gpio[0] vccd sky130_ef_io__gpiov2_pad_wrapped
Xsky130_ef_io__gpiov2_pad_wrapped_6 gpio_in_h[31] analog_noesd_io[31] analog_io[31]
+ sky130_ef_io__gpiov2_pad_wrapped_6/PAD_A_ESD_1_H gpio_dm2[31] gpio_dm1[31] gpio_dm0[31]
+ gpio_in[31] gpio_inp_dis[31] gpio_ib_mode_sel[31] porb_h porb_h sky130_ef_io__gpiov2_pad_wrapped_6/TIE_LO_ESD
+ gpio_oeb[31] sky130_ef_io__gpiov2_pad_wrapped_6/HLD_H_N sky130_ef_io__gpiov2_pad_wrapped_6/TIE_LO_ESD
+ gpio_slow_sel[31] gpio_vtrip_sel[31] gpio_holdover[31] gpio_analog_en[31] gpio_analog_sel[31]
+ gpio_loopback_one[31] sky130_ef_io__gpiov2_pad_wrapped_6/TIE_LO_ESD gpio_analog_pol[31]
+ gpio_out[31] FILLER_9/VDDIO_Q w_21151_534874# sky130_ef_io__gpiov2_pad_wrapped_6/HLD_H_N
+ FILLER_9/VSSIO_Q w_21253_537965# vccd FILLER_9/AMUXBUS_B FILLER_9/AMUXBUS_A vssio
+ vddio vdda2 w_23367_537965# vddio vssa2 w_23367_534874# vssd gpio[31] vccd sky130_ef_io__gpiov2_pad_wrapped
Xconstant_value_inst[27] vccd gpio_loopback_zero[27] gpio_loopback_one[27] vssd constant_block
Xuser1_vssa_hvclamp_pad\[0\] vssd vssa1 vddio vssa1_pad vccd vddio vssio FILLER_9/VDDIO_Q
+ vdda1 FILLER_9/VSSIO_Q vccd FILLER_9/AMUXBUS_B FILLER_9/AMUXBUS_A sky130_ef_io__vssa_hvc_clamped_pad
Xsky130_ef_io__gpiov2_pad_wrapped_7 gpio_in_h[30] analog_noesd_io[30] analog_io[30]
+ sky130_ef_io__gpiov2_pad_wrapped_7/PAD_A_ESD_1_H gpio_dm2[30] gpio_dm1[30] gpio_dm0[30]
+ gpio_in[30] gpio_inp_dis[30] gpio_ib_mode_sel[30] porb_h porb_h sky130_ef_io__gpiov2_pad_wrapped_7/TIE_LO_ESD
+ gpio_oeb[30] sky130_ef_io__gpiov2_pad_wrapped_7/HLD_H_N sky130_ef_io__gpiov2_pad_wrapped_7/TIE_LO_ESD
+ gpio_slow_sel[30] gpio_vtrip_sel[30] gpio_holdover[30] gpio_analog_en[30] gpio_analog_sel[30]
+ gpio_loopback_one[30] sky130_ef_io__gpiov2_pad_wrapped_7/TIE_LO_ESD gpio_analog_pol[30]
+ gpio_out[30] FILLER_9/VDDIO_Q w_21151_578074# sky130_ef_io__gpiov2_pad_wrapped_7/HLD_H_N
+ FILLER_9/VSSIO_Q w_21253_581165# vccd FILLER_9/AMUXBUS_B FILLER_9/AMUXBUS_A vssio
+ vddio vdda2 w_23367_581165# vddio vssa2 w_23367_578074# vssd gpio[30] vccd sky130_ef_io__gpiov2_pad_wrapped
Xconstant_value_inst[43] vccd gpio_loopback_zero[43] gpio_loopback_one[43] vssd constant_block
Xconstant_value_inst[26] vccd gpio_loopback_zero[26] gpio_loopback_one[26] vssd constant_block
Xuser1_vccd_lvclamp_pad vdda1 vccd vssd1 vddio vddio FILLER_9/AMUXBUS_B vssio FILLER_9/AMUXBUS_A
+ vccd vccd1_pad vccd1 vssd FILLER_9/VDDIO_Q vssa1 FILLER_9/VSSIO_Q sky130_ef_io__vccd_lvc_clamped3_pad
Xsky130_ef_io__gpiov2_pad_wrapped_8 gpio_in_h[29] analog_noesd_io[29] analog_io[29]
+ sky130_ef_io__gpiov2_pad_wrapped_8/PAD_A_ESD_1_H gpio_dm2[29] gpio_dm1[29] gpio_dm0[29]
+ gpio_in[29] gpio_inp_dis[29] gpio_ib_mode_sel[29] porb_h porb_h sky130_ef_io__gpiov2_pad_wrapped_8/TIE_LO_ESD
+ gpio_oeb[29] sky130_ef_io__gpiov2_pad_wrapped_8/HLD_H_N sky130_ef_io__gpiov2_pad_wrapped_8/TIE_LO_ESD
+ gpio_slow_sel[29] gpio_vtrip_sel[29] gpio_holdover[29] gpio_analog_en[29] gpio_analog_sel[29]
+ gpio_loopback_one[29] sky130_ef_io__gpiov2_pad_wrapped_8/TIE_LO_ESD gpio_analog_pol[29]
+ gpio_out[29] FILLER_9/VDDIO_Q w_21151_621274# sky130_ef_io__gpiov2_pad_wrapped_8/HLD_H_N
+ FILLER_9/VSSIO_Q w_21253_624365# vccd FILLER_9/AMUXBUS_B FILLER_9/AMUXBUS_A vssio
+ vddio vdda2 w_23367_624365# vddio vssa2 w_23367_621274# vssd gpio[29] vccd sky130_ef_io__gpiov2_pad_wrapped
Xconstant_value_inst[42] vccd gpio_loopback_zero[42] gpio_loopback_one[42] vssd constant_block
Xconstant_value_inst[25] vccd gpio_loopback_zero[25] gpio_loopback_one[25] vssd constant_block
.ends

.subckt caravel_openframe vddio vddio_2 vssio vssio_2 vdda vssa vccd vssd vdda1 vdda1_2
+ vssa1 vssa1_2 vssa2 vccd1 vccd2 vssd1 vssd2 gpio[0] gpio[1] gpio[2] gpio[3] gpio[4]
+ gpio[5] gpio[6] gpio[7] gpio[8] gpio[9] gpio[10] gpio[11] gpio[12] gpio[13] gpio[14]
+ gpio[15] gpio[16] gpio[17] gpio[18] gpio[19] gpio[20] gpio[21] gpio[22] gpio[23]
+ gpio[24] gpio[25] gpio[26] gpio[27] gpio[28] gpio[29] gpio[30] gpio[31] gpio[32]
+ gpio[33] gpio[34] gpio[35] gpio[36] gpio[37] gpio[38] gpio[39] gpio[40] gpio[41]
+ gpio[42] gpio[43] resetb vdda2
Xchip_io_openframe_0 vddio vssio vdda1_2 vccd2 chip_io_openframe_0/vddio chip_io_openframe_0/vccd
+ chip_io_openframe_0/vdda chip_io_openframe_0/vdda1 chip_io_openframe_0/vdda2 chip_io_openframe_0/vccd1
+ chip_io_openframe_0/vccd2 chip_io_openframe_0/porb_l chip_io_openframe_0/por_l chip_io_openframe_0/resetb_h
+ chip_io_openframe_0/resetb_l chip_io_openframe_0/mask_rev[31] chip_io_openframe_0/mask_rev[30]
+ chip_io_openframe_0/mask_rev[29] chip_io_openframe_0/mask_rev[28] chip_io_openframe_0/mask_rev[27]
+ chip_io_openframe_0/mask_rev[26] chip_io_openframe_0/mask_rev[25] chip_io_openframe_0/mask_rev[24]
+ chip_io_openframe_0/mask_rev[23] chip_io_openframe_0/mask_rev[22] chip_io_openframe_0/mask_rev[21]
+ chip_io_openframe_0/mask_rev[20] chip_io_openframe_0/mask_rev[19] chip_io_openframe_0/mask_rev[18]
+ chip_io_openframe_0/mask_rev[17] chip_io_openframe_0/mask_rev[16] chip_io_openframe_0/mask_rev[15]
+ chip_io_openframe_0/mask_rev[14] chip_io_openframe_0/mask_rev[13] chip_io_openframe_0/mask_rev[12]
+ chip_io_openframe_0/mask_rev[11] chip_io_openframe_0/mask_rev[10] chip_io_openframe_0/mask_rev[9]
+ chip_io_openframe_0/mask_rev[8] chip_io_openframe_0/mask_rev[7] chip_io_openframe_0/mask_rev[6]
+ chip_io_openframe_0/mask_rev[5] chip_io_openframe_0/mask_rev[4] chip_io_openframe_0/mask_rev[3]
+ chip_io_openframe_0/mask_rev[2] chip_io_openframe_0/mask_rev[1] chip_io_openframe_0/mask_rev[0]
+ gpio[36] chip_io_openframe_0/gpio_out[41] chip_io_openframe_0/gpio_out[39] chip_io_openframe_0/gpio_out[38]
+ chip_io_openframe_0/gpio_out[37] chip_io_openframe_0/gpio_out[36] chip_io_openframe_0/gpio_out[35]
+ chip_io_openframe_0/gpio_out[33] chip_io_openframe_0/gpio_out[32] chip_io_openframe_0/gpio_out[30]
+ chip_io_openframe_0/gpio_out[26] chip_io_openframe_0/gpio_out[23] chip_io_openframe_0/gpio_out[18]
+ chip_io_openframe_0/gpio_out[17] chip_io_openframe_0/gpio_out[16] chip_io_openframe_0/gpio_out[15]
+ chip_io_openframe_0/gpio_out[13] chip_io_openframe_0/gpio_out[12] chip_io_openframe_0/gpio_oeb[43]
+ chip_io_openframe_0/gpio_oeb[42] chip_io_openframe_0/gpio_oeb[41] chip_io_openframe_0/gpio_oeb[37]
+ chip_io_openframe_0/gpio_oeb[34] chip_io_openframe_0/gpio_oeb[29] chip_io_openframe_0/gpio_oeb[28]
+ chip_io_openframe_0/gpio_oeb[27] chip_io_openframe_0/gpio_oeb[26] chip_io_openframe_0/gpio_oeb[25]
+ chip_io_openframe_0/gpio_oeb[24] chip_io_openframe_0/gpio_oeb[23] chip_io_openframe_0/gpio_oeb[22]
+ chip_io_openframe_0/gpio_oeb[21] chip_io_openframe_0/gpio_oeb[20] chip_io_openframe_0/gpio_oeb[18]
+ chip_io_openframe_0/gpio_oeb[17] chip_io_openframe_0/gpio_oeb[16] chip_io_openframe_0/gpio_oeb[15]
+ chip_io_openframe_0/gpio_oeb[14] chip_io_openframe_0/gpio_oeb[13] chip_io_openframe_0/gpio_oeb[6]
+ chip_io_openframe_0/gpio_oeb[3] chip_io_openframe_0/gpio_oeb[0] chip_io_openframe_0/gpio_inp_dis[39]
+ chip_io_openframe_0/gpio_inp_dis[37] chip_io_openframe_0/gpio_inp_dis[36] chip_io_openframe_0/gpio_inp_dis[33]
+ chip_io_openframe_0/gpio_inp_dis[32] chip_io_openframe_0/gpio_inp_dis[22] chip_io_openframe_0/gpio_inp_dis[21]
+ chip_io_openframe_0/gpio_inp_dis[20] chip_io_openframe_0/gpio_inp_dis[18] chip_io_openframe_0/gpio_inp_dis[15]
+ chip_io_openframe_0/gpio_inp_dis[14] chip_io_openframe_0/gpio_inp_dis[12] chip_io_openframe_0/gpio_inp_dis[11]
+ chip_io_openframe_0/gpio_inp_dis[8] chip_io_openframe_0/gpio_inp_dis[4] chip_io_openframe_0/gpio_ib_mode_sel[43]
+ chip_io_openframe_0/gpio_ib_mode_sel[42] chip_io_openframe_0/gpio_ib_mode_sel[40]
+ chip_io_openframe_0/gpio_ib_mode_sel[39] chip_io_openframe_0/gpio_ib_mode_sel[38]
+ chip_io_openframe_0/gpio_ib_mode_sel[37] chip_io_openframe_0/gpio_ib_mode_sel[36]
+ chip_io_openframe_0/gpio_ib_mode_sel[35] chip_io_openframe_0/gpio_ib_mode_sel[34]
+ chip_io_openframe_0/gpio_ib_mode_sel[33] chip_io_openframe_0/gpio_ib_mode_sel[32]
+ chip_io_openframe_0/gpio_ib_mode_sel[31] chip_io_openframe_0/gpio_ib_mode_sel[30]
+ chip_io_openframe_0/gpio_ib_mode_sel[26] chip_io_openframe_0/gpio_ib_mode_sel[25]
+ chip_io_openframe_0/gpio_ib_mode_sel[24] chip_io_openframe_0/gpio_ib_mode_sel[23]
+ chip_io_openframe_0/gpio_ib_mode_sel[22] chip_io_openframe_0/gpio_ib_mode_sel[21]
+ chip_io_openframe_0/gpio_ib_mode_sel[20] chip_io_openframe_0/gpio_ib_mode_sel[18]
+ chip_io_openframe_0/gpio_ib_mode_sel[15] chip_io_openframe_0/gpio_ib_mode_sel[14]
+ chip_io_openframe_0/gpio_ib_mode_sel[10] chip_io_openframe_0/gpio_ib_mode_sel[8]
+ chip_io_openframe_0/gpio_ib_mode_sel[7] chip_io_openframe_0/gpio_ib_mode_sel[6]
+ chip_io_openframe_0/gpio_ib_mode_sel[5] chip_io_openframe_0/gpio_ib_mode_sel[4]
+ chip_io_openframe_0/gpio_vtrip_sel[42] chip_io_openframe_0/gpio_vtrip_sel[41] chip_io_openframe_0/gpio_vtrip_sel[40]
+ chip_io_openframe_0/gpio_vtrip_sel[37] chip_io_openframe_0/gpio_vtrip_sel[36] chip_io_openframe_0/gpio_vtrip_sel[34]
+ chip_io_openframe_0/gpio_vtrip_sel[33] chip_io_openframe_0/gpio_vtrip_sel[32] chip_io_openframe_0/gpio_vtrip_sel[30]
+ chip_io_openframe_0/gpio_vtrip_sel[29] chip_io_openframe_0/gpio_vtrip_sel[19] chip_io_openframe_0/gpio_vtrip_sel[18]
+ chip_io_openframe_0/gpio_vtrip_sel[17] chip_io_openframe_0/gpio_vtrip_sel[16] chip_io_openframe_0/gpio_vtrip_sel[15]
+ chip_io_openframe_0/gpio_vtrip_sel[14] chip_io_openframe_0/gpio_vtrip_sel[13] chip_io_openframe_0/gpio_vtrip_sel[12]
+ chip_io_openframe_0/gpio_vtrip_sel[5] chip_io_openframe_0/gpio_vtrip_sel[4] chip_io_openframe_0/gpio_vtrip_sel[3]
+ chip_io_openframe_0/gpio_vtrip_sel[2] chip_io_openframe_0/gpio_vtrip_sel[1] chip_io_openframe_0/gpio_vtrip_sel[0]
+ chip_io_openframe_0/gpio_slow_sel[34] chip_io_openframe_0/gpio_slow_sel[33] chip_io_openframe_0/gpio_slow_sel[32]
+ chip_io_openframe_0/gpio_slow_sel[31] chip_io_openframe_0/gpio_slow_sel[30] chip_io_openframe_0/gpio_slow_sel[29]
+ chip_io_openframe_0/gpio_slow_sel[24] chip_io_openframe_0/gpio_slow_sel[23] chip_io_openframe_0/gpio_slow_sel[22]
+ chip_io_openframe_0/gpio_slow_sel[21] chip_io_openframe_0/gpio_slow_sel[20] chip_io_openframe_0/gpio_slow_sel[17]
+ chip_io_openframe_0/gpio_slow_sel[16] chip_io_openframe_0/gpio_slow_sel[15] chip_io_openframe_0/gpio_slow_sel[14]
+ chip_io_openframe_0/gpio_slow_sel[13] chip_io_openframe_0/gpio_slow_sel[12] chip_io_openframe_0/gpio_slow_sel[11]
+ chip_io_openframe_0/gpio_slow_sel[10] chip_io_openframe_0/gpio_slow_sel[9] chip_io_openframe_0/gpio_slow_sel[8]
+ chip_io_openframe_0/gpio_slow_sel[5] chip_io_openframe_0/gpio_holdover[43] chip_io_openframe_0/gpio_holdover[42]
+ chip_io_openframe_0/gpio_holdover[32] chip_io_openframe_0/gpio_holdover[31] chip_io_openframe_0/gpio_holdover[29]
+ chip_io_openframe_0/gpio_holdover[28] chip_io_openframe_0/gpio_holdover[27] chip_io_openframe_0/gpio_holdover[24]
+ chip_io_openframe_0/gpio_holdover[21] chip_io_openframe_0/gpio_holdover[20] chip_io_openframe_0/gpio_holdover[15]
+ chip_io_openframe_0/gpio_holdover[14] chip_io_openframe_0/gpio_holdover[13] chip_io_openframe_0/gpio_holdover[12]
+ chip_io_openframe_0/gpio_holdover[11] chip_io_openframe_0/gpio_holdover[10] chip_io_openframe_0/gpio_holdover[9]
+ chip_io_openframe_0/gpio_holdover[8] chip_io_openframe_0/gpio_holdover[7] chip_io_openframe_0/gpio_holdover[6]
+ chip_io_openframe_0/gpio_holdover[4] chip_io_openframe_0/gpio_holdover[3] chip_io_openframe_0/gpio_holdover[2]
+ chip_io_openframe_0/gpio_holdover[0] chip_io_openframe_0/gpio_analog_en[38] chip_io_openframe_0/gpio_analog_en[37]
+ chip_io_openframe_0/gpio_analog_en[36] chip_io_openframe_0/gpio_analog_en[35] chip_io_openframe_0/gpio_analog_en[34]
+ chip_io_openframe_0/gpio_analog_en[33] chip_io_openframe_0/gpio_analog_en[31] chip_io_openframe_0/gpio_analog_en[30]
+ chip_io_openframe_0/gpio_analog_en[26] chip_io_openframe_0/gpio_analog_en[25] chip_io_openframe_0/gpio_analog_en[19]
+ chip_io_openframe_0/gpio_analog_en[17] chip_io_openframe_0/gpio_analog_en[16] chip_io_openframe_0/gpio_analog_en[15]
+ chip_io_openframe_0/gpio_analog_en[14] chip_io_openframe_0/gpio_analog_en[13] chip_io_openframe_0/gpio_analog_en[12]
+ chip_io_openframe_0/gpio_analog_en[11] chip_io_openframe_0/gpio_analog_en[10] chip_io_openframe_0/gpio_analog_en[7]
+ chip_io_openframe_0/gpio_analog_en[6] chip_io_openframe_0/gpio_analog_en[5] chip_io_openframe_0/gpio_analog_en[3]
+ chip_io_openframe_0/gpio_analog_en[2] chip_io_openframe_0/gpio_analog_en[1] chip_io_openframe_0/gpio_analog_sel[36]
+ chip_io_openframe_0/gpio_analog_sel[35] chip_io_openframe_0/gpio_analog_sel[34]
+ chip_io_openframe_0/gpio_analog_sel[33] chip_io_openframe_0/gpio_analog_sel[32]
+ chip_io_openframe_0/gpio_analog_sel[31] chip_io_openframe_0/gpio_analog_sel[30]
+ chip_io_openframe_0/gpio_analog_sel[19] chip_io_openframe_0/gpio_analog_sel[18]
+ chip_io_openframe_0/gpio_analog_sel[17] chip_io_openframe_0/gpio_analog_sel[16]
+ chip_io_openframe_0/gpio_analog_sel[8] chip_io_openframe_0/gpio_analog_sel[7] chip_io_openframe_0/gpio_analog_sel[6]
+ chip_io_openframe_0/gpio_analog_pol[39] chip_io_openframe_0/gpio_analog_pol[38]
+ chip_io_openframe_0/gpio_analog_pol[37] chip_io_openframe_0/gpio_analog_pol[36]
+ chip_io_openframe_0/gpio_analog_pol[32] chip_io_openframe_0/gpio_analog_pol[31]
+ chip_io_openframe_0/gpio_analog_pol[30] chip_io_openframe_0/gpio_analog_pol[27]
+ chip_io_openframe_0/gpio_analog_pol[26] chip_io_openframe_0/gpio_analog_pol[25]
+ chip_io_openframe_0/gpio_analog_pol[19] chip_io_openframe_0/gpio_analog_pol[9] chip_io_openframe_0/gpio_analog_pol[6]
+ chip_io_openframe_0/gpio_analog_pol[5] chip_io_openframe_0/gpio_analog_pol[4] chip_io_openframe_0/gpio_analog_pol[3]
+ chip_io_openframe_0/gpio_analog_pol[2] chip_io_openframe_0/gpio_dm0[43] chip_io_openframe_0/gpio_dm0[42]
+ chip_io_openframe_0/gpio_dm0[39] chip_io_openframe_0/gpio_dm0[30] chip_io_openframe_0/gpio_dm0[27]
+ chip_io_openframe_0/gpio_dm0[23] chip_io_openframe_0/gpio_dm0[22] chip_io_openframe_0/gpio_dm0[13]
+ chip_io_openframe_0/gpio_dm0[12] chip_io_openframe_0/gpio_dm0[10] chip_io_openframe_0/gpio_dm0[9]
+ chip_io_openframe_0/gpio_dm0[8] chip_io_openframe_0/gpio_dm0[7] chip_io_openframe_0/gpio_dm0[6]
+ chip_io_openframe_0/gpio_dm0[5] chip_io_openframe_0/gpio_dm0[4] chip_io_openframe_0/gpio_dm0[3]
+ chip_io_openframe_0/gpio_dm1[43] chip_io_openframe_0/gpio_dm1[42] chip_io_openframe_0/gpio_dm1[41]
+ chip_io_openframe_0/gpio_dm1[39] chip_io_openframe_0/gpio_dm1[38] chip_io_openframe_0/gpio_dm1[29]
+ chip_io_openframe_0/gpio_dm1[28] chip_io_openframe_0/gpio_dm1[27] chip_io_openframe_0/gpio_dm1[26]
+ chip_io_openframe_0/gpio_dm1[25] chip_io_openframe_0/gpio_dm1[24] chip_io_openframe_0/gpio_dm1[23]
+ chip_io_openframe_0/gpio_dm1[22] chip_io_openframe_0/gpio_dm1[21] chip_io_openframe_0/gpio_dm1[20]
+ chip_io_openframe_0/gpio_dm1[16] chip_io_openframe_0/gpio_dm1[15] chip_io_openframe_0/gpio_dm1[11]
+ chip_io_openframe_0/gpio_dm1[10] chip_io_openframe_0/gpio_dm1[2] chip_io_openframe_0/gpio_dm1[1]
+ chip_io_openframe_0/gpio_dm1[0] chip_io_openframe_0/gpio_dm2[39] chip_io_openframe_0/gpio_dm2[38]
+ chip_io_openframe_0/gpio_dm2[37] chip_io_openframe_0/gpio_dm2[36] chip_io_openframe_0/gpio_dm2[24]
+ chip_io_openframe_0/gpio_dm2[16] chip_io_openframe_0/gpio_dm2[15] chip_io_openframe_0/gpio_dm2[14]
+ chip_io_openframe_0/gpio_dm2[11] chip_io_openframe_0/gpio_dm2[10] chip_io_openframe_0/gpio_dm2[9]
+ chip_io_openframe_0/gpio_dm2[8] chip_io_openframe_0/gpio_dm2[7] chip_io_openframe_0/gpio_dm2[6]
+ chip_io_openframe_0/gpio_dm2[5] chip_io_openframe_0/gpio_dm2[4] chip_io_openframe_0/gpio_dm2[3]
+ chip_io_openframe_0/gpio_dm2[2] chip_io_openframe_0/gpio_dm2[1] chip_io_openframe_0/gpio_dm2[0]
+ chip_io_openframe_0/gpio_in[42] chip_io_openframe_0/gpio_in[39] chip_io_openframe_0/gpio_in[38]
+ chip_io_openframe_0/gpio_in[37] chip_io_openframe_0/gpio_in[35] chip_io_openframe_0/gpio_in[34]
+ chip_io_openframe_0/gpio_in[32] chip_io_openframe_0/gpio_in[31] chip_io_openframe_0/gpio_in[28]
+ chip_io_openframe_0/gpio_in[25] chip_io_openframe_0/gpio_in[22] chip_io_openframe_0/gpio_in[19]
+ chip_io_openframe_0/gpio_in[18] chip_io_openframe_0/gpio_in[17] chip_io_openframe_0/gpio_in[16]
+ chip_io_openframe_0/gpio_in[14] chip_io_openframe_0/gpio_in[13] chip_io_openframe_0/gpio_in[11]
+ chip_io_openframe_0/gpio_in[10] chip_io_openframe_0/gpio_in[9] chip_io_openframe_0/gpio_in[7]
+ chip_io_openframe_0/gpio_in[4] chip_io_openframe_0/gpio_in[1] chip_io_openframe_0/gpio_in_h[40]
+ chip_io_openframe_0/gpio_in_h[39] chip_io_openframe_0/gpio_in_h[38] chip_io_openframe_0/gpio_in_h[37]
+ chip_io_openframe_0/gpio_in_h[36] chip_io_openframe_0/gpio_in_h[34] chip_io_openframe_0/gpio_in_h[33]
+ chip_io_openframe_0/gpio_in_h[31] chip_io_openframe_0/gpio_in_h[30] chip_io_openframe_0/gpio_in_h[20]
+ chip_io_openframe_0/gpio_in_h[19] chip_io_openframe_0/gpio_in_h[18] chip_io_openframe_0/gpio_in_h[17]
+ chip_io_openframe_0/gpio_in_h[16] chip_io_openframe_0/gpio_in_h[15] chip_io_openframe_0/gpio_in_h[14]
+ chip_io_openframe_0/gpio_in_h[13] chip_io_openframe_0/gpio_in_h[12] chip_io_openframe_0/gpio_in_h[11]
+ chip_io_openframe_0/gpio_in_h[10] chip_io_openframe_0/gpio_in_h[6] chip_io_openframe_0/gpio_in_h[3]
+ chip_io_openframe_0/gpio_in_h[0] chip_io_openframe_0/gpio_loopback_zero[43] chip_io_openframe_0/gpio_loopback_zero[42]
+ chip_io_openframe_0/gpio_loopback_zero[41] chip_io_openframe_0/gpio_loopback_zero[40]
+ chip_io_openframe_0/gpio_loopback_zero[39] chip_io_openframe_0/gpio_loopback_zero[38]
+ chip_io_openframe_0/gpio_loopback_zero[37] chip_io_openframe_0/gpio_loopback_zero[36]
+ chip_io_openframe_0/gpio_loopback_zero[35] chip_io_openframe_0/gpio_loopback_zero[34]
+ chip_io_openframe_0/gpio_loopback_zero[33] chip_io_openframe_0/gpio_loopback_zero[32]
+ chip_io_openframe_0/gpio_loopback_zero[31] chip_io_openframe_0/gpio_loopback_zero[30]
+ chip_io_openframe_0/gpio_loopback_zero[29] chip_io_openframe_0/gpio_loopback_zero[28]
+ chip_io_openframe_0/gpio_loopback_zero[27] chip_io_openframe_0/gpio_loopback_zero[26]
+ chip_io_openframe_0/gpio_loopback_zero[25] chip_io_openframe_0/gpio_loopback_zero[24]
+ chip_io_openframe_0/gpio_loopback_zero[23] chip_io_openframe_0/gpio_loopback_zero[22]
+ chip_io_openframe_0/gpio_loopback_zero[21] chip_io_openframe_0/gpio_loopback_zero[20]
+ chip_io_openframe_0/gpio_loopback_zero[19] chip_io_openframe_0/gpio_loopback_zero[18]
+ chip_io_openframe_0/gpio_loopback_zero[17] chip_io_openframe_0/gpio_loopback_zero[16]
+ chip_io_openframe_0/gpio_loopback_zero[15] chip_io_openframe_0/gpio_loopback_zero[14]
+ chip_io_openframe_0/gpio_loopback_zero[13] chip_io_openframe_0/gpio_loopback_zero[12]
+ chip_io_openframe_0/gpio_loopback_zero[11] chip_io_openframe_0/gpio_loopback_zero[10]
+ chip_io_openframe_0/gpio_loopback_zero[9] chip_io_openframe_0/gpio_loopback_zero[8]
+ chip_io_openframe_0/gpio_loopback_zero[7] chip_io_openframe_0/gpio_loopback_zero[6]
+ chip_io_openframe_0/gpio_loopback_zero[5] chip_io_openframe_0/gpio_loopback_zero[4]
+ chip_io_openframe_0/gpio_loopback_zero[3] chip_io_openframe_0/gpio_loopback_zero[2]
+ chip_io_openframe_0/gpio_loopback_zero[1] chip_io_openframe_0/gpio_loopback_zero[0]
+ chip_io_openframe_0/gpio_loopback_one[43] chip_io_openframe_0/gpio_loopback_one[42]
+ chip_io_openframe_0/gpio_loopback_one[41] chip_io_openframe_0/gpio_loopback_one[38]
+ chip_io_openframe_0/gpio_loopback_one[36] chip_io_openframe_0/gpio_loopback_one[35]
+ chip_io_openframe_0/gpio_loopback_one[31] chip_io_openframe_0/gpio_loopback_one[30]
+ chip_io_openframe_0/gpio_loopback_one[29] chip_io_openframe_0/gpio_loopback_one[28]
+ chip_io_openframe_0/gpio_loopback_one[27] chip_io_openframe_0/gpio_loopback_one[26]
+ chip_io_openframe_0/gpio_loopback_one[25] chip_io_openframe_0/gpio_loopback_one[24]
+ chip_io_openframe_0/gpio_loopback_one[22] chip_io_openframe_0/gpio_loopback_one[21]
+ chip_io_openframe_0/gpio_loopback_one[14] chip_io_openframe_0/gpio_loopback_one[11]
+ chip_io_openframe_0/gpio_loopback_one[8] chip_io_openframe_0/gpio_loopback_one[3]
+ chip_io_openframe_0/analog_io[39] chip_io_openframe_0/analog_io[36] chip_io_openframe_0/analog_io[35]
+ chip_io_openframe_0/analog_io[33] chip_io_openframe_0/analog_io[30] chip_io_openframe_0/analog_io[28]
+ chip_io_openframe_0/analog_io[26] chip_io_openframe_0/analog_io[20] chip_io_openframe_0/analog_io[19]
+ chip_io_openframe_0/analog_io[18] chip_io_openframe_0/analog_io[17] chip_io_openframe_0/analog_io[15]
+ chip_io_openframe_0/analog_io[14] chip_io_openframe_0/analog_io[13] chip_io_openframe_0/analog_io[10]
+ chip_io_openframe_0/analog_io[7] chip_io_openframe_0/analog_io[5] chip_io_openframe_0/analog_io[2]
+ chip_io_openframe_0/analog_noesd_io[43] chip_io_openframe_0/analog_noesd_io[42]
+ chip_io_openframe_0/analog_noesd_io[41] chip_io_openframe_0/analog_noesd_io[40]
+ chip_io_openframe_0/analog_noesd_io[39] chip_io_openframe_0/analog_noesd_io[38]
+ chip_io_openframe_0/analog_noesd_io[37] chip_io_openframe_0/analog_noesd_io[34]
+ chip_io_openframe_0/analog_noesd_io[28] chip_io_openframe_0/analog_noesd_io[27]
+ chip_io_openframe_0/analog_noesd_io[26] chip_io_openframe_0/analog_noesd_io[25]
+ chip_io_openframe_0/analog_noesd_io[23] chip_io_openframe_0/analog_noesd_io[22]
+ chip_io_openframe_0/analog_noesd_io[21] chip_io_openframe_0/analog_noesd_io[16]
+ chip_io_openframe_0/analog_noesd_io[12] chip_io_openframe_0/analog_noesd_io[6] chip_io_openframe_0/analog_noesd_io[1]
+ chip_io_openframe_0/analog_noesd_io[0] w_694469_865869# chip_io_openframe_0/gpio_analog_pol[20]
+ w_23367_407274# w_694469_100152# w_23367_534874# chip_io_openframe_0/gpio_out[0]
+ w_137274_1012253# chip_io_openframe_0/area1_gpio_pad[11]/PAD_A_ESD_1_H chip_io_openframe_0/sky130_ef_io__gpiov2_pad_wrapped_17/PAD_A_ESD_1_H
+ chip_io_openframe_0/sky130_ef_io__gpiov2_pad_wrapped_2/PAD_A_ESD_1_H w_188674_1014469#
+ w_404752_21253# w_459552_23367# chip_io_openframe_0/gpio_vtrip_sel[39] chip_io_openframe_0/gpio_analog_pol[21]
+ chip_io_openframe_0/area1_gpio_pad[5]/PAD_A_ESD_1_H w_485565_1014469# w_291674_1014469#
+ w_638765_1014469# w_23367_280765# chip_io_openframe_0/gpio_inp_dis[0] chip_io_openframe_0/analog_noesd_io[29]
+ chip_io_openframe_0/gpio_analog_pol[22] chip_io_openframe_0/gpio_dm0[16] w_692253_776670#
+ w_23367_710765# w_692355_547952# chip_io_openframe_0/gpio_analog_pol[23] w_23367_537965#
+ chip_io_openframe_0/area1_gpio_pad[15]/PAD_A_ESD_1_H w_21151_364074# chip_io_openframe_0/analog_noesd_io[3]
+ w_21253_966965# chip_io_openframe_0/gpio_out[3] chip_io_openframe_0/gpio_in_h[41]
+ chip_io_openframe_0/area1_gpio_pad[9]/PAD_A_ESD_1_H chip_io_openframe_0/gpio_analog_pol[24]
+ chip_io_openframe_0/gpio_inp_dis[42] w_459552_21253# w_694469_145352# w_692355_593152#
+ w_485565_1012355# w_694469_951752# w_694469_190352# w_638765_1012355# chip_io_openframe_0/gpio_vtrip_sel[6]
+ w_349952_23367# chip_io_openframe_0/gpio_inp_dis[27] w_692355_325552# chip_io_openframe_0/gpio_in_h[42]
+ chip_io_openframe_0/gpio_dm1[8] chip_io_openframe_0/sky130_ef_io__gpiov2_pad_wrapped_5/PAD_A_ESD_1_H
+ w_189869_23367# chip_io_openframe_0/gpio_slow_sel[36] w_694469_235552# w_21151_794074#
+ w_692355_683352# w_21253_194365# chip_io_openframe_0/gpio_holdover[37] w_694469_280552#
+ w_85874_1014469# chip_io_openframe_0/sky130_ef_io__gpiov2_pad_wrapped_5/HLD_H_N
+ chip_io_openframe_0/gpio_inp_dis[29] chip_io_openframe_0/gpio_in_h[43] chip_io_openframe_0/gpio_dm1[7]
+ chip_io_openframe_0/sky130_ef_io__gpiov2_pad_wrapped_12/PAD_A_ESD_1_H chip_io_openframe_0/gpio_out[6]
+ w_21253_624365# w_482474_1012253# chip_io_openframe_0/gpio_ib_mode_sel[27] chip_io_openframe_0/gpio_holdover[33]
+ w_295152_23367# w_635674_1012253# chip_io_openframe_0/gpio_dm2[23] w_349952_21253#
+ w_23367_578074# chip_io_openframe_0/analog_io[43] w_692253_551270# chip_io_openframe_0/gpio_dm1[6]
+ w_694469_370752# chip_io_openframe_0/area0_gpio_pad[3]/PAD_A_ESD_1_H w_189869_21253#
+ chip_io_openframe_0/gpio_holdover[18] chip_io_openframe_0/gpio_ib_mode_sel[29] chip_io_openframe_0/gpio_inp_dis[24]
+ chip_io_openframe_0/area1_gpio_pad[3]/HLD_H_N chip_io_openframe_0/gpio_vtrip_sel[20]
+ chip_io_openframe_0/sky130_ef_io__gpiov2_pad_wrapped_12/HLD_H_N chip_io_openframe_0/analog_io[23]
+ w_21151_277674# chip_io_openframe_0/area1_gpio_pad[2]/PAD_A_ESD_1_H chip_io_openframe_0/gpio_dm0[15]
+ chip_io_openframe_0/gpio_oeb[30] chip_io_openframe_0/gpio_dm1[5] chip_io_openframe_0/analog_noesd_io[8]
+ chip_io_openframe_0/gpio_slow_sel[19] chip_io_openframe_0/gpio_ib_mode_sel[28] chip_io_openframe_0/gpio_holdover[39]
+ w_692253_641470# chip_io_openframe_0/sky130_ef_io__gpiov2_pad_wrapped_8/PAD_A_ESD_1_H
+ w_692253_955070# w_295152_21253# w_294765_1014469# chip_io_openframe_0/gpio_dm0[38]
+ chip_io_openframe_0/sky130_ef_io__gpiov2_pad_wrapped_6/HLD_H_N w_21151_707674# chip_io_openframe_0/gpio_inp_dis[7]
+ w_23367_234474# chip_io_openframe_0/gpio_dm1[9] w_692355_100152# w_694469_776669#
+ chip_io_openframe_0/gpio_analog_pol[29] w_393474_1014469# w_21151_963874# chip_io_openframe_0/gpio_dm1[4]
+ chip_io_openframe_0/gpio_out[20] chip_io_openframe_0/sky130_ef_io__gpiov2_pad_wrapped_15/PAD_A_ESD_1_H
+ chip_io_openframe_0/gpio_inp_dis[3] chip_io_openframe_0/area1_gpio_pad[12]/PAD_A_ESD_1_H
+ w_692253_596470# chip_io_openframe_0/gpio_analog_en[9] chip_io_openframe_0/analog_io[27]
+ chip_io_openframe_0/sky130_ef_io__gpiov2_pad_wrapped_0/PAD_A_ESD_1_H w_692253_731670#
+ chip_io_openframe_0/gpio_loopback_one[4] w_21253_280765# chip_io_openframe_0/area1_gpio_pad[6]/PAD_A_ESD_1_H
+ w_692253_328870# chip_io_openframe_0/gpio_dm1[3] chip_io_openframe_0/analog_noesd_io[31]
+ w_23367_410365# chip_io_openframe_0/gpio_vtrip_sel[21] chip_io_openframe_0/gpio_oeb[33]
+ w_21253_710765# chip_io_openframe_0/area1_gpio_pad[0]/HLD_H_N chip_io_openframe_0/gpio_dm0[2]
+ w_294765_1012355# w_462869_23367# w_23367_237565# w_21253_537965# chip_io_openframe_0/sky130_ef_io__gpiov2_pad_wrapped_6/TIE_LO_ESD
+ chip_io_openframe_0/gpio_in[2] w_23367_664474# w_692253_686670# w_21151_191274#
+ w_692253_374070# chip_io_openframe_0/area1_gpio_pad[5]/TIE_LO_ESD chip_io_openframe_0/area1_gpio_pad[16]/PAD_A_ESD_1_H
+ chip_io_openframe_0/analog_noesd_io[5] chip_io_openframe_0/gpio_in[5] w_692355_145352#
+ w_21151_621274# chip_io_openframe_0/gpio_dm0[1] chip_io_openframe_0/analog_noesd_io[13]
+ chip_io_openframe_0/area1_gpio_pad[9]/HLD_H_N chip_io_openframe_0/gpio_analog_pol[28]
+ chip_io_openframe_0/sky130_ef_io__gpiov2_pad_wrapped_13/HLD_H_N w_692355_951752#
+ w_692355_190352# chip_io_openframe_0/gpio_dm2[22] chip_io_openframe_0/gpio_analog_sel[20]
+ chip_io_openframe_0/gpio_analog_en[39] chip_io_openframe_0/analog_io[4] w_694469_862552#
+ chip_io_openframe_0/gpio_in[8] w_88965_1014469# chip_io_openframe_0/gpio_loopback_one[12]
+ chip_io_openframe_0/area1_gpio_pad[0]/TIE_LO_ESD w_188674_1012253# chip_io_openframe_0/gpio_analog_sel[21]
+ chip_io_openframe_0/gpio_dm2[43] chip_io_openframe_0/gpio_oeb[36] chip_io_openframe_0/gpio_dm0[0]
+ chip_io_openframe_0/sky130_ef_io__gpiov2_pad_wrapped_18/PAD_A_ESD_1_H chip_io_openframe_0/gpio_loopback_one[32]
+ w_291674_1012253# chip_io_openframe_0/gpio_vtrip_sel[43] chip_io_openframe_0/gpio_out[42]
+ chip_io_openframe_0/sky130_ef_io__gpiov2_pad_wrapped_3/PAD_A_ESD_1_H w_462869_21253#
+ w_23367_667565# chip_io_openframe_0/analog_io[40] chip_io_openframe_0/gpio_out[2]
+ chip_io_openframe_0/gpio_inp_dis[43] w_692355_235552# w_694469_551269# chip_io_openframe_0/gpio_oeb[2]
+ chip_io_openframe_0/gpio_vtrip_sel[22] w_23367_320874# chip_io_openframe_0/gpio_loopback_one[37]
+ chip_io_openframe_0/area1_gpio_pad[8]/TIE_LO_ESD chip_io_openframe_0/gpio_analog_sel[22]
+ chip_io_openframe_0/area1_gpio_pad[7]/HLD_H_N w_692355_280552# chip_io_openframe_0/area0_gpio_pad[0]/PAD_A_ESD_1_H
+ chip_io_openframe_0/gpio_holdover[36] chip_io_openframe_0/gpio_dm0[14] chip_io_openframe_0/analog_noesd_io[17]
+ chip_io_openframe_0/gpio_inp_dis[9] chip_io_openframe_0/gpio_in[26] chip_io_openframe_0/gpio_inp_dis[28]
+ chip_io_openframe_0/gpio_analog_sel[23] chip_io_openframe_0/sky130_ef_io__gpiov2_pad_wrapped_10/PAD_A_ESD_1_H
+ chip_io_openframe_0/gpio_out[29] chip_io_openframe_0/gpio_out[27] chip_io_openframe_0/gpio_ib_mode_sel[3]
+ w_88965_1012355# chip_io_openframe_0/gpio_dm1[14] w_692253_103470# chip_io_openframe_0/sky130_ef_io__gpiov2_pad_wrapped_13/TIE_LO_ESD
+ w_140365_1014469# chip_io_openframe_0/sky130_ef_io__gpiov2_pad_wrapped_10/TIE_LO_ESD
+ w_694469_641469# w_694469_955069# chip_io_openframe_0/area1_gpio_pad[2]/TIE_LO_ESD
+ chip_io_openframe_0/gpio_analog_sel[24] chip_io_openframe_0/gpio_slow_sel[35] chip_io_openframe_0/gpio_slow_sel[25]
+ chip_io_openframe_0/gpio_analog_en[40] chip_io_openframe_0/analog_noesd_io[2] w_692355_370752#
+ chip_io_openframe_0/gpio_ib_mode_sel[2] chip_io_openframe_0/analog_noesd_io[36]
+ w_23367_323965# chip_io_openframe_0/gpio_dm2[27] chip_io_openframe_0/gpio_slow_sel[1]
+ chip_io_openframe_0/analog_io[11] w_23367_750874# chip_io_openframe_0/area0_gpio_pad[4]/PAD_A_ESD_1_H
+ chip_io_openframe_0/sky130_ef_io__gpiov2_pad_wrapped_3/HLD_H_N chip_io_openframe_0/analog_io[1]
+ chip_io_openframe_0/gpio_analog_sel[25] chip_io_openframe_0/gpio_oeb[5] chip_io_openframe_0/gpio_loopback_one[0]
+ chip_io_openframe_0/gpio_ib_mode_sel[13] chip_io_openframe_0/gpio_out[5] chip_io_openframe_0/gpio_loopback_one[15]
+ w_396565_1014469# chip_io_openframe_0/gpio_ib_mode_sel[1] chip_io_openframe_0/gpio_oeb[19]
+ chip_io_openframe_0/gpio_dm0[21] w_240074_1014469# chip_io_openframe_0/analog_io[24]
+ w_694469_596469# chip_io_openframe_0/gpio_slow_sel[26] w_23367_581165# chip_io_openframe_0/gpio_loopback_one[5]
+ chip_io_openframe_0/gpio_vtrip_sel[23] chip_io_openframe_0/gpio_analog_pol[10] chip_io_openframe_0/gpio_in[23]
+ w_694469_731669# chip_io_openframe_0/sky130_ef_io__gpiov2_pad_wrapped_7/HLD_H_N
+ chip_io_openframe_0/gpio_analog_sel[26] chip_io_openframe_0/gpio_analog_sel[5] chip_io_openframe_0/area1_gpio_pad[3]/PAD_A_ESD_1_H
+ chip_io_openframe_0/gpio_inp_dis[40] chip_io_openframe_0/sky130_ef_io__gpiov2_pad_wrapped_6/PAD_A_ESD_1_H
+ chip_io_openframe_0/gpio_in_h[2] chip_io_openframe_0/gpio_ib_mode_sel[0] w_21151_407274#
+ w_186552_23367# w_517669_23367# w_21151_534874# chip_io_openframe_0/gpio_analog_pol[1]
+ chip_io_openframe_0/gpio_out[24] w_85874_1012253# chip_io_openframe_0/gpio_inp_dis[6]
+ chip_io_openframe_0/analog_noesd_io[19] chip_io_openframe_0/gpio_analog_pol[40]
+ chip_io_openframe_0/gpio_in[29] w_694469_328869# w_140365_1012355# chip_io_openframe_0/gpio_analog_pol[11]
+ chip_io_openframe_0/gpio_inp_dis[25] chip_io_openframe_0/gpio_analog_sel[27] chip_io_openframe_0/gpio_slow_sel[27]
+ chip_io_openframe_0/sky130_ef_io__gpiov2_pad_wrapped_9/HLD_H_N w_692253_148670#
+ chip_io_openframe_0/gpio_analog_pol[41] chip_io_openframe_0/gpio_inp_dis[2] w_23367_753965#
+ chip_io_openframe_0/gpio_in[43] w_694469_686669# chip_io_openframe_0/gpio_dm2[21]
+ chip_io_openframe_0/gpio_analog_pol[12] chip_io_openframe_0/gpio_holdover[40] chip_io_openframe_0/sky130_ef_io__gpiov2_pad_wrapped_13/PAD_A_ESD_1_H
+ w_692253_193670# chip_io_openframe_0/gpio_analog_sel[9] chip_io_openframe_0/gpio_slow_sel[4]
+ chip_io_openframe_0/gpio_analog_en[41] chip_io_openframe_0/area1_gpio_pad[13]/PAD_A_ESD_1_H
+ w_694469_374069# chip_io_openframe_0/analog_io[9] chip_io_openframe_0/gpio_oeb[8]
+ w_396565_1012355# chip_io_openframe_0/gpio_analog_en[20] chip_io_openframe_0/analog_noesd_io[10]
+ chip_io_openframe_0/gpio_out[8] chip_io_openframe_0/gpio_analog_pol[42] chip_io_openframe_0/gpio_holdover[25]
+ chip_io_openframe_0/gpio_analog_pol[13] chip_io_openframe_0/area1_gpio_pad[7]/PAD_A_ESD_1_H
+ chip_io_openframe_0/gpio_dm2[42] w_21253_410365# w_694469_638152# chip_io_openframe_0/analog_noesd_io[33]
+ chip_io_openframe_0/sky130_ef_io__gpiov2_pad_wrapped_15/TIE_LO_ESD chip_io_openframe_0/gpio_inp_dis[16]
+ chip_io_openframe_0/gpio_in[20] w_186552_21253# chip_io_openframe_0/gpio_in_h[5]
+ w_517669_21253# w_21253_237565# chip_io_openframe_0/gpio_analog_pol[43] w_692253_238870#
+ w_23367_364074# chip_io_openframe_0/gpio_dm0[37] chip_io_openframe_0/gpio_analog_pol[14]
+ chip_io_openframe_0/gpio_vtrip_sel[24] chip_io_openframe_0/gpio_out[21] chip_io_openframe_0/sky130_ef_io__gpiov2_pad_wrapped_16/HLD_H_N
+ chip_io_openframe_0/analog_io[32] w_692253_283870# chip_io_openframe_0/gpio_loopback_one[18]
+ chip_io_openframe_0/sky130_ef_io__gpiov2_pad_wrapped_10/HLD_H_N chip_io_openframe_0/gpio_analog_sel[4]
+ chip_io_openframe_0/gpio_dm0[26] w_533874_1014469# chip_io_openframe_0/gpio_loopback_one[33]
+ chip_io_openframe_0/gpio_vtrip_sel[28] chip_io_openframe_0/gpio_analog_pol[0] chip_io_openframe_0/gpio_analog_pol[15]
+ chip_io_openframe_0/area1_gpio_pad[17]/PAD_A_ESD_1_H chip_io_openframe_0/analog_noesd_io[7]
+ chip_io_openframe_0/sky130_ef_io__gpiov2_pad_wrapped_9/PAD_A_ESD_1_H chip_io_openframe_0/gpio_holdover[16]
+ chip_io_openframe_0/gpio_out[10] chip_io_openframe_0/gpio_dm1[37] chip_io_openframe_0/gpio_slow_sel[28]
+ chip_io_openframe_0/sky130_ef_io__gpiov2_pad_wrapped_14/HLD_H_N w_694469_728352#
+ chip_io_openframe_0/gpio_in[40] chip_io_openframe_0/gpio_slow_sel[7] chip_io_openframe_0/analog_noesd_io[14]
+ w_692355_862552# chip_io_openframe_0/gpio_dm0[36] chip_io_openframe_0/gpio_dm1[13]
+ chip_io_openframe_0/gpio_oeb[32] chip_io_openframe_0/gpio_analog_sel[29] w_393474_1012253#
+ chip_io_openframe_0/gpio_vtrip_sel[8] w_694469_773352# chip_io_openframe_0/analog_io[6]
+ chip_io_openframe_0/gpio_inp_dis[35] chip_io_openframe_0/gpio_analog_pol[16] chip_io_openframe_0/gpio_loopback_one[10]
+ chip_io_openframe_0/area0_gpio_pad[0]/HLD_H_N chip_io_openframe_0/gpio_analog_en[42]
+ chip_io_openframe_0/gpio_slow_sel[38] w_23367_367165# chip_io_openframe_0/sky130_ef_io__gpiov2_pad_wrapped_12/TIE_LO_ESD
+ chip_io_openframe_0/gpio_dm2[26] w_21253_667565# chip_io_openframe_0/gpio_analog_en[21]
+ chip_io_openframe_0/gpio_dm1[36] chip_io_openframe_0/gpio_in_h[29] chip_io_openframe_0/gpio_dm2[13]
+ chip_io_openframe_0/sky130_ef_io__gpiov2_pad_wrapped_16/PAD_A_ESD_1_H w_23367_794074#
+ w_694469_103469# chip_io_openframe_0/gpio_in[0] chip_io_openframe_0/gpio_analog_pol[17]
+ chip_io_openframe_0/gpio_inp_dis[31] chip_io_openframe_0/gpio_in_h[8] chip_io_openframe_0/sky130_ef_io__gpiov2_pad_wrapped_1/PAD_A_ESD_1_H
+ chip_io_openframe_0/gpio_in_h[21] chip_io_openframe_0/gpio_dm0[35] w_137274_1014469#
+ w_353269_23367# chip_io_openframe_0/gpio_holdover[22] chip_io_openframe_0/gpio_dm0[20]
+ chip_io_openframe_0/area1_gpio_pad[10]/HLD_H_N chip_io_openframe_0/analog_io[41]
+ chip_io_openframe_0/gpio_ib_mode_sel[17] chip_io_openframe_0/gpio_holdover[35] chip_io_openframe_0/gpio_in[3]
+ chip_io_openframe_0/gpio_analog_pol[18] chip_io_openframe_0/gpio_inp_dis[13] chip_io_openframe_0/area0_gpio_pad[1]/PAD_A_ESD_1_H
+ chip_io_openframe_0/sky130_ef_io__gpiov2_pad_wrapped_17/HLD_H_N chip_io_openframe_0/analog_noesd_io[30]
+ chip_io_openframe_0/gpio_slow_sel[39] chip_io_openframe_0/analog_noesd_io[18] chip_io_openframe_0/gpio_loopback_one[1]
+ chip_io_openframe_0/area0_gpio_pad[2]/HLD_H_N chip_io_openframe_0/gpio_ib_mode_sel[12]
+ chip_io_openframe_0/gpio_analog_sel[3] chip_io_openframe_0/gpio_dm1[35] chip_io_openframe_0/area1_gpio_pad[11]/HLD_H_N
+ w_21151_578074# chip_io_openframe_0/gpio_dm0[41] chip_io_openframe_0/area1_gpio_pad[4]/HLD_H_N
+ chip_io_openframe_0/gpio_in[6] chip_io_openframe_0/gpio_in_h[22] chip_io_openframe_0/gpio_dm0[34]
+ chip_io_openframe_0/analog_io[21] chip_io_openframe_0/gpio_analog_en[29] vccd chip_io_openframe_0/gpio_oeb[35]
+ chip_io_openframe_0/analog_io[29] chip_io_openframe_0/gpio_loopback_one[6] w_243165_1014469#
+ chip_io_openframe_0/gpio_dm0[18] chip_io_openframe_0/gpio_out[43] chip_io_openframe_0/area0_gpio_pad[3]/HLD_H_N
+ chip_io_openframe_0/gpio_out[1] chip_io_openframe_0/area1_gpio_pad[0]/PAD_A_ESD_1_H
+ chip_io_openframe_0/area1_gpio_pad[8]/HLD_H_N chip_io_openframe_0/sky130_ef_io__gpiov2_pad_wrapped_0/HLD_H_N
+ chip_io_openframe_0/gpio_oeb[1] chip_io_openframe_0/gpio_dm2[35] chip_io_openframe_0/area0_gpio_pad[0]/TIE_LO_ESD
+ chip_io_openframe_0/gpio_analog_sel[28] w_23367_797165# chip_io_openframe_0/gpio_slow_sel[40]
+ chip_io_openframe_0/analog_noesd_io[4] chip_io_openframe_0/gpio_dm2[20] chip_io_openframe_0/gpio_dm1[34]
+ resetb w_21253_323965# chip_io_openframe_0/gpio_analog_pol[35] chip_io_openframe_0/gpio_in_h[32]
+ chip_io_openframe_0/gpio_in[27] chip_io_openframe_0/gpio_inp_dis[19] chip_io_openframe_0/gpio_in_h[23]
+ chip_io_openframe_0/area0_gpio_pad[4]/HLD_H_N chip_io_openframe_0/gpio_dm0[33] chip_io_openframe_0/sky130_ef_io__gpiov2_pad_wrapped_8/TIE_LO_ESD
+ chip_io_openframe_0/gpio_analog_en[43] chip_io_openframe_0/gpio_dm1[18] w_353269_21253#
+ chip_io_openframe_0/sky130_ef_io__gpiov2_pad_wrapped_4/HLD_H_N chip_io_openframe_0/area1_gpio_pad[13]/HLD_H_N
+ chip_io_openframe_0/area0_gpio_pad[1]/TIE_LO_ESD chip_io_openframe_0/analog_io[3]
+ chip_io_openframe_0/analog_io[12] chip_io_openframe_0/area0_gpio_pad[5]/PAD_A_ESD_1_H
+ w_23367_277674# chip_io_openframe_0/gpio_analog_en[22] w_694469_148669# chip_io_openframe_0/gpio_out[28]
+ chip_io_openframe_0/analog_io[37] chip_io_openframe_0/gpio_loopback_one[13] chip_io_openframe_0/gpio_dm2[41]
+ chip_io_openframe_0/sky130_ef_io__gpiov2_pad_wrapped_3/TIE_LO_ESD chip_io_openframe_0/gpio_out[9]
+ w_21253_581165# chip_io_openframe_0/gpio_dm2[34] w_694469_193669# chip_io_openframe_0/area0_gpio_pad[5]/HLD_H_N
+ vdda1 chip_io_openframe_0/area1_gpio_pad[10]/PAD_A_ESD_1_H chip_io_openframe_0/gpio_slow_sel[41]
+ chip_io_openframe_0/area1_gpio_pad[14]/HLD_H_N chip_io_openframe_0/sky130_ef_io__gpiov2_pad_wrapped_17/TIE_LO_ESD
+ chip_io_openframe_0/sky130_ef_io__gpiov2_pad_wrapped_8/HLD_H_N chip_io_openframe_0/analog_io[25]
+ chip_io_openframe_0/gpio_dm1[33] chip_io_openframe_0/gpio_loopback_one[9] w_23367_707674#
+ chip_io_openframe_0/gpio_dm2[18] w_21151_234474# chip_io_openframe_0/gpio_in_h[24]
+ chip_io_openframe_0/gpio_dm0[32] chip_io_openframe_0/gpio_holdover[19] chip_io_openframe_0/sky130_ef_io__gpiov2_pad_wrapped_4/PAD_A_ESD_1_H
+ chip_io_openframe_0/area1_gpio_pad[4]/PAD_A_ESD_1_H chip_io_openframe_0/gpio_vtrip_sel[26]
+ chip_io_openframe_0/sky130_ef_io__gpiov2_pad_wrapped_18/HLD_H_N vddio_2 chip_io_openframe_0/gpio_inp_dis[5]
+ chip_io_openframe_0/gpio_dm0[25] w_243165_1012355# vdda w_23367_963874# chip_io_openframe_0/gpio_analog_sel[2]
+ chip_io_openframe_0/gpio_out[40] chip_io_openframe_0/gpio_inp_dis[10] chip_io_openframe_0/gpio_slow_sel[0]
+ chip_io_openframe_0/analog_noesd_io[20] chip_io_openframe_0/area0_gpio_pad[3]/TIE_LO_ESD
+ chip_io_openframe_0/area1_gpio_pad[9]/TIE_LO_ESD chip_io_openframe_0/gpio_loopback_one[19]
+ chip_io_openframe_0/gpio_dm2[33] chip_io_openframe_0/area1_gpio_pad[12]/TIE_LO_ESD
+ chip_io_openframe_0/sky130_ef_io__gpiov2_pad_wrapped_0/TIE_LO_ESD gpio[23] chip_io_openframe_0/gpio_oeb[4]
+ chip_io_openframe_0/area1_gpio_pad[6]/HLD_H_N chip_io_openframe_0/gpio_slow_sel[42]
+ w_694469_238869# w_21253_753965# chip_io_openframe_0/gpio_dm1[32] chip_io_openframe_0/gpio_loopback_one[39]
+ chip_io_openframe_0/vssd1 chip_io_openframe_0/area0_gpio_pad[1]/HLD_H_N chip_io_openframe_0/gpio_inp_dis[1]
+ chip_io_openframe_0/gpio_analog_en[27] chip_io_openframe_0/area1_gpio_pad[10]/TIE_LO_ESD
+ chip_io_openframe_0/gpio_loopback_one[34] w_694469_283869# chip_io_openframe_0/gpio_in_h[35]
+ chip_io_openframe_0/gpio_in_h[25] chip_io_openframe_0/area1_gpio_pad[16]/HLD_H_N
+ chip_io_openframe_0/gpio_dm0[31] chip_io_openframe_0/analog_io[16] chip_io_openframe_0/gpio_loopback_one[20]
+ chip_io_openframe_0/vssd2 chip_io_openframe_0/gpio_dm1[12] w_692253_865870# chip_io_openframe_0/gpio_inp_dis[41]
+ chip_io_openframe_0/sky130_ef_io__gpiov2_pad_wrapped_11/PAD_A_ESD_1_H chip_io_openframe_0/gpio_in[24]
+ chip_io_openframe_0/gpio_oeb[9] chip_io_openframe_0/gpio_ib_mode_sel[19] chip_io_openframe_0/gpio_in[15]
+ chip_io_openframe_0/area1_gpio_pad[13]/TIE_LO_ESD w_536965_1014469# chip_io_openframe_0/gpio_holdover[5]
+ chip_io_openframe_0/area1_gpio_pad[5]/HLD_H_N chip_io_openframe_0/area1_gpio_pad[14]/PAD_A_ESD_1_H
+ chip_io_openframe_0/gpio_in_h[1] chip_io_openframe_0/gpio_analog_pol[34] w_298469_23367#
+ w_191765_1014469# chip_io_openframe_0/gpio_dm2[32] chip_io_openframe_0/gpio_inp_dis[26]
+ w_694469_547952# w_482474_1014469# chip_io_openframe_0/gpio_out[25] chip_io_openframe_0/area1_gpio_pad[17]/HLD_H_N
+ chip_io_openframe_0/area0_gpio_pad[2]/TIE_LO_ESD chip_io_openframe_0/gpio_out[31]
+ w_692355_638152# vssa2 chip_io_openframe_0/gpio_slow_sel[43] chip_io_openframe_0/analog_noesd_io[11]
+ gpio[8] chip_io_openframe_0/gpio_analog_sel[38] w_635674_1014469# chip_io_openframe_0/gpio_dm1[31]
+ chip_io_openframe_0/gpio_dm2[25] chip_io_openframe_0/gpio_dm2[12] chip_io_openframe_0/area1_gpio_pad[14]/TIE_LO_ESD
+ w_21151_664474# chip_io_openframe_0/area1_gpio_pad[8]/PAD_A_ESD_1_H chip_io_openframe_0/gpio_analog_en[23]
+ chip_io_openframe_0/gpio_loopback_one[17] vdda2 chip_io_openframe_0/gpio_holdover[1]
+ chip_io_openframe_0/area1_gpio_pad[3]/TIE_LO_ESD chip_io_openframe_0/analog_noesd_io[35]
+ chip_io_openframe_0/area1_gpio_pad[1]/HLD_H_N gpio[2] chip_io_openframe_0/gpio_in_h[26]
+ chip_io_openframe_0/sky130_ef_io__gpiov2_pad_wrapped_16/TIE_LO_ESD chip_io_openframe_0/area1_gpio_pad[1]/TIE_LO_ESD
+ chip_io_openframe_0/sky130_ef_io__gpiov2_pad_wrapped_5/TIE_LO_ESD w_23367_191274#
+ w_23367_966965# chip_io_openframe_0/gpio_slow_sel[37] vssd chip_io_openframe_0/gpio_holdover[41]
+ chip_io_openframe_0/analog_noesd_io[24] w_240074_1012253# chip_io_openframe_0/gpio_dm0[19]
+ gpio[40] w_408069_23367# chip_io_openframe_0/area1_gpio_pad[18]/HLD_H_N chip_io_openframe_0/gpio_vtrip_sel[10]
+ chip_io_openframe_0/sky130_ef_io__gpiov2_pad_wrapped_18/TIE_LO_ESD chip_io_openframe_0/analog_io[0]
+ chip_io_openframe_0/gpio_analog_sel[39] chip_io_openframe_0/gpio_out[14] chip_io_openframe_0/sky130_ef_io__gpiov2_pad_wrapped_11/HLD_H_N
+ chip_io_openframe_0/analog_io[34] chip_io_openframe_0/gpio_analog_sel[10] w_694469_593152#
+ chip_io_openframe_0/sky130_ef_io__gpiov2_pad_wrapped_11/TIE_LO_ESD chip_io_openframe_0/gpio_in[30]
+ chip_io_openframe_0/gpio_slow_sel[3] chip_io_openframe_0/gpio_dm2[31] gpio[30] w_23367_621274#
+ chip_io_openframe_0/gpio_slow_sel[2] gpio[35] chip_io_openframe_0/area1_gpio_pad[4]/TIE_LO_ESD
+ chip_io_openframe_0/gpio_holdover[26] chip_io_openframe_0/gpio_vtrip_sel[27] gpio[3]
+ chip_io_openframe_0/gpio_oeb[7] chip_io_openframe_0/gpio_dm1[30] gpio[17] chip_io_openframe_0/area1_gpio_pad[15]/HLD_H_N
+ chip_io_openframe_0/gpio_out[7] chip_io_openframe_0/gpio_analog_sel[1] vssd1 chip_io_openframe_0/gpio_dm0[40]
+ chip_io_openframe_0/analog_io[38] chip_io_openframe_0/gpio_vtrip_sel[7] chip_io_openframe_0/gpio_ib_mode_sel[16]
+ chip_io_openframe_0/gpio_analog_sel[40] gpio[29] chip_io_openframe_0/gpio_dm1[19]
+ chip_io_openframe_0/gpio_in_h[27] chip_io_openframe_0/gpio_dm0[29] w_692355_728352#
+ chip_io_openframe_0/sky130_ef_io__gpiov2_pad_wrapped_15/HLD_H_N chip_io_openframe_0/gpio_vtrip_sel[31]
+ chip_io_openframe_0/gpio_in[33] chip_io_openframe_0/gpio_loopback_one[40] gpio[27]
+ chip_io_openframe_0/gpio_inp_dis[17] chip_io_openframe_0/gpio_analog_sel[11] chip_io_openframe_0/sky130_ef_io__gpiov2_pad_wrapped_7/PAD_A_ESD_1_H
+ chip_io_openframe_0/gpio_analog_pol[8] chip_io_openframe_0/area1_gpio_pad[16]/TIE_LO_ESD
+ chip_io_openframe_0/area1_gpio_pad[18]/PAD_A_ESD_1_H chip_io_openframe_0/sky130_ef_io__gpiov2_pad_wrapped_1/TIE_LO_ESD
+ w_514352_23367# chip_io_openframe_0/sky130_ef_io__gpiov2_pad_wrapped_9/TIE_LO_ESD
+ w_694469_325552# chip_io_openframe_0/gpio_oeb[10] w_536965_1012355# w_692355_773352#
+ vssio_2 chip_io_openframe_0/gpio_dm0[17] chip_io_openframe_0/gpio_in[21] gpio[26]
+ chip_io_openframe_0/gpio_loopback_one[2] w_298469_21253# chip_io_openframe_0/gpio_inp_dis[34]
+ chip_io_openframe_0/gpio_in[12] w_191765_1012355# chip_io_openframe_0/analog_noesd_io[15]
+ chip_io_openframe_0/gpio_ib_mode_sel[11] chip_io_openframe_0/gpio_oeb[38] chip_io_openframe_0/gpio_in_h[4]
+ chip_io_openframe_0/area1_gpio_pad[15]/TIE_LO_ESD chip_io_openframe_0/sky130_ef_io__gpiov2_pad_wrapped_4/TIE_LO_ESD
+ chip_io_openframe_0/analog_io[8] chip_io_openframe_0/gpio_dm2[30] chip_io_openframe_0/gpio_in[36]
+ chip_io_openframe_0/sky130_ef_io__gpiov2_pad_wrapped_2/HLD_H_N chip_io_openframe_0/gpio_analog_sel[41]
+ chip_io_openframe_0/gpio_dm1[40] chip_io_openframe_0/gpio_out[22] chip_io_openframe_0/gpio_analog_sel[37]
+ chip_io_openframe_0/gpio_analog_sel[12] gpio[18] chip_io_openframe_0/area1_gpio_pad[17]/TIE_LO_ESD
+ gpio[14] chip_io_openframe_0/gpio_dm2[19] gpio[16] vccd1 w_694469_683352# chip_io_openframe_0/gpio_vtrip_sel[35]
+ w_21253_367165# chip_io_openframe_0/area0_gpio_pad[4]/TIE_LO_ESD chip_io_openframe_0/gpio_out[34]
+ chip_io_openframe_0/gpio_loopback_one[7] w_23367_194365# chip_io_openframe_0/analog_noesd_io[9]
+ gpio[39] w_21151_320874# chip_io_openframe_0/gpio_inp_dis[38] chip_io_openframe_0/gpio_analog_pol[33]
+ chip_io_openframe_0/gpio_analog_en[0] chip_io_openframe_0/gpio_in_h[9] chip_io_openframe_0/gpio_dm0[28]
+ chip_io_openframe_0/gpio_analog_en[18] chip_io_openframe_0/gpio_loopback_one[23]
+ chip_io_openframe_0/gpio_inp_dis[30] chip_io_openframe_0/gpio_dm1[17] vssd2 gpio[37]
+ gpio[38] chip_io_openframe_0/sky130_ef_io__gpiov2_pad_wrapped_14/PAD_A_ESD_1_H chip_io_openframe_0/gpio_holdover[17]
+ gpio[15] chip_io_openframe_0/gpio_vtrip_sel[25] chip_io_openframe_0/gpio_oeb[11]
+ chip_io_openframe_0/area1_gpio_pad[2]/HLD_H_N gpio[10] w_408069_21253# chip_io_openframe_0/gpio_analog_sel[42]
+ chip_io_openframe_0/gpio_analog_sel[13] chip_io_openframe_0/area1_gpio_pad[18]/TIE_LO_ESD
+ w_23367_624365# chip_io_openframe_0/gpio_slow_sel[18] chip_io_openframe_0/gpio_out[11]
+ gpio[6] vssa1 chip_io_openframe_0/gpio_inp_dis[23] chip_io_openframe_0/gpio_oeb[39]
+ chip_io_openframe_0/gpio_analog_en[24] chip_io_openframe_0/gpio_dm2[40] chip_io_openframe_0/gpio_holdover[34]
+ chip_io_openframe_0/gpio_in[41] gpio[20] chip_io_openframe_0/gpio_dm2[29] chip_io_openframe_0/area1_gpio_pad[6]/TIE_LO_ESD
+ chip_io_openframe_0/gpio_loopback_one[16] chip_io_openframe_0/gpio_slow_sel[6] chip_io_openframe_0/analog_io[42]
+ chip_io_openframe_0/gpio_out[4] chip_io_openframe_0/area0_gpio_pad[5]/TIE_LO_ESD
+ chip_io_openframe_0/gpio_oeb[31] chip_io_openframe_0/sky130_ef_io__gpiov2_pad_wrapped_7/TIE_LO_ESD
+ chip_io_openframe_0/gpio_analog_en[4] gpio[0] gpio[1] gpio[7] chip_io_openframe_0/gpio_ib_mode_sel[41]
+ chip_io_openframe_0/gpio_vtrip_sel[11] chip_io_openframe_0/gpio_dm2[17] chip_io_openframe_0/gpio_analog_en[28]
+ gpio[43] chip_io_openframe_0/gpio_analog_sel[43] gpio[34] chip_io_openframe_0/gpio_vtrip_sel[38]
+ chip_io_openframe_0/vssa chip_io_openframe_0/gpio_analog_sel[14] gpio[19] chip_io_openframe_0/analog_noesd_io[32]
+ chip_io_openframe_0/area0_gpio_pad[2]/PAD_A_ESD_1_H chip_io_openframe_0/gpio_holdover[38]
+ gpio[41] w_514352_21253# chip_io_openframe_0/gpio_holdover[30] w_533874_1012253#
+ chip_io_openframe_0/gpio_oeb[12] gpio[32] chip_io_openframe_0/gpio_dm0[24] chip_io_openframe_0/gpio_vtrip_sel[9]
+ chip_io_openframe_0/gpio_dm0[11] gpio[25] gpio[33] chip_io_openframe_0/area1_gpio_pad[11]/TIE_LO_ESD
+ chip_io_openframe_0/gpio_analog_sel[0] chip_io_openframe_0/gpio_oeb[40] chip_io_openframe_0/gpio_in_h[28]
+ chip_io_openframe_0/sky130_ef_io__gpiov2_pad_wrapped_14/TIE_LO_ESD w_404752_23367#
+ chip_io_openframe_0/analog_io[22] vssa1_2 chip_io_openframe_0/analog_io[31] gpio[22]
+ chip_io_openframe_0/gpio_holdover[23] chip_io_openframe_0/gpio_analog_en[8] chip_io_openframe_0/gpio_dm2[28]
+ chip_io_openframe_0/gpio_in_h[7] chip_io_openframe_0/sky130_ef_io__gpiov2_pad_wrapped_1/HLD_H_N
+ chip_io_openframe_0/gpio_analog_sel[15] gpio[4] VSUBS chip_io_openframe_0/porb_h
+ chip_io_openframe_0/gpio_analog_en[32] chip_io_openframe_0/gpio_analog_pol[7] gpio[24]
+ vssa chip_io_openframe_0/sky130_ef_io__gpiov2_pad_wrapped_2/TIE_LO_ESD gpio[11]
+ chip_io_openframe_0/area1_gpio_pad[7]/TIE_LO_ESD chip_io_openframe_0/vssio chip_io_openframe_0/area1_gpio_pad[12]/HLD_H_N
+ gpio[31] gpio[9] gpio[42] w_21253_797165# chip_io_openframe_0/FILLER_9/VSSIO_Q chip_io_openframe_0/gpio_out[19]
+ gpio[5] chip_io_openframe_0/vssa2 w_21151_750874# chip_io_openframe_0/vssa1 chip_io_openframe_0/area1_gpio_pad[1]/PAD_A_ESD_1_H
+ gpio[28] gpio[13] gpio[21] chip_io_openframe_0/gpio_ib_mode_sel[9] gpio[12] chip_io_openframe
.ends

