magic
tech sky130A
magscale 1 2
timestamp 1677507641
<< viali >>
rect 2145 7361 2179 7395
rect 7113 7361 7147 7395
rect 1593 6817 1627 6851
rect 3341 6817 3375 6851
rect 3985 6817 4019 6851
rect 5733 6817 5767 6851
rect 2145 6749 2179 6783
rect 3433 6749 3467 6783
rect 6653 6749 6687 6783
rect 7113 6749 7147 6783
rect 7205 6613 7239 6647
rect 4905 6341 4939 6375
rect 1869 6273 1903 6307
rect 2145 6273 2179 6307
rect 4537 6273 4571 6307
rect 4721 6273 4755 6307
rect 6561 6273 6595 6307
rect 1777 6205 1811 6239
rect 2605 6205 2639 6239
rect 3341 6205 3375 6239
rect 6469 5865 6503 5899
rect 2697 5729 2731 5763
rect 6101 5729 6135 5763
rect 1593 5661 1627 5695
rect 3985 5661 4019 5695
rect 5917 5661 5951 5695
rect 6009 5525 6043 5559
rect 1593 5185 1627 5219
rect 7113 4981 7147 5015
rect 2697 4709 2731 4743
rect 2237 4641 2271 4675
rect 2145 4573 2179 4607
rect 2237 4437 2271 4471
rect 2329 4097 2363 4131
rect 5273 4097 5307 4131
rect 5457 4097 5491 4131
rect 6745 4097 6779 4131
rect 5089 4029 5123 4063
rect 2973 3145 3007 3179
rect 2053 3009 2087 3043
rect 3157 3009 3191 3043
rect 5549 3009 5583 3043
rect 5733 3009 5767 3043
rect 4629 2941 4663 2975
rect 4997 2941 5031 2975
rect 2697 2805 2731 2839
rect 5549 2805 5583 2839
rect 6561 2805 6595 2839
rect 2881 2601 2915 2635
rect 2237 2465 2271 2499
rect 1593 2397 1627 2431
rect 5457 2397 5491 2431
rect 4077 2057 4111 2091
rect 3893 1921 3927 1955
rect 4905 1921 4939 1955
rect 2053 1853 2087 1887
rect 2421 1853 2455 1887
rect 4997 1853 5031 1887
rect 4353 1785 4387 1819
rect 5733 1717 5767 1751
rect 7297 1717 7331 1751
rect 1593 1513 1627 1547
rect 2605 1445 2639 1479
rect 3985 1377 4019 1411
rect 3065 1309 3099 1343
rect 7297 1309 7331 1343
rect 7205 1173 7239 1207
<< metal1 >>
rect 1104 7642 7820 7664
rect 1104 7590 3150 7642
rect 3202 7590 3214 7642
rect 3266 7590 3278 7642
rect 3330 7590 3342 7642
rect 3394 7590 3406 7642
rect 3458 7590 7150 7642
rect 7202 7590 7214 7642
rect 7266 7590 7278 7642
rect 7330 7590 7342 7642
rect 7394 7590 7406 7642
rect 7458 7590 7820 7642
rect 1104 7568 7820 7590
rect 2130 7392 2136 7404
rect 2091 7364 2136 7392
rect 2130 7352 2136 7364
rect 2188 7352 2194 7404
rect 6086 7352 6092 7404
rect 6144 7392 6150 7404
rect 7101 7395 7159 7401
rect 7101 7392 7113 7395
rect 6144 7364 7113 7392
rect 6144 7352 6150 7364
rect 7101 7361 7113 7364
rect 7147 7392 7159 7395
rect 7558 7392 7564 7404
rect 7147 7364 7564 7392
rect 7147 7361 7159 7364
rect 7101 7355 7159 7361
rect 7558 7352 7564 7364
rect 7616 7352 7622 7404
rect 1104 7098 7820 7120
rect 1104 7046 1150 7098
rect 1202 7046 1214 7098
rect 1266 7046 1278 7098
rect 1330 7046 1342 7098
rect 1394 7046 1406 7098
rect 1458 7046 5150 7098
rect 5202 7046 5214 7098
rect 5266 7046 5278 7098
rect 5330 7046 5342 7098
rect 5394 7046 5406 7098
rect 5458 7046 7820 7098
rect 1104 7024 7820 7046
rect 14 6876 20 6928
rect 72 6916 78 6928
rect 72 6888 2636 6916
rect 72 6876 78 6888
rect 1578 6848 1584 6860
rect 1539 6820 1584 6848
rect 1578 6808 1584 6820
rect 1636 6808 1642 6860
rect 2608 6848 2636 6888
rect 3329 6851 3387 6857
rect 3329 6848 3341 6851
rect 2608 6820 3341 6848
rect 3329 6817 3341 6820
rect 3375 6817 3387 6851
rect 3329 6811 3387 6817
rect 3602 6808 3608 6860
rect 3660 6848 3666 6860
rect 3973 6851 4031 6857
rect 3973 6848 3985 6851
rect 3660 6820 3985 6848
rect 3660 6808 3666 6820
rect 3973 6817 3985 6820
rect 4019 6817 4031 6851
rect 3973 6811 4031 6817
rect 5721 6851 5779 6857
rect 5721 6817 5733 6851
rect 5767 6848 5779 6851
rect 8386 6848 8392 6860
rect 5767 6820 8392 6848
rect 5767 6817 5779 6820
rect 5721 6811 5779 6817
rect 2130 6780 2136 6792
rect 2091 6752 2136 6780
rect 2130 6740 2136 6752
rect 2188 6740 2194 6792
rect 3421 6783 3479 6789
rect 3421 6749 3433 6783
rect 3467 6780 3479 6783
rect 5736 6780 5764 6811
rect 8386 6808 8392 6820
rect 8444 6808 8450 6860
rect 3467 6752 5764 6780
rect 6641 6783 6699 6789
rect 3467 6749 3479 6752
rect 3421 6743 3479 6749
rect 6641 6749 6653 6783
rect 6687 6780 6699 6783
rect 6822 6780 6828 6792
rect 6687 6752 6828 6780
rect 6687 6749 6699 6752
rect 6641 6743 6699 6749
rect 6822 6740 6828 6752
rect 6880 6780 6886 6792
rect 7101 6783 7159 6789
rect 7101 6780 7113 6783
rect 6880 6752 7113 6780
rect 6880 6740 6886 6752
rect 7101 6749 7113 6752
rect 7147 6749 7159 6783
rect 7101 6743 7159 6749
rect 7193 6647 7251 6653
rect 7193 6613 7205 6647
rect 7239 6644 7251 6647
rect 7558 6644 7564 6656
rect 7239 6616 7564 6644
rect 7239 6613 7251 6616
rect 7193 6607 7251 6613
rect 7558 6604 7564 6616
rect 7616 6604 7622 6656
rect 1104 6554 7820 6576
rect 1104 6502 3150 6554
rect 3202 6502 3214 6554
rect 3266 6502 3278 6554
rect 3330 6502 3342 6554
rect 3394 6502 3406 6554
rect 3458 6502 7150 6554
rect 7202 6502 7214 6554
rect 7266 6502 7278 6554
rect 7330 6502 7342 6554
rect 7394 6502 7406 6554
rect 7458 6502 7820 6554
rect 1104 6480 7820 6502
rect 3602 6332 3608 6384
rect 3660 6372 3666 6384
rect 4890 6372 4896 6384
rect 3660 6344 4752 6372
rect 4851 6344 4896 6372
rect 3660 6332 3666 6344
rect 1578 6264 1584 6316
rect 1636 6304 1642 6316
rect 1857 6307 1915 6313
rect 1857 6304 1869 6307
rect 1636 6276 1869 6304
rect 1636 6264 1642 6276
rect 1857 6273 1869 6276
rect 1903 6273 1915 6307
rect 1857 6267 1915 6273
rect 2133 6307 2191 6313
rect 2133 6273 2145 6307
rect 2179 6304 2191 6307
rect 4522 6304 4528 6316
rect 2179 6276 2774 6304
rect 4483 6276 4528 6304
rect 2179 6273 2191 6276
rect 2133 6267 2191 6273
rect 1762 6236 1768 6248
rect 1723 6208 1768 6236
rect 1762 6196 1768 6208
rect 1820 6196 1826 6248
rect 1946 6196 1952 6248
rect 2004 6236 2010 6248
rect 2593 6239 2651 6245
rect 2593 6236 2605 6239
rect 2004 6208 2605 6236
rect 2004 6196 2010 6208
rect 2593 6205 2605 6208
rect 2639 6205 2651 6239
rect 2746 6236 2774 6276
rect 4522 6264 4528 6276
rect 4580 6264 4586 6316
rect 4724 6313 4752 6344
rect 4890 6332 4896 6344
rect 4948 6332 4954 6384
rect 4709 6307 4767 6313
rect 4709 6273 4721 6307
rect 4755 6273 4767 6307
rect 6546 6304 6552 6316
rect 6459 6276 6552 6304
rect 4709 6267 4767 6273
rect 6546 6264 6552 6276
rect 6604 6304 6610 6316
rect 7742 6304 7748 6316
rect 6604 6276 7748 6304
rect 6604 6264 6610 6276
rect 7742 6264 7748 6276
rect 7800 6264 7806 6316
rect 3329 6239 3387 6245
rect 3329 6236 3341 6239
rect 2746 6208 3341 6236
rect 2593 6199 2651 6205
rect 3329 6205 3341 6208
rect 3375 6236 3387 6239
rect 5074 6236 5080 6248
rect 3375 6208 5080 6236
rect 3375 6205 3387 6208
rect 3329 6199 3387 6205
rect 5074 6196 5080 6208
rect 5132 6196 5138 6248
rect 1104 6010 7820 6032
rect 1104 5958 1150 6010
rect 1202 5958 1214 6010
rect 1266 5958 1278 6010
rect 1330 5958 1342 6010
rect 1394 5958 1406 6010
rect 1458 5958 5150 6010
rect 5202 5958 5214 6010
rect 5266 5958 5278 6010
rect 5330 5958 5342 6010
rect 5394 5958 5406 6010
rect 5458 5958 7820 6010
rect 1104 5936 7820 5958
rect 6457 5899 6515 5905
rect 6457 5865 6469 5899
rect 6503 5896 6515 5899
rect 7006 5896 7012 5908
rect 6503 5868 7012 5896
rect 6503 5865 6515 5868
rect 6457 5859 6515 5865
rect 7006 5856 7012 5868
rect 7064 5856 7070 5908
rect 2685 5763 2743 5769
rect 2685 5729 2697 5763
rect 2731 5760 2743 5763
rect 2774 5760 2780 5772
rect 2731 5732 2780 5760
rect 2731 5729 2743 5732
rect 2685 5723 2743 5729
rect 2774 5720 2780 5732
rect 2832 5760 2838 5772
rect 5534 5760 5540 5772
rect 2832 5732 5540 5760
rect 2832 5720 2838 5732
rect 5534 5720 5540 5732
rect 5592 5720 5598 5772
rect 6086 5760 6092 5772
rect 6047 5732 6092 5760
rect 6086 5720 6092 5732
rect 6144 5720 6150 5772
rect 1578 5692 1584 5704
rect 1539 5664 1584 5692
rect 1578 5652 1584 5664
rect 1636 5652 1642 5704
rect 3970 5692 3976 5704
rect 3931 5664 3976 5692
rect 3970 5652 3976 5664
rect 4028 5652 4034 5704
rect 5905 5695 5963 5701
rect 5905 5661 5917 5695
rect 5951 5692 5963 5695
rect 6822 5692 6828 5704
rect 5951 5664 6828 5692
rect 5951 5661 5963 5664
rect 5905 5655 5963 5661
rect 6822 5652 6828 5664
rect 6880 5652 6886 5704
rect 5994 5556 6000 5568
rect 5955 5528 6000 5556
rect 5994 5516 6000 5528
rect 6052 5516 6058 5568
rect 1104 5466 7820 5488
rect 1104 5414 3150 5466
rect 3202 5414 3214 5466
rect 3266 5414 3278 5466
rect 3330 5414 3342 5466
rect 3394 5414 3406 5466
rect 3458 5414 7150 5466
rect 7202 5414 7214 5466
rect 7266 5414 7278 5466
rect 7330 5414 7342 5466
rect 7394 5414 7406 5466
rect 7458 5414 7820 5466
rect 1104 5392 7820 5414
rect 2958 5312 2964 5364
rect 3016 5352 3022 5364
rect 3970 5352 3976 5364
rect 3016 5324 3976 5352
rect 3016 5312 3022 5324
rect 3970 5312 3976 5324
rect 4028 5352 4034 5364
rect 5810 5352 5816 5364
rect 4028 5324 5816 5352
rect 4028 5312 4034 5324
rect 5810 5312 5816 5324
rect 5868 5312 5874 5364
rect 658 5176 664 5228
rect 716 5216 722 5228
rect 1581 5219 1639 5225
rect 1581 5216 1593 5219
rect 716 5188 1593 5216
rect 716 5176 722 5188
rect 1581 5185 1593 5188
rect 1627 5216 1639 5219
rect 2130 5216 2136 5228
rect 1627 5188 2136 5216
rect 1627 5185 1639 5188
rect 1581 5179 1639 5185
rect 2130 5176 2136 5188
rect 2188 5176 2194 5228
rect 6822 4972 6828 5024
rect 6880 5012 6886 5024
rect 7101 5015 7159 5021
rect 7101 5012 7113 5015
rect 6880 4984 7113 5012
rect 6880 4972 6886 4984
rect 7101 4981 7113 4984
rect 7147 4981 7159 5015
rect 7101 4975 7159 4981
rect 1104 4922 7820 4944
rect 1104 4870 1150 4922
rect 1202 4870 1214 4922
rect 1266 4870 1278 4922
rect 1330 4870 1342 4922
rect 1394 4870 1406 4922
rect 1458 4870 5150 4922
rect 5202 4870 5214 4922
rect 5266 4870 5278 4922
rect 5330 4870 5342 4922
rect 5394 4870 5406 4922
rect 5458 4870 7820 4922
rect 1104 4848 7820 4870
rect 2685 4743 2743 4749
rect 2685 4709 2697 4743
rect 2731 4740 2743 4743
rect 5074 4740 5080 4752
rect 2731 4712 5080 4740
rect 2731 4709 2743 4712
rect 2685 4703 2743 4709
rect 5074 4700 5080 4712
rect 5132 4700 5138 4752
rect 1946 4632 1952 4684
rect 2004 4672 2010 4684
rect 2225 4675 2283 4681
rect 2225 4672 2237 4675
rect 2004 4644 2237 4672
rect 2004 4632 2010 4644
rect 2225 4641 2237 4644
rect 2271 4641 2283 4675
rect 2225 4635 2283 4641
rect 2130 4604 2136 4616
rect 2091 4576 2136 4604
rect 2130 4564 2136 4576
rect 2188 4564 2194 4616
rect 1578 4428 1584 4480
rect 1636 4468 1642 4480
rect 2225 4471 2283 4477
rect 2225 4468 2237 4471
rect 1636 4440 2237 4468
rect 1636 4428 1642 4440
rect 2225 4437 2237 4440
rect 2271 4437 2283 4471
rect 2225 4431 2283 4437
rect 1104 4378 7820 4400
rect 1104 4326 3150 4378
rect 3202 4326 3214 4378
rect 3266 4326 3278 4378
rect 3330 4326 3342 4378
rect 3394 4326 3406 4378
rect 3458 4326 7150 4378
rect 7202 4326 7214 4378
rect 7266 4326 7278 4378
rect 7330 4326 7342 4378
rect 7394 4326 7406 4378
rect 7458 4326 7820 4378
rect 1104 4304 7820 4326
rect 2317 4131 2375 4137
rect 2317 4097 2329 4131
rect 2363 4128 2375 4131
rect 2866 4128 2872 4140
rect 2363 4100 2872 4128
rect 2363 4097 2375 4100
rect 2317 4091 2375 4097
rect 2866 4088 2872 4100
rect 2924 4128 2930 4140
rect 4522 4128 4528 4140
rect 2924 4100 4528 4128
rect 2924 4088 2930 4100
rect 4522 4088 4528 4100
rect 4580 4088 4586 4140
rect 5261 4131 5319 4137
rect 5261 4097 5273 4131
rect 5307 4097 5319 4131
rect 5261 4091 5319 4097
rect 5445 4131 5503 4137
rect 5445 4097 5457 4131
rect 5491 4128 5503 4131
rect 6730 4128 6736 4140
rect 5491 4100 6736 4128
rect 5491 4097 5503 4100
rect 5445 4091 5503 4097
rect 1026 4020 1032 4072
rect 1084 4060 1090 4072
rect 5077 4063 5135 4069
rect 5077 4060 5089 4063
rect 1084 4032 5089 4060
rect 1084 4020 1090 4032
rect 5077 4029 5089 4032
rect 5123 4029 5135 4063
rect 5276 4060 5304 4091
rect 6730 4088 6736 4100
rect 6788 4088 6794 4140
rect 6546 4060 6552 4072
rect 5276 4032 6552 4060
rect 5077 4023 5135 4029
rect 6546 4020 6552 4032
rect 6604 4020 6610 4072
rect 1104 3834 7820 3856
rect 1104 3782 1150 3834
rect 1202 3782 1214 3834
rect 1266 3782 1278 3834
rect 1330 3782 1342 3834
rect 1394 3782 1406 3834
rect 1458 3782 5150 3834
rect 5202 3782 5214 3834
rect 5266 3782 5278 3834
rect 5330 3782 5342 3834
rect 5394 3782 5406 3834
rect 5458 3782 7820 3834
rect 1104 3760 7820 3782
rect 3050 3680 3056 3732
rect 3108 3720 3114 3732
rect 5994 3720 6000 3732
rect 3108 3692 6000 3720
rect 3108 3680 3114 3692
rect 5994 3680 6000 3692
rect 6052 3680 6058 3732
rect 1104 3290 7820 3312
rect 1104 3238 3150 3290
rect 3202 3238 3214 3290
rect 3266 3238 3278 3290
rect 3330 3238 3342 3290
rect 3394 3238 3406 3290
rect 3458 3238 7150 3290
rect 7202 3238 7214 3290
rect 7266 3238 7278 3290
rect 7330 3238 7342 3290
rect 7394 3238 7406 3290
rect 7458 3238 7820 3290
rect 1104 3216 7820 3238
rect 2961 3179 3019 3185
rect 2961 3145 2973 3179
rect 3007 3176 3019 3179
rect 4338 3176 4344 3188
rect 3007 3148 4344 3176
rect 3007 3145 3019 3148
rect 2961 3139 3019 3145
rect 4338 3136 4344 3148
rect 4396 3136 4402 3188
rect 3602 3068 3608 3120
rect 3660 3068 3666 3120
rect 2041 3043 2099 3049
rect 2041 3009 2053 3043
rect 2087 3040 2099 3043
rect 2774 3040 2780 3052
rect 2087 3012 2780 3040
rect 2087 3009 2099 3012
rect 2041 3003 2099 3009
rect 2774 3000 2780 3012
rect 2832 3000 2838 3052
rect 3145 3043 3203 3049
rect 3145 3009 3157 3043
rect 3191 3009 3203 3043
rect 5534 3040 5540 3052
rect 5495 3012 5540 3040
rect 3145 3003 3203 3009
rect 14 2864 20 2916
rect 72 2904 78 2916
rect 3050 2904 3056 2916
rect 72 2876 3056 2904
rect 72 2864 78 2876
rect 3050 2864 3056 2876
rect 3108 2864 3114 2916
rect 2685 2839 2743 2845
rect 2685 2805 2697 2839
rect 2731 2836 2743 2839
rect 2774 2836 2780 2848
rect 2731 2808 2780 2836
rect 2731 2805 2743 2808
rect 2685 2799 2743 2805
rect 2774 2796 2780 2808
rect 2832 2796 2838 2848
rect 3160 2836 3188 3003
rect 5534 3000 5540 3012
rect 5592 3000 5598 3052
rect 5721 3043 5779 3049
rect 5721 3009 5733 3043
rect 5767 3040 5779 3043
rect 5810 3040 5816 3052
rect 5767 3012 5816 3040
rect 5767 3009 5779 3012
rect 5721 3003 5779 3009
rect 5810 3000 5816 3012
rect 5868 3000 5874 3052
rect 3970 2932 3976 2984
rect 4028 2972 4034 2984
rect 4617 2975 4675 2981
rect 4617 2972 4629 2975
rect 4028 2944 4629 2972
rect 4028 2932 4034 2944
rect 4617 2941 4629 2944
rect 4663 2941 4675 2975
rect 4982 2972 4988 2984
rect 4943 2944 4988 2972
rect 4617 2935 4675 2941
rect 4982 2932 4988 2944
rect 5040 2932 5046 2984
rect 5000 2876 6592 2904
rect 5000 2836 5028 2876
rect 6564 2848 6592 2876
rect 5534 2836 5540 2848
rect 3160 2808 5028 2836
rect 5495 2808 5540 2836
rect 5534 2796 5540 2808
rect 5592 2796 5598 2848
rect 6546 2836 6552 2848
rect 6507 2808 6552 2836
rect 6546 2796 6552 2808
rect 6604 2796 6610 2848
rect 1104 2746 7820 2768
rect 1104 2694 1150 2746
rect 1202 2694 1214 2746
rect 1266 2694 1278 2746
rect 1330 2694 1342 2746
rect 1394 2694 1406 2746
rect 1458 2694 5150 2746
rect 5202 2694 5214 2746
rect 5266 2694 5278 2746
rect 5330 2694 5342 2746
rect 5394 2694 5406 2746
rect 5458 2694 7820 2746
rect 1104 2672 7820 2694
rect 2869 2635 2927 2641
rect 2869 2601 2881 2635
rect 2915 2632 2927 2635
rect 3050 2632 3056 2644
rect 2915 2604 3056 2632
rect 2915 2601 2927 2604
rect 2869 2595 2927 2601
rect 3050 2592 3056 2604
rect 3108 2592 3114 2644
rect 1302 2456 1308 2508
rect 1360 2496 1366 2508
rect 2225 2499 2283 2505
rect 2225 2496 2237 2499
rect 1360 2468 2237 2496
rect 1360 2456 1366 2468
rect 2225 2465 2237 2468
rect 2271 2465 2283 2499
rect 2225 2459 2283 2465
rect 1578 2428 1584 2440
rect 1539 2400 1584 2428
rect 1578 2388 1584 2400
rect 1636 2388 1642 2440
rect 4982 2388 4988 2440
rect 5040 2428 5046 2440
rect 5442 2428 5448 2440
rect 5040 2400 5448 2428
rect 5040 2388 5046 2400
rect 5442 2388 5448 2400
rect 5500 2388 5506 2440
rect 1104 2202 7820 2224
rect 1104 2150 3150 2202
rect 3202 2150 3214 2202
rect 3266 2150 3278 2202
rect 3330 2150 3342 2202
rect 3394 2150 3406 2202
rect 3458 2150 7150 2202
rect 7202 2150 7214 2202
rect 7266 2150 7278 2202
rect 7330 2150 7342 2202
rect 7394 2150 7406 2202
rect 7458 2150 7820 2202
rect 1104 2128 7820 2150
rect 2866 2048 2872 2100
rect 2924 2088 2930 2100
rect 2924 2060 4016 2088
rect 2924 2048 2930 2060
rect 3050 1980 3056 2032
rect 3108 1980 3114 2032
rect 3878 1952 3884 1964
rect 3839 1924 3884 1952
rect 3878 1912 3884 1924
rect 3936 1912 3942 1964
rect 3988 1952 4016 2060
rect 4062 2048 4068 2100
rect 4120 2088 4126 2100
rect 4120 2060 4165 2088
rect 4120 2048 4126 2060
rect 4893 1955 4951 1961
rect 4893 1952 4905 1955
rect 3988 1924 4905 1952
rect 4893 1921 4905 1924
rect 4939 1921 4951 1955
rect 4893 1915 4951 1921
rect 658 1844 664 1896
rect 716 1884 722 1896
rect 1302 1884 1308 1896
rect 716 1856 1308 1884
rect 716 1844 722 1856
rect 1302 1844 1308 1856
rect 1360 1884 1366 1896
rect 2041 1887 2099 1893
rect 2041 1884 2053 1887
rect 1360 1856 2053 1884
rect 1360 1844 1366 1856
rect 2041 1853 2053 1856
rect 2087 1853 2099 1887
rect 2041 1847 2099 1853
rect 2409 1887 2467 1893
rect 2409 1853 2421 1887
rect 2455 1884 2467 1887
rect 2958 1884 2964 1896
rect 2455 1856 2964 1884
rect 2455 1853 2467 1856
rect 2409 1847 2467 1853
rect 2958 1844 2964 1856
rect 3016 1844 3022 1896
rect 4985 1887 5043 1893
rect 4985 1853 4997 1887
rect 5031 1884 5043 1887
rect 8386 1884 8392 1896
rect 5031 1856 8392 1884
rect 5031 1853 5043 1856
rect 4985 1847 5043 1853
rect 8386 1844 8392 1856
rect 8444 1844 8450 1896
rect 4341 1819 4399 1825
rect 4341 1785 4353 1819
rect 4387 1816 4399 1819
rect 6454 1816 6460 1828
rect 4387 1788 6460 1816
rect 4387 1785 4399 1788
rect 4341 1779 4399 1785
rect 6454 1776 6460 1788
rect 6512 1776 6518 1828
rect 5721 1751 5779 1757
rect 5721 1717 5733 1751
rect 5767 1748 5779 1751
rect 5810 1748 5816 1760
rect 5767 1720 5816 1748
rect 5767 1717 5779 1720
rect 5721 1711 5779 1717
rect 5810 1708 5816 1720
rect 5868 1708 5874 1760
rect 7282 1748 7288 1760
rect 7243 1720 7288 1748
rect 7282 1708 7288 1720
rect 7340 1708 7346 1760
rect 1104 1658 7820 1680
rect 1104 1606 1150 1658
rect 1202 1606 1214 1658
rect 1266 1606 1278 1658
rect 1330 1606 1342 1658
rect 1394 1606 1406 1658
rect 1458 1606 5150 1658
rect 5202 1606 5214 1658
rect 5266 1606 5278 1658
rect 5330 1606 5342 1658
rect 5394 1606 5406 1658
rect 5458 1606 7820 1658
rect 1104 1584 7820 1606
rect 1486 1504 1492 1556
rect 1544 1544 1550 1556
rect 1581 1547 1639 1553
rect 1581 1544 1593 1547
rect 1544 1516 1593 1544
rect 1544 1504 1550 1516
rect 1581 1513 1593 1516
rect 1627 1544 1639 1547
rect 3970 1544 3976 1556
rect 1627 1516 3976 1544
rect 1627 1513 1639 1516
rect 1581 1507 1639 1513
rect 3970 1504 3976 1516
rect 4028 1504 4034 1556
rect 2593 1479 2651 1485
rect 2593 1445 2605 1479
rect 2639 1476 2651 1479
rect 3050 1476 3056 1488
rect 2639 1448 3056 1476
rect 2639 1445 2651 1448
rect 2593 1439 2651 1445
rect 3050 1436 3056 1448
rect 3108 1436 3114 1488
rect 2682 1368 2688 1420
rect 2740 1408 2746 1420
rect 3602 1408 3608 1420
rect 2740 1380 3608 1408
rect 2740 1368 2746 1380
rect 3068 1349 3096 1380
rect 3602 1368 3608 1380
rect 3660 1368 3666 1420
rect 3878 1368 3884 1420
rect 3936 1408 3942 1420
rect 3973 1411 4031 1417
rect 3973 1408 3985 1411
rect 3936 1380 3985 1408
rect 3936 1368 3942 1380
rect 3973 1377 3985 1380
rect 4019 1377 4031 1411
rect 3973 1371 4031 1377
rect 3053 1343 3111 1349
rect 3053 1309 3065 1343
rect 3099 1309 3111 1343
rect 7282 1340 7288 1352
rect 7195 1312 7288 1340
rect 3053 1303 3111 1309
rect 7282 1300 7288 1312
rect 7340 1340 7346 1352
rect 7742 1340 7748 1352
rect 7340 1312 7748 1340
rect 7340 1300 7346 1312
rect 7742 1300 7748 1312
rect 7800 1300 7806 1352
rect 7193 1207 7251 1213
rect 7193 1173 7205 1207
rect 7239 1204 7251 1207
rect 7834 1204 7840 1216
rect 7239 1176 7840 1204
rect 7239 1173 7251 1176
rect 7193 1167 7251 1173
rect 7834 1164 7840 1176
rect 7892 1164 7898 1216
rect 1104 1114 7820 1136
rect 1104 1062 3150 1114
rect 3202 1062 3214 1114
rect 3266 1062 3278 1114
rect 3330 1062 3342 1114
rect 3394 1062 3406 1114
rect 3458 1062 7150 1114
rect 7202 1062 7214 1114
rect 7266 1062 7278 1114
rect 7330 1062 7342 1114
rect 7394 1062 7406 1114
rect 7458 1062 7820 1114
rect 1104 1040 7820 1062
<< via1 >>
rect 3150 7590 3202 7642
rect 3214 7590 3266 7642
rect 3278 7590 3330 7642
rect 3342 7590 3394 7642
rect 3406 7590 3458 7642
rect 7150 7590 7202 7642
rect 7214 7590 7266 7642
rect 7278 7590 7330 7642
rect 7342 7590 7394 7642
rect 7406 7590 7458 7642
rect 2136 7395 2188 7404
rect 2136 7361 2145 7395
rect 2145 7361 2179 7395
rect 2179 7361 2188 7395
rect 2136 7352 2188 7361
rect 6092 7352 6144 7404
rect 7564 7352 7616 7404
rect 1150 7046 1202 7098
rect 1214 7046 1266 7098
rect 1278 7046 1330 7098
rect 1342 7046 1394 7098
rect 1406 7046 1458 7098
rect 5150 7046 5202 7098
rect 5214 7046 5266 7098
rect 5278 7046 5330 7098
rect 5342 7046 5394 7098
rect 5406 7046 5458 7098
rect 20 6876 72 6928
rect 1584 6851 1636 6860
rect 1584 6817 1593 6851
rect 1593 6817 1627 6851
rect 1627 6817 1636 6851
rect 1584 6808 1636 6817
rect 3608 6808 3660 6860
rect 2136 6783 2188 6792
rect 2136 6749 2145 6783
rect 2145 6749 2179 6783
rect 2179 6749 2188 6783
rect 2136 6740 2188 6749
rect 8392 6808 8444 6860
rect 6828 6740 6880 6792
rect 7564 6604 7616 6656
rect 3150 6502 3202 6554
rect 3214 6502 3266 6554
rect 3278 6502 3330 6554
rect 3342 6502 3394 6554
rect 3406 6502 3458 6554
rect 7150 6502 7202 6554
rect 7214 6502 7266 6554
rect 7278 6502 7330 6554
rect 7342 6502 7394 6554
rect 7406 6502 7458 6554
rect 3608 6332 3660 6384
rect 4896 6375 4948 6384
rect 1584 6264 1636 6316
rect 4528 6307 4580 6316
rect 1768 6239 1820 6248
rect 1768 6205 1777 6239
rect 1777 6205 1811 6239
rect 1811 6205 1820 6239
rect 1768 6196 1820 6205
rect 1952 6196 2004 6248
rect 4528 6273 4537 6307
rect 4537 6273 4571 6307
rect 4571 6273 4580 6307
rect 4528 6264 4580 6273
rect 4896 6341 4905 6375
rect 4905 6341 4939 6375
rect 4939 6341 4948 6375
rect 4896 6332 4948 6341
rect 6552 6307 6604 6316
rect 6552 6273 6561 6307
rect 6561 6273 6595 6307
rect 6595 6273 6604 6307
rect 6552 6264 6604 6273
rect 7748 6264 7800 6316
rect 5080 6196 5132 6248
rect 1150 5958 1202 6010
rect 1214 5958 1266 6010
rect 1278 5958 1330 6010
rect 1342 5958 1394 6010
rect 1406 5958 1458 6010
rect 5150 5958 5202 6010
rect 5214 5958 5266 6010
rect 5278 5958 5330 6010
rect 5342 5958 5394 6010
rect 5406 5958 5458 6010
rect 7012 5856 7064 5908
rect 2780 5720 2832 5772
rect 5540 5720 5592 5772
rect 6092 5763 6144 5772
rect 6092 5729 6101 5763
rect 6101 5729 6135 5763
rect 6135 5729 6144 5763
rect 6092 5720 6144 5729
rect 1584 5695 1636 5704
rect 1584 5661 1593 5695
rect 1593 5661 1627 5695
rect 1627 5661 1636 5695
rect 1584 5652 1636 5661
rect 3976 5695 4028 5704
rect 3976 5661 3985 5695
rect 3985 5661 4019 5695
rect 4019 5661 4028 5695
rect 3976 5652 4028 5661
rect 6828 5652 6880 5704
rect 6000 5559 6052 5568
rect 6000 5525 6009 5559
rect 6009 5525 6043 5559
rect 6043 5525 6052 5559
rect 6000 5516 6052 5525
rect 3150 5414 3202 5466
rect 3214 5414 3266 5466
rect 3278 5414 3330 5466
rect 3342 5414 3394 5466
rect 3406 5414 3458 5466
rect 7150 5414 7202 5466
rect 7214 5414 7266 5466
rect 7278 5414 7330 5466
rect 7342 5414 7394 5466
rect 7406 5414 7458 5466
rect 2964 5312 3016 5364
rect 3976 5312 4028 5364
rect 5816 5312 5868 5364
rect 664 5176 716 5228
rect 2136 5176 2188 5228
rect 6828 4972 6880 5024
rect 1150 4870 1202 4922
rect 1214 4870 1266 4922
rect 1278 4870 1330 4922
rect 1342 4870 1394 4922
rect 1406 4870 1458 4922
rect 5150 4870 5202 4922
rect 5214 4870 5266 4922
rect 5278 4870 5330 4922
rect 5342 4870 5394 4922
rect 5406 4870 5458 4922
rect 5080 4700 5132 4752
rect 1952 4632 2004 4684
rect 2136 4607 2188 4616
rect 2136 4573 2145 4607
rect 2145 4573 2179 4607
rect 2179 4573 2188 4607
rect 2136 4564 2188 4573
rect 1584 4428 1636 4480
rect 3150 4326 3202 4378
rect 3214 4326 3266 4378
rect 3278 4326 3330 4378
rect 3342 4326 3394 4378
rect 3406 4326 3458 4378
rect 7150 4326 7202 4378
rect 7214 4326 7266 4378
rect 7278 4326 7330 4378
rect 7342 4326 7394 4378
rect 7406 4326 7458 4378
rect 2872 4088 2924 4140
rect 4528 4088 4580 4140
rect 6736 4131 6788 4140
rect 1032 4020 1084 4072
rect 6736 4097 6745 4131
rect 6745 4097 6779 4131
rect 6779 4097 6788 4131
rect 6736 4088 6788 4097
rect 6552 4020 6604 4072
rect 1150 3782 1202 3834
rect 1214 3782 1266 3834
rect 1278 3782 1330 3834
rect 1342 3782 1394 3834
rect 1406 3782 1458 3834
rect 5150 3782 5202 3834
rect 5214 3782 5266 3834
rect 5278 3782 5330 3834
rect 5342 3782 5394 3834
rect 5406 3782 5458 3834
rect 3056 3680 3108 3732
rect 6000 3680 6052 3732
rect 3150 3238 3202 3290
rect 3214 3238 3266 3290
rect 3278 3238 3330 3290
rect 3342 3238 3394 3290
rect 3406 3238 3458 3290
rect 7150 3238 7202 3290
rect 7214 3238 7266 3290
rect 7278 3238 7330 3290
rect 7342 3238 7394 3290
rect 7406 3238 7458 3290
rect 4344 3136 4396 3188
rect 3608 3068 3660 3120
rect 2780 3000 2832 3052
rect 5540 3043 5592 3052
rect 20 2864 72 2916
rect 3056 2864 3108 2916
rect 2780 2796 2832 2848
rect 5540 3009 5549 3043
rect 5549 3009 5583 3043
rect 5583 3009 5592 3043
rect 5540 3000 5592 3009
rect 5816 3000 5868 3052
rect 3976 2932 4028 2984
rect 4988 2975 5040 2984
rect 4988 2941 4997 2975
rect 4997 2941 5031 2975
rect 5031 2941 5040 2975
rect 4988 2932 5040 2941
rect 5540 2839 5592 2848
rect 5540 2805 5549 2839
rect 5549 2805 5583 2839
rect 5583 2805 5592 2839
rect 5540 2796 5592 2805
rect 6552 2839 6604 2848
rect 6552 2805 6561 2839
rect 6561 2805 6595 2839
rect 6595 2805 6604 2839
rect 6552 2796 6604 2805
rect 1150 2694 1202 2746
rect 1214 2694 1266 2746
rect 1278 2694 1330 2746
rect 1342 2694 1394 2746
rect 1406 2694 1458 2746
rect 5150 2694 5202 2746
rect 5214 2694 5266 2746
rect 5278 2694 5330 2746
rect 5342 2694 5394 2746
rect 5406 2694 5458 2746
rect 3056 2592 3108 2644
rect 1308 2456 1360 2508
rect 1584 2431 1636 2440
rect 1584 2397 1593 2431
rect 1593 2397 1627 2431
rect 1627 2397 1636 2431
rect 1584 2388 1636 2397
rect 4988 2388 5040 2440
rect 5448 2431 5500 2440
rect 5448 2397 5457 2431
rect 5457 2397 5491 2431
rect 5491 2397 5500 2431
rect 5448 2388 5500 2397
rect 3150 2150 3202 2202
rect 3214 2150 3266 2202
rect 3278 2150 3330 2202
rect 3342 2150 3394 2202
rect 3406 2150 3458 2202
rect 7150 2150 7202 2202
rect 7214 2150 7266 2202
rect 7278 2150 7330 2202
rect 7342 2150 7394 2202
rect 7406 2150 7458 2202
rect 2872 2048 2924 2100
rect 3056 1980 3108 2032
rect 3884 1955 3936 1964
rect 3884 1921 3893 1955
rect 3893 1921 3927 1955
rect 3927 1921 3936 1955
rect 3884 1912 3936 1921
rect 4068 2091 4120 2100
rect 4068 2057 4077 2091
rect 4077 2057 4111 2091
rect 4111 2057 4120 2091
rect 4068 2048 4120 2057
rect 664 1844 716 1896
rect 1308 1844 1360 1896
rect 2964 1844 3016 1896
rect 8392 1844 8444 1896
rect 6460 1776 6512 1828
rect 5816 1708 5868 1760
rect 7288 1751 7340 1760
rect 7288 1717 7297 1751
rect 7297 1717 7331 1751
rect 7331 1717 7340 1751
rect 7288 1708 7340 1717
rect 1150 1606 1202 1658
rect 1214 1606 1266 1658
rect 1278 1606 1330 1658
rect 1342 1606 1394 1658
rect 1406 1606 1458 1658
rect 5150 1606 5202 1658
rect 5214 1606 5266 1658
rect 5278 1606 5330 1658
rect 5342 1606 5394 1658
rect 5406 1606 5458 1658
rect 1492 1504 1544 1556
rect 3976 1504 4028 1556
rect 3056 1436 3108 1488
rect 2688 1368 2740 1420
rect 3608 1368 3660 1420
rect 3884 1368 3936 1420
rect 7288 1343 7340 1352
rect 7288 1309 7297 1343
rect 7297 1309 7331 1343
rect 7331 1309 7340 1343
rect 7288 1300 7340 1309
rect 7748 1300 7800 1352
rect 7840 1164 7892 1216
rect 3150 1062 3202 1114
rect 3214 1062 3266 1114
rect 3278 1062 3330 1114
rect 3342 1062 3394 1114
rect 3406 1062 3458 1114
rect 7150 1062 7202 1114
rect 7214 1062 7266 1114
rect 7278 1062 7330 1114
rect 7342 1062 7394 1114
rect 7406 1062 7458 1114
<< metal2 >>
rect 18 8200 74 9000
rect 662 8200 718 9000
rect 1950 8200 2006 9000
rect 2148 8214 2544 8242
rect 32 6934 60 8200
rect 20 6928 72 6934
rect 20 6870 72 6876
rect 676 5234 704 8200
rect 1582 7576 1638 7585
rect 1582 7511 1638 7520
rect 1150 7100 1458 7109
rect 1150 7098 1156 7100
rect 1212 7098 1236 7100
rect 1292 7098 1316 7100
rect 1372 7098 1396 7100
rect 1452 7098 1458 7100
rect 1212 7046 1214 7098
rect 1394 7046 1396 7098
rect 1150 7044 1156 7046
rect 1212 7044 1236 7046
rect 1292 7044 1316 7046
rect 1372 7044 1396 7046
rect 1452 7044 1458 7046
rect 1150 7035 1458 7044
rect 1596 6866 1624 7511
rect 1584 6860 1636 6866
rect 1584 6802 1636 6808
rect 1584 6316 1636 6322
rect 1584 6258 1636 6264
rect 1150 6012 1458 6021
rect 1150 6010 1156 6012
rect 1212 6010 1236 6012
rect 1292 6010 1316 6012
rect 1372 6010 1396 6012
rect 1452 6010 1458 6012
rect 1212 5958 1214 6010
rect 1394 5958 1396 6010
rect 1150 5956 1156 5958
rect 1212 5956 1236 5958
rect 1292 5956 1316 5958
rect 1372 5956 1396 5958
rect 1452 5956 1458 5958
rect 1150 5947 1458 5956
rect 1596 5710 1624 6258
rect 1964 6254 1992 8200
rect 2148 7410 2176 8214
rect 2516 8106 2544 8214
rect 2594 8200 2650 9000
rect 2778 8936 2834 8945
rect 2778 8871 2834 8880
rect 2608 8106 2636 8200
rect 2516 8078 2636 8106
rect 2136 7404 2188 7410
rect 2136 7346 2188 7352
rect 2148 6798 2176 7346
rect 2136 6792 2188 6798
rect 2136 6734 2188 6740
rect 1768 6248 1820 6254
rect 1766 6216 1768 6225
rect 1952 6248 2004 6254
rect 1820 6216 1822 6225
rect 1952 6190 2004 6196
rect 1766 6151 1822 6160
rect 1584 5704 1636 5710
rect 1584 5646 1636 5652
rect 664 5228 716 5234
rect 664 5170 716 5176
rect 1596 5137 1624 5646
rect 1582 5128 1638 5137
rect 1582 5063 1638 5072
rect 1150 4924 1458 4933
rect 1150 4922 1156 4924
rect 1212 4922 1236 4924
rect 1292 4922 1316 4924
rect 1372 4922 1396 4924
rect 1452 4922 1458 4924
rect 1212 4870 1214 4922
rect 1394 4870 1396 4922
rect 1150 4868 1156 4870
rect 1212 4868 1236 4870
rect 1292 4868 1316 4870
rect 1372 4868 1396 4870
rect 1452 4868 1458 4870
rect 1150 4859 1458 4868
rect 1964 4690 1992 6190
rect 2792 5778 2820 8871
rect 3238 8200 3294 9000
rect 3344 8214 3648 8242
rect 3252 8106 3280 8200
rect 3344 8106 3372 8214
rect 3252 8078 3372 8106
rect 3150 7644 3458 7653
rect 3150 7642 3156 7644
rect 3212 7642 3236 7644
rect 3292 7642 3316 7644
rect 3372 7642 3396 7644
rect 3452 7642 3458 7644
rect 3212 7590 3214 7642
rect 3394 7590 3396 7642
rect 3150 7588 3156 7590
rect 3212 7588 3236 7590
rect 3292 7588 3316 7590
rect 3372 7588 3396 7590
rect 3452 7588 3458 7590
rect 3150 7579 3458 7588
rect 3620 6866 3648 8214
rect 4526 8200 4582 9000
rect 5170 8200 5226 9000
rect 5814 8200 5870 9000
rect 6826 8256 6882 8265
rect 7102 8200 7158 9000
rect 7746 8200 7802 9000
rect 8390 8200 8446 9000
rect 4066 6896 4122 6905
rect 3608 6860 3660 6866
rect 4066 6831 4122 6840
rect 3608 6802 3660 6808
rect 3150 6556 3458 6565
rect 3150 6554 3156 6556
rect 3212 6554 3236 6556
rect 3292 6554 3316 6556
rect 3372 6554 3396 6556
rect 3452 6554 3458 6556
rect 3212 6502 3214 6554
rect 3394 6502 3396 6554
rect 3150 6500 3156 6502
rect 3212 6500 3236 6502
rect 3292 6500 3316 6502
rect 3372 6500 3396 6502
rect 3452 6500 3458 6502
rect 3150 6491 3458 6500
rect 3620 6390 3648 6802
rect 3608 6384 3660 6390
rect 3608 6326 3660 6332
rect 2780 5772 2832 5778
rect 2780 5714 2832 5720
rect 3976 5704 4028 5710
rect 3976 5646 4028 5652
rect 3150 5468 3458 5477
rect 3150 5466 3156 5468
rect 3212 5466 3236 5468
rect 3292 5466 3316 5468
rect 3372 5466 3396 5468
rect 3452 5466 3458 5468
rect 3212 5414 3214 5466
rect 3394 5414 3396 5466
rect 3150 5412 3156 5414
rect 3212 5412 3236 5414
rect 3292 5412 3316 5414
rect 3372 5412 3396 5414
rect 3452 5412 3458 5414
rect 3150 5403 3458 5412
rect 3988 5370 4016 5646
rect 2964 5364 3016 5370
rect 2964 5306 3016 5312
rect 3976 5364 4028 5370
rect 3976 5306 4028 5312
rect 2136 5228 2188 5234
rect 2136 5170 2188 5176
rect 1952 4684 2004 4690
rect 1952 4626 2004 4632
rect 2148 4622 2176 5170
rect 2136 4616 2188 4622
rect 2136 4558 2188 4564
rect 1584 4480 1636 4486
rect 1584 4422 1636 4428
rect 1032 4072 1084 4078
rect 1032 4014 1084 4020
rect 20 2916 72 2922
rect 20 2858 72 2864
rect 32 800 60 2858
rect 664 1896 716 1902
rect 664 1838 716 1844
rect 676 800 704 1838
rect 18 0 74 800
rect 662 0 718 800
rect 1044 762 1072 4014
rect 1150 3836 1458 3845
rect 1150 3834 1156 3836
rect 1212 3834 1236 3836
rect 1292 3834 1316 3836
rect 1372 3834 1396 3836
rect 1452 3834 1458 3836
rect 1212 3782 1214 3834
rect 1394 3782 1396 3834
rect 1150 3780 1156 3782
rect 1212 3780 1236 3782
rect 1292 3780 1316 3782
rect 1372 3780 1396 3782
rect 1452 3780 1458 3782
rect 1150 3771 1458 3780
rect 1150 2748 1458 2757
rect 1150 2746 1156 2748
rect 1212 2746 1236 2748
rect 1292 2746 1316 2748
rect 1372 2746 1396 2748
rect 1452 2746 1458 2748
rect 1212 2694 1214 2746
rect 1394 2694 1396 2746
rect 1150 2692 1156 2694
rect 1212 2692 1236 2694
rect 1292 2692 1316 2694
rect 1372 2692 1396 2694
rect 1452 2692 1458 2694
rect 1150 2683 1458 2692
rect 1308 2508 1360 2514
rect 1308 2450 1360 2456
rect 1320 1902 1348 2450
rect 1596 2446 1624 4422
rect 2778 4176 2834 4185
rect 2778 4111 2834 4120
rect 2872 4140 2924 4146
rect 2792 3058 2820 4111
rect 2872 4082 2924 4088
rect 2884 3505 2912 4082
rect 2870 3496 2926 3505
rect 2870 3431 2926 3440
rect 2780 3052 2832 3058
rect 2780 2994 2832 3000
rect 2792 2938 2820 2994
rect 2792 2910 2912 2938
rect 2780 2848 2832 2854
rect 2780 2790 2832 2796
rect 1584 2440 1636 2446
rect 1584 2382 1636 2388
rect 1308 1896 1360 1902
rect 1308 1838 1360 1844
rect 1150 1660 1458 1669
rect 1150 1658 1156 1660
rect 1212 1658 1236 1660
rect 1292 1658 1316 1660
rect 1372 1658 1396 1660
rect 1452 1658 1458 1660
rect 1212 1606 1214 1658
rect 1394 1606 1396 1658
rect 1150 1604 1156 1606
rect 1212 1604 1236 1606
rect 1292 1604 1316 1606
rect 1372 1604 1396 1606
rect 1452 1604 1458 1606
rect 1150 1595 1458 1604
rect 1492 1556 1544 1562
rect 1492 1498 1544 1504
rect 1228 870 1348 898
rect 1228 762 1256 870
rect 1320 800 1348 870
rect 1044 734 1256 762
rect 1306 0 1362 800
rect 1504 785 1532 1498
rect 1596 1465 1624 2382
rect 2792 2145 2820 2790
rect 2778 2136 2834 2145
rect 2884 2106 2912 2910
rect 2778 2071 2834 2080
rect 2872 2100 2924 2106
rect 2872 2042 2924 2048
rect 2976 1902 3004 5306
rect 3150 4380 3458 4389
rect 3150 4378 3156 4380
rect 3212 4378 3236 4380
rect 3292 4378 3316 4380
rect 3372 4378 3396 4380
rect 3452 4378 3458 4380
rect 3212 4326 3214 4378
rect 3394 4326 3396 4378
rect 3150 4324 3156 4326
rect 3212 4324 3236 4326
rect 3292 4324 3316 4326
rect 3372 4324 3396 4326
rect 3452 4324 3458 4326
rect 3150 4315 3458 4324
rect 3056 3732 3108 3738
rect 3056 3674 3108 3680
rect 3068 2922 3096 3674
rect 3150 3292 3458 3301
rect 3150 3290 3156 3292
rect 3212 3290 3236 3292
rect 3292 3290 3316 3292
rect 3372 3290 3396 3292
rect 3452 3290 3458 3292
rect 3212 3238 3214 3290
rect 3394 3238 3396 3290
rect 3150 3236 3156 3238
rect 3212 3236 3236 3238
rect 3292 3236 3316 3238
rect 3372 3236 3396 3238
rect 3452 3236 3458 3238
rect 3150 3227 3458 3236
rect 3608 3120 3660 3126
rect 3608 3062 3660 3068
rect 3056 2916 3108 2922
rect 3056 2858 3108 2864
rect 3068 2650 3096 2858
rect 3056 2644 3108 2650
rect 3056 2586 3108 2592
rect 3150 2204 3458 2213
rect 3150 2202 3156 2204
rect 3212 2202 3236 2204
rect 3292 2202 3316 2204
rect 3372 2202 3396 2204
rect 3452 2202 3458 2204
rect 3212 2150 3214 2202
rect 3394 2150 3396 2202
rect 3150 2148 3156 2150
rect 3212 2148 3236 2150
rect 3292 2148 3316 2150
rect 3372 2148 3396 2150
rect 3452 2148 3458 2150
rect 3150 2139 3458 2148
rect 3056 2032 3108 2038
rect 3056 1974 3108 1980
rect 2964 1896 3016 1902
rect 2964 1838 3016 1844
rect 3068 1494 3096 1974
rect 3056 1488 3108 1494
rect 1582 1456 1638 1465
rect 3056 1430 3108 1436
rect 1582 1391 1638 1400
rect 2688 1420 2740 1426
rect 2688 1362 2740 1368
rect 2700 1306 2728 1362
rect 2608 1278 2728 1306
rect 2608 800 2636 1278
rect 3068 898 3096 1430
rect 3620 1426 3648 3062
rect 3976 2984 4028 2990
rect 3976 2926 4028 2932
rect 3884 1964 3936 1970
rect 3884 1906 3936 1912
rect 3896 1426 3924 1906
rect 3988 1562 4016 2926
rect 4080 2106 4108 6831
rect 4540 6474 4568 8200
rect 5184 7290 5212 8200
rect 5092 7262 5212 7290
rect 4894 6896 4950 6905
rect 4894 6831 4950 6840
rect 4356 6446 4568 6474
rect 4356 3194 4384 6446
rect 4908 6390 4936 6831
rect 4896 6384 4948 6390
rect 4896 6326 4948 6332
rect 4528 6316 4580 6322
rect 4528 6258 4580 6264
rect 4540 4146 4568 6258
rect 5092 6254 5120 7262
rect 5150 7100 5458 7109
rect 5150 7098 5156 7100
rect 5212 7098 5236 7100
rect 5292 7098 5316 7100
rect 5372 7098 5396 7100
rect 5452 7098 5458 7100
rect 5212 7046 5214 7098
rect 5394 7046 5396 7098
rect 5150 7044 5156 7046
rect 5212 7044 5236 7046
rect 5292 7044 5316 7046
rect 5372 7044 5396 7046
rect 5452 7044 5458 7046
rect 5150 7035 5458 7044
rect 5080 6248 5132 6254
rect 5080 6190 5132 6196
rect 5150 6012 5458 6021
rect 5150 6010 5156 6012
rect 5212 6010 5236 6012
rect 5292 6010 5316 6012
rect 5372 6010 5396 6012
rect 5452 6010 5458 6012
rect 5212 5958 5214 6010
rect 5394 5958 5396 6010
rect 5150 5956 5156 5958
rect 5212 5956 5236 5958
rect 5292 5956 5316 5958
rect 5372 5956 5396 5958
rect 5452 5956 5458 5958
rect 5150 5947 5458 5956
rect 5540 5772 5592 5778
rect 5540 5714 5592 5720
rect 5150 4924 5458 4933
rect 5150 4922 5156 4924
rect 5212 4922 5236 4924
rect 5292 4922 5316 4924
rect 5372 4922 5396 4924
rect 5452 4922 5458 4924
rect 5212 4870 5214 4922
rect 5394 4870 5396 4922
rect 5150 4868 5156 4870
rect 5212 4868 5236 4870
rect 5292 4868 5316 4870
rect 5372 4868 5396 4870
rect 5452 4868 5458 4870
rect 5150 4859 5458 4868
rect 5080 4752 5132 4758
rect 5080 4694 5132 4700
rect 4528 4140 4580 4146
rect 4528 4082 4580 4088
rect 4344 3188 4396 3194
rect 4344 3130 4396 3136
rect 4988 2984 5040 2990
rect 4988 2926 5040 2932
rect 5000 2446 5028 2926
rect 4988 2440 5040 2446
rect 4988 2382 5040 2388
rect 4068 2100 4120 2106
rect 4068 2042 4120 2048
rect 3976 1556 4028 1562
rect 3976 1498 4028 1504
rect 5092 1442 5120 4694
rect 5150 3836 5458 3845
rect 5150 3834 5156 3836
rect 5212 3834 5236 3836
rect 5292 3834 5316 3836
rect 5372 3834 5396 3836
rect 5452 3834 5458 3836
rect 5212 3782 5214 3834
rect 5394 3782 5396 3834
rect 5150 3780 5156 3782
rect 5212 3780 5236 3782
rect 5292 3780 5316 3782
rect 5372 3780 5396 3782
rect 5452 3780 5458 3782
rect 5150 3771 5458 3780
rect 5552 3058 5580 5714
rect 5828 5370 5856 8200
rect 6826 8191 6882 8200
rect 6092 7404 6144 7410
rect 6092 7346 6144 7352
rect 6104 5778 6132 7346
rect 6840 6798 6868 8191
rect 7116 7834 7144 8200
rect 7024 7806 7144 7834
rect 6828 6792 6880 6798
rect 6828 6734 6880 6740
rect 6552 6316 6604 6322
rect 6552 6258 6604 6264
rect 6092 5772 6144 5778
rect 6092 5714 6144 5720
rect 6000 5568 6052 5574
rect 6000 5510 6052 5516
rect 5816 5364 5868 5370
rect 5816 5306 5868 5312
rect 6012 3738 6040 5510
rect 6564 4078 6592 6258
rect 7024 5914 7052 7806
rect 7150 7644 7458 7653
rect 7150 7642 7156 7644
rect 7212 7642 7236 7644
rect 7292 7642 7316 7644
rect 7372 7642 7396 7644
rect 7452 7642 7458 7644
rect 7212 7590 7214 7642
rect 7394 7590 7396 7642
rect 7150 7588 7156 7590
rect 7212 7588 7236 7590
rect 7292 7588 7316 7590
rect 7372 7588 7396 7590
rect 7452 7588 7458 7590
rect 7150 7579 7458 7588
rect 7562 7576 7618 7585
rect 7562 7511 7618 7520
rect 7576 7410 7604 7511
rect 7564 7404 7616 7410
rect 7564 7346 7616 7352
rect 7564 6656 7616 6662
rect 7564 6598 7616 6604
rect 7150 6556 7458 6565
rect 7150 6554 7156 6556
rect 7212 6554 7236 6556
rect 7292 6554 7316 6556
rect 7372 6554 7396 6556
rect 7452 6554 7458 6556
rect 7212 6502 7214 6554
rect 7394 6502 7396 6554
rect 7150 6500 7156 6502
rect 7212 6500 7236 6502
rect 7292 6500 7316 6502
rect 7372 6500 7396 6502
rect 7452 6500 7458 6502
rect 7150 6491 7458 6500
rect 7012 5908 7064 5914
rect 7012 5850 7064 5856
rect 6828 5704 6880 5710
rect 6828 5646 6880 5652
rect 6840 5030 6868 5646
rect 7576 5545 7604 6598
rect 7760 6322 7788 8200
rect 8404 6866 8432 8200
rect 8392 6860 8444 6866
rect 8392 6802 8444 6808
rect 7748 6316 7800 6322
rect 7748 6258 7800 6264
rect 7562 5536 7618 5545
rect 7150 5468 7458 5477
rect 7562 5471 7618 5480
rect 7150 5466 7156 5468
rect 7212 5466 7236 5468
rect 7292 5466 7316 5468
rect 7372 5466 7396 5468
rect 7452 5466 7458 5468
rect 7212 5414 7214 5466
rect 7394 5414 7396 5466
rect 7150 5412 7156 5414
rect 7212 5412 7236 5414
rect 7292 5412 7316 5414
rect 7372 5412 7396 5414
rect 7452 5412 7458 5414
rect 7150 5403 7458 5412
rect 6828 5024 6880 5030
rect 6828 4966 6880 4972
rect 6840 4865 6868 4966
rect 6826 4856 6882 4865
rect 6826 4791 6882 4800
rect 7150 4380 7458 4389
rect 7150 4378 7156 4380
rect 7212 4378 7236 4380
rect 7292 4378 7316 4380
rect 7372 4378 7396 4380
rect 7452 4378 7458 4380
rect 7212 4326 7214 4378
rect 7394 4326 7396 4378
rect 7150 4324 7156 4326
rect 7212 4324 7236 4326
rect 7292 4324 7316 4326
rect 7372 4324 7396 4326
rect 7452 4324 7458 4326
rect 7150 4315 7458 4324
rect 6734 4176 6790 4185
rect 6734 4111 6736 4120
rect 6788 4111 6790 4120
rect 6736 4082 6788 4088
rect 6552 4072 6604 4078
rect 6552 4014 6604 4020
rect 6000 3732 6052 3738
rect 6000 3674 6052 3680
rect 7150 3292 7458 3301
rect 7150 3290 7156 3292
rect 7212 3290 7236 3292
rect 7292 3290 7316 3292
rect 7372 3290 7396 3292
rect 7452 3290 7458 3292
rect 7212 3238 7214 3290
rect 7394 3238 7396 3290
rect 7150 3236 7156 3238
rect 7212 3236 7236 3238
rect 7292 3236 7316 3238
rect 7372 3236 7396 3238
rect 7452 3236 7458 3238
rect 7150 3227 7458 3236
rect 5540 3052 5592 3058
rect 5540 2994 5592 3000
rect 5816 3052 5868 3058
rect 5816 2994 5868 3000
rect 5540 2848 5592 2854
rect 5540 2790 5592 2796
rect 5150 2748 5458 2757
rect 5150 2746 5156 2748
rect 5212 2746 5236 2748
rect 5292 2746 5316 2748
rect 5372 2746 5396 2748
rect 5452 2746 5458 2748
rect 5212 2694 5214 2746
rect 5394 2694 5396 2746
rect 5150 2692 5156 2694
rect 5212 2692 5236 2694
rect 5292 2692 5316 2694
rect 5372 2692 5396 2694
rect 5452 2692 5458 2694
rect 5150 2683 5458 2692
rect 5448 2440 5500 2446
rect 5446 2408 5448 2417
rect 5500 2408 5502 2417
rect 5446 2343 5502 2352
rect 5150 1660 5458 1669
rect 5150 1658 5156 1660
rect 5212 1658 5236 1660
rect 5292 1658 5316 1660
rect 5372 1658 5396 1660
rect 5452 1658 5458 1660
rect 5212 1606 5214 1658
rect 5394 1606 5396 1658
rect 5150 1604 5156 1606
rect 5212 1604 5236 1606
rect 5292 1604 5316 1606
rect 5372 1604 5396 1606
rect 5452 1604 5458 1606
rect 5150 1595 5458 1604
rect 5552 1465 5580 2790
rect 5828 1766 5856 2994
rect 6552 2848 6604 2854
rect 6550 2816 6552 2825
rect 6604 2816 6606 2825
rect 6550 2751 6606 2760
rect 7150 2204 7458 2213
rect 7150 2202 7156 2204
rect 7212 2202 7236 2204
rect 7292 2202 7316 2204
rect 7372 2202 7396 2204
rect 7452 2202 7458 2204
rect 7212 2150 7214 2202
rect 7394 2150 7396 2202
rect 7150 2148 7156 2150
rect 7212 2148 7236 2150
rect 7292 2148 7316 2150
rect 7372 2148 7396 2150
rect 7452 2148 7458 2150
rect 7150 2139 7458 2148
rect 8392 1896 8444 1902
rect 8392 1838 8444 1844
rect 6460 1828 6512 1834
rect 6460 1770 6512 1776
rect 5816 1760 5868 1766
rect 5816 1702 5868 1708
rect 5538 1456 5594 1465
rect 3608 1420 3660 1426
rect 3608 1362 3660 1368
rect 3884 1420 3936 1426
rect 5092 1414 5212 1442
rect 3884 1362 3936 1368
rect 3150 1116 3458 1125
rect 3150 1114 3156 1116
rect 3212 1114 3236 1116
rect 3292 1114 3316 1116
rect 3372 1114 3396 1116
rect 3452 1114 3458 1116
rect 3212 1062 3214 1114
rect 3394 1062 3396 1114
rect 3150 1060 3156 1062
rect 3212 1060 3236 1062
rect 3292 1060 3316 1062
rect 3372 1060 3396 1062
rect 3452 1060 3458 1062
rect 3150 1051 3458 1060
rect 3068 870 3280 898
rect 3252 800 3280 870
rect 3896 800 3924 1362
rect 5184 800 5212 1414
rect 5538 1391 5594 1400
rect 5828 800 5856 1702
rect 6472 800 6500 1770
rect 7288 1760 7340 1766
rect 7288 1702 7340 1708
rect 7300 1358 7328 1702
rect 7288 1352 7340 1358
rect 7288 1294 7340 1300
rect 7748 1352 7800 1358
rect 7748 1294 7800 1300
rect 7150 1116 7458 1125
rect 7150 1114 7156 1116
rect 7212 1114 7236 1116
rect 7292 1114 7316 1116
rect 7372 1114 7396 1116
rect 7452 1114 7458 1116
rect 7212 1062 7214 1114
rect 7394 1062 7396 1114
rect 7150 1060 7156 1062
rect 7212 1060 7236 1062
rect 7292 1060 7316 1062
rect 7372 1060 7396 1062
rect 7452 1060 7458 1062
rect 7150 1051 7458 1060
rect 7760 800 7788 1294
rect 7840 1216 7892 1222
rect 7840 1158 7892 1164
rect 1490 776 1546 785
rect 1490 711 1546 720
rect 2594 0 2650 800
rect 3238 0 3294 800
rect 3882 0 3938 800
rect 5170 0 5226 800
rect 5814 0 5870 800
rect 6458 0 6514 800
rect 7746 0 7802 800
rect 7852 105 7880 1158
rect 8404 800 8432 1838
rect 7838 96 7894 105
rect 7838 31 7894 40
rect 8390 0 8446 800
<< via2 >>
rect 1582 7520 1638 7576
rect 1156 7098 1212 7100
rect 1236 7098 1292 7100
rect 1316 7098 1372 7100
rect 1396 7098 1452 7100
rect 1156 7046 1202 7098
rect 1202 7046 1212 7098
rect 1236 7046 1266 7098
rect 1266 7046 1278 7098
rect 1278 7046 1292 7098
rect 1316 7046 1330 7098
rect 1330 7046 1342 7098
rect 1342 7046 1372 7098
rect 1396 7046 1406 7098
rect 1406 7046 1452 7098
rect 1156 7044 1212 7046
rect 1236 7044 1292 7046
rect 1316 7044 1372 7046
rect 1396 7044 1452 7046
rect 1156 6010 1212 6012
rect 1236 6010 1292 6012
rect 1316 6010 1372 6012
rect 1396 6010 1452 6012
rect 1156 5958 1202 6010
rect 1202 5958 1212 6010
rect 1236 5958 1266 6010
rect 1266 5958 1278 6010
rect 1278 5958 1292 6010
rect 1316 5958 1330 6010
rect 1330 5958 1342 6010
rect 1342 5958 1372 6010
rect 1396 5958 1406 6010
rect 1406 5958 1452 6010
rect 1156 5956 1212 5958
rect 1236 5956 1292 5958
rect 1316 5956 1372 5958
rect 1396 5956 1452 5958
rect 2778 8880 2834 8936
rect 1766 6196 1768 6216
rect 1768 6196 1820 6216
rect 1820 6196 1822 6216
rect 1766 6160 1822 6196
rect 1582 5072 1638 5128
rect 1156 4922 1212 4924
rect 1236 4922 1292 4924
rect 1316 4922 1372 4924
rect 1396 4922 1452 4924
rect 1156 4870 1202 4922
rect 1202 4870 1212 4922
rect 1236 4870 1266 4922
rect 1266 4870 1278 4922
rect 1278 4870 1292 4922
rect 1316 4870 1330 4922
rect 1330 4870 1342 4922
rect 1342 4870 1372 4922
rect 1396 4870 1406 4922
rect 1406 4870 1452 4922
rect 1156 4868 1212 4870
rect 1236 4868 1292 4870
rect 1316 4868 1372 4870
rect 1396 4868 1452 4870
rect 3156 7642 3212 7644
rect 3236 7642 3292 7644
rect 3316 7642 3372 7644
rect 3396 7642 3452 7644
rect 3156 7590 3202 7642
rect 3202 7590 3212 7642
rect 3236 7590 3266 7642
rect 3266 7590 3278 7642
rect 3278 7590 3292 7642
rect 3316 7590 3330 7642
rect 3330 7590 3342 7642
rect 3342 7590 3372 7642
rect 3396 7590 3406 7642
rect 3406 7590 3452 7642
rect 3156 7588 3212 7590
rect 3236 7588 3292 7590
rect 3316 7588 3372 7590
rect 3396 7588 3452 7590
rect 6826 8200 6882 8256
rect 4066 6840 4122 6896
rect 3156 6554 3212 6556
rect 3236 6554 3292 6556
rect 3316 6554 3372 6556
rect 3396 6554 3452 6556
rect 3156 6502 3202 6554
rect 3202 6502 3212 6554
rect 3236 6502 3266 6554
rect 3266 6502 3278 6554
rect 3278 6502 3292 6554
rect 3316 6502 3330 6554
rect 3330 6502 3342 6554
rect 3342 6502 3372 6554
rect 3396 6502 3406 6554
rect 3406 6502 3452 6554
rect 3156 6500 3212 6502
rect 3236 6500 3292 6502
rect 3316 6500 3372 6502
rect 3396 6500 3452 6502
rect 3156 5466 3212 5468
rect 3236 5466 3292 5468
rect 3316 5466 3372 5468
rect 3396 5466 3452 5468
rect 3156 5414 3202 5466
rect 3202 5414 3212 5466
rect 3236 5414 3266 5466
rect 3266 5414 3278 5466
rect 3278 5414 3292 5466
rect 3316 5414 3330 5466
rect 3330 5414 3342 5466
rect 3342 5414 3372 5466
rect 3396 5414 3406 5466
rect 3406 5414 3452 5466
rect 3156 5412 3212 5414
rect 3236 5412 3292 5414
rect 3316 5412 3372 5414
rect 3396 5412 3452 5414
rect 1156 3834 1212 3836
rect 1236 3834 1292 3836
rect 1316 3834 1372 3836
rect 1396 3834 1452 3836
rect 1156 3782 1202 3834
rect 1202 3782 1212 3834
rect 1236 3782 1266 3834
rect 1266 3782 1278 3834
rect 1278 3782 1292 3834
rect 1316 3782 1330 3834
rect 1330 3782 1342 3834
rect 1342 3782 1372 3834
rect 1396 3782 1406 3834
rect 1406 3782 1452 3834
rect 1156 3780 1212 3782
rect 1236 3780 1292 3782
rect 1316 3780 1372 3782
rect 1396 3780 1452 3782
rect 1156 2746 1212 2748
rect 1236 2746 1292 2748
rect 1316 2746 1372 2748
rect 1396 2746 1452 2748
rect 1156 2694 1202 2746
rect 1202 2694 1212 2746
rect 1236 2694 1266 2746
rect 1266 2694 1278 2746
rect 1278 2694 1292 2746
rect 1316 2694 1330 2746
rect 1330 2694 1342 2746
rect 1342 2694 1372 2746
rect 1396 2694 1406 2746
rect 1406 2694 1452 2746
rect 1156 2692 1212 2694
rect 1236 2692 1292 2694
rect 1316 2692 1372 2694
rect 1396 2692 1452 2694
rect 2778 4120 2834 4176
rect 2870 3440 2926 3496
rect 1156 1658 1212 1660
rect 1236 1658 1292 1660
rect 1316 1658 1372 1660
rect 1396 1658 1452 1660
rect 1156 1606 1202 1658
rect 1202 1606 1212 1658
rect 1236 1606 1266 1658
rect 1266 1606 1278 1658
rect 1278 1606 1292 1658
rect 1316 1606 1330 1658
rect 1330 1606 1342 1658
rect 1342 1606 1372 1658
rect 1396 1606 1406 1658
rect 1406 1606 1452 1658
rect 1156 1604 1212 1606
rect 1236 1604 1292 1606
rect 1316 1604 1372 1606
rect 1396 1604 1452 1606
rect 2778 2080 2834 2136
rect 3156 4378 3212 4380
rect 3236 4378 3292 4380
rect 3316 4378 3372 4380
rect 3396 4378 3452 4380
rect 3156 4326 3202 4378
rect 3202 4326 3212 4378
rect 3236 4326 3266 4378
rect 3266 4326 3278 4378
rect 3278 4326 3292 4378
rect 3316 4326 3330 4378
rect 3330 4326 3342 4378
rect 3342 4326 3372 4378
rect 3396 4326 3406 4378
rect 3406 4326 3452 4378
rect 3156 4324 3212 4326
rect 3236 4324 3292 4326
rect 3316 4324 3372 4326
rect 3396 4324 3452 4326
rect 3156 3290 3212 3292
rect 3236 3290 3292 3292
rect 3316 3290 3372 3292
rect 3396 3290 3452 3292
rect 3156 3238 3202 3290
rect 3202 3238 3212 3290
rect 3236 3238 3266 3290
rect 3266 3238 3278 3290
rect 3278 3238 3292 3290
rect 3316 3238 3330 3290
rect 3330 3238 3342 3290
rect 3342 3238 3372 3290
rect 3396 3238 3406 3290
rect 3406 3238 3452 3290
rect 3156 3236 3212 3238
rect 3236 3236 3292 3238
rect 3316 3236 3372 3238
rect 3396 3236 3452 3238
rect 3156 2202 3212 2204
rect 3236 2202 3292 2204
rect 3316 2202 3372 2204
rect 3396 2202 3452 2204
rect 3156 2150 3202 2202
rect 3202 2150 3212 2202
rect 3236 2150 3266 2202
rect 3266 2150 3278 2202
rect 3278 2150 3292 2202
rect 3316 2150 3330 2202
rect 3330 2150 3342 2202
rect 3342 2150 3372 2202
rect 3396 2150 3406 2202
rect 3406 2150 3452 2202
rect 3156 2148 3212 2150
rect 3236 2148 3292 2150
rect 3316 2148 3372 2150
rect 3396 2148 3452 2150
rect 1582 1400 1638 1456
rect 4894 6840 4950 6896
rect 5156 7098 5212 7100
rect 5236 7098 5292 7100
rect 5316 7098 5372 7100
rect 5396 7098 5452 7100
rect 5156 7046 5202 7098
rect 5202 7046 5212 7098
rect 5236 7046 5266 7098
rect 5266 7046 5278 7098
rect 5278 7046 5292 7098
rect 5316 7046 5330 7098
rect 5330 7046 5342 7098
rect 5342 7046 5372 7098
rect 5396 7046 5406 7098
rect 5406 7046 5452 7098
rect 5156 7044 5212 7046
rect 5236 7044 5292 7046
rect 5316 7044 5372 7046
rect 5396 7044 5452 7046
rect 5156 6010 5212 6012
rect 5236 6010 5292 6012
rect 5316 6010 5372 6012
rect 5396 6010 5452 6012
rect 5156 5958 5202 6010
rect 5202 5958 5212 6010
rect 5236 5958 5266 6010
rect 5266 5958 5278 6010
rect 5278 5958 5292 6010
rect 5316 5958 5330 6010
rect 5330 5958 5342 6010
rect 5342 5958 5372 6010
rect 5396 5958 5406 6010
rect 5406 5958 5452 6010
rect 5156 5956 5212 5958
rect 5236 5956 5292 5958
rect 5316 5956 5372 5958
rect 5396 5956 5452 5958
rect 5156 4922 5212 4924
rect 5236 4922 5292 4924
rect 5316 4922 5372 4924
rect 5396 4922 5452 4924
rect 5156 4870 5202 4922
rect 5202 4870 5212 4922
rect 5236 4870 5266 4922
rect 5266 4870 5278 4922
rect 5278 4870 5292 4922
rect 5316 4870 5330 4922
rect 5330 4870 5342 4922
rect 5342 4870 5372 4922
rect 5396 4870 5406 4922
rect 5406 4870 5452 4922
rect 5156 4868 5212 4870
rect 5236 4868 5292 4870
rect 5316 4868 5372 4870
rect 5396 4868 5452 4870
rect 5156 3834 5212 3836
rect 5236 3834 5292 3836
rect 5316 3834 5372 3836
rect 5396 3834 5452 3836
rect 5156 3782 5202 3834
rect 5202 3782 5212 3834
rect 5236 3782 5266 3834
rect 5266 3782 5278 3834
rect 5278 3782 5292 3834
rect 5316 3782 5330 3834
rect 5330 3782 5342 3834
rect 5342 3782 5372 3834
rect 5396 3782 5406 3834
rect 5406 3782 5452 3834
rect 5156 3780 5212 3782
rect 5236 3780 5292 3782
rect 5316 3780 5372 3782
rect 5396 3780 5452 3782
rect 7156 7642 7212 7644
rect 7236 7642 7292 7644
rect 7316 7642 7372 7644
rect 7396 7642 7452 7644
rect 7156 7590 7202 7642
rect 7202 7590 7212 7642
rect 7236 7590 7266 7642
rect 7266 7590 7278 7642
rect 7278 7590 7292 7642
rect 7316 7590 7330 7642
rect 7330 7590 7342 7642
rect 7342 7590 7372 7642
rect 7396 7590 7406 7642
rect 7406 7590 7452 7642
rect 7156 7588 7212 7590
rect 7236 7588 7292 7590
rect 7316 7588 7372 7590
rect 7396 7588 7452 7590
rect 7562 7520 7618 7576
rect 7156 6554 7212 6556
rect 7236 6554 7292 6556
rect 7316 6554 7372 6556
rect 7396 6554 7452 6556
rect 7156 6502 7202 6554
rect 7202 6502 7212 6554
rect 7236 6502 7266 6554
rect 7266 6502 7278 6554
rect 7278 6502 7292 6554
rect 7316 6502 7330 6554
rect 7330 6502 7342 6554
rect 7342 6502 7372 6554
rect 7396 6502 7406 6554
rect 7406 6502 7452 6554
rect 7156 6500 7212 6502
rect 7236 6500 7292 6502
rect 7316 6500 7372 6502
rect 7396 6500 7452 6502
rect 7562 5480 7618 5536
rect 7156 5466 7212 5468
rect 7236 5466 7292 5468
rect 7316 5466 7372 5468
rect 7396 5466 7452 5468
rect 7156 5414 7202 5466
rect 7202 5414 7212 5466
rect 7236 5414 7266 5466
rect 7266 5414 7278 5466
rect 7278 5414 7292 5466
rect 7316 5414 7330 5466
rect 7330 5414 7342 5466
rect 7342 5414 7372 5466
rect 7396 5414 7406 5466
rect 7406 5414 7452 5466
rect 7156 5412 7212 5414
rect 7236 5412 7292 5414
rect 7316 5412 7372 5414
rect 7396 5412 7452 5414
rect 6826 4800 6882 4856
rect 7156 4378 7212 4380
rect 7236 4378 7292 4380
rect 7316 4378 7372 4380
rect 7396 4378 7452 4380
rect 7156 4326 7202 4378
rect 7202 4326 7212 4378
rect 7236 4326 7266 4378
rect 7266 4326 7278 4378
rect 7278 4326 7292 4378
rect 7316 4326 7330 4378
rect 7330 4326 7342 4378
rect 7342 4326 7372 4378
rect 7396 4326 7406 4378
rect 7406 4326 7452 4378
rect 7156 4324 7212 4326
rect 7236 4324 7292 4326
rect 7316 4324 7372 4326
rect 7396 4324 7452 4326
rect 6734 4140 6790 4176
rect 6734 4120 6736 4140
rect 6736 4120 6788 4140
rect 6788 4120 6790 4140
rect 7156 3290 7212 3292
rect 7236 3290 7292 3292
rect 7316 3290 7372 3292
rect 7396 3290 7452 3292
rect 7156 3238 7202 3290
rect 7202 3238 7212 3290
rect 7236 3238 7266 3290
rect 7266 3238 7278 3290
rect 7278 3238 7292 3290
rect 7316 3238 7330 3290
rect 7330 3238 7342 3290
rect 7342 3238 7372 3290
rect 7396 3238 7406 3290
rect 7406 3238 7452 3290
rect 7156 3236 7212 3238
rect 7236 3236 7292 3238
rect 7316 3236 7372 3238
rect 7396 3236 7452 3238
rect 5156 2746 5212 2748
rect 5236 2746 5292 2748
rect 5316 2746 5372 2748
rect 5396 2746 5452 2748
rect 5156 2694 5202 2746
rect 5202 2694 5212 2746
rect 5236 2694 5266 2746
rect 5266 2694 5278 2746
rect 5278 2694 5292 2746
rect 5316 2694 5330 2746
rect 5330 2694 5342 2746
rect 5342 2694 5372 2746
rect 5396 2694 5406 2746
rect 5406 2694 5452 2746
rect 5156 2692 5212 2694
rect 5236 2692 5292 2694
rect 5316 2692 5372 2694
rect 5396 2692 5452 2694
rect 5446 2388 5448 2408
rect 5448 2388 5500 2408
rect 5500 2388 5502 2408
rect 5446 2352 5502 2388
rect 5156 1658 5212 1660
rect 5236 1658 5292 1660
rect 5316 1658 5372 1660
rect 5396 1658 5452 1660
rect 5156 1606 5202 1658
rect 5202 1606 5212 1658
rect 5236 1606 5266 1658
rect 5266 1606 5278 1658
rect 5278 1606 5292 1658
rect 5316 1606 5330 1658
rect 5330 1606 5342 1658
rect 5342 1606 5372 1658
rect 5396 1606 5406 1658
rect 5406 1606 5452 1658
rect 5156 1604 5212 1606
rect 5236 1604 5292 1606
rect 5316 1604 5372 1606
rect 5396 1604 5452 1606
rect 6550 2796 6552 2816
rect 6552 2796 6604 2816
rect 6604 2796 6606 2816
rect 6550 2760 6606 2796
rect 7156 2202 7212 2204
rect 7236 2202 7292 2204
rect 7316 2202 7372 2204
rect 7396 2202 7452 2204
rect 7156 2150 7202 2202
rect 7202 2150 7212 2202
rect 7236 2150 7266 2202
rect 7266 2150 7278 2202
rect 7278 2150 7292 2202
rect 7316 2150 7330 2202
rect 7330 2150 7342 2202
rect 7342 2150 7372 2202
rect 7396 2150 7406 2202
rect 7406 2150 7452 2202
rect 7156 2148 7212 2150
rect 7236 2148 7292 2150
rect 7316 2148 7372 2150
rect 7396 2148 7452 2150
rect 3156 1114 3212 1116
rect 3236 1114 3292 1116
rect 3316 1114 3372 1116
rect 3396 1114 3452 1116
rect 3156 1062 3202 1114
rect 3202 1062 3212 1114
rect 3236 1062 3266 1114
rect 3266 1062 3278 1114
rect 3278 1062 3292 1114
rect 3316 1062 3330 1114
rect 3330 1062 3342 1114
rect 3342 1062 3372 1114
rect 3396 1062 3406 1114
rect 3406 1062 3452 1114
rect 3156 1060 3212 1062
rect 3236 1060 3292 1062
rect 3316 1060 3372 1062
rect 3396 1060 3452 1062
rect 5538 1400 5594 1456
rect 7156 1114 7212 1116
rect 7236 1114 7292 1116
rect 7316 1114 7372 1116
rect 7396 1114 7452 1116
rect 7156 1062 7202 1114
rect 7202 1062 7212 1114
rect 7236 1062 7266 1114
rect 7266 1062 7278 1114
rect 7278 1062 7292 1114
rect 7316 1062 7330 1114
rect 7330 1062 7342 1114
rect 7342 1062 7372 1114
rect 7396 1062 7406 1114
rect 7406 1062 7452 1114
rect 7156 1060 7212 1062
rect 7236 1060 7292 1062
rect 7316 1060 7372 1062
rect 7396 1060 7452 1062
rect 1490 720 1546 776
rect 7838 40 7894 96
<< metal3 >>
rect 0 8938 800 8968
rect 2773 8938 2839 8941
rect 0 8936 2839 8938
rect 0 8880 2778 8936
rect 2834 8880 2839 8936
rect 0 8878 2839 8880
rect 0 8848 800 8878
rect 2773 8875 2839 8878
rect 6821 8258 6887 8261
rect 8200 8258 9000 8288
rect 6821 8256 9000 8258
rect 6821 8200 6826 8256
rect 6882 8200 9000 8256
rect 6821 8198 9000 8200
rect 6821 8195 6887 8198
rect 8200 8168 9000 8198
rect 3146 7648 3462 7649
rect 0 7578 800 7608
rect 3146 7584 3152 7648
rect 3216 7584 3232 7648
rect 3296 7584 3312 7648
rect 3376 7584 3392 7648
rect 3456 7584 3462 7648
rect 3146 7583 3462 7584
rect 7146 7648 7462 7649
rect 7146 7584 7152 7648
rect 7216 7584 7232 7648
rect 7296 7584 7312 7648
rect 7376 7584 7392 7648
rect 7456 7584 7462 7648
rect 7146 7583 7462 7584
rect 1577 7578 1643 7581
rect 0 7576 1643 7578
rect 0 7520 1582 7576
rect 1638 7520 1643 7576
rect 0 7518 1643 7520
rect 0 7488 800 7518
rect 1577 7515 1643 7518
rect 7557 7578 7623 7581
rect 8200 7578 9000 7608
rect 7557 7576 9000 7578
rect 7557 7520 7562 7576
rect 7618 7520 9000 7576
rect 7557 7518 9000 7520
rect 7557 7515 7623 7518
rect 8200 7488 9000 7518
rect 1146 7104 1462 7105
rect 1146 7040 1152 7104
rect 1216 7040 1232 7104
rect 1296 7040 1312 7104
rect 1376 7040 1392 7104
rect 1456 7040 1462 7104
rect 1146 7039 1462 7040
rect 5146 7104 5462 7105
rect 5146 7040 5152 7104
rect 5216 7040 5232 7104
rect 5296 7040 5312 7104
rect 5376 7040 5392 7104
rect 5456 7040 5462 7104
rect 5146 7039 5462 7040
rect 0 6898 800 6928
rect 4061 6898 4127 6901
rect 0 6896 4127 6898
rect 0 6840 4066 6896
rect 4122 6840 4127 6896
rect 0 6838 4127 6840
rect 0 6808 800 6838
rect 4061 6835 4127 6838
rect 4889 6898 4955 6901
rect 8200 6898 9000 6928
rect 4889 6896 9000 6898
rect 4889 6840 4894 6896
rect 4950 6840 9000 6896
rect 4889 6838 9000 6840
rect 4889 6835 4955 6838
rect 8200 6808 9000 6838
rect 3146 6560 3462 6561
rect 3146 6496 3152 6560
rect 3216 6496 3232 6560
rect 3296 6496 3312 6560
rect 3376 6496 3392 6560
rect 3456 6496 3462 6560
rect 3146 6495 3462 6496
rect 7146 6560 7462 6561
rect 7146 6496 7152 6560
rect 7216 6496 7232 6560
rect 7296 6496 7312 6560
rect 7376 6496 7392 6560
rect 7456 6496 7462 6560
rect 7146 6495 7462 6496
rect 0 6218 800 6248
rect 1761 6218 1827 6221
rect 0 6216 1827 6218
rect 0 6160 1766 6216
rect 1822 6160 1827 6216
rect 0 6158 1827 6160
rect 0 6128 800 6158
rect 1761 6155 1827 6158
rect 1146 6016 1462 6017
rect 1146 5952 1152 6016
rect 1216 5952 1232 6016
rect 1296 5952 1312 6016
rect 1376 5952 1392 6016
rect 1456 5952 1462 6016
rect 1146 5951 1462 5952
rect 5146 6016 5462 6017
rect 5146 5952 5152 6016
rect 5216 5952 5232 6016
rect 5296 5952 5312 6016
rect 5376 5952 5392 6016
rect 5456 5952 5462 6016
rect 5146 5951 5462 5952
rect 7557 5538 7623 5541
rect 8200 5538 9000 5568
rect 7557 5536 9000 5538
rect 7557 5480 7562 5536
rect 7618 5480 9000 5536
rect 7557 5478 9000 5480
rect 7557 5475 7623 5478
rect 3146 5472 3462 5473
rect 3146 5408 3152 5472
rect 3216 5408 3232 5472
rect 3296 5408 3312 5472
rect 3376 5408 3392 5472
rect 3456 5408 3462 5472
rect 3146 5407 3462 5408
rect 7146 5472 7462 5473
rect 7146 5408 7152 5472
rect 7216 5408 7232 5472
rect 7296 5408 7312 5472
rect 7376 5408 7392 5472
rect 7456 5408 7462 5472
rect 8200 5448 9000 5478
rect 7146 5407 7462 5408
rect 1577 5130 1643 5133
rect 982 5128 1643 5130
rect 982 5072 1582 5128
rect 1638 5072 1643 5128
rect 982 5070 1643 5072
rect 0 4858 800 4888
rect 982 4858 1042 5070
rect 1577 5067 1643 5070
rect 1146 4928 1462 4929
rect 1146 4864 1152 4928
rect 1216 4864 1232 4928
rect 1296 4864 1312 4928
rect 1376 4864 1392 4928
rect 1456 4864 1462 4928
rect 1146 4863 1462 4864
rect 5146 4928 5462 4929
rect 5146 4864 5152 4928
rect 5216 4864 5232 4928
rect 5296 4864 5312 4928
rect 5376 4864 5392 4928
rect 5456 4864 5462 4928
rect 5146 4863 5462 4864
rect 0 4798 1042 4858
rect 6821 4858 6887 4861
rect 8200 4858 9000 4888
rect 6821 4856 9000 4858
rect 6821 4800 6826 4856
rect 6882 4800 9000 4856
rect 6821 4798 9000 4800
rect 0 4768 800 4798
rect 6821 4795 6887 4798
rect 8200 4768 9000 4798
rect 3146 4384 3462 4385
rect 3146 4320 3152 4384
rect 3216 4320 3232 4384
rect 3296 4320 3312 4384
rect 3376 4320 3392 4384
rect 3456 4320 3462 4384
rect 3146 4319 3462 4320
rect 7146 4384 7462 4385
rect 7146 4320 7152 4384
rect 7216 4320 7232 4384
rect 7296 4320 7312 4384
rect 7376 4320 7392 4384
rect 7456 4320 7462 4384
rect 7146 4319 7462 4320
rect 0 4178 800 4208
rect 2773 4178 2839 4181
rect 0 4176 2839 4178
rect 0 4120 2778 4176
rect 2834 4120 2839 4176
rect 0 4118 2839 4120
rect 0 4088 800 4118
rect 2773 4115 2839 4118
rect 6729 4178 6795 4181
rect 8200 4178 9000 4208
rect 6729 4176 9000 4178
rect 6729 4120 6734 4176
rect 6790 4120 9000 4176
rect 6729 4118 9000 4120
rect 6729 4115 6795 4118
rect 8200 4088 9000 4118
rect 1146 3840 1462 3841
rect 1146 3776 1152 3840
rect 1216 3776 1232 3840
rect 1296 3776 1312 3840
rect 1376 3776 1392 3840
rect 1456 3776 1462 3840
rect 1146 3775 1462 3776
rect 5146 3840 5462 3841
rect 5146 3776 5152 3840
rect 5216 3776 5232 3840
rect 5296 3776 5312 3840
rect 5376 3776 5392 3840
rect 5456 3776 5462 3840
rect 5146 3775 5462 3776
rect 0 3498 800 3528
rect 2865 3498 2931 3501
rect 0 3496 2931 3498
rect 0 3440 2870 3496
rect 2926 3440 2931 3496
rect 0 3438 2931 3440
rect 0 3408 800 3438
rect 2865 3435 2931 3438
rect 3146 3296 3462 3297
rect 3146 3232 3152 3296
rect 3216 3232 3232 3296
rect 3296 3232 3312 3296
rect 3376 3232 3392 3296
rect 3456 3232 3462 3296
rect 3146 3231 3462 3232
rect 7146 3296 7462 3297
rect 7146 3232 7152 3296
rect 7216 3232 7232 3296
rect 7296 3232 7312 3296
rect 7376 3232 7392 3296
rect 7456 3232 7462 3296
rect 7146 3231 7462 3232
rect 6545 2818 6611 2821
rect 8200 2818 9000 2848
rect 6545 2816 9000 2818
rect 6545 2760 6550 2816
rect 6606 2760 9000 2816
rect 6545 2758 9000 2760
rect 6545 2755 6611 2758
rect 1146 2752 1462 2753
rect 1146 2688 1152 2752
rect 1216 2688 1232 2752
rect 1296 2688 1312 2752
rect 1376 2688 1392 2752
rect 1456 2688 1462 2752
rect 1146 2687 1462 2688
rect 5146 2752 5462 2753
rect 5146 2688 5152 2752
rect 5216 2688 5232 2752
rect 5296 2688 5312 2752
rect 5376 2688 5392 2752
rect 5456 2688 5462 2752
rect 8200 2728 9000 2758
rect 5146 2687 5462 2688
rect 5441 2410 5507 2413
rect 5441 2408 7666 2410
rect 5441 2352 5446 2408
rect 5502 2352 7666 2408
rect 5441 2350 7666 2352
rect 5441 2347 5507 2350
rect 3146 2208 3462 2209
rect 0 2138 800 2168
rect 3146 2144 3152 2208
rect 3216 2144 3232 2208
rect 3296 2144 3312 2208
rect 3376 2144 3392 2208
rect 3456 2144 3462 2208
rect 3146 2143 3462 2144
rect 7146 2208 7462 2209
rect 7146 2144 7152 2208
rect 7216 2144 7232 2208
rect 7296 2144 7312 2208
rect 7376 2144 7392 2208
rect 7456 2144 7462 2208
rect 7146 2143 7462 2144
rect 2773 2138 2839 2141
rect 0 2136 2839 2138
rect 0 2080 2778 2136
rect 2834 2080 2839 2136
rect 0 2078 2839 2080
rect 7606 2138 7666 2350
rect 8200 2138 9000 2168
rect 7606 2078 9000 2138
rect 0 2048 800 2078
rect 2773 2075 2839 2078
rect 8200 2048 9000 2078
rect 1146 1664 1462 1665
rect 1146 1600 1152 1664
rect 1216 1600 1232 1664
rect 1296 1600 1312 1664
rect 1376 1600 1392 1664
rect 1456 1600 1462 1664
rect 1146 1599 1462 1600
rect 5146 1664 5462 1665
rect 5146 1600 5152 1664
rect 5216 1600 5232 1664
rect 5296 1600 5312 1664
rect 5376 1600 5392 1664
rect 5456 1600 5462 1664
rect 5146 1599 5462 1600
rect 0 1458 800 1488
rect 1577 1458 1643 1461
rect 0 1456 1643 1458
rect 0 1400 1582 1456
rect 1638 1400 1643 1456
rect 0 1398 1643 1400
rect 0 1368 800 1398
rect 1577 1395 1643 1398
rect 5533 1458 5599 1461
rect 8200 1458 9000 1488
rect 5533 1456 9000 1458
rect 5533 1400 5538 1456
rect 5594 1400 9000 1456
rect 5533 1398 9000 1400
rect 5533 1395 5599 1398
rect 8200 1368 9000 1398
rect 3146 1120 3462 1121
rect 3146 1056 3152 1120
rect 3216 1056 3232 1120
rect 3296 1056 3312 1120
rect 3376 1056 3392 1120
rect 3456 1056 3462 1120
rect 3146 1055 3462 1056
rect 7146 1120 7462 1121
rect 7146 1056 7152 1120
rect 7216 1056 7232 1120
rect 7296 1056 7312 1120
rect 7376 1056 7392 1120
rect 7456 1056 7462 1120
rect 7146 1055 7462 1056
rect 0 778 800 808
rect 1485 778 1551 781
rect 0 776 1551 778
rect 0 720 1490 776
rect 1546 720 1551 776
rect 0 718 1551 720
rect 0 688 800 718
rect 1485 715 1551 718
rect 7833 98 7899 101
rect 8200 98 9000 128
rect 7833 96 9000 98
rect 7833 40 7838 96
rect 7894 40 9000 96
rect 7833 38 9000 40
rect 7833 35 7899 38
rect 8200 8 9000 38
<< via3 >>
rect 3152 7644 3216 7648
rect 3152 7588 3156 7644
rect 3156 7588 3212 7644
rect 3212 7588 3216 7644
rect 3152 7584 3216 7588
rect 3232 7644 3296 7648
rect 3232 7588 3236 7644
rect 3236 7588 3292 7644
rect 3292 7588 3296 7644
rect 3232 7584 3296 7588
rect 3312 7644 3376 7648
rect 3312 7588 3316 7644
rect 3316 7588 3372 7644
rect 3372 7588 3376 7644
rect 3312 7584 3376 7588
rect 3392 7644 3456 7648
rect 3392 7588 3396 7644
rect 3396 7588 3452 7644
rect 3452 7588 3456 7644
rect 3392 7584 3456 7588
rect 7152 7644 7216 7648
rect 7152 7588 7156 7644
rect 7156 7588 7212 7644
rect 7212 7588 7216 7644
rect 7152 7584 7216 7588
rect 7232 7644 7296 7648
rect 7232 7588 7236 7644
rect 7236 7588 7292 7644
rect 7292 7588 7296 7644
rect 7232 7584 7296 7588
rect 7312 7644 7376 7648
rect 7312 7588 7316 7644
rect 7316 7588 7372 7644
rect 7372 7588 7376 7644
rect 7312 7584 7376 7588
rect 7392 7644 7456 7648
rect 7392 7588 7396 7644
rect 7396 7588 7452 7644
rect 7452 7588 7456 7644
rect 7392 7584 7456 7588
rect 1152 7100 1216 7104
rect 1152 7044 1156 7100
rect 1156 7044 1212 7100
rect 1212 7044 1216 7100
rect 1152 7040 1216 7044
rect 1232 7100 1296 7104
rect 1232 7044 1236 7100
rect 1236 7044 1292 7100
rect 1292 7044 1296 7100
rect 1232 7040 1296 7044
rect 1312 7100 1376 7104
rect 1312 7044 1316 7100
rect 1316 7044 1372 7100
rect 1372 7044 1376 7100
rect 1312 7040 1376 7044
rect 1392 7100 1456 7104
rect 1392 7044 1396 7100
rect 1396 7044 1452 7100
rect 1452 7044 1456 7100
rect 1392 7040 1456 7044
rect 5152 7100 5216 7104
rect 5152 7044 5156 7100
rect 5156 7044 5212 7100
rect 5212 7044 5216 7100
rect 5152 7040 5216 7044
rect 5232 7100 5296 7104
rect 5232 7044 5236 7100
rect 5236 7044 5292 7100
rect 5292 7044 5296 7100
rect 5232 7040 5296 7044
rect 5312 7100 5376 7104
rect 5312 7044 5316 7100
rect 5316 7044 5372 7100
rect 5372 7044 5376 7100
rect 5312 7040 5376 7044
rect 5392 7100 5456 7104
rect 5392 7044 5396 7100
rect 5396 7044 5452 7100
rect 5452 7044 5456 7100
rect 5392 7040 5456 7044
rect 3152 6556 3216 6560
rect 3152 6500 3156 6556
rect 3156 6500 3212 6556
rect 3212 6500 3216 6556
rect 3152 6496 3216 6500
rect 3232 6556 3296 6560
rect 3232 6500 3236 6556
rect 3236 6500 3292 6556
rect 3292 6500 3296 6556
rect 3232 6496 3296 6500
rect 3312 6556 3376 6560
rect 3312 6500 3316 6556
rect 3316 6500 3372 6556
rect 3372 6500 3376 6556
rect 3312 6496 3376 6500
rect 3392 6556 3456 6560
rect 3392 6500 3396 6556
rect 3396 6500 3452 6556
rect 3452 6500 3456 6556
rect 3392 6496 3456 6500
rect 7152 6556 7216 6560
rect 7152 6500 7156 6556
rect 7156 6500 7212 6556
rect 7212 6500 7216 6556
rect 7152 6496 7216 6500
rect 7232 6556 7296 6560
rect 7232 6500 7236 6556
rect 7236 6500 7292 6556
rect 7292 6500 7296 6556
rect 7232 6496 7296 6500
rect 7312 6556 7376 6560
rect 7312 6500 7316 6556
rect 7316 6500 7372 6556
rect 7372 6500 7376 6556
rect 7312 6496 7376 6500
rect 7392 6556 7456 6560
rect 7392 6500 7396 6556
rect 7396 6500 7452 6556
rect 7452 6500 7456 6556
rect 7392 6496 7456 6500
rect 1152 6012 1216 6016
rect 1152 5956 1156 6012
rect 1156 5956 1212 6012
rect 1212 5956 1216 6012
rect 1152 5952 1216 5956
rect 1232 6012 1296 6016
rect 1232 5956 1236 6012
rect 1236 5956 1292 6012
rect 1292 5956 1296 6012
rect 1232 5952 1296 5956
rect 1312 6012 1376 6016
rect 1312 5956 1316 6012
rect 1316 5956 1372 6012
rect 1372 5956 1376 6012
rect 1312 5952 1376 5956
rect 1392 6012 1456 6016
rect 1392 5956 1396 6012
rect 1396 5956 1452 6012
rect 1452 5956 1456 6012
rect 1392 5952 1456 5956
rect 5152 6012 5216 6016
rect 5152 5956 5156 6012
rect 5156 5956 5212 6012
rect 5212 5956 5216 6012
rect 5152 5952 5216 5956
rect 5232 6012 5296 6016
rect 5232 5956 5236 6012
rect 5236 5956 5292 6012
rect 5292 5956 5296 6012
rect 5232 5952 5296 5956
rect 5312 6012 5376 6016
rect 5312 5956 5316 6012
rect 5316 5956 5372 6012
rect 5372 5956 5376 6012
rect 5312 5952 5376 5956
rect 5392 6012 5456 6016
rect 5392 5956 5396 6012
rect 5396 5956 5452 6012
rect 5452 5956 5456 6012
rect 5392 5952 5456 5956
rect 3152 5468 3216 5472
rect 3152 5412 3156 5468
rect 3156 5412 3212 5468
rect 3212 5412 3216 5468
rect 3152 5408 3216 5412
rect 3232 5468 3296 5472
rect 3232 5412 3236 5468
rect 3236 5412 3292 5468
rect 3292 5412 3296 5468
rect 3232 5408 3296 5412
rect 3312 5468 3376 5472
rect 3312 5412 3316 5468
rect 3316 5412 3372 5468
rect 3372 5412 3376 5468
rect 3312 5408 3376 5412
rect 3392 5468 3456 5472
rect 3392 5412 3396 5468
rect 3396 5412 3452 5468
rect 3452 5412 3456 5468
rect 3392 5408 3456 5412
rect 7152 5468 7216 5472
rect 7152 5412 7156 5468
rect 7156 5412 7212 5468
rect 7212 5412 7216 5468
rect 7152 5408 7216 5412
rect 7232 5468 7296 5472
rect 7232 5412 7236 5468
rect 7236 5412 7292 5468
rect 7292 5412 7296 5468
rect 7232 5408 7296 5412
rect 7312 5468 7376 5472
rect 7312 5412 7316 5468
rect 7316 5412 7372 5468
rect 7372 5412 7376 5468
rect 7312 5408 7376 5412
rect 7392 5468 7456 5472
rect 7392 5412 7396 5468
rect 7396 5412 7452 5468
rect 7452 5412 7456 5468
rect 7392 5408 7456 5412
rect 1152 4924 1216 4928
rect 1152 4868 1156 4924
rect 1156 4868 1212 4924
rect 1212 4868 1216 4924
rect 1152 4864 1216 4868
rect 1232 4924 1296 4928
rect 1232 4868 1236 4924
rect 1236 4868 1292 4924
rect 1292 4868 1296 4924
rect 1232 4864 1296 4868
rect 1312 4924 1376 4928
rect 1312 4868 1316 4924
rect 1316 4868 1372 4924
rect 1372 4868 1376 4924
rect 1312 4864 1376 4868
rect 1392 4924 1456 4928
rect 1392 4868 1396 4924
rect 1396 4868 1452 4924
rect 1452 4868 1456 4924
rect 1392 4864 1456 4868
rect 5152 4924 5216 4928
rect 5152 4868 5156 4924
rect 5156 4868 5212 4924
rect 5212 4868 5216 4924
rect 5152 4864 5216 4868
rect 5232 4924 5296 4928
rect 5232 4868 5236 4924
rect 5236 4868 5292 4924
rect 5292 4868 5296 4924
rect 5232 4864 5296 4868
rect 5312 4924 5376 4928
rect 5312 4868 5316 4924
rect 5316 4868 5372 4924
rect 5372 4868 5376 4924
rect 5312 4864 5376 4868
rect 5392 4924 5456 4928
rect 5392 4868 5396 4924
rect 5396 4868 5452 4924
rect 5452 4868 5456 4924
rect 5392 4864 5456 4868
rect 3152 4380 3216 4384
rect 3152 4324 3156 4380
rect 3156 4324 3212 4380
rect 3212 4324 3216 4380
rect 3152 4320 3216 4324
rect 3232 4380 3296 4384
rect 3232 4324 3236 4380
rect 3236 4324 3292 4380
rect 3292 4324 3296 4380
rect 3232 4320 3296 4324
rect 3312 4380 3376 4384
rect 3312 4324 3316 4380
rect 3316 4324 3372 4380
rect 3372 4324 3376 4380
rect 3312 4320 3376 4324
rect 3392 4380 3456 4384
rect 3392 4324 3396 4380
rect 3396 4324 3452 4380
rect 3452 4324 3456 4380
rect 3392 4320 3456 4324
rect 7152 4380 7216 4384
rect 7152 4324 7156 4380
rect 7156 4324 7212 4380
rect 7212 4324 7216 4380
rect 7152 4320 7216 4324
rect 7232 4380 7296 4384
rect 7232 4324 7236 4380
rect 7236 4324 7292 4380
rect 7292 4324 7296 4380
rect 7232 4320 7296 4324
rect 7312 4380 7376 4384
rect 7312 4324 7316 4380
rect 7316 4324 7372 4380
rect 7372 4324 7376 4380
rect 7312 4320 7376 4324
rect 7392 4380 7456 4384
rect 7392 4324 7396 4380
rect 7396 4324 7452 4380
rect 7452 4324 7456 4380
rect 7392 4320 7456 4324
rect 1152 3836 1216 3840
rect 1152 3780 1156 3836
rect 1156 3780 1212 3836
rect 1212 3780 1216 3836
rect 1152 3776 1216 3780
rect 1232 3836 1296 3840
rect 1232 3780 1236 3836
rect 1236 3780 1292 3836
rect 1292 3780 1296 3836
rect 1232 3776 1296 3780
rect 1312 3836 1376 3840
rect 1312 3780 1316 3836
rect 1316 3780 1372 3836
rect 1372 3780 1376 3836
rect 1312 3776 1376 3780
rect 1392 3836 1456 3840
rect 1392 3780 1396 3836
rect 1396 3780 1452 3836
rect 1452 3780 1456 3836
rect 1392 3776 1456 3780
rect 5152 3836 5216 3840
rect 5152 3780 5156 3836
rect 5156 3780 5212 3836
rect 5212 3780 5216 3836
rect 5152 3776 5216 3780
rect 5232 3836 5296 3840
rect 5232 3780 5236 3836
rect 5236 3780 5292 3836
rect 5292 3780 5296 3836
rect 5232 3776 5296 3780
rect 5312 3836 5376 3840
rect 5312 3780 5316 3836
rect 5316 3780 5372 3836
rect 5372 3780 5376 3836
rect 5312 3776 5376 3780
rect 5392 3836 5456 3840
rect 5392 3780 5396 3836
rect 5396 3780 5452 3836
rect 5452 3780 5456 3836
rect 5392 3776 5456 3780
rect 3152 3292 3216 3296
rect 3152 3236 3156 3292
rect 3156 3236 3212 3292
rect 3212 3236 3216 3292
rect 3152 3232 3216 3236
rect 3232 3292 3296 3296
rect 3232 3236 3236 3292
rect 3236 3236 3292 3292
rect 3292 3236 3296 3292
rect 3232 3232 3296 3236
rect 3312 3292 3376 3296
rect 3312 3236 3316 3292
rect 3316 3236 3372 3292
rect 3372 3236 3376 3292
rect 3312 3232 3376 3236
rect 3392 3292 3456 3296
rect 3392 3236 3396 3292
rect 3396 3236 3452 3292
rect 3452 3236 3456 3292
rect 3392 3232 3456 3236
rect 7152 3292 7216 3296
rect 7152 3236 7156 3292
rect 7156 3236 7212 3292
rect 7212 3236 7216 3292
rect 7152 3232 7216 3236
rect 7232 3292 7296 3296
rect 7232 3236 7236 3292
rect 7236 3236 7292 3292
rect 7292 3236 7296 3292
rect 7232 3232 7296 3236
rect 7312 3292 7376 3296
rect 7312 3236 7316 3292
rect 7316 3236 7372 3292
rect 7372 3236 7376 3292
rect 7312 3232 7376 3236
rect 7392 3292 7456 3296
rect 7392 3236 7396 3292
rect 7396 3236 7452 3292
rect 7452 3236 7456 3292
rect 7392 3232 7456 3236
rect 1152 2748 1216 2752
rect 1152 2692 1156 2748
rect 1156 2692 1212 2748
rect 1212 2692 1216 2748
rect 1152 2688 1216 2692
rect 1232 2748 1296 2752
rect 1232 2692 1236 2748
rect 1236 2692 1292 2748
rect 1292 2692 1296 2748
rect 1232 2688 1296 2692
rect 1312 2748 1376 2752
rect 1312 2692 1316 2748
rect 1316 2692 1372 2748
rect 1372 2692 1376 2748
rect 1312 2688 1376 2692
rect 1392 2748 1456 2752
rect 1392 2692 1396 2748
rect 1396 2692 1452 2748
rect 1452 2692 1456 2748
rect 1392 2688 1456 2692
rect 5152 2748 5216 2752
rect 5152 2692 5156 2748
rect 5156 2692 5212 2748
rect 5212 2692 5216 2748
rect 5152 2688 5216 2692
rect 5232 2748 5296 2752
rect 5232 2692 5236 2748
rect 5236 2692 5292 2748
rect 5292 2692 5296 2748
rect 5232 2688 5296 2692
rect 5312 2748 5376 2752
rect 5312 2692 5316 2748
rect 5316 2692 5372 2748
rect 5372 2692 5376 2748
rect 5312 2688 5376 2692
rect 5392 2748 5456 2752
rect 5392 2692 5396 2748
rect 5396 2692 5452 2748
rect 5452 2692 5456 2748
rect 5392 2688 5456 2692
rect 3152 2204 3216 2208
rect 3152 2148 3156 2204
rect 3156 2148 3212 2204
rect 3212 2148 3216 2204
rect 3152 2144 3216 2148
rect 3232 2204 3296 2208
rect 3232 2148 3236 2204
rect 3236 2148 3292 2204
rect 3292 2148 3296 2204
rect 3232 2144 3296 2148
rect 3312 2204 3376 2208
rect 3312 2148 3316 2204
rect 3316 2148 3372 2204
rect 3372 2148 3376 2204
rect 3312 2144 3376 2148
rect 3392 2204 3456 2208
rect 3392 2148 3396 2204
rect 3396 2148 3452 2204
rect 3452 2148 3456 2204
rect 3392 2144 3456 2148
rect 7152 2204 7216 2208
rect 7152 2148 7156 2204
rect 7156 2148 7212 2204
rect 7212 2148 7216 2204
rect 7152 2144 7216 2148
rect 7232 2204 7296 2208
rect 7232 2148 7236 2204
rect 7236 2148 7292 2204
rect 7292 2148 7296 2204
rect 7232 2144 7296 2148
rect 7312 2204 7376 2208
rect 7312 2148 7316 2204
rect 7316 2148 7372 2204
rect 7372 2148 7376 2204
rect 7312 2144 7376 2148
rect 7392 2204 7456 2208
rect 7392 2148 7396 2204
rect 7396 2148 7452 2204
rect 7452 2148 7456 2204
rect 7392 2144 7456 2148
rect 1152 1660 1216 1664
rect 1152 1604 1156 1660
rect 1156 1604 1212 1660
rect 1212 1604 1216 1660
rect 1152 1600 1216 1604
rect 1232 1660 1296 1664
rect 1232 1604 1236 1660
rect 1236 1604 1292 1660
rect 1292 1604 1296 1660
rect 1232 1600 1296 1604
rect 1312 1660 1376 1664
rect 1312 1604 1316 1660
rect 1316 1604 1372 1660
rect 1372 1604 1376 1660
rect 1312 1600 1376 1604
rect 1392 1660 1456 1664
rect 1392 1604 1396 1660
rect 1396 1604 1452 1660
rect 1452 1604 1456 1660
rect 1392 1600 1456 1604
rect 5152 1660 5216 1664
rect 5152 1604 5156 1660
rect 5156 1604 5212 1660
rect 5212 1604 5216 1660
rect 5152 1600 5216 1604
rect 5232 1660 5296 1664
rect 5232 1604 5236 1660
rect 5236 1604 5292 1660
rect 5292 1604 5296 1660
rect 5232 1600 5296 1604
rect 5312 1660 5376 1664
rect 5312 1604 5316 1660
rect 5316 1604 5372 1660
rect 5372 1604 5376 1660
rect 5312 1600 5376 1604
rect 5392 1660 5456 1664
rect 5392 1604 5396 1660
rect 5396 1604 5452 1660
rect 5452 1604 5456 1660
rect 5392 1600 5456 1604
rect 3152 1116 3216 1120
rect 3152 1060 3156 1116
rect 3156 1060 3212 1116
rect 3212 1060 3216 1116
rect 3152 1056 3216 1060
rect 3232 1116 3296 1120
rect 3232 1060 3236 1116
rect 3236 1060 3292 1116
rect 3292 1060 3296 1116
rect 3232 1056 3296 1060
rect 3312 1116 3376 1120
rect 3312 1060 3316 1116
rect 3316 1060 3372 1116
rect 3372 1060 3376 1116
rect 3312 1056 3376 1060
rect 3392 1116 3456 1120
rect 3392 1060 3396 1116
rect 3396 1060 3452 1116
rect 3452 1060 3456 1116
rect 3392 1056 3456 1060
rect 7152 1116 7216 1120
rect 7152 1060 7156 1116
rect 7156 1060 7212 1116
rect 7212 1060 7216 1116
rect 7152 1056 7216 1060
rect 7232 1116 7296 1120
rect 7232 1060 7236 1116
rect 7236 1060 7292 1116
rect 7292 1060 7296 1116
rect 7232 1056 7296 1060
rect 7312 1116 7376 1120
rect 7312 1060 7316 1116
rect 7316 1060 7372 1116
rect 7372 1060 7376 1116
rect 7312 1056 7376 1060
rect 7392 1116 7456 1120
rect 7392 1060 7396 1116
rect 7396 1060 7452 1116
rect 7452 1060 7456 1116
rect 7392 1056 7456 1060
<< metal4 >>
rect 1144 7104 1464 7664
rect 1144 7040 1152 7104
rect 1216 7040 1232 7104
rect 1296 7040 1312 7104
rect 1376 7040 1392 7104
rect 1456 7040 1464 7104
rect 1144 6016 1464 7040
rect 1144 5952 1152 6016
rect 1216 5952 1232 6016
rect 1296 5952 1312 6016
rect 1376 5952 1392 6016
rect 1456 5952 1464 6016
rect 1144 4928 1464 5952
rect 1144 4864 1152 4928
rect 1216 4864 1232 4928
rect 1296 4864 1312 4928
rect 1376 4864 1392 4928
rect 1456 4864 1464 4928
rect 1144 3840 1464 4864
rect 1144 3776 1152 3840
rect 1216 3776 1232 3840
rect 1296 3776 1312 3840
rect 1376 3776 1392 3840
rect 1456 3776 1464 3840
rect 1144 2752 1464 3776
rect 1144 2688 1152 2752
rect 1216 2688 1232 2752
rect 1296 2688 1312 2752
rect 1376 2688 1392 2752
rect 1456 2688 1464 2752
rect 1144 1664 1464 2688
rect 1144 1600 1152 1664
rect 1216 1600 1232 1664
rect 1296 1600 1312 1664
rect 1376 1600 1392 1664
rect 1456 1600 1464 1664
rect 1144 1040 1464 1600
rect 3144 7648 3464 7664
rect 3144 7584 3152 7648
rect 3216 7584 3232 7648
rect 3296 7584 3312 7648
rect 3376 7584 3392 7648
rect 3456 7584 3464 7648
rect 3144 6560 3464 7584
rect 3144 6496 3152 6560
rect 3216 6496 3232 6560
rect 3296 6496 3312 6560
rect 3376 6496 3392 6560
rect 3456 6496 3464 6560
rect 3144 5472 3464 6496
rect 3144 5408 3152 5472
rect 3216 5408 3232 5472
rect 3296 5408 3312 5472
rect 3376 5408 3392 5472
rect 3456 5408 3464 5472
rect 3144 4384 3464 5408
rect 3144 4320 3152 4384
rect 3216 4320 3232 4384
rect 3296 4320 3312 4384
rect 3376 4320 3392 4384
rect 3456 4320 3464 4384
rect 3144 3296 3464 4320
rect 3144 3232 3152 3296
rect 3216 3232 3232 3296
rect 3296 3232 3312 3296
rect 3376 3232 3392 3296
rect 3456 3232 3464 3296
rect 3144 2208 3464 3232
rect 3144 2144 3152 2208
rect 3216 2144 3232 2208
rect 3296 2144 3312 2208
rect 3376 2144 3392 2208
rect 3456 2144 3464 2208
rect 3144 1120 3464 2144
rect 3144 1056 3152 1120
rect 3216 1056 3232 1120
rect 3296 1056 3312 1120
rect 3376 1056 3392 1120
rect 3456 1056 3464 1120
rect 3144 1040 3464 1056
rect 5144 7104 5464 7664
rect 5144 7040 5152 7104
rect 5216 7040 5232 7104
rect 5296 7040 5312 7104
rect 5376 7040 5392 7104
rect 5456 7040 5464 7104
rect 5144 6016 5464 7040
rect 5144 5952 5152 6016
rect 5216 5952 5232 6016
rect 5296 5952 5312 6016
rect 5376 5952 5392 6016
rect 5456 5952 5464 6016
rect 5144 4928 5464 5952
rect 5144 4864 5152 4928
rect 5216 4864 5232 4928
rect 5296 4864 5312 4928
rect 5376 4864 5392 4928
rect 5456 4864 5464 4928
rect 5144 3840 5464 4864
rect 5144 3776 5152 3840
rect 5216 3776 5232 3840
rect 5296 3776 5312 3840
rect 5376 3776 5392 3840
rect 5456 3776 5464 3840
rect 5144 2752 5464 3776
rect 5144 2688 5152 2752
rect 5216 2688 5232 2752
rect 5296 2688 5312 2752
rect 5376 2688 5392 2752
rect 5456 2688 5464 2752
rect 5144 1664 5464 2688
rect 5144 1600 5152 1664
rect 5216 1600 5232 1664
rect 5296 1600 5312 1664
rect 5376 1600 5392 1664
rect 5456 1600 5464 1664
rect 5144 1040 5464 1600
rect 7144 7648 7464 7664
rect 7144 7584 7152 7648
rect 7216 7584 7232 7648
rect 7296 7584 7312 7648
rect 7376 7584 7392 7648
rect 7456 7584 7464 7648
rect 7144 6560 7464 7584
rect 7144 6496 7152 6560
rect 7216 6496 7232 6560
rect 7296 6496 7312 6560
rect 7376 6496 7392 6560
rect 7456 6496 7464 6560
rect 7144 5472 7464 6496
rect 7144 5408 7152 5472
rect 7216 5408 7232 5472
rect 7296 5408 7312 5472
rect 7376 5408 7392 5472
rect 7456 5408 7464 5472
rect 7144 4384 7464 5408
rect 7144 4320 7152 4384
rect 7216 4320 7232 4384
rect 7296 4320 7312 4384
rect 7376 4320 7392 4384
rect 7456 4320 7464 4384
rect 7144 3296 7464 4320
rect 7144 3232 7152 3296
rect 7216 3232 7232 3296
rect 7296 3232 7312 3296
rect 7376 3232 7392 3296
rect 7456 3232 7464 3296
rect 7144 2208 7464 3232
rect 7144 2144 7152 2208
rect 7216 2144 7232 2208
rect 7296 2144 7312 2208
rect 7376 2144 7392 2208
rect 7456 2144 7464 2208
rect 7144 1120 7464 2144
rect 7144 1056 7152 1120
rect 7216 1056 7232 1120
rect 7296 1056 7312 1120
rect 7376 1056 7392 1120
rect 7456 1056 7464 1120
rect 7144 1040 7464 1056
use sky130_fd_sc_hd__fill_2  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 1380 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 1840 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 2668 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24
timestamp 1673029049
transform 1 0 3312 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1673029049
transform 1 0 3772 0 1 1088
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 4232 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 5336 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1673029049
transform 1 0 6072 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57
timestamp 1673029049
transform 1 0 6348 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68
timestamp 1673029049
transform 1 0 7360 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3
timestamp 1673029049
transform 1 0 1380 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 1932 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_36
timestamp 1673029049
transform 1 0 4416 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_40
timestamp 1673029049
transform 1 0 4784 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_44
timestamp 1673029049
transform 1 0 5152 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1673029049
transform 1 0 5796 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1673029049
transform 1 0 6164 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_57
timestamp 1673029049
transform 1 0 6348 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_68
timestamp 1673029049
transform 1 0 7360 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1673029049
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_8
timestamp 1673029049
transform 1 0 1840 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_15
timestamp 1673029049
transform 1 0 2484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_22
timestamp 1673029049
transform 1 0 3128 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1673029049
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_41
timestamp 1673029049
transform 1 0 4876 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_50
timestamp 1673029049
transform 1 0 5704 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_62
timestamp 1673029049
transform 1 0 6808 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3
timestamp 1673029049
transform 1 0 1380 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_9
timestamp 1673029049
transform 1 0 1932 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_13
timestamp 1673029049
transform 1 0 2300 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_43
timestamp 1673029049
transform 1 0 5060 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_52
timestamp 1673029049
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp 1673029049
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_62
timestamp 1673029049
transform 1 0 6808 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1673029049
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1673029049
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1673029049
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1673029049
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1673029049
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1673029049
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_65
timestamp 1673029049
transform 1 0 7084 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_69
timestamp 1673029049
transform 1 0 7452 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_3
timestamp 1673029049
transform 1 0 1380 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_11
timestamp 1673029049
transform 1 0 2116 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_16
timestamp 1673029049
transform 1 0 2576 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_28
timestamp 1673029049
transform 1 0 3680 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_40 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 4784 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_48
timestamp 1673029049
transform 1 0 5520 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_57
timestamp 1673029049
transform 1 0 6348 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_64
timestamp 1673029049
transform 1 0 6992 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3
timestamp 1673029049
transform 1 0 1380 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_9
timestamp 1673029049
transform 1 0 1932 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_19
timestamp 1673029049
transform 1 0 2852 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1673029049
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1673029049
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1673029049
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1673029049
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_65
timestamp 1673029049
transform 1 0 7084 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_69
timestamp 1673029049
transform 1 0 7452 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1673029049
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_8
timestamp 1673029049
transform 1 0 1840 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_20
timestamp 1673029049
transform 1 0 2944 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_32
timestamp 1673029049
transform 1 0 4048 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_44
timestamp 1673029049
transform 1 0 5152 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_57
timestamp 1673029049
transform 1 0 6348 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_68
timestamp 1673029049
transform 1 0 7360 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1673029049
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_8
timestamp 1673029049
transform 1 0 1840 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_16
timestamp 1673029049
transform 1 0 2576 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_20
timestamp 1673029049
transform 1 0 2944 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1673029049
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_34
timestamp 1673029049
transform 1 0 4232 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_46
timestamp 1673029049
transform 1 0 5336 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_50
timestamp 1673029049
transform 1 0 5704 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_60
timestamp 1673029049
transform 1 0 6624 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_68
timestamp 1673029049
transform 1 0 7360 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_3
timestamp 1673029049
transform 1 0 1380 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_12
timestamp 1673029049
transform 1 0 2208 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_19
timestamp 1673029049
transform 1 0 2852 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_23
timestamp 1673029049
transform 1 0 3220 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_27
timestamp 1673029049
transform 1 0 3588 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_35
timestamp 1673029049
transform 1 0 4324 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_42
timestamp 1673029049
transform 1 0 4968 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1673029049
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1673029049
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_62
timestamp 1673029049
transform 1 0 6808 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1673029049
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_14
timestamp 1673029049
transform 1 0 2392 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_22
timestamp 1673029049
transform 1 0 3128 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_26
timestamp 1673029049
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1673029049
transform 1 0 3772 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_34
timestamp 1673029049
transform 1 0 4232 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_46
timestamp 1673029049
transform 1 0 5336 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_53
timestamp 1673029049
transform 1 0 5980 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_57
timestamp 1673029049
transform 1 0 6348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_61
timestamp 1673029049
transform 1 0 6716 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_68
timestamp 1673029049
transform 1 0 7360 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_3
timestamp 1673029049
transform 1 0 1380 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_11_14
timestamp 1673029049
transform 1 0 2392 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_26
timestamp 1673029049
transform 1 0 3496 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_29
timestamp 1673029049
transform 1 0 3772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_41
timestamp 1673029049
transform 1 0 4876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_53
timestamp 1673029049
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_57
timestamp 1673029049
transform 1 0 6348 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_68
timestamp 1673029049
transform 1 0 7360 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1673029049
transform 1 0 1104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1673029049
transform -1 0 7820 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1673029049
transform 1 0 1104 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1673029049
transform -1 0 7820 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1673029049
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1673029049
transform -1 0 7820 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1673029049
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1673029049
transform -1 0 7820 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1673029049
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1673029049
transform -1 0 7820 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1673029049
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1673029049
transform -1 0 7820 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1673029049
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1673029049
transform -1 0 7820 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1673029049
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1673029049
transform -1 0 7820 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1673029049
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1673029049
transform -1 0 7820 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1673029049
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1673029049
transform -1 0 7820 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1673029049
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1673029049
transform -1 0 7820 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1673029049
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1673029049
transform -1 0 7820 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_24 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 3680 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_25
timestamp 1673029049
transform 1 0 6256 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_26
timestamp 1673029049
transform 1 0 6256 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_27
timestamp 1673029049
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28
timestamp 1673029049
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1673029049
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1673029049
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 1673029049
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 1673029049
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 1673029049
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 1673029049
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1673029049
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1673029049
transform 1 0 3680 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1673029049
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  spare_logic_biginv $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 1564 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[0\] $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 2300 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[1\]
timestamp 1673029049
transform 1 0 7084 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[2\]
timestamp 1673029049
transform 1 0 6440 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[3\]
timestamp 1673029049
transform -1 0 5980 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[4\]
timestamp 1673029049
transform -1 0 2392 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[5\]
timestamp 1673029049
transform -1 0 4232 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[6\]
timestamp 1673029049
transform 1 0 5520 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[7\]
timestamp 1673029049
transform -1 0 2576 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[8\]
timestamp 1673029049
transform -1 0 2944 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[9\]
timestamp 1673029049
transform -1 0 6992 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[10\]
timestamp 1673029049
transform -1 0 3588 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[11\]
timestamp 1673029049
transform -1 0 6808 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[12\]
timestamp 1673029049
transform -1 0 1840 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[13\]
timestamp 1673029049
transform -1 0 7360 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[14\]
timestamp 1673029049
transform -1 0 2852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[15\]
timestamp 1673029049
transform -1 0 3128 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[16\]
timestamp 1673029049
transform -1 0 1840 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[17\]
timestamp 1673029049
transform -1 0 7360 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[18\]
timestamp 1673029049
transform -1 0 1840 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[19\]
timestamp 1673029049
transform -1 0 1840 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[20\]
timestamp 1673029049
transform -1 0 4232 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[21\]
timestamp 1673029049
transform -1 0 5704 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[22\]
timestamp 1673029049
transform -1 0 2484 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[23\]
timestamp 1673029049
transform -1 0 3312 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[24\]
timestamp 1673029049
transform 1 0 2392 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[25\]
timestamp 1673029049
transform -1 0 6808 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spare_logic_const\[26\]
timestamp 1673029049
transform -1 0 4232 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__dfbbp_1  spare_logic_flop\[0\] $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 5060 0 -1 3264
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbp_1  spare_logic_flop\[1\]
timestamp 1673029049
transform 1 0 2024 0 -1 2176
box -38 -48 2430 592
use sky130_fd_sc_hd__inv_2  spare_logic_inv\[0\] $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 4876 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  spare_logic_inv\[1\]
timestamp 1673029049
transform -1 0 7360 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  spare_logic_inv\[2\]
timestamp 1673029049
transform 1 0 7084 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  spare_logic_inv\[3\]
timestamp 1673029049
transform -1 0 3496 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  spare_logic_mux\[0\] $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 6624 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  spare_logic_mux\[1\]
timestamp 1673029049
transform -1 0 2852 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  spare_logic_nand\[0\] $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 4508 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  spare_logic_nand\[1\]
timestamp 1673029049
transform 1 0 5428 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  spare_logic_nor\[0\] $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform -1 0 5520 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  spare_logic_nor\[1\]
timestamp 1673029049
transform -1 0 2208 0 -1 6528
box -38 -48 498 592
<< labels >>
flabel metal3 s 0 2048 800 2168 0 FreeSans 480 0 0 0 spare_xfq[0]
port 0 nsew signal tristate
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 spare_xfq[1]
port 1 nsew signal tristate
flabel metal2 s 4526 8200 4582 9000 0 FreeSans 224 90 0 0 spare_xfqn[0]
port 2 nsew signal tristate
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 spare_xfqn[1]
port 3 nsew signal tristate
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 spare_xi[0]
port 4 nsew signal tristate
flabel metal3 s 8200 8 9000 128 0 FreeSans 480 0 0 0 spare_xi[1]
port 5 nsew signal tristate
flabel metal3 s 8200 5448 9000 5568 0 FreeSans 480 0 0 0 spare_xi[2]
port 6 nsew signal tristate
flabel metal2 s 18 8200 74 9000 0 FreeSans 224 90 0 0 spare_xi[3]
port 7 nsew signal tristate
flabel metal3 s 0 7488 800 7608 0 FreeSans 480 0 0 0 spare_xib
port 8 nsew signal tristate
flabel metal2 s 7102 8200 7158 9000 0 FreeSans 224 90 0 0 spare_xmx[0]
port 9 nsew signal tristate
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 spare_xmx[1]
port 10 nsew signal tristate
flabel metal3 s 8200 6808 9000 6928 0 FreeSans 480 0 0 0 spare_xna[0]
port 11 nsew signal tristate
flabel metal3 s 8200 1368 9000 1488 0 FreeSans 480 0 0 0 spare_xna[1]
port 12 nsew signal tristate
flabel metal2 s 1306 0 1362 800 0 FreeSans 224 90 0 0 spare_xno[0]
port 13 nsew signal tristate
flabel metal3 s 0 6128 800 6248 0 FreeSans 480 0 0 0 spare_xno[1]
port 14 nsew signal tristate
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 spare_xz[0]
port 15 nsew signal tristate
flabel metal2 s 5170 8200 5226 9000 0 FreeSans 224 90 0 0 spare_xz[10]
port 16 nsew signal tristate
flabel metal2 s 7746 8200 7802 9000 0 FreeSans 224 90 0 0 spare_xz[11]
port 17 nsew signal tristate
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 spare_xz[12]
port 18 nsew signal tristate
flabel metal3 s 8200 7488 9000 7608 0 FreeSans 480 0 0 0 spare_xz[13]
port 19 nsew signal tristate
flabel metal2 s 1950 8200 2006 9000 0 FreeSans 224 90 0 0 spare_xz[14]
port 20 nsew signal tristate
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 spare_xz[15]
port 21 nsew signal tristate
flabel metal3 s 0 1368 800 1488 0 FreeSans 480 0 0 0 spare_xz[16]
port 22 nsew signal tristate
flabel metal3 s 8200 4768 9000 4888 0 FreeSans 480 0 0 0 spare_xz[17]
port 23 nsew signal tristate
flabel metal2 s 662 8200 718 9000 0 FreeSans 224 90 0 0 spare_xz[18]
port 24 nsew signal tristate
flabel metal3 s 0 688 800 808 0 FreeSans 480 0 0 0 spare_xz[19]
port 25 nsew signal tristate
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 spare_xz[1]
port 26 nsew signal tristate
flabel metal2 s 5814 8200 5870 9000 0 FreeSans 224 90 0 0 spare_xz[20]
port 27 nsew signal tristate
flabel metal3 s 8200 2048 9000 2168 0 FreeSans 480 0 0 0 spare_xz[21]
port 28 nsew signal tristate
flabel metal2 s 662 0 718 800 0 FreeSans 224 90 0 0 spare_xz[22]
port 29 nsew signal tristate
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 spare_xz[23]
port 30 nsew signal tristate
flabel metal2 s 3238 0 3294 800 0 FreeSans 224 90 0 0 spare_xz[24]
port 31 nsew signal tristate
flabel metal3 s 8200 2728 9000 2848 0 FreeSans 480 0 0 0 spare_xz[25]
port 32 nsew signal tristate
flabel metal2 s 3882 0 3938 800 0 FreeSans 224 90 0 0 spare_xz[26]
port 33 nsew signal tristate
flabel metal3 s 8200 8168 9000 8288 0 FreeSans 480 0 0 0 spare_xz[2]
port 34 nsew signal tristate
flabel metal2 s 8390 8200 8446 9000 0 FreeSans 224 90 0 0 spare_xz[3]
port 35 nsew signal tristate
flabel metal2 s 2594 8200 2650 9000 0 FreeSans 224 90 0 0 spare_xz[4]
port 36 nsew signal tristate
flabel metal2 s 3238 8200 3294 9000 0 FreeSans 224 90 0 0 spare_xz[5]
port 37 nsew signal tristate
flabel metal2 s 5814 0 5870 800 0 FreeSans 224 90 0 0 spare_xz[6]
port 38 nsew signal tristate
flabel metal3 s 0 3408 800 3528 0 FreeSans 480 0 0 0 spare_xz[7]
port 39 nsew signal tristate
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 spare_xz[8]
port 40 nsew signal tristate
flabel metal3 s 8200 4088 9000 4208 0 FreeSans 480 0 0 0 spare_xz[9]
port 41 nsew signal tristate
flabel metal4 s 1144 1040 1464 7664 0 FreeSans 1920 90 0 0 vccd
port 42 nsew power bidirectional
flabel metal4 s 5144 1040 5464 7664 0 FreeSans 1920 90 0 0 vccd
port 42 nsew power bidirectional
flabel metal4 s 3144 1040 3464 7664 0 FreeSans 1920 90 0 0 vssd
port 43 nsew ground bidirectional
flabel metal4 s 7144 1040 7464 7664 0 FreeSans 1920 90 0 0 vssd
port 43 nsew ground bidirectional
rlabel metal1 4462 7072 4462 7072 0 vccd
rlabel metal1 4462 7616 4462 7616 0 vssd
rlabel metal3 1740 2108 1740 2108 0 spare_xfq[0]
rlabel metal2 6486 1282 6486 1282 0 spare_xfq[1]
rlabel metal1 3680 3162 3680 3162 0 spare_xfqn[0]
rlabel metal3 2384 6868 2384 6868 0 spare_xfqn[1]
rlabel metal2 8418 1316 8418 1316 0 spare_xi[0]
rlabel metal1 7544 1190 7544 1190 0 spare_xi[1]
rlabel metal1 7406 6630 7406 6630 0 spare_xi[2]
rlabel metal1 1334 6902 1334 6902 0 spare_xi[3]
rlabel metal3 1142 7548 1142 7548 0 spare_xib
rlabel metal1 6762 5882 6762 5882 0 spare_xmx[0]
rlabel metal2 5198 1095 5198 1095 0 spare_xmx[1]
rlabel metal2 4922 6613 4922 6613 0 spare_xna[0]
rlabel metal3 6954 1428 6954 1428 0 spare_xna[1]
rlabel metal2 1334 823 1334 823 0 spare_xno[0]
rlabel metal3 1234 6188 1234 6188 0 spare_xno[1]
rlabel metal1 4462 1938 4462 1938 0 spare_xz[0]
rlabel metal1 2461 6290 2461 6290 0 spare_xz[10]
rlabel metal1 7176 6290 7176 6290 0 spare_xz[11]
rlabel metal2 1610 5389 1610 5389 0 spare_xz[12]
rlabel metal1 7360 7378 7360 7378 0 spare_xz[13]
rlabel metal1 2300 6222 2300 6222 0 spare_xz[14]
rlabel metal1 2990 2618 2990 2618 0 spare_xz[15]
rlabel metal2 1610 1921 1610 1921 0 spare_xz[16]
rlabel metal1 6992 4998 6992 4998 0 spare_xz[17]
rlabel metal1 1150 5202 1150 5202 0 spare_xz[18]
rlabel metal1 2806 1530 2806 1530 0 spare_xz[19]
rlabel metal1 7544 1326 7544 1326 0 spare_xz[1]
rlabel metal1 2714 1870 2714 1870 0 spare_xz[20]
rlabel via2 5474 2397 5474 2397 0 spare_xz[21]
rlabel metal1 1380 1870 1380 1870 0 spare_xz[22]
rlabel metal1 3082 1360 3082 1360 0 spare_xz[23]
rlabel via1 3082 1445 3082 1445 0 spare_xz[24]
rlabel via2 6578 2805 6578 2805 0 spare_xz[25]
rlabel metal1 3956 1394 3956 1394 0 spare_xz[26]
rlabel metal1 6992 6766 6992 6766 0 spare_xz[2]
rlabel metal1 7084 6834 7084 6834 0 spare_xz[3]
rlabel metal2 2346 8228 2346 8228 0 spare_xz[4]
rlabel metal1 3818 6834 3818 6834 0 spare_xz[5]
rlabel metal1 5796 1734 5796 1734 0 spare_xz[6]
rlabel metal2 4554 5202 4554 5202 0 spare_xz[7]
rlabel metal2 5566 4386 5566 4386 0 spare_xz[8]
rlabel via2 6762 4131 6762 4131 0 spare_xz[9]
<< properties >>
string FIXED_BBOX 0 0 9000 9000
<< end >>
