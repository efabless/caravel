magic
tech sky130A
magscale 1 2
timestamp 1637846189
<< locali >>
rect 5273 10115 5307 10217
rect 10367 9537 10459 9571
rect 1501 9435 1535 9537
rect 10425 9367 10459 9537
rect 2789 8347 2823 8517
rect 7849 6647 7883 6817
rect 9413 6715 9447 6885
rect 6561 6171 6595 6273
rect 5365 2839 5399 2941
rect 14105 1751 14139 1921
rect 9965 663 9999 969
rect 10425 663 10459 765
<< viali >>
rect 6929 10761 6963 10795
rect 7205 10761 7239 10795
rect 10977 10761 11011 10795
rect 2329 10693 2363 10727
rect 8094 10693 8128 10727
rect 1317 10625 1351 10659
rect 5457 10625 5491 10659
rect 6745 10625 6779 10659
rect 7021 10625 7055 10659
rect 7389 10625 7423 10659
rect 9321 10625 9355 10659
rect 10425 10625 10459 10659
rect 11161 10625 11195 10659
rect 12265 10625 12299 10659
rect 13277 10625 13311 10659
rect 17923 10625 17957 10659
rect 18153 10625 18187 10659
rect 18337 10625 18371 10659
rect 2697 10557 2731 10591
rect 3065 10557 3099 10591
rect 5549 10557 5583 10591
rect 7849 10557 7883 10591
rect 12357 10557 12391 10591
rect 12449 10557 12483 10591
rect 13645 10557 13679 10591
rect 16129 10557 16163 10591
rect 16497 10557 16531 10591
rect 11897 10489 11931 10523
rect 4491 10421 4525 10455
rect 5825 10421 5859 10455
rect 7481 10421 7515 10455
rect 9229 10421 9263 10455
rect 9965 10421 9999 10455
rect 10701 10421 10735 10455
rect 10885 10421 10919 10455
rect 15071 10421 15105 10455
rect 18153 10421 18187 10455
rect 3525 10217 3559 10251
rect 5273 10217 5307 10251
rect 6009 10217 6043 10251
rect 7941 10217 7975 10251
rect 10885 10217 10919 10251
rect 13093 10217 13127 10251
rect 13645 10217 13679 10251
rect 16635 10217 16669 10251
rect 18337 10217 18371 10251
rect 305 10081 339 10115
rect 2053 10081 2087 10115
rect 3065 10081 3099 10115
rect 5273 10081 5307 10115
rect 5457 10081 5491 10115
rect 8401 10081 8435 10115
rect 14841 10081 14875 10115
rect 15209 10081 15243 10115
rect 2329 10013 2363 10047
rect 2697 10013 2731 10047
rect 3249 10013 3283 10047
rect 3341 10013 3375 10047
rect 3617 10013 3651 10047
rect 3893 10013 3927 10047
rect 4261 10013 4295 10047
rect 4813 10013 4847 10047
rect 4997 10013 5031 10047
rect 5549 10013 5583 10047
rect 6009 10013 6043 10047
rect 6193 10013 6227 10047
rect 8953 10013 8987 10047
rect 9137 10013 9171 10047
rect 9597 10013 9631 10047
rect 12081 10013 12115 10047
rect 13277 10013 13311 10047
rect 17969 10013 18003 10047
rect 18521 10013 18555 10047
rect 581 9945 615 9979
rect 2789 9945 2823 9979
rect 2973 9945 3007 9979
rect 3065 9945 3099 9979
rect 3801 9945 3835 9979
rect 8401 9945 8435 9979
rect 8493 9945 8527 9979
rect 11897 9945 11931 9979
rect 2237 9877 2271 9911
rect 2697 9877 2731 9911
rect 4997 9877 5031 9911
rect 5917 9877 5951 9911
rect 9045 9877 9079 9911
rect 17785 9877 17819 9911
rect 1133 9673 1167 9707
rect 5917 9673 5951 9707
rect 12449 9673 12483 9707
rect 4813 9605 4847 9639
rect 6009 9605 6043 9639
rect 9965 9605 9999 9639
rect 17693 9605 17727 9639
rect 1409 9537 1443 9571
rect 1501 9537 1535 9571
rect 1593 9537 1627 9571
rect 1777 9537 1811 9571
rect 2973 9537 3007 9571
rect 3157 9537 3191 9571
rect 4721 9537 4755 9571
rect 6745 9537 6779 9571
rect 10241 9537 10275 9571
rect 10333 9537 10367 9571
rect 12817 9537 12851 9571
rect 1133 9469 1167 9503
rect 1685 9469 1719 9503
rect 4997 9469 5031 9503
rect 6193 9469 6227 9503
rect 6837 9469 6871 9503
rect 6929 9469 6963 9503
rect 1317 9401 1351 9435
rect 1501 9401 1535 9435
rect 4353 9401 4387 9435
rect 5549 9401 5583 9435
rect 10609 9469 10643 9503
rect 10885 9469 10919 9503
rect 12909 9469 12943 9503
rect 13001 9469 13035 9503
rect 13277 9469 13311 9503
rect 15025 9469 15059 9503
rect 15301 9469 15335 9503
rect 17969 9469 18003 9503
rect 12357 9401 12391 9435
rect 16221 9401 16255 9435
rect 3065 9333 3099 9367
rect 6377 9333 6411 9367
rect 8493 9333 8527 9367
rect 10425 9333 10459 9367
rect 2053 9129 2087 9163
rect 5549 9129 5583 9163
rect 9229 9129 9263 9163
rect 9597 9129 9631 9163
rect 10701 9129 10735 9163
rect 18337 9129 18371 9163
rect 2237 9061 2271 9095
rect 2329 9061 2363 9095
rect 305 8993 339 9027
rect 581 8993 615 9027
rect 2145 8993 2179 9027
rect 3157 8993 3191 9027
rect 4445 8993 4479 9027
rect 6101 8993 6135 9027
rect 10057 8993 10091 9027
rect 10241 8993 10275 9027
rect 10793 8993 10827 9027
rect 12817 8993 12851 9027
rect 15761 8993 15795 9027
rect 2421 8925 2455 8959
rect 2881 8925 2915 8959
rect 5917 8925 5951 8959
rect 6653 8925 6687 8959
rect 7849 8925 7883 8959
rect 8116 8925 8150 8959
rect 9413 8925 9447 8959
rect 10333 8925 10367 8959
rect 13369 8925 13403 8959
rect 13553 8925 13587 8959
rect 15393 8925 15427 8959
rect 15853 8925 15887 8959
rect 16221 8925 16255 8959
rect 18153 8925 18187 8959
rect 4169 8857 4203 8891
rect 12541 8857 12575 8891
rect 3801 8789 3835 8823
rect 4261 8789 4295 8823
rect 6009 8789 6043 8823
rect 6561 8789 6595 8823
rect 9873 8789 9907 8823
rect 13461 8789 13495 8823
rect 13967 8789 14001 8823
rect 17969 8789 18003 8823
rect 2329 8585 2363 8619
rect 2513 8585 2547 8619
rect 3249 8585 3283 8619
rect 3341 8585 3375 8619
rect 4629 8585 4663 8619
rect 2789 8517 2823 8551
rect 5457 8517 5491 8551
rect 5733 8517 5767 8551
rect 6193 8517 6227 8551
rect 10241 8517 10275 8551
rect 11989 8517 12023 8551
rect 12173 8517 12207 8551
rect 13553 8517 13587 8551
rect 14473 8517 14507 8551
rect 15807 8517 15841 8551
rect 2421 8449 2455 8483
rect 2513 8449 2547 8483
rect 2697 8449 2731 8483
rect 3709 8449 3743 8483
rect 3893 8449 3927 8483
rect 4353 8449 4387 8483
rect 4537 8449 4571 8483
rect 4813 8449 4847 8483
rect 5273 8449 5307 8483
rect 5547 8471 5581 8505
rect 5641 8449 5675 8483
rect 5917 8449 5951 8483
rect 6377 8449 6411 8483
rect 8677 8449 8711 8483
rect 10425 8449 10459 8483
rect 10692 8449 10726 8483
rect 13645 8449 13679 8483
rect 14381 8449 14415 8483
rect 14565 8449 14599 8483
rect 14841 8449 14875 8483
rect 17601 8449 17635 8483
rect 18521 8449 18555 8483
rect 3525 8381 3559 8415
rect 6745 8381 6779 8415
rect 13461 8381 13495 8415
rect 17233 8381 17267 8415
rect 2789 8313 2823 8347
rect 3801 8313 3835 8347
rect 5365 8313 5399 8347
rect 5825 8313 5859 8347
rect 6009 8313 6043 8347
rect 18337 8313 18371 8347
rect 2881 8245 2915 8279
rect 8171 8245 8205 8279
rect 11805 8245 11839 8279
rect 14013 8245 14047 8279
rect 14933 8245 14967 8279
rect 4537 8041 4571 8075
rect 4629 8041 4663 8075
rect 5549 8041 5583 8075
rect 7941 8041 7975 8075
rect 8309 8041 8343 8075
rect 10149 8041 10183 8075
rect 10333 8041 10367 8075
rect 11621 8041 11655 8075
rect 14381 8041 14415 8075
rect 15025 8041 15059 8075
rect 9781 7973 9815 8007
rect 10885 7973 10919 8007
rect 11437 7973 11471 8007
rect 12725 7973 12759 8007
rect 13277 7973 13311 8007
rect 305 7905 339 7939
rect 3341 7905 3375 7939
rect 4353 7905 4387 7939
rect 4905 7905 4939 7939
rect 5089 7905 5123 7939
rect 9689 7905 9723 7939
rect 10241 7905 10275 7939
rect 10701 7905 10735 7939
rect 10793 7905 10827 7939
rect 11253 7905 11287 7939
rect 12265 7905 12299 7939
rect 15945 7905 15979 7939
rect 2881 7837 2915 7871
rect 3249 7837 3283 7871
rect 3433 7837 3467 7871
rect 3617 7837 3651 7871
rect 4077 7837 4111 7871
rect 4445 7837 4479 7871
rect 4721 7837 4755 7871
rect 4813 7837 4847 7871
rect 4997 7837 5031 7871
rect 8033 7837 8067 7871
rect 9965 7837 9999 7871
rect 10517 7837 10551 7871
rect 10885 7837 10919 7871
rect 10977 7837 11011 7871
rect 11161 7837 11195 7871
rect 11528 7815 11562 7849
rect 11621 7837 11655 7871
rect 12357 7837 12391 7871
rect 13001 7837 13035 7871
rect 13185 7837 13219 7871
rect 13829 7837 13863 7871
rect 14013 7837 14047 7871
rect 14611 7837 14645 7871
rect 14841 7837 14875 7871
rect 14933 7837 14967 7871
rect 15209 7837 15243 7871
rect 15485 7837 15519 7871
rect 581 7769 615 7803
rect 5825 7769 5859 7803
rect 6193 7769 6227 7803
rect 6377 7769 6411 7803
rect 9444 7769 9478 7803
rect 11253 7769 11287 7803
rect 11713 7769 11747 7803
rect 11897 7769 11931 7803
rect 15117 7769 15151 7803
rect 15393 7769 15427 7803
rect 16221 7769 16255 7803
rect 17969 7769 18003 7803
rect 2053 7701 2087 7735
rect 2789 7701 2823 7735
rect 3709 7701 3743 7735
rect 3893 7701 3927 7735
rect 5917 7701 5951 7735
rect 14749 7701 14783 7735
rect 1685 7497 1719 7531
rect 2973 7497 3007 7531
rect 9965 7497 9999 7531
rect 15577 7497 15611 7531
rect 17785 7497 17819 7531
rect 1869 7429 1903 7463
rect 6469 7429 6503 7463
rect 17049 7429 17083 7463
rect 1409 7361 1443 7395
rect 1961 7361 1995 7395
rect 2329 7361 2363 7395
rect 2513 7361 2547 7395
rect 2789 7361 2823 7395
rect 3157 7361 3191 7395
rect 3249 7361 3283 7395
rect 3341 7361 3375 7395
rect 3709 7361 3743 7395
rect 4813 7361 4847 7395
rect 4997 7361 5031 7395
rect 5273 7361 5307 7395
rect 5733 7361 5767 7395
rect 5917 7361 5951 7395
rect 6377 7361 6411 7395
rect 6745 7361 6779 7395
rect 7849 7361 7883 7395
rect 8953 7361 8987 7395
rect 9045 7361 9079 7395
rect 9597 7361 9631 7395
rect 9689 7361 9723 7395
rect 9781 7361 9815 7395
rect 10609 7361 10643 7395
rect 12403 7361 12437 7395
rect 12541 7361 12575 7395
rect 15117 7361 15151 7395
rect 17325 7361 17359 7395
rect 2421 7293 2455 7327
rect 5089 7293 5123 7327
rect 6009 7293 6043 7327
rect 6837 7293 6871 7327
rect 7941 7293 7975 7327
rect 10977 7293 11011 7327
rect 17877 7293 17911 7327
rect 17969 7293 18003 7327
rect 8217 7225 8251 7259
rect 1501 7157 1535 7191
rect 2697 7157 2731 7191
rect 3617 7157 3651 7191
rect 9229 7157 9263 7191
rect 12633 7157 12667 7191
rect 15025 7157 15059 7191
rect 17417 7157 17451 7191
rect 10149 6953 10183 6987
rect 10425 6953 10459 6987
rect 15209 6953 15243 6987
rect 17785 6953 17819 6987
rect 18337 6953 18371 6987
rect 2421 6885 2455 6919
rect 9413 6885 9447 6919
rect 1961 6817 1995 6851
rect 6377 6817 6411 6851
rect 7573 6817 7607 6851
rect 7849 6817 7883 6851
rect 8493 6817 8527 6851
rect 8677 6817 8711 6851
rect 1501 6749 1535 6783
rect 1593 6749 1627 6783
rect 2789 6749 2823 6783
rect 3065 6749 3099 6783
rect 3249 6749 3283 6783
rect 3341 6749 3375 6783
rect 3525 6749 3559 6783
rect 4077 6749 4111 6783
rect 6469 6749 6503 6783
rect 2053 6681 2087 6715
rect 3433 6681 3467 6715
rect 4353 6681 4387 6715
rect 7297 6681 7331 6715
rect 8401 6749 8435 6783
rect 11345 6817 11379 6851
rect 13921 6817 13955 6851
rect 15025 6817 15059 6851
rect 15577 6817 15611 6851
rect 17325 6817 17359 6851
rect 9505 6749 9539 6783
rect 9965 6749 9999 6783
rect 10149 6749 10183 6783
rect 11161 6749 11195 6783
rect 11621 6749 11655 6783
rect 14749 6749 14783 6783
rect 15393 6749 15427 6783
rect 15485 6749 15519 6783
rect 17141 6749 17175 6783
rect 17785 6749 17819 6783
rect 18521 6749 18555 6783
rect 9413 6681 9447 6715
rect 13645 6681 13679 6715
rect 17233 6681 17267 6715
rect 1317 6613 1351 6647
rect 2513 6613 2547 6647
rect 2973 6613 3007 6647
rect 5825 6613 5859 6647
rect 6193 6613 6227 6647
rect 6837 6613 6871 6647
rect 6929 6613 6963 6647
rect 7389 6613 7423 6647
rect 7849 6613 7883 6647
rect 8033 6613 8067 6647
rect 9597 6613 9631 6647
rect 10793 6613 10827 6647
rect 11253 6613 11287 6647
rect 11805 6613 11839 6647
rect 13277 6613 13311 6647
rect 13737 6613 13771 6647
rect 14381 6613 14415 6647
rect 14841 6613 14875 6647
rect 16773 6613 16807 6647
rect 2053 6409 2087 6443
rect 4445 6409 4479 6443
rect 5089 6409 5123 6443
rect 6193 6409 6227 6443
rect 6837 6409 6871 6443
rect 8033 6409 8067 6443
rect 8493 6409 8527 6443
rect 10241 6409 10275 6443
rect 10425 6409 10459 6443
rect 11161 6409 11195 6443
rect 11529 6409 11563 6443
rect 11621 6409 11655 6443
rect 14013 6409 14047 6443
rect 14657 6409 14691 6443
rect 16589 6409 16623 6443
rect 18475 6409 18509 6443
rect 581 6341 615 6375
rect 5641 6341 5675 6375
rect 15025 6341 15059 6375
rect 2329 6273 2363 6307
rect 2421 6273 2455 6307
rect 4629 6273 4663 6307
rect 5733 6273 5767 6307
rect 6101 6273 6135 6307
rect 6285 6273 6319 6307
rect 6377 6273 6411 6307
rect 6561 6273 6595 6307
rect 6653 6273 6687 6307
rect 6745 6273 6779 6307
rect 6929 6273 6963 6307
rect 8401 6273 8435 6307
rect 9965 6273 9999 6307
rect 10149 6273 10183 6307
rect 10241 6273 10275 6307
rect 10793 6273 10827 6307
rect 12265 6273 12299 6307
rect 14289 6273 14323 6307
rect 14749 6273 14783 6307
rect 16405 6273 16439 6307
rect 17049 6273 17083 6307
rect 305 6205 339 6239
rect 2605 6205 2639 6239
rect 4721 6205 4755 6239
rect 5825 6205 5859 6239
rect 8677 6205 8711 6239
rect 10885 6205 10919 6239
rect 11713 6205 11747 6239
rect 12541 6205 12575 6239
rect 14381 6205 14415 6239
rect 14841 6205 14875 6239
rect 16681 6205 16715 6239
rect 5273 6137 5307 6171
rect 6561 6137 6595 6171
rect 2513 6069 2547 6103
rect 11069 6069 11103 6103
rect 14933 6069 14967 6103
rect 4491 5865 4525 5899
rect 7619 5865 7653 5899
rect 10057 5865 10091 5899
rect 13001 5865 13035 5899
rect 15117 5865 15151 5899
rect 16693 5865 16727 5899
rect 5825 5729 5859 5763
rect 6193 5729 6227 5763
rect 14841 5729 14875 5763
rect 15209 5729 15243 5763
rect 16957 5729 16991 5763
rect 2329 5661 2363 5695
rect 2421 5661 2455 5695
rect 2697 5661 2731 5695
rect 3065 5661 3099 5695
rect 9873 5661 9907 5695
rect 11805 5661 11839 5695
rect 13185 5661 13219 5695
rect 14749 5661 14783 5695
rect 18521 5661 18555 5695
rect 11529 5593 11563 5627
rect 8585 5525 8619 5559
rect 18337 5525 18371 5559
rect 9321 5321 9355 5355
rect 10885 5321 10919 5355
rect 8585 5253 8619 5287
rect 8769 5253 8803 5287
rect 9045 5253 9079 5287
rect 10793 5253 10827 5287
rect 5733 5185 5767 5219
rect 7573 5185 7607 5219
rect 7757 5185 7791 5219
rect 8033 5185 8067 5219
rect 8859 5185 8893 5219
rect 8953 5175 8987 5209
rect 9229 5185 9263 5219
rect 9781 5185 9815 5219
rect 12357 5185 12391 5219
rect 18521 5185 18555 5219
rect 7665 5117 7699 5151
rect 7941 5117 7975 5151
rect 8401 5117 8435 5151
rect 12265 5117 12299 5151
rect 12725 5117 12759 5151
rect 14289 5117 14323 5151
rect 14565 5117 14599 5151
rect 18245 5117 18279 5151
rect 8677 5049 8711 5083
rect 12817 5049 12851 5083
rect 5825 4981 5859 5015
rect 9965 4981 9999 5015
rect 16773 4981 16807 5015
rect 5089 4777 5123 4811
rect 12265 4777 12299 4811
rect 14105 4777 14139 4811
rect 9689 4641 9723 4675
rect 9781 4641 9815 4675
rect 15853 4641 15887 4675
rect 17693 4641 17727 4675
rect 2329 4573 2363 4607
rect 2421 4573 2455 4607
rect 2697 4573 2731 4607
rect 3065 4573 3099 4607
rect 4491 4573 4525 4607
rect 4813 4573 4847 4607
rect 6837 4573 6871 4607
rect 7205 4573 7239 4607
rect 7849 4573 7883 4607
rect 8217 4573 8251 4607
rect 12357 4573 12391 4607
rect 12443 4573 12477 4607
rect 12547 4573 12581 4607
rect 12725 4573 12759 4607
rect 17969 4573 18003 4607
rect 18521 4573 18555 4607
rect 6561 4505 6595 4539
rect 7021 4505 7055 4539
rect 10057 4505 10091 4539
rect 12173 4505 12207 4539
rect 15577 4505 15611 4539
rect 15945 4505 15979 4539
rect 4721 4437 4755 4471
rect 11529 4437 11563 4471
rect 12633 4437 12667 4471
rect 18337 4437 18371 4471
rect 3249 4233 3283 4267
rect 8033 4233 8067 4267
rect 8769 4233 8803 4267
rect 9229 4233 9263 4267
rect 10425 4233 10459 4267
rect 10793 4233 10827 4267
rect 11253 4233 11287 4267
rect 9597 4165 9631 4199
rect 11621 4165 11655 4199
rect 16313 4165 16347 4199
rect 3525 4097 3559 4131
rect 4905 4097 4939 4131
rect 5089 4097 5123 4131
rect 6745 4097 6779 4131
rect 6929 4097 6963 4131
rect 7205 4097 7239 4131
rect 7481 4097 7515 4131
rect 7849 4097 7883 4131
rect 8861 4097 8895 4131
rect 10885 4097 10919 4131
rect 12081 4097 12115 4131
rect 12265 4097 12299 4131
rect 12449 4097 12483 4131
rect 12541 4097 12575 4131
rect 12629 4097 12663 4131
rect 13369 4097 13403 4131
rect 14381 4097 14415 4131
rect 14565 4097 14599 4131
rect 16129 4097 16163 4131
rect 3249 4029 3283 4063
rect 6377 4029 6411 4063
rect 6653 4029 6687 4063
rect 7113 4029 7147 4063
rect 8953 4029 8987 4063
rect 9689 4029 9723 4063
rect 9873 4029 9907 4063
rect 10977 4029 11011 4063
rect 11713 4029 11747 4063
rect 11805 4029 11839 4063
rect 12817 4029 12851 4063
rect 13277 4029 13311 4063
rect 17877 4029 17911 4063
rect 18521 4029 18555 4063
rect 8401 3961 8435 3995
rect 12173 3961 12207 3995
rect 3433 3893 3467 3927
rect 4905 3893 4939 3927
rect 6837 3893 6871 3927
rect 13645 3893 13679 3927
rect 14381 3893 14415 3927
rect 17417 3893 17451 3927
rect 18061 3893 18095 3927
rect 4169 3689 4203 3723
rect 5641 3689 5675 3723
rect 5733 3689 5767 3723
rect 7941 3689 7975 3723
rect 9597 3689 9631 3723
rect 10885 3689 10919 3723
rect 3893 3621 3927 3655
rect 5917 3621 5951 3655
rect 6285 3621 6319 3655
rect 8585 3621 8619 3655
rect 18153 3621 18187 3655
rect 765 3553 799 3587
rect 2513 3553 2547 3587
rect 3341 3553 3375 3587
rect 6929 3553 6963 3587
rect 7113 3553 7147 3587
rect 9045 3553 9079 3587
rect 10517 3553 10551 3587
rect 13829 3553 13863 3587
rect 15853 3553 15887 3587
rect 17601 3553 17635 3587
rect 2881 3485 2915 3519
rect 2973 3485 3007 3519
rect 3617 3485 3651 3519
rect 3893 3485 3927 3519
rect 4077 3485 4111 3519
rect 4353 3485 4387 3519
rect 4445 3485 4479 3519
rect 4537 3485 4571 3519
rect 4997 3485 5031 3519
rect 5273 3485 5307 3519
rect 5825 3485 5859 3519
rect 5917 3485 5951 3519
rect 6101 3485 6135 3519
rect 8033 3485 8067 3519
rect 8217 3485 8251 3519
rect 9137 3485 9171 3519
rect 9781 3485 9815 3519
rect 10609 3485 10643 3519
rect 14197 3485 14231 3519
rect 16221 3485 16255 3519
rect 18337 3485 18371 3519
rect 1041 3417 1075 3451
rect 2697 3417 2731 3451
rect 7849 3417 7883 3451
rect 4813 3349 4847 3383
rect 5365 3349 5399 3383
rect 6653 3349 6687 3383
rect 6745 3349 6779 3383
rect 7573 3349 7607 3383
rect 9229 3349 9263 3383
rect 15623 3349 15657 3383
rect 3433 3145 3467 3179
rect 3617 3145 3651 3179
rect 5549 3145 5583 3179
rect 14565 3145 14599 3179
rect 15991 3145 16025 3179
rect 18337 3145 18371 3179
rect 2973 3077 3007 3111
rect 8125 3077 8159 3111
rect 8309 3077 8343 3111
rect 12909 3077 12943 3111
rect 14473 3077 14507 3111
rect 3709 3009 3743 3043
rect 4813 3009 4847 3043
rect 5549 3009 5583 3043
rect 5917 3009 5951 3043
rect 6009 3009 6043 3043
rect 6193 3009 6227 3043
rect 7113 3009 7147 3043
rect 7389 3009 7423 3043
rect 7573 3009 7607 3043
rect 7665 3009 7699 3043
rect 7849 3009 7883 3043
rect 8401 3009 8435 3043
rect 12541 3009 12575 3043
rect 12817 3009 12851 3043
rect 13185 3009 13219 3043
rect 14013 3009 14047 3043
rect 17785 3009 17819 3043
rect 4905 2941 4939 2975
rect 5365 2941 5399 2975
rect 5641 2941 5675 2975
rect 5825 2941 5859 2975
rect 8769 2941 8803 2975
rect 10425 2941 10459 2975
rect 10793 2941 10827 2975
rect 14657 2941 14691 2975
rect 17417 2941 17451 2975
rect 17877 2941 17911 2975
rect 3341 2873 3375 2907
rect 6101 2873 6135 2907
rect 7757 2873 7791 2907
rect 13553 2873 13587 2907
rect 13737 2873 13771 2907
rect 14105 2873 14139 2907
rect 5365 2805 5399 2839
rect 7205 2805 7239 2839
rect 10195 2805 10229 2839
rect 12219 2805 12253 2839
rect 6837 2601 6871 2635
rect 12265 2601 12299 2635
rect 3157 2533 3191 2567
rect 3249 2533 3283 2567
rect 5825 2533 5859 2567
rect 12173 2533 12207 2567
rect 765 2465 799 2499
rect 1041 2465 1075 2499
rect 3065 2465 3099 2499
rect 4169 2465 4203 2499
rect 4997 2465 5031 2499
rect 5181 2465 5215 2499
rect 10149 2465 10183 2499
rect 11713 2465 11747 2499
rect 15393 2465 15427 2499
rect 15761 2465 15795 2499
rect 17969 2465 18003 2499
rect 3341 2397 3375 2431
rect 4445 2397 4479 2431
rect 5641 2397 5675 2431
rect 5825 2397 5859 2431
rect 6101 2397 6135 2431
rect 6745 2397 6779 2431
rect 6837 2397 6871 2431
rect 7481 2397 7515 2431
rect 8585 2397 8619 2431
rect 8677 2397 8711 2431
rect 10241 2397 10275 2431
rect 11805 2397 11839 2431
rect 12265 2397 12299 2431
rect 12633 2397 12667 2431
rect 15485 2397 15519 2431
rect 15577 2397 15611 2431
rect 18521 2397 18555 2431
rect 4905 2329 4939 2363
rect 6561 2329 6595 2363
rect 8861 2329 8895 2363
rect 12357 2329 12391 2363
rect 12541 2329 12575 2363
rect 15148 2329 15182 2363
rect 15945 2329 15979 2363
rect 17693 2329 17727 2363
rect 2513 2261 2547 2295
rect 4537 2261 4571 2295
rect 7573 2261 7607 2295
rect 8769 2261 8803 2295
rect 12725 2261 12759 2295
rect 14013 2261 14047 2295
rect 15761 2261 15795 2295
rect 18337 2261 18371 2295
rect 3525 2057 3559 2091
rect 3709 2057 3743 2091
rect 4353 2057 4387 2091
rect 6469 2057 6503 2091
rect 9137 2057 9171 2091
rect 9873 2057 9907 2091
rect 10517 2057 10551 2091
rect 10977 2057 11011 2091
rect 12265 2057 12299 2091
rect 13093 2057 13127 2091
rect 14289 2057 14323 2091
rect 14841 2057 14875 2091
rect 17417 2057 17451 2091
rect 15945 1989 15979 2023
rect 3617 1921 3651 1955
rect 3709 1921 3743 1955
rect 3893 1921 3927 1955
rect 5457 1921 5491 1955
rect 6377 1921 6411 1955
rect 7389 1921 7423 1955
rect 10885 1921 10919 1955
rect 12437 1921 12471 1955
rect 12541 1921 12575 1955
rect 12633 1921 12667 1955
rect 12817 1921 12851 1955
rect 13001 1921 13035 1955
rect 13277 1921 13311 1955
rect 14105 1921 14139 1955
rect 14197 1921 14231 1955
rect 14381 1921 14415 1955
rect 14657 1921 14691 1955
rect 15117 1921 15151 1955
rect 15669 1921 15703 1955
rect 4445 1853 4479 1887
rect 4537 1853 4571 1887
rect 5549 1853 5583 1887
rect 5825 1853 5859 1887
rect 6561 1853 6595 1887
rect 7665 1853 7699 1887
rect 9965 1853 9999 1887
rect 10149 1853 10183 1887
rect 11161 1853 11195 1887
rect 3985 1785 4019 1819
rect 14473 1853 14507 1887
rect 15393 1853 15427 1887
rect 14933 1785 14967 1819
rect 6009 1717 6043 1751
rect 9505 1717 9539 1751
rect 14105 1717 14139 1751
rect 15301 1717 15335 1751
rect 2973 1513 3007 1547
rect 5549 1513 5583 1547
rect 10609 1513 10643 1547
rect 2881 1445 2915 1479
rect 3525 1445 3559 1479
rect 765 1377 799 1411
rect 1041 1377 1075 1411
rect 2789 1377 2823 1411
rect 3985 1377 4019 1411
rect 6101 1377 6135 1411
rect 6285 1377 6319 1411
rect 8769 1377 8803 1411
rect 10149 1377 10183 1411
rect 14105 1377 14139 1411
rect 16497 1377 16531 1411
rect 16589 1377 16623 1411
rect 3065 1309 3099 1343
rect 3525 1309 3559 1343
rect 3709 1309 3743 1343
rect 3801 1309 3835 1343
rect 3893 1309 3927 1343
rect 4077 1309 4111 1343
rect 4445 1309 4479 1343
rect 4997 1309 5031 1343
rect 5181 1309 5215 1343
rect 5365 1309 5399 1343
rect 5549 1309 5583 1343
rect 6009 1309 6043 1343
rect 6469 1309 6503 1343
rect 8493 1309 8527 1343
rect 8677 1309 8711 1343
rect 9137 1309 9171 1343
rect 10241 1309 10275 1343
rect 11161 1309 11195 1343
rect 11253 1309 11287 1343
rect 12633 1309 12667 1343
rect 12725 1309 12759 1343
rect 14013 1309 14047 1343
rect 18245 1309 18279 1343
rect 18337 1309 18371 1343
rect 3249 1241 3283 1275
rect 3433 1241 3467 1275
rect 10885 1241 10919 1275
rect 11069 1241 11103 1275
rect 11345 1241 11379 1275
rect 14473 1241 14507 1275
rect 16221 1241 16255 1275
rect 16834 1241 16868 1275
rect 2513 1173 2547 1207
rect 5181 1173 5215 1207
rect 5641 1173 5675 1207
rect 6929 1173 6963 1207
rect 11161 1173 11195 1207
rect 13553 1173 13587 1207
rect 13921 1173 13955 1207
rect 17969 1173 18003 1207
rect 5825 969 5859 1003
rect 6377 969 6411 1003
rect 6469 969 6503 1003
rect 9597 969 9631 1003
rect 9965 969 9999 1003
rect 10149 969 10183 1003
rect 10517 969 10551 1003
rect 11437 969 11471 1003
rect 12449 969 12483 1003
rect 12541 969 12575 1003
rect 13645 969 13679 1003
rect 13737 969 13771 1003
rect 14197 969 14231 1003
rect 16037 969 16071 1003
rect 17325 969 17359 1003
rect 9505 901 9539 935
rect 3249 833 3283 867
rect 3801 833 3835 867
rect 3893 833 3927 867
rect 3985 833 4019 867
rect 4169 833 4203 867
rect 5457 833 5491 867
rect 2973 765 3007 799
rect 4077 765 4111 799
rect 5549 765 5583 799
rect 6561 765 6595 799
rect 7205 765 7239 799
rect 7573 765 7607 799
rect 9781 765 9815 799
rect 3157 697 3191 731
rect 8999 697 9033 731
rect 12357 901 12391 935
rect 17233 901 17267 935
rect 10057 833 10091 867
rect 10241 833 10275 867
rect 10885 833 10919 867
rect 11345 833 11379 867
rect 12173 833 12207 867
rect 12449 833 12483 867
rect 14197 833 14231 867
rect 15853 833 15887 867
rect 16957 833 16991 867
rect 17049 833 17083 867
rect 17785 833 17819 867
rect 18337 833 18371 867
rect 3065 629 3099 663
rect 6009 629 6043 663
rect 9137 629 9171 663
rect 9965 629 9999 663
rect 10425 765 10459 799
rect 10977 765 11011 799
rect 11161 765 11195 799
rect 12909 765 12943 799
rect 13001 765 13035 799
rect 13875 765 13909 799
rect 15577 765 15611 799
rect 17877 765 17911 799
rect 13277 697 13311 731
rect 15669 697 15703 731
rect 16957 697 16991 731
rect 10425 629 10459 663
rect 13185 629 13219 663
rect 17693 629 17727 663
rect 18061 629 18095 663
rect 5641 425 5675 459
rect 8125 425 8159 459
rect 10885 425 10919 459
rect 14749 425 14783 459
rect 17509 425 17543 459
rect 18337 425 18371 459
rect 4491 357 4525 391
rect 3065 289 3099 323
rect 6101 289 6135 323
rect 6285 289 6319 323
rect 8309 289 8343 323
rect 8401 289 8435 323
rect 10701 289 10735 323
rect 13001 289 13035 323
rect 16129 289 16163 323
rect 2329 221 2363 255
rect 2421 221 2455 255
rect 2697 221 2731 255
rect 6009 221 6043 255
rect 8861 221 8895 255
rect 8953 221 8987 255
rect 10609 221 10643 255
rect 18521 221 18555 255
rect 9137 153 9171 187
rect 13277 153 13311 187
rect 16374 153 16408 187
rect 8769 85 8803 119
rect 8861 85 8895 119
<< metal1 >>
rect 0 10906 18860 10928
rect 0 10854 4660 10906
rect 4712 10854 4724 10906
rect 4776 10854 4788 10906
rect 4840 10854 4852 10906
rect 4904 10854 4916 10906
rect 4968 10854 7760 10906
rect 7812 10854 7824 10906
rect 7876 10854 7888 10906
rect 7940 10854 7952 10906
rect 8004 10854 8016 10906
rect 8068 10854 10860 10906
rect 10912 10854 10924 10906
rect 10976 10854 10988 10906
rect 11040 10854 11052 10906
rect 11104 10854 11116 10906
rect 11168 10854 13960 10906
rect 14012 10854 14024 10906
rect 14076 10854 14088 10906
rect 14140 10854 14152 10906
rect 14204 10854 14216 10906
rect 14268 10854 17060 10906
rect 17112 10854 17124 10906
rect 17176 10854 17188 10906
rect 17240 10854 17252 10906
rect 17304 10854 17316 10906
rect 17368 10854 18860 10906
rect 0 10832 18860 10854
rect 3786 10792 3792 10804
rect 2332 10764 3792 10792
rect 2130 10684 2136 10736
rect 2188 10724 2194 10736
rect 2332 10733 2360 10764
rect 2317 10727 2375 10733
rect 2317 10724 2329 10727
rect 2188 10696 2329 10724
rect 2188 10684 2194 10696
rect 2317 10693 2329 10696
rect 2363 10693 2375 10727
rect 3436 10710 3464 10764
rect 3786 10752 3792 10764
rect 3844 10752 3850 10804
rect 6917 10795 6975 10801
rect 6917 10761 6929 10795
rect 6963 10792 6975 10795
rect 7098 10792 7104 10804
rect 6963 10764 7104 10792
rect 6963 10761 6975 10764
rect 6917 10755 6975 10761
rect 7098 10752 7104 10764
rect 7156 10752 7162 10804
rect 7193 10795 7251 10801
rect 7193 10761 7205 10795
rect 7239 10761 7251 10795
rect 7193 10755 7251 10761
rect 7208 10724 7236 10755
rect 9950 10752 9956 10804
rect 10008 10792 10014 10804
rect 10965 10795 11023 10801
rect 10965 10792 10977 10795
rect 10008 10764 10977 10792
rect 10008 10752 10014 10764
rect 10965 10761 10977 10764
rect 11011 10761 11023 10795
rect 10965 10755 11023 10761
rect 15948 10764 16896 10792
rect 15948 10736 15976 10764
rect 8082 10727 8140 10733
rect 8082 10724 8094 10727
rect 7208 10696 8094 10724
rect 2317 10687 2375 10693
rect 8082 10693 8094 10696
rect 8128 10693 8140 10727
rect 13354 10724 13360 10736
rect 8082 10687 8140 10693
rect 10796 10696 13360 10724
rect 1302 10656 1308 10668
rect 1263 10628 1308 10656
rect 1302 10616 1308 10628
rect 1360 10616 1366 10668
rect 5445 10659 5503 10665
rect 5445 10656 5457 10659
rect 4356 10628 5457 10656
rect 2682 10588 2688 10600
rect 2643 10560 2688 10588
rect 2682 10548 2688 10560
rect 2740 10548 2746 10600
rect 2958 10548 2964 10600
rect 3016 10588 3022 10600
rect 3053 10591 3111 10597
rect 3053 10588 3065 10591
rect 3016 10560 3065 10588
rect 3016 10548 3022 10560
rect 3053 10557 3065 10560
rect 3099 10557 3111 10591
rect 3053 10551 3111 10557
rect 4356 10464 4384 10628
rect 5445 10625 5457 10628
rect 5491 10625 5503 10659
rect 6730 10656 6736 10668
rect 6691 10628 6736 10656
rect 5445 10619 5503 10625
rect 6730 10616 6736 10628
rect 6788 10616 6794 10668
rect 7006 10656 7012 10668
rect 6967 10628 7012 10656
rect 7006 10616 7012 10628
rect 7064 10616 7070 10668
rect 7377 10659 7435 10665
rect 7377 10625 7389 10659
rect 7423 10656 7435 10659
rect 9214 10656 9220 10668
rect 7423 10628 9220 10656
rect 7423 10625 7435 10628
rect 7377 10619 7435 10625
rect 9214 10616 9220 10628
rect 9272 10616 9278 10668
rect 9309 10659 9367 10665
rect 9309 10625 9321 10659
rect 9355 10625 9367 10659
rect 10410 10656 10416 10668
rect 10371 10628 10416 10656
rect 9309 10619 9367 10625
rect 5537 10591 5595 10597
rect 5537 10557 5549 10591
rect 5583 10588 5595 10591
rect 5994 10588 6000 10600
rect 5583 10560 6000 10588
rect 5583 10557 5595 10560
rect 5537 10551 5595 10557
rect 5994 10548 6000 10560
rect 6052 10548 6058 10600
rect 7650 10548 7656 10600
rect 7708 10588 7714 10600
rect 7837 10591 7895 10597
rect 7837 10588 7849 10591
rect 7708 10560 7849 10588
rect 7708 10548 7714 10560
rect 7837 10557 7849 10560
rect 7883 10557 7895 10591
rect 9324 10588 9352 10619
rect 10410 10616 10416 10628
rect 10468 10616 10474 10668
rect 7837 10551 7895 10557
rect 9232 10560 9352 10588
rect 2314 10412 2320 10464
rect 2372 10452 2378 10464
rect 4338 10452 4344 10464
rect 2372 10424 4344 10452
rect 2372 10412 2378 10424
rect 4338 10412 4344 10424
rect 4396 10412 4402 10464
rect 4430 10412 4436 10464
rect 4488 10461 4494 10464
rect 4488 10455 4537 10461
rect 4488 10421 4491 10455
rect 4525 10421 4537 10455
rect 5810 10452 5816 10464
rect 5771 10424 5816 10452
rect 4488 10415 4537 10421
rect 4488 10412 4494 10415
rect 5810 10412 5816 10424
rect 5868 10412 5874 10464
rect 7466 10452 7472 10464
rect 7427 10424 7472 10452
rect 7466 10412 7472 10424
rect 7524 10412 7530 10464
rect 9030 10412 9036 10464
rect 9088 10452 9094 10464
rect 9232 10461 9260 10560
rect 9674 10480 9680 10532
rect 9732 10520 9738 10532
rect 10796 10520 10824 10696
rect 13354 10684 13360 10696
rect 13412 10684 13418 10736
rect 15930 10724 15936 10736
rect 14674 10696 15936 10724
rect 15930 10684 15936 10696
rect 15988 10684 15994 10736
rect 16868 10710 16896 10764
rect 11149 10659 11207 10665
rect 11149 10625 11161 10659
rect 11195 10656 11207 10659
rect 11195 10628 11928 10656
rect 11195 10625 11207 10628
rect 11149 10619 11207 10625
rect 11900 10529 11928 10628
rect 12158 10616 12164 10668
rect 12216 10656 12222 10668
rect 12253 10659 12311 10665
rect 12253 10656 12265 10659
rect 12216 10628 12265 10656
rect 12216 10616 12222 10628
rect 12253 10625 12265 10628
rect 12299 10625 12311 10659
rect 13262 10656 13268 10668
rect 13175 10628 13268 10656
rect 12253 10619 12311 10625
rect 13262 10616 13268 10628
rect 13320 10656 13326 10668
rect 17911 10659 17969 10665
rect 13320 10628 13768 10656
rect 13320 10616 13326 10628
rect 12345 10591 12403 10597
rect 12345 10557 12357 10591
rect 12391 10557 12403 10591
rect 12345 10551 12403 10557
rect 12437 10591 12495 10597
rect 12437 10557 12449 10591
rect 12483 10557 12495 10591
rect 13630 10588 13636 10600
rect 13591 10560 13636 10588
rect 12437 10551 12495 10557
rect 9732 10492 10824 10520
rect 11885 10523 11943 10529
rect 9732 10480 9738 10492
rect 9217 10455 9275 10461
rect 9217 10452 9229 10455
rect 9088 10424 9229 10452
rect 9088 10412 9094 10424
rect 9217 10421 9229 10424
rect 9263 10421 9275 10455
rect 9950 10452 9956 10464
rect 9911 10424 9956 10452
rect 9217 10415 9275 10421
rect 9950 10412 9956 10424
rect 10008 10412 10014 10464
rect 10704 10461 10732 10492
rect 11885 10489 11897 10523
rect 11931 10489 11943 10523
rect 11885 10483 11943 10489
rect 12250 10480 12256 10532
rect 12308 10520 12314 10532
rect 12360 10520 12388 10551
rect 12308 10492 12388 10520
rect 12308 10480 12314 10492
rect 10689 10455 10747 10461
rect 10689 10421 10701 10455
rect 10735 10421 10747 10455
rect 10689 10415 10747 10421
rect 10778 10412 10784 10464
rect 10836 10452 10842 10464
rect 10873 10455 10931 10461
rect 10873 10452 10885 10455
rect 10836 10424 10885 10452
rect 10836 10412 10842 10424
rect 10873 10421 10885 10424
rect 10919 10421 10931 10455
rect 10873 10415 10931 10421
rect 12066 10412 12072 10464
rect 12124 10452 12130 10464
rect 12452 10452 12480 10551
rect 13630 10548 13636 10560
rect 13688 10548 13694 10600
rect 13740 10588 13768 10628
rect 17911 10625 17923 10659
rect 17957 10656 17969 10659
rect 18141 10659 18199 10665
rect 18141 10656 18153 10659
rect 17957 10628 18153 10656
rect 17957 10625 17969 10628
rect 17911 10619 17969 10625
rect 18141 10625 18153 10628
rect 18187 10625 18199 10659
rect 18322 10656 18328 10668
rect 18283 10628 18328 10656
rect 18141 10619 18199 10625
rect 18322 10616 18328 10628
rect 18380 10616 18386 10668
rect 14826 10588 14832 10600
rect 13740 10560 14832 10588
rect 14826 10548 14832 10560
rect 14884 10588 14890 10600
rect 16117 10591 16175 10597
rect 16117 10588 16129 10591
rect 14884 10560 16129 10588
rect 14884 10548 14890 10560
rect 16117 10557 16129 10560
rect 16163 10557 16175 10591
rect 16482 10588 16488 10600
rect 16443 10560 16488 10588
rect 16117 10551 16175 10557
rect 16482 10548 16488 10560
rect 16540 10548 16546 10600
rect 12124 10424 12480 10452
rect 15059 10455 15117 10461
rect 12124 10412 12130 10424
rect 15059 10421 15071 10455
rect 15105 10452 15117 10455
rect 15194 10452 15200 10464
rect 15105 10424 15200 10452
rect 15105 10421 15117 10424
rect 15059 10415 15117 10421
rect 15194 10412 15200 10424
rect 15252 10412 15258 10464
rect 15286 10412 15292 10464
rect 15344 10452 15350 10464
rect 18141 10455 18199 10461
rect 18141 10452 18153 10455
rect 15344 10424 18153 10452
rect 15344 10412 15350 10424
rect 18141 10421 18153 10424
rect 18187 10421 18199 10455
rect 18141 10415 18199 10421
rect 0 10362 18860 10384
rect 0 10310 3110 10362
rect 3162 10310 3174 10362
rect 3226 10310 3238 10362
rect 3290 10310 3302 10362
rect 3354 10310 3366 10362
rect 3418 10310 6210 10362
rect 6262 10310 6274 10362
rect 6326 10310 6338 10362
rect 6390 10310 6402 10362
rect 6454 10310 6466 10362
rect 6518 10310 9310 10362
rect 9362 10310 9374 10362
rect 9426 10310 9438 10362
rect 9490 10310 9502 10362
rect 9554 10310 9566 10362
rect 9618 10310 12410 10362
rect 12462 10310 12474 10362
rect 12526 10310 12538 10362
rect 12590 10310 12602 10362
rect 12654 10310 12666 10362
rect 12718 10310 15510 10362
rect 15562 10310 15574 10362
rect 15626 10310 15638 10362
rect 15690 10310 15702 10362
rect 15754 10310 15766 10362
rect 15818 10310 18860 10362
rect 0 10288 18860 10310
rect 2682 10208 2688 10260
rect 2740 10248 2746 10260
rect 3513 10251 3571 10257
rect 3513 10248 3525 10251
rect 2740 10220 3525 10248
rect 2740 10208 2746 10220
rect 3513 10217 3525 10220
rect 3559 10217 3571 10251
rect 5261 10251 5319 10257
rect 5261 10248 5273 10251
rect 3513 10211 3571 10217
rect 4172 10220 5273 10248
rect 1596 10152 3648 10180
rect 290 10112 296 10124
rect 203 10084 296 10112
rect 290 10072 296 10084
rect 348 10112 354 10124
rect 1596 10112 1624 10152
rect 348 10084 1624 10112
rect 2041 10115 2099 10121
rect 348 10072 354 10084
rect 2041 10081 2053 10115
rect 2087 10112 2099 10115
rect 2087 10084 2360 10112
rect 2087 10081 2099 10084
rect 2041 10075 2099 10081
rect 2332 10056 2360 10084
rect 2958 10072 2964 10124
rect 3016 10072 3022 10124
rect 3053 10115 3111 10121
rect 3053 10081 3065 10115
rect 3099 10112 3111 10115
rect 3418 10112 3424 10124
rect 3099 10084 3424 10112
rect 3099 10081 3111 10084
rect 3053 10075 3111 10081
rect 3418 10072 3424 10084
rect 3476 10072 3482 10124
rect 2314 10044 2320 10056
rect 2275 10016 2320 10044
rect 2314 10004 2320 10016
rect 2372 10004 2378 10056
rect 2685 10047 2743 10053
rect 2685 10013 2697 10047
rect 2731 10013 2743 10047
rect 2976 10044 3004 10072
rect 3234 10044 3240 10056
rect 2976 10016 3096 10044
rect 3195 10016 3240 10044
rect 2685 10007 2743 10013
rect 566 9976 572 9988
rect 527 9948 572 9976
rect 566 9936 572 9948
rect 624 9936 630 9988
rect 2130 9976 2136 9988
rect 1794 9948 2136 9976
rect 2130 9936 2136 9948
rect 2188 9936 2194 9988
rect 2700 9976 2728 10007
rect 2240 9948 2728 9976
rect 2777 9979 2835 9985
rect 2240 9920 2268 9948
rect 2777 9945 2789 9979
rect 2823 9945 2835 9979
rect 2777 9939 2835 9945
rect 2222 9908 2228 9920
rect 2183 9880 2228 9908
rect 2222 9868 2228 9880
rect 2280 9868 2286 9920
rect 2682 9908 2688 9920
rect 2643 9880 2688 9908
rect 2682 9868 2688 9880
rect 2740 9868 2746 9920
rect 2792 9908 2820 9939
rect 2866 9936 2872 9988
rect 2924 9976 2930 9988
rect 3068 9985 3096 10016
rect 3234 10004 3240 10016
rect 3292 10004 3298 10056
rect 3620 10053 3648 10152
rect 3329 10047 3387 10053
rect 3329 10013 3341 10047
rect 3375 10013 3387 10047
rect 3329 10007 3387 10013
rect 3605 10047 3663 10053
rect 3605 10013 3617 10047
rect 3651 10013 3663 10047
rect 3605 10007 3663 10013
rect 3881 10047 3939 10053
rect 3881 10013 3893 10047
rect 3927 10013 3939 10047
rect 3881 10007 3939 10013
rect 2961 9979 3019 9985
rect 2961 9976 2973 9979
rect 2924 9948 2973 9976
rect 2924 9936 2930 9948
rect 2961 9945 2973 9948
rect 3007 9945 3019 9979
rect 2961 9939 3019 9945
rect 3053 9979 3111 9985
rect 3053 9945 3065 9979
rect 3099 9945 3111 9979
rect 3053 9939 3111 9945
rect 3344 9976 3372 10007
rect 3789 9979 3847 9985
rect 3789 9976 3801 9979
rect 3344 9948 3801 9976
rect 3344 9908 3372 9948
rect 3789 9945 3801 9948
rect 3835 9945 3847 9979
rect 3896 9976 3924 10007
rect 4062 10004 4068 10056
rect 4120 10044 4126 10056
rect 4172 10044 4200 10220
rect 5261 10217 5273 10220
rect 5307 10217 5319 10251
rect 5994 10248 6000 10260
rect 5955 10220 6000 10248
rect 5261 10211 5319 10217
rect 5994 10208 6000 10220
rect 6052 10208 6058 10260
rect 7006 10208 7012 10260
rect 7064 10248 7070 10260
rect 7929 10251 7987 10257
rect 7929 10248 7941 10251
rect 7064 10220 7941 10248
rect 7064 10208 7070 10220
rect 7929 10217 7941 10220
rect 7975 10217 7987 10251
rect 7929 10211 7987 10217
rect 9214 10208 9220 10260
rect 9272 10248 9278 10260
rect 10873 10251 10931 10257
rect 10873 10248 10885 10251
rect 9272 10220 10885 10248
rect 9272 10208 9278 10220
rect 10873 10217 10885 10220
rect 10919 10217 10931 10251
rect 10873 10211 10931 10217
rect 4246 10140 4252 10192
rect 4304 10180 4310 10192
rect 4304 10152 9628 10180
rect 4304 10140 4310 10152
rect 4338 10072 4344 10124
rect 4396 10112 4402 10124
rect 5261 10115 5319 10121
rect 4396 10084 5028 10112
rect 4396 10072 4402 10084
rect 5000 10053 5028 10084
rect 5261 10081 5273 10115
rect 5307 10112 5319 10115
rect 5445 10115 5503 10121
rect 5445 10112 5457 10115
rect 5307 10084 5457 10112
rect 5307 10081 5319 10084
rect 5261 10075 5319 10081
rect 5445 10081 5457 10084
rect 5491 10112 5503 10115
rect 8389 10115 8447 10121
rect 5491 10084 6040 10112
rect 5491 10081 5503 10084
rect 5445 10075 5503 10081
rect 6012 10053 6040 10084
rect 8389 10081 8401 10115
rect 8435 10112 8447 10115
rect 9030 10112 9036 10124
rect 8435 10084 9036 10112
rect 8435 10081 8447 10084
rect 8389 10075 8447 10081
rect 9030 10072 9036 10084
rect 9088 10072 9094 10124
rect 4249 10047 4307 10053
rect 4249 10044 4261 10047
rect 4120 10016 4261 10044
rect 4120 10004 4126 10016
rect 4249 10013 4261 10016
rect 4295 10013 4307 10047
rect 4249 10007 4307 10013
rect 4801 10047 4859 10053
rect 4801 10013 4813 10047
rect 4847 10013 4859 10047
rect 4801 10007 4859 10013
rect 4985 10047 5043 10053
rect 4985 10013 4997 10047
rect 5031 10013 5043 10047
rect 4985 10007 5043 10013
rect 5537 10047 5595 10053
rect 5537 10013 5549 10047
rect 5583 10013 5595 10047
rect 5537 10007 5595 10013
rect 5997 10047 6055 10053
rect 5997 10013 6009 10047
rect 6043 10013 6055 10047
rect 5997 10007 6055 10013
rect 6181 10047 6239 10053
rect 6181 10013 6193 10047
rect 6227 10013 6239 10047
rect 6181 10007 6239 10013
rect 4430 9976 4436 9988
rect 3896 9948 4436 9976
rect 3789 9939 3847 9945
rect 4430 9936 4436 9948
rect 4488 9976 4494 9988
rect 4816 9976 4844 10007
rect 5552 9976 5580 10007
rect 6196 9976 6224 10007
rect 7466 10004 7472 10056
rect 7524 10044 7530 10056
rect 8938 10044 8944 10056
rect 7524 10016 8432 10044
rect 8899 10016 8944 10044
rect 7524 10004 7530 10016
rect 8404 9985 8432 10016
rect 8938 10004 8944 10016
rect 8996 10004 9002 10056
rect 9122 10044 9128 10056
rect 9083 10016 9128 10044
rect 9122 10004 9128 10016
rect 9180 10004 9186 10056
rect 9600 10053 9628 10152
rect 9585 10047 9643 10053
rect 9585 10013 9597 10047
rect 9631 10013 9643 10047
rect 10888 10044 10916 10211
rect 12802 10208 12808 10260
rect 12860 10248 12866 10260
rect 13081 10251 13139 10257
rect 13081 10248 13093 10251
rect 12860 10220 13093 10248
rect 12860 10208 12866 10220
rect 13081 10217 13093 10220
rect 13127 10217 13139 10251
rect 13630 10248 13636 10260
rect 13591 10220 13636 10248
rect 13081 10211 13139 10217
rect 13630 10208 13636 10220
rect 13688 10208 13694 10260
rect 16482 10208 16488 10260
rect 16540 10248 16546 10260
rect 16623 10251 16681 10257
rect 16623 10248 16635 10251
rect 16540 10220 16635 10248
rect 16540 10208 16546 10220
rect 16623 10217 16635 10220
rect 16669 10217 16681 10251
rect 18322 10248 18328 10260
rect 18283 10220 18328 10248
rect 16623 10211 16681 10217
rect 18322 10208 18328 10220
rect 18380 10208 18386 10260
rect 14826 10112 14832 10124
rect 14787 10084 14832 10112
rect 14826 10072 14832 10084
rect 14884 10072 14890 10124
rect 15194 10112 15200 10124
rect 15155 10084 15200 10112
rect 15194 10072 15200 10084
rect 15252 10072 15258 10124
rect 12069 10047 12127 10053
rect 12069 10044 12081 10047
rect 10888 10016 12081 10044
rect 9585 10007 9643 10013
rect 12069 10013 12081 10016
rect 12115 10013 12127 10047
rect 12069 10007 12127 10013
rect 13265 10047 13323 10053
rect 13265 10013 13277 10047
rect 13311 10044 13323 10047
rect 15286 10044 15292 10056
rect 13311 10016 15292 10044
rect 13311 10013 13323 10016
rect 13265 10007 13323 10013
rect 15286 10004 15292 10016
rect 15344 10004 15350 10056
rect 17954 10044 17960 10056
rect 17915 10016 17960 10044
rect 17954 10004 17960 10016
rect 18012 10004 18018 10056
rect 18509 10047 18567 10053
rect 18509 10013 18521 10047
rect 18555 10044 18567 10047
rect 18782 10044 18788 10056
rect 18555 10016 18788 10044
rect 18555 10013 18567 10016
rect 18509 10007 18567 10013
rect 18782 10004 18788 10016
rect 18840 10004 18846 10056
rect 4488 9948 6224 9976
rect 8389 9979 8447 9985
rect 4488 9936 4494 9948
rect 8389 9945 8401 9979
rect 8435 9945 8447 9979
rect 8389 9939 8447 9945
rect 8481 9979 8539 9985
rect 8481 9945 8493 9979
rect 8527 9945 8539 9979
rect 8481 9939 8539 9945
rect 4982 9908 4988 9920
rect 2792 9880 3372 9908
rect 4943 9880 4988 9908
rect 4982 9868 4988 9880
rect 5040 9868 5046 9920
rect 5902 9908 5908 9920
rect 5863 9880 5908 9908
rect 5902 9868 5908 9880
rect 5960 9868 5966 9920
rect 8294 9868 8300 9920
rect 8352 9908 8358 9920
rect 8496 9908 8524 9939
rect 11238 9936 11244 9988
rect 11296 9976 11302 9988
rect 11885 9979 11943 9985
rect 11885 9976 11897 9979
rect 11296 9948 11897 9976
rect 11296 9936 11302 9948
rect 11885 9945 11897 9948
rect 11931 9945 11943 9979
rect 11885 9939 11943 9945
rect 15930 9936 15936 9988
rect 15988 9936 15994 9988
rect 8352 9880 8524 9908
rect 9033 9911 9091 9917
rect 8352 9868 8358 9880
rect 9033 9877 9045 9911
rect 9079 9908 9091 9911
rect 11514 9908 11520 9920
rect 9079 9880 11520 9908
rect 9079 9877 9091 9880
rect 9033 9871 9091 9877
rect 11514 9868 11520 9880
rect 11572 9868 11578 9920
rect 17770 9908 17776 9920
rect 17731 9880 17776 9908
rect 17770 9868 17776 9880
rect 17828 9868 17834 9920
rect 0 9818 18860 9840
rect 0 9766 4660 9818
rect 4712 9766 4724 9818
rect 4776 9766 4788 9818
rect 4840 9766 4852 9818
rect 4904 9766 4916 9818
rect 4968 9766 7760 9818
rect 7812 9766 7824 9818
rect 7876 9766 7888 9818
rect 7940 9766 7952 9818
rect 8004 9766 8016 9818
rect 8068 9766 10860 9818
rect 10912 9766 10924 9818
rect 10976 9766 10988 9818
rect 11040 9766 11052 9818
rect 11104 9766 11116 9818
rect 11168 9766 13960 9818
rect 14012 9766 14024 9818
rect 14076 9766 14088 9818
rect 14140 9766 14152 9818
rect 14204 9766 14216 9818
rect 14268 9766 17060 9818
rect 17112 9766 17124 9818
rect 17176 9766 17188 9818
rect 17240 9766 17252 9818
rect 17304 9766 17316 9818
rect 17368 9766 18860 9818
rect 0 9744 18860 9766
rect 566 9664 572 9716
rect 624 9704 630 9716
rect 1121 9707 1179 9713
rect 1121 9704 1133 9707
rect 624 9676 1133 9704
rect 624 9664 630 9676
rect 1121 9673 1133 9676
rect 1167 9673 1179 9707
rect 1121 9667 1179 9673
rect 2774 9664 2780 9716
rect 2832 9704 2838 9716
rect 4338 9704 4344 9716
rect 2832 9676 4344 9704
rect 2832 9664 2838 9676
rect 4338 9664 4344 9676
rect 4396 9664 4402 9716
rect 5810 9664 5816 9716
rect 5868 9704 5874 9716
rect 5905 9707 5963 9713
rect 5905 9704 5917 9707
rect 5868 9676 5917 9704
rect 5868 9664 5874 9676
rect 5905 9673 5917 9676
rect 5951 9673 5963 9707
rect 5905 9667 5963 9673
rect 6730 9664 6736 9716
rect 6788 9704 6794 9716
rect 12437 9707 12495 9713
rect 12437 9704 12449 9707
rect 6788 9676 12449 9704
rect 6788 9664 6794 9676
rect 12437 9673 12449 9676
rect 12483 9704 12495 9707
rect 13262 9704 13268 9716
rect 12483 9676 13268 9704
rect 12483 9673 12495 9676
rect 12437 9667 12495 9673
rect 13262 9664 13268 9676
rect 13320 9664 13326 9716
rect 2222 9636 2228 9648
rect 1412 9608 2228 9636
rect 1412 9577 1440 9608
rect 2222 9596 2228 9608
rect 2280 9596 2286 9648
rect 3234 9636 3240 9648
rect 2976 9608 3240 9636
rect 2976 9577 3004 9608
rect 3234 9596 3240 9608
rect 3292 9596 3298 9648
rect 4801 9639 4859 9645
rect 4801 9605 4813 9639
rect 4847 9636 4859 9639
rect 5626 9636 5632 9648
rect 4847 9608 5632 9636
rect 4847 9605 4859 9608
rect 4801 9599 4859 9605
rect 5626 9596 5632 9608
rect 5684 9636 5690 9648
rect 5997 9639 6055 9645
rect 5997 9636 6009 9639
rect 5684 9608 6009 9636
rect 5684 9596 5690 9608
rect 5997 9605 6009 9608
rect 6043 9605 6055 9639
rect 5997 9599 6055 9605
rect 8294 9596 8300 9648
rect 8352 9636 8358 9648
rect 9950 9636 9956 9648
rect 8352 9622 8786 9636
rect 8352 9608 8800 9622
rect 9911 9608 9956 9636
rect 8352 9596 8358 9608
rect 1397 9571 1455 9577
rect 1397 9537 1409 9571
rect 1443 9537 1455 9571
rect 1397 9531 1455 9537
rect 1489 9571 1547 9577
rect 1489 9537 1501 9571
rect 1535 9568 1547 9571
rect 1581 9571 1639 9577
rect 1581 9568 1593 9571
rect 1535 9540 1593 9568
rect 1535 9537 1547 9540
rect 1489 9531 1547 9537
rect 1581 9537 1593 9540
rect 1627 9537 1639 9571
rect 1581 9531 1639 9537
rect 1765 9571 1823 9577
rect 1765 9537 1777 9571
rect 1811 9537 1823 9571
rect 1765 9531 1823 9537
rect 2961 9571 3019 9577
rect 2961 9537 2973 9571
rect 3007 9537 3019 9571
rect 2961 9531 3019 9537
rect 3145 9571 3203 9577
rect 3145 9537 3157 9571
rect 3191 9568 3203 9571
rect 4614 9568 4620 9580
rect 3191 9540 4620 9568
rect 3191 9537 3203 9540
rect 3145 9531 3203 9537
rect 1121 9503 1179 9509
rect 1121 9469 1133 9503
rect 1167 9500 1179 9503
rect 1673 9503 1731 9509
rect 1673 9500 1685 9503
rect 1167 9472 1685 9500
rect 1167 9469 1179 9472
rect 1121 9463 1179 9469
rect 1673 9469 1685 9472
rect 1719 9469 1731 9503
rect 1780 9500 1808 9531
rect 4614 9528 4620 9540
rect 4672 9528 4678 9580
rect 4709 9571 4767 9577
rect 4709 9537 4721 9571
rect 4755 9568 4767 9571
rect 4755 9540 5580 9568
rect 4755 9537 4767 9540
rect 4709 9531 4767 9537
rect 4985 9503 5043 9509
rect 1780 9472 4384 9500
rect 1673 9463 1731 9469
rect 1305 9435 1363 9441
rect 1305 9401 1317 9435
rect 1351 9432 1363 9435
rect 1489 9435 1547 9441
rect 1489 9432 1501 9435
rect 1351 9404 1501 9432
rect 1351 9401 1363 9404
rect 1305 9395 1363 9401
rect 1489 9401 1501 9404
rect 1535 9432 1547 9435
rect 2958 9432 2964 9444
rect 1535 9404 2964 9432
rect 1535 9401 1547 9404
rect 1489 9395 1547 9401
rect 2958 9392 2964 9404
rect 3016 9432 3022 9444
rect 3234 9432 3240 9444
rect 3016 9404 3240 9432
rect 3016 9392 3022 9404
rect 3234 9392 3240 9404
rect 3292 9392 3298 9444
rect 3418 9392 3424 9444
rect 3476 9392 3482 9444
rect 4356 9441 4384 9472
rect 4985 9469 4997 9503
rect 5031 9500 5043 9503
rect 5442 9500 5448 9512
rect 5031 9472 5448 9500
rect 5031 9469 5043 9472
rect 4985 9463 5043 9469
rect 5442 9460 5448 9472
rect 5500 9460 5506 9512
rect 5552 9441 5580 9540
rect 5902 9528 5908 9580
rect 5960 9568 5966 9580
rect 6733 9571 6791 9577
rect 6733 9568 6745 9571
rect 5960 9540 6745 9568
rect 5960 9528 5966 9540
rect 6733 9537 6745 9540
rect 6779 9537 6791 9571
rect 6733 9531 6791 9537
rect 6181 9503 6239 9509
rect 6181 9469 6193 9503
rect 6227 9469 6239 9503
rect 6822 9500 6828 9512
rect 6783 9472 6828 9500
rect 6181 9463 6239 9469
rect 4341 9435 4399 9441
rect 4341 9401 4353 9435
rect 4387 9401 4399 9435
rect 4341 9395 4399 9401
rect 5537 9435 5595 9441
rect 5537 9401 5549 9435
rect 5583 9401 5595 9435
rect 6196 9432 6224 9463
rect 6822 9460 6828 9472
rect 6880 9460 6886 9512
rect 6917 9503 6975 9509
rect 6917 9469 6929 9503
rect 6963 9469 6975 9503
rect 8772 9500 8800 9608
rect 9950 9596 9956 9608
rect 10008 9596 10014 9648
rect 11330 9636 11336 9648
rect 10520 9608 11336 9636
rect 10229 9571 10287 9577
rect 10229 9537 10241 9571
rect 10275 9568 10287 9571
rect 10321 9571 10379 9577
rect 10321 9568 10333 9571
rect 10275 9540 10333 9568
rect 10275 9537 10287 9540
rect 10229 9531 10287 9537
rect 10321 9537 10333 9540
rect 10367 9537 10379 9571
rect 10321 9531 10379 9537
rect 10520 9500 10548 9608
rect 11330 9596 11336 9608
rect 11388 9596 11394 9648
rect 12526 9596 12532 9648
rect 12584 9636 12590 9648
rect 17681 9639 17739 9645
rect 12584 9622 13846 9636
rect 12584 9608 13860 9622
rect 12584 9596 12590 9608
rect 12158 9528 12164 9580
rect 12216 9568 12222 9580
rect 12805 9571 12863 9577
rect 12805 9568 12817 9571
rect 12216 9540 12817 9568
rect 12216 9528 12222 9540
rect 12805 9537 12817 9540
rect 12851 9537 12863 9571
rect 12805 9531 12863 9537
rect 8772 9472 10548 9500
rect 10597 9503 10655 9509
rect 6917 9463 6975 9469
rect 10597 9469 10609 9503
rect 10643 9500 10655 9503
rect 10870 9500 10876 9512
rect 10643 9472 10723 9500
rect 10783 9472 10876 9500
rect 10643 9469 10655 9472
rect 10597 9463 10655 9469
rect 6932 9432 6960 9463
rect 5537 9395 5595 9401
rect 5644 9404 6960 9432
rect 3053 9367 3111 9373
rect 3053 9333 3065 9367
rect 3099 9364 3111 9367
rect 3436 9364 3464 9392
rect 3099 9336 3464 9364
rect 3099 9333 3111 9336
rect 3053 9327 3111 9333
rect 4982 9324 4988 9376
rect 5040 9364 5046 9376
rect 5644 9364 5672 9404
rect 5040 9336 5672 9364
rect 5040 9324 5046 9336
rect 5902 9324 5908 9376
rect 5960 9364 5966 9376
rect 6365 9367 6423 9373
rect 6365 9364 6377 9367
rect 5960 9336 6377 9364
rect 5960 9324 5966 9336
rect 6365 9333 6377 9336
rect 6411 9333 6423 9367
rect 6365 9327 6423 9333
rect 8481 9367 8539 9373
rect 8481 9333 8493 9367
rect 8527 9364 8539 9367
rect 10226 9364 10232 9376
rect 8527 9336 10232 9364
rect 8527 9333 8539 9336
rect 8481 9327 8539 9333
rect 10226 9324 10232 9336
rect 10284 9324 10290 9376
rect 10413 9367 10471 9373
rect 10413 9333 10425 9367
rect 10459 9364 10471 9367
rect 10594 9364 10600 9376
rect 10459 9336 10600 9364
rect 10459 9333 10471 9336
rect 10413 9327 10471 9333
rect 10594 9324 10600 9336
rect 10652 9364 10658 9376
rect 10695 9364 10723 9472
rect 10870 9460 10876 9472
rect 10928 9500 10934 9512
rect 12526 9500 12532 9512
rect 10928 9472 11928 9500
rect 10928 9460 10934 9472
rect 10652 9336 10723 9364
rect 11900 9364 11928 9472
rect 11992 9472 12532 9500
rect 11992 9444 12020 9472
rect 12526 9460 12532 9472
rect 12584 9460 12590 9512
rect 12894 9500 12900 9512
rect 12855 9472 12900 9500
rect 12894 9460 12900 9472
rect 12952 9460 12958 9512
rect 12989 9503 13047 9509
rect 12989 9469 13001 9503
rect 13035 9469 13047 9503
rect 12989 9463 13047 9469
rect 13265 9503 13323 9509
rect 13265 9469 13277 9503
rect 13311 9500 13323 9503
rect 13538 9500 13544 9512
rect 13311 9472 13544 9500
rect 13311 9469 13323 9472
rect 13265 9463 13323 9469
rect 11974 9392 11980 9444
rect 12032 9392 12038 9444
rect 12066 9392 12072 9444
rect 12124 9432 12130 9444
rect 12345 9435 12403 9441
rect 12345 9432 12357 9435
rect 12124 9404 12357 9432
rect 12124 9392 12130 9404
rect 12345 9401 12357 9404
rect 12391 9432 12403 9435
rect 13004 9432 13032 9463
rect 13538 9460 13544 9472
rect 13596 9460 13602 9512
rect 13832 9500 13860 9608
rect 17681 9605 17693 9639
rect 17727 9636 17739 9639
rect 17770 9636 17776 9648
rect 17727 9608 17776 9636
rect 17727 9605 17739 9608
rect 17681 9599 17739 9605
rect 17770 9596 17776 9608
rect 17828 9596 17834 9648
rect 15930 9528 15936 9580
rect 15988 9568 15994 9580
rect 15988 9540 16606 9568
rect 15988 9528 15994 9540
rect 16500 9512 16528 9540
rect 14366 9500 14372 9512
rect 13832 9472 14372 9500
rect 14366 9460 14372 9472
rect 14424 9460 14430 9512
rect 15013 9503 15071 9509
rect 15013 9469 15025 9503
rect 15059 9500 15071 9503
rect 15289 9503 15347 9509
rect 15059 9472 15240 9500
rect 15059 9469 15071 9472
rect 15013 9463 15071 9469
rect 12391 9404 13032 9432
rect 15212 9432 15240 9472
rect 15289 9469 15301 9503
rect 15335 9500 15347 9503
rect 15838 9500 15844 9512
rect 15335 9472 15844 9500
rect 15335 9469 15347 9472
rect 15289 9463 15347 9469
rect 15838 9460 15844 9472
rect 15896 9460 15902 9512
rect 16482 9460 16488 9512
rect 16540 9460 16546 9512
rect 17954 9500 17960 9512
rect 17915 9472 17960 9500
rect 17954 9460 17960 9472
rect 18012 9460 18018 9512
rect 16209 9435 16267 9441
rect 16209 9432 16221 9435
rect 15212 9404 16221 9432
rect 12391 9401 12403 9404
rect 12345 9395 12403 9401
rect 16209 9401 16221 9404
rect 16255 9401 16267 9435
rect 16209 9395 16267 9401
rect 14458 9364 14464 9376
rect 11900 9336 14464 9364
rect 10652 9324 10658 9336
rect 14458 9324 14464 9336
rect 14516 9324 14522 9376
rect 0 9274 18860 9296
rect 0 9222 3110 9274
rect 3162 9222 3174 9274
rect 3226 9222 3238 9274
rect 3290 9222 3302 9274
rect 3354 9222 3366 9274
rect 3418 9222 6210 9274
rect 6262 9222 6274 9274
rect 6326 9222 6338 9274
rect 6390 9222 6402 9274
rect 6454 9222 6466 9274
rect 6518 9222 9310 9274
rect 9362 9222 9374 9274
rect 9426 9222 9438 9274
rect 9490 9222 9502 9274
rect 9554 9222 9566 9274
rect 9618 9222 12410 9274
rect 12462 9222 12474 9274
rect 12526 9222 12538 9274
rect 12590 9222 12602 9274
rect 12654 9222 12666 9274
rect 12718 9222 15510 9274
rect 15562 9222 15574 9274
rect 15626 9222 15638 9274
rect 15690 9222 15702 9274
rect 15754 9222 15766 9274
rect 15818 9222 18860 9274
rect 0 9200 18860 9222
rect 2041 9163 2099 9169
rect 2041 9129 2053 9163
rect 2087 9160 2099 9163
rect 2866 9160 2872 9172
rect 2087 9132 2872 9160
rect 2087 9129 2099 9132
rect 2041 9123 2099 9129
rect 2866 9120 2872 9132
rect 2924 9160 2930 9172
rect 4062 9160 4068 9172
rect 2924 9132 4068 9160
rect 2924 9120 2930 9132
rect 4062 9120 4068 9132
rect 4120 9120 4126 9172
rect 4614 9120 4620 9172
rect 4672 9160 4678 9172
rect 5537 9163 5595 9169
rect 5537 9160 5549 9163
rect 4672 9132 5549 9160
rect 4672 9120 4678 9132
rect 5537 9129 5549 9132
rect 5583 9129 5595 9163
rect 5537 9123 5595 9129
rect 9217 9163 9275 9169
rect 9217 9129 9229 9163
rect 9263 9160 9275 9163
rect 9585 9163 9643 9169
rect 9585 9160 9597 9163
rect 9263 9132 9597 9160
rect 9263 9129 9275 9132
rect 9217 9123 9275 9129
rect 9585 9129 9597 9132
rect 9631 9160 9643 9163
rect 10410 9160 10416 9172
rect 9631 9132 10416 9160
rect 9631 9129 9643 9132
rect 9585 9123 9643 9129
rect 10410 9120 10416 9132
rect 10468 9120 10474 9172
rect 10689 9163 10747 9169
rect 10689 9129 10701 9163
rect 10735 9160 10747 9163
rect 12158 9160 12164 9172
rect 10735 9132 12164 9160
rect 10735 9129 10747 9132
rect 10689 9123 10747 9129
rect 12158 9120 12164 9132
rect 12216 9120 12222 9172
rect 13354 9120 13360 9172
rect 13412 9160 13418 9172
rect 17954 9160 17960 9172
rect 13412 9132 17960 9160
rect 13412 9120 13418 9132
rect 17954 9120 17960 9132
rect 18012 9160 18018 9172
rect 18325 9163 18383 9169
rect 18325 9160 18337 9163
rect 18012 9132 18337 9160
rect 18012 9120 18018 9132
rect 18325 9129 18337 9132
rect 18371 9129 18383 9163
rect 18325 9123 18383 9129
rect 2225 9095 2283 9101
rect 2225 9092 2237 9095
rect 1596 9064 2237 9092
rect 290 9024 296 9036
rect 251 8996 296 9024
rect 290 8984 296 8996
rect 348 8984 354 9036
rect 569 9027 627 9033
rect 569 8993 581 9027
rect 615 9024 627 9027
rect 1596 9024 1624 9064
rect 2225 9061 2237 9064
rect 2271 9061 2283 9095
rect 2225 9055 2283 9061
rect 2317 9095 2375 9101
rect 2317 9061 2329 9095
rect 2363 9092 2375 9095
rect 10870 9092 10876 9104
rect 2363 9064 2774 9092
rect 2363 9061 2375 9064
rect 2317 9055 2375 9061
rect 615 8996 1624 9024
rect 2133 9027 2191 9033
rect 615 8993 627 8996
rect 569 8987 627 8993
rect 2133 8993 2145 9027
rect 2179 9024 2191 9027
rect 2498 9024 2504 9036
rect 2179 8996 2504 9024
rect 2179 8993 2191 8996
rect 2133 8987 2191 8993
rect 2498 8984 2504 8996
rect 2556 8984 2562 9036
rect 2746 9024 2774 9064
rect 10060 9064 10876 9092
rect 2958 9024 2964 9036
rect 2746 8996 2964 9024
rect 2958 8984 2964 8996
rect 3016 9024 3022 9036
rect 3145 9027 3203 9033
rect 3145 9024 3157 9027
rect 3016 8996 3157 9024
rect 3016 8984 3022 8996
rect 3145 8993 3157 8996
rect 3191 8993 3203 9027
rect 3145 8987 3203 8993
rect 4433 9027 4491 9033
rect 4433 8993 4445 9027
rect 4479 9024 4491 9027
rect 4982 9024 4988 9036
rect 4479 8996 4988 9024
rect 4479 8993 4491 8996
rect 4433 8987 4491 8993
rect 4982 8984 4988 8996
rect 5040 8984 5046 9036
rect 5534 8984 5540 9036
rect 5592 9024 5598 9036
rect 6086 9024 6092 9036
rect 5592 8996 6092 9024
rect 5592 8984 5598 8996
rect 6086 8984 6092 8996
rect 6144 8984 6150 9036
rect 6178 8984 6184 9036
rect 6236 9024 6242 9036
rect 6822 9024 6828 9036
rect 6236 8996 6828 9024
rect 6236 8984 6242 8996
rect 6822 8984 6828 8996
rect 6880 8984 6886 9036
rect 9674 9024 9680 9036
rect 9324 8996 9680 9024
rect 2409 8959 2467 8965
rect 2409 8925 2421 8959
rect 2455 8925 2467 8959
rect 2409 8919 2467 8925
rect 1854 8888 1860 8900
rect 1794 8860 1860 8888
rect 1854 8848 1860 8860
rect 1912 8848 1918 8900
rect 2424 8888 2452 8919
rect 2774 8916 2780 8968
rect 2832 8956 2838 8968
rect 2869 8959 2927 8965
rect 2869 8956 2881 8959
rect 2832 8928 2881 8956
rect 2832 8916 2838 8928
rect 2869 8925 2881 8928
rect 2915 8925 2927 8959
rect 2869 8919 2927 8925
rect 3602 8916 3608 8968
rect 3660 8956 3666 8968
rect 5552 8956 5580 8984
rect 5902 8956 5908 8968
rect 3660 8928 5580 8956
rect 5863 8928 5908 8956
rect 3660 8916 3666 8928
rect 5902 8916 5908 8928
rect 5960 8916 5966 8968
rect 5994 8916 6000 8968
rect 6052 8956 6058 8968
rect 8110 8965 8116 8968
rect 6641 8959 6699 8965
rect 6641 8956 6653 8959
rect 6052 8928 6653 8956
rect 6052 8916 6058 8928
rect 6641 8925 6653 8928
rect 6687 8956 6699 8959
rect 7837 8959 7895 8965
rect 7837 8956 7849 8959
rect 6687 8928 7849 8956
rect 6687 8925 6699 8928
rect 6641 8919 6699 8925
rect 7837 8925 7849 8928
rect 7883 8925 7895 8959
rect 8104 8956 8116 8965
rect 8023 8928 8116 8956
rect 7837 8919 7895 8925
rect 8104 8919 8116 8928
rect 8168 8956 8174 8968
rect 9324 8956 9352 8996
rect 9674 8984 9680 8996
rect 9732 8984 9738 9036
rect 10060 9033 10088 9064
rect 10870 9052 10876 9064
rect 10928 9052 10934 9104
rect 10045 9027 10103 9033
rect 10045 8993 10057 9027
rect 10091 8993 10103 9027
rect 10226 9024 10232 9036
rect 10187 8996 10232 9024
rect 10045 8987 10103 8993
rect 10226 8984 10232 8996
rect 10284 8984 10290 9036
rect 10410 8984 10416 9036
rect 10468 9024 10474 9036
rect 10781 9027 10839 9033
rect 10781 9024 10793 9027
rect 10468 8996 10793 9024
rect 10468 8984 10474 8996
rect 10781 8993 10793 8996
rect 10827 8993 10839 9027
rect 10781 8987 10839 8993
rect 11330 8984 11336 9036
rect 11388 9024 11394 9036
rect 11974 9024 11980 9036
rect 11388 8996 11980 9024
rect 11388 8984 11394 8996
rect 11974 8984 11980 8996
rect 12032 8984 12038 9036
rect 12158 8984 12164 9036
rect 12216 9024 12222 9036
rect 12805 9027 12863 9033
rect 12805 9024 12817 9027
rect 12216 8996 12817 9024
rect 12216 8984 12222 8996
rect 12805 8993 12817 8996
rect 12851 8993 12863 9027
rect 12805 8987 12863 8993
rect 13722 8984 13728 9036
rect 13780 9024 13786 9036
rect 15749 9027 15807 9033
rect 15749 9024 15761 9027
rect 13780 8996 15761 9024
rect 13780 8984 13786 8996
rect 15749 8993 15761 8996
rect 15795 9024 15807 9027
rect 16666 9024 16672 9036
rect 15795 8996 16672 9024
rect 15795 8993 15807 8996
rect 15749 8987 15807 8993
rect 16666 8984 16672 8996
rect 16724 8984 16730 9036
rect 8168 8928 9352 8956
rect 9401 8959 9459 8965
rect 8110 8916 8116 8919
rect 8168 8916 8174 8928
rect 9401 8925 9413 8959
rect 9447 8956 9459 8959
rect 10321 8959 10379 8965
rect 9447 8928 10272 8956
rect 9447 8925 9459 8928
rect 9401 8919 9459 8925
rect 4157 8891 4215 8897
rect 4157 8888 4169 8891
rect 2424 8860 4169 8888
rect 2314 8780 2320 8832
rect 2372 8820 2378 8832
rect 2424 8820 2452 8860
rect 4157 8857 4169 8860
rect 4203 8857 4215 8891
rect 4157 8851 4215 8857
rect 5442 8848 5448 8900
rect 5500 8888 5506 8900
rect 6914 8888 6920 8900
rect 5500 8860 6920 8888
rect 5500 8848 5506 8860
rect 6914 8848 6920 8860
rect 6972 8848 6978 8900
rect 2372 8792 2452 8820
rect 2372 8780 2378 8792
rect 3234 8780 3240 8832
rect 3292 8820 3298 8832
rect 3789 8823 3847 8829
rect 3789 8820 3801 8823
rect 3292 8792 3801 8820
rect 3292 8780 3298 8792
rect 3789 8789 3801 8792
rect 3835 8789 3847 8823
rect 4246 8820 4252 8832
rect 4207 8792 4252 8820
rect 3789 8783 3847 8789
rect 4246 8780 4252 8792
rect 4304 8780 4310 8832
rect 5997 8823 6055 8829
rect 5997 8789 6009 8823
rect 6043 8820 6055 8823
rect 6178 8820 6184 8832
rect 6043 8792 6184 8820
rect 6043 8789 6055 8792
rect 5997 8783 6055 8789
rect 6178 8780 6184 8792
rect 6236 8780 6242 8832
rect 6362 8780 6368 8832
rect 6420 8820 6426 8832
rect 6549 8823 6607 8829
rect 6549 8820 6561 8823
rect 6420 8792 6561 8820
rect 6420 8780 6426 8792
rect 6549 8789 6561 8792
rect 6595 8789 6607 8823
rect 6549 8783 6607 8789
rect 6822 8780 6828 8832
rect 6880 8820 6886 8832
rect 9416 8820 9444 8919
rect 10244 8900 10272 8928
rect 10321 8925 10333 8959
rect 10367 8956 10379 8959
rect 11238 8956 11244 8968
rect 10367 8928 11244 8956
rect 10367 8925 10379 8928
rect 10321 8919 10379 8925
rect 11238 8916 11244 8928
rect 11296 8916 11302 8968
rect 11348 8956 11376 8984
rect 13354 8956 13360 8968
rect 11348 8928 11454 8956
rect 13315 8928 13360 8956
rect 13354 8916 13360 8928
rect 13412 8916 13418 8968
rect 13538 8956 13544 8968
rect 13499 8928 13544 8956
rect 13538 8916 13544 8928
rect 13596 8916 13602 8968
rect 15286 8916 15292 8968
rect 15344 8956 15350 8968
rect 15381 8959 15439 8965
rect 15381 8956 15393 8959
rect 15344 8928 15393 8956
rect 15344 8916 15350 8928
rect 15381 8925 15393 8928
rect 15427 8925 15439 8959
rect 15381 8919 15439 8925
rect 15838 8916 15844 8968
rect 15896 8956 15902 8968
rect 15896 8928 15941 8956
rect 15896 8916 15902 8928
rect 16114 8916 16120 8968
rect 16172 8956 16178 8968
rect 16209 8959 16267 8965
rect 16209 8956 16221 8959
rect 16172 8928 16221 8956
rect 16172 8916 16178 8928
rect 16209 8925 16221 8928
rect 16255 8925 16267 8959
rect 18141 8959 18199 8965
rect 18141 8956 18153 8959
rect 16209 8919 16267 8925
rect 17972 8928 18153 8956
rect 10226 8848 10232 8900
rect 10284 8888 10290 8900
rect 10284 8860 10548 8888
rect 10284 8848 10290 8860
rect 9858 8820 9864 8832
rect 6880 8792 9444 8820
rect 9819 8792 9864 8820
rect 6880 8780 6886 8792
rect 9858 8780 9864 8792
rect 9916 8780 9922 8832
rect 10520 8820 10548 8860
rect 12434 8848 12440 8900
rect 12492 8888 12498 8900
rect 12529 8891 12587 8897
rect 12529 8888 12541 8891
rect 12492 8860 12541 8888
rect 12492 8848 12498 8860
rect 12529 8857 12541 8860
rect 12575 8857 12587 8891
rect 12529 8851 12587 8857
rect 13280 8860 14320 8888
rect 13280 8820 13308 8860
rect 13446 8820 13452 8832
rect 10520 8792 13308 8820
rect 13407 8792 13452 8820
rect 13446 8780 13452 8792
rect 13504 8780 13510 8832
rect 13814 8780 13820 8832
rect 13872 8820 13878 8832
rect 13955 8823 14013 8829
rect 13955 8820 13967 8823
rect 13872 8792 13967 8820
rect 13872 8780 13878 8792
rect 13955 8789 13967 8792
rect 14001 8789 14013 8823
rect 14292 8820 14320 8860
rect 14366 8848 14372 8900
rect 14424 8848 14430 8900
rect 16482 8848 16488 8900
rect 16540 8888 16546 8900
rect 16540 8860 16606 8888
rect 16540 8848 16546 8860
rect 17972 8829 18000 8928
rect 18141 8925 18153 8928
rect 18187 8925 18199 8959
rect 18141 8919 18199 8925
rect 17957 8823 18015 8829
rect 17957 8820 17969 8823
rect 14292 8792 17969 8820
rect 13955 8783 14013 8789
rect 17957 8789 17969 8792
rect 18003 8789 18015 8823
rect 17957 8783 18015 8789
rect 0 8730 18860 8752
rect 0 8678 4660 8730
rect 4712 8678 4724 8730
rect 4776 8678 4788 8730
rect 4840 8678 4852 8730
rect 4904 8678 4916 8730
rect 4968 8678 7760 8730
rect 7812 8678 7824 8730
rect 7876 8678 7888 8730
rect 7940 8678 7952 8730
rect 8004 8678 8016 8730
rect 8068 8678 10860 8730
rect 10912 8678 10924 8730
rect 10976 8678 10988 8730
rect 11040 8678 11052 8730
rect 11104 8678 11116 8730
rect 11168 8678 13960 8730
rect 14012 8678 14024 8730
rect 14076 8678 14088 8730
rect 14140 8678 14152 8730
rect 14204 8678 14216 8730
rect 14268 8678 17060 8730
rect 17112 8678 17124 8730
rect 17176 8678 17188 8730
rect 17240 8678 17252 8730
rect 17304 8678 17316 8730
rect 17368 8678 18860 8730
rect 0 8656 18860 8678
rect 2314 8616 2320 8628
rect 2275 8588 2320 8616
rect 2314 8576 2320 8588
rect 2372 8576 2378 8628
rect 2498 8616 2504 8628
rect 2459 8588 2504 8616
rect 2498 8576 2504 8588
rect 2556 8576 2562 8628
rect 3234 8616 3240 8628
rect 3195 8588 3240 8616
rect 3234 8576 3240 8588
rect 3292 8576 3298 8628
rect 3329 8619 3387 8625
rect 3329 8585 3341 8619
rect 3375 8616 3387 8619
rect 4246 8616 4252 8628
rect 3375 8588 4252 8616
rect 3375 8585 3387 8588
rect 3329 8579 3387 8585
rect 4246 8576 4252 8588
rect 4304 8576 4310 8628
rect 4617 8619 4675 8625
rect 4617 8585 4629 8619
rect 4663 8616 4675 8619
rect 18506 8616 18512 8628
rect 4663 8588 5764 8616
rect 4663 8585 4675 8588
rect 4617 8579 4675 8585
rect 2774 8548 2780 8560
rect 2516 8520 2780 8548
rect 2516 8489 2544 8520
rect 2774 8508 2780 8520
rect 2832 8548 2838 8560
rect 5442 8548 5448 8560
rect 2832 8520 2925 8548
rect 4816 8520 5448 8548
rect 2832 8508 2838 8520
rect 2409 8483 2467 8489
rect 2409 8449 2421 8483
rect 2455 8449 2467 8483
rect 2409 8443 2467 8449
rect 2501 8483 2559 8489
rect 2501 8449 2513 8483
rect 2547 8449 2559 8483
rect 2501 8443 2559 8449
rect 2685 8483 2743 8489
rect 2685 8449 2697 8483
rect 2731 8480 2743 8483
rect 2958 8480 2964 8492
rect 2731 8452 2964 8480
rect 2731 8449 2743 8452
rect 2685 8443 2743 8449
rect 2424 8412 2452 8443
rect 2958 8440 2964 8452
rect 3016 8440 3022 8492
rect 3694 8480 3700 8492
rect 3655 8452 3700 8480
rect 3694 8440 3700 8452
rect 3752 8440 3758 8492
rect 3881 8483 3939 8489
rect 3881 8449 3893 8483
rect 3927 8449 3939 8483
rect 4338 8480 4344 8492
rect 4299 8452 4344 8480
rect 3881 8443 3939 8449
rect 2866 8412 2872 8424
rect 2424 8384 2872 8412
rect 2866 8372 2872 8384
rect 2924 8372 2930 8424
rect 3513 8415 3571 8421
rect 3513 8381 3525 8415
rect 3559 8412 3571 8415
rect 3602 8412 3608 8424
rect 3559 8384 3608 8412
rect 3559 8381 3571 8384
rect 3513 8375 3571 8381
rect 3602 8372 3608 8384
rect 3660 8372 3666 8424
rect 3896 8412 3924 8443
rect 4338 8440 4344 8452
rect 4396 8440 4402 8492
rect 4522 8480 4528 8492
rect 4483 8452 4528 8480
rect 4522 8440 4528 8452
rect 4580 8440 4586 8492
rect 4816 8489 4844 8520
rect 5442 8508 5448 8520
rect 5500 8508 5506 8560
rect 5736 8557 5764 8588
rect 6196 8588 8708 8616
rect 6196 8557 6224 8588
rect 5721 8551 5779 8557
rect 4801 8483 4859 8489
rect 4801 8449 4813 8483
rect 4847 8449 4859 8483
rect 4801 8443 4859 8449
rect 4982 8440 4988 8492
rect 5040 8480 5046 8492
rect 5261 8483 5319 8489
rect 5261 8480 5273 8483
rect 5040 8452 5273 8480
rect 5040 8440 5046 8452
rect 5261 8449 5273 8452
rect 5307 8449 5319 8483
rect 5534 8474 5540 8526
rect 5592 8474 5598 8526
rect 5721 8517 5733 8551
rect 5767 8517 5779 8551
rect 5721 8511 5779 8517
rect 6181 8551 6239 8557
rect 6181 8517 6193 8551
rect 6227 8517 6239 8551
rect 8294 8548 8300 8560
rect 7774 8520 8300 8548
rect 6181 8511 6239 8517
rect 8294 8508 8300 8520
rect 8352 8508 8358 8560
rect 5629 8483 5687 8489
rect 5535 8471 5547 8474
rect 5581 8471 5593 8474
rect 5535 8465 5593 8471
rect 5261 8443 5319 8449
rect 5629 8449 5641 8483
rect 5675 8449 5687 8483
rect 5902 8480 5908 8492
rect 5863 8452 5908 8480
rect 5629 8443 5687 8449
rect 4540 8412 4568 8440
rect 3896 8384 4568 8412
rect 2777 8347 2835 8353
rect 2777 8313 2789 8347
rect 2823 8344 2835 8347
rect 3789 8347 3847 8353
rect 3789 8344 3801 8347
rect 2823 8316 3801 8344
rect 2823 8313 2835 8316
rect 2777 8307 2835 8313
rect 3789 8313 3801 8316
rect 3835 8313 3847 8347
rect 3789 8307 3847 8313
rect 5353 8347 5411 8353
rect 5353 8313 5365 8347
rect 5399 8344 5411 8347
rect 5644 8344 5672 8443
rect 5902 8440 5908 8452
rect 5960 8440 5966 8492
rect 6362 8480 6368 8492
rect 6323 8452 6368 8480
rect 6362 8440 6368 8452
rect 6420 8440 6426 8492
rect 8680 8489 8708 8588
rect 10244 8588 18512 8616
rect 10244 8557 10272 8588
rect 18506 8576 18512 8588
rect 18564 8576 18570 8628
rect 10229 8551 10287 8557
rect 10229 8517 10241 8551
rect 10275 8517 10287 8551
rect 11977 8551 12035 8557
rect 11977 8548 11989 8551
rect 10229 8511 10287 8517
rect 10336 8520 11989 8548
rect 8665 8483 8723 8489
rect 8665 8449 8677 8483
rect 8711 8480 8723 8483
rect 10336 8480 10364 8520
rect 11977 8517 11989 8520
rect 12023 8517 12035 8551
rect 11977 8511 12035 8517
rect 12158 8508 12164 8560
rect 12216 8548 12222 8560
rect 13541 8551 13599 8557
rect 13541 8548 13553 8551
rect 12216 8520 13553 8548
rect 12216 8508 12222 8520
rect 13541 8517 13553 8520
rect 13587 8548 13599 8551
rect 13722 8548 13728 8560
rect 13587 8520 13728 8548
rect 13587 8517 13599 8520
rect 13541 8511 13599 8517
rect 13722 8508 13728 8520
rect 13780 8508 13786 8560
rect 14461 8551 14519 8557
rect 14461 8517 14473 8551
rect 14507 8548 14519 8551
rect 15286 8548 15292 8560
rect 14507 8520 15292 8548
rect 14507 8517 14519 8520
rect 14461 8511 14519 8517
rect 15286 8508 15292 8520
rect 15344 8508 15350 8560
rect 15795 8551 15853 8557
rect 15795 8517 15807 8551
rect 15841 8548 15853 8551
rect 16022 8548 16028 8560
rect 15841 8520 16028 8548
rect 15841 8517 15853 8520
rect 15795 8511 15853 8517
rect 16022 8508 16028 8520
rect 16080 8508 16086 8560
rect 16298 8508 16304 8560
rect 16356 8508 16362 8560
rect 10686 8489 10692 8492
rect 8711 8452 10364 8480
rect 10413 8483 10471 8489
rect 8711 8449 8723 8452
rect 8665 8443 8723 8449
rect 10413 8449 10425 8483
rect 10459 8449 10471 8483
rect 10680 8480 10692 8489
rect 10647 8452 10692 8480
rect 10413 8443 10471 8449
rect 10680 8443 10692 8452
rect 6733 8415 6791 8421
rect 6733 8412 6745 8415
rect 5828 8384 6745 8412
rect 5828 8353 5856 8384
rect 6733 8381 6745 8384
rect 6779 8381 6791 8415
rect 6733 8375 6791 8381
rect 5399 8316 5672 8344
rect 5813 8347 5871 8353
rect 5399 8313 5411 8316
rect 5353 8307 5411 8313
rect 5813 8313 5825 8347
rect 5859 8313 5871 8347
rect 5994 8344 6000 8356
rect 5955 8316 6000 8344
rect 5813 8307 5871 8313
rect 5994 8304 6000 8316
rect 6052 8304 6058 8356
rect 2869 8279 2927 8285
rect 2869 8245 2881 8279
rect 2915 8276 2927 8279
rect 2958 8276 2964 8288
rect 2915 8248 2964 8276
rect 2915 8245 2927 8248
rect 2869 8239 2927 8245
rect 2958 8236 2964 8248
rect 3016 8236 3022 8288
rect 4614 8236 4620 8288
rect 4672 8276 4678 8288
rect 5626 8276 5632 8288
rect 4672 8248 5632 8276
rect 4672 8236 4678 8248
rect 5626 8236 5632 8248
rect 5684 8236 5690 8288
rect 8018 8236 8024 8288
rect 8076 8276 8082 8288
rect 8159 8279 8217 8285
rect 8159 8276 8171 8279
rect 8076 8248 8171 8276
rect 8076 8236 8082 8248
rect 8159 8245 8171 8248
rect 8205 8245 8217 8279
rect 8159 8239 8217 8245
rect 9858 8236 9864 8288
rect 9916 8276 9922 8288
rect 10428 8276 10456 8443
rect 10686 8440 10692 8443
rect 10744 8440 10750 8492
rect 13633 8483 13691 8489
rect 13633 8449 13645 8483
rect 13679 8449 13691 8483
rect 14366 8480 14372 8492
rect 14327 8452 14372 8480
rect 13633 8443 13691 8449
rect 13446 8412 13452 8424
rect 13407 8384 13452 8412
rect 13446 8372 13452 8384
rect 13504 8372 13510 8424
rect 13648 8412 13676 8443
rect 14366 8440 14372 8452
rect 14424 8440 14430 8492
rect 14550 8480 14556 8492
rect 14511 8452 14556 8480
rect 14550 8440 14556 8452
rect 14608 8440 14614 8492
rect 14829 8483 14887 8489
rect 14829 8449 14841 8483
rect 14875 8449 14887 8483
rect 17494 8480 17500 8492
rect 14829 8443 14887 8449
rect 17144 8452 17500 8480
rect 13814 8412 13820 8424
rect 13648 8384 13820 8412
rect 13814 8372 13820 8384
rect 13872 8412 13878 8424
rect 14844 8412 14872 8443
rect 13872 8384 14872 8412
rect 13872 8372 13878 8384
rect 15838 8372 15844 8424
rect 15896 8412 15902 8424
rect 17144 8412 17172 8452
rect 17494 8440 17500 8452
rect 17552 8480 17558 8492
rect 17589 8483 17647 8489
rect 17589 8480 17601 8483
rect 17552 8452 17601 8480
rect 17552 8440 17558 8452
rect 17589 8449 17601 8452
rect 17635 8480 17647 8483
rect 17862 8480 17868 8492
rect 17635 8452 17868 8480
rect 17635 8449 17647 8452
rect 17589 8443 17647 8449
rect 17862 8440 17868 8452
rect 17920 8440 17926 8492
rect 18506 8480 18512 8492
rect 18467 8452 18512 8480
rect 18506 8440 18512 8452
rect 18564 8440 18570 8492
rect 15896 8384 17172 8412
rect 17221 8415 17279 8421
rect 15896 8372 15902 8384
rect 17221 8381 17233 8415
rect 17267 8412 17279 8415
rect 17267 8384 18368 8412
rect 17267 8381 17279 8384
rect 17221 8375 17279 8381
rect 12158 8344 12164 8356
rect 11348 8316 12164 8344
rect 11348 8288 11376 8316
rect 12158 8304 12164 8316
rect 12216 8304 12222 8356
rect 18340 8353 18368 8384
rect 18325 8347 18383 8353
rect 18325 8313 18337 8347
rect 18371 8313 18383 8347
rect 18325 8307 18383 8313
rect 11330 8276 11336 8288
rect 9916 8248 11336 8276
rect 9916 8236 9922 8248
rect 11330 8236 11336 8248
rect 11388 8236 11394 8288
rect 11422 8236 11428 8288
rect 11480 8276 11486 8288
rect 11793 8279 11851 8285
rect 11793 8276 11805 8279
rect 11480 8248 11805 8276
rect 11480 8236 11486 8248
rect 11793 8245 11805 8248
rect 11839 8245 11851 8279
rect 11793 8239 11851 8245
rect 13814 8236 13820 8288
rect 13872 8276 13878 8288
rect 14001 8279 14059 8285
rect 14001 8276 14013 8279
rect 13872 8248 14013 8276
rect 13872 8236 13878 8248
rect 14001 8245 14013 8248
rect 14047 8245 14059 8279
rect 14918 8276 14924 8288
rect 14879 8248 14924 8276
rect 14001 8239 14059 8245
rect 14918 8236 14924 8248
rect 14976 8236 14982 8288
rect 0 8186 18860 8208
rect 0 8134 3110 8186
rect 3162 8134 3174 8186
rect 3226 8134 3238 8186
rect 3290 8134 3302 8186
rect 3354 8134 3366 8186
rect 3418 8134 6210 8186
rect 6262 8134 6274 8186
rect 6326 8134 6338 8186
rect 6390 8134 6402 8186
rect 6454 8134 6466 8186
rect 6518 8134 9310 8186
rect 9362 8134 9374 8186
rect 9426 8134 9438 8186
rect 9490 8134 9502 8186
rect 9554 8134 9566 8186
rect 9618 8134 12410 8186
rect 12462 8134 12474 8186
rect 12526 8134 12538 8186
rect 12590 8134 12602 8186
rect 12654 8134 12666 8186
rect 12718 8134 15510 8186
rect 15562 8134 15574 8186
rect 15626 8134 15638 8186
rect 15690 8134 15702 8186
rect 15754 8134 15766 8186
rect 15818 8134 18860 8186
rect 0 8112 18860 8134
rect 4522 8072 4528 8084
rect 4483 8044 4528 8072
rect 4522 8032 4528 8044
rect 4580 8032 4586 8084
rect 4614 8032 4620 8084
rect 4672 8072 4678 8084
rect 5534 8072 5540 8084
rect 4672 8044 4717 8072
rect 5495 8044 5540 8072
rect 4672 8032 4678 8044
rect 5534 8032 5540 8044
rect 5592 8032 5598 8084
rect 6914 8032 6920 8084
rect 6972 8072 6978 8084
rect 7929 8075 7987 8081
rect 7929 8072 7941 8075
rect 6972 8044 7941 8072
rect 6972 8032 6978 8044
rect 7929 8041 7941 8044
rect 7975 8041 7987 8075
rect 7929 8035 7987 8041
rect 8297 8075 8355 8081
rect 8297 8041 8309 8075
rect 8343 8072 8355 8075
rect 8938 8072 8944 8084
rect 8343 8044 8944 8072
rect 8343 8041 8355 8044
rect 8297 8035 8355 8041
rect 8938 8032 8944 8044
rect 8996 8032 9002 8084
rect 10134 8072 10140 8084
rect 10095 8044 10140 8072
rect 10134 8032 10140 8044
rect 10192 8032 10198 8084
rect 10321 8075 10379 8081
rect 10321 8041 10333 8075
rect 10367 8072 10379 8075
rect 10502 8072 10508 8084
rect 10367 8044 10508 8072
rect 10367 8041 10379 8044
rect 10321 8035 10379 8041
rect 10502 8032 10508 8044
rect 10560 8032 10566 8084
rect 10686 8032 10692 8084
rect 10744 8032 10750 8084
rect 10778 8032 10784 8084
rect 10836 8072 10842 8084
rect 11609 8075 11667 8081
rect 11609 8072 11621 8075
rect 10836 8044 11621 8072
rect 10836 8032 10842 8044
rect 11609 8041 11621 8044
rect 11655 8041 11667 8075
rect 11609 8035 11667 8041
rect 12250 8032 12256 8084
rect 12308 8072 12314 8084
rect 14366 8072 14372 8084
rect 12308 8044 13308 8072
rect 14327 8044 14372 8072
rect 12308 8032 12314 8044
rect 6822 8004 6828 8016
rect 4816 7976 6828 8004
rect 290 7936 296 7948
rect 251 7908 296 7936
rect 290 7896 296 7908
rect 348 7896 354 7948
rect 3329 7939 3387 7945
rect 3329 7905 3341 7939
rect 3375 7936 3387 7939
rect 4341 7939 4399 7945
rect 4341 7936 4353 7939
rect 3375 7908 4353 7936
rect 3375 7905 3387 7908
rect 3329 7899 3387 7905
rect 4341 7905 4353 7908
rect 4387 7905 4399 7939
rect 4816 7936 4844 7976
rect 6822 7964 6828 7976
rect 6880 7964 6886 8016
rect 9766 8004 9772 8016
rect 9727 7976 9772 8004
rect 9766 7964 9772 7976
rect 9824 7964 9830 8016
rect 10704 8004 10732 8032
rect 9968 7976 10732 8004
rect 10873 8007 10931 8013
rect 4341 7899 4399 7905
rect 4724 7908 4844 7936
rect 4893 7939 4951 7945
rect 2869 7871 2927 7877
rect 2869 7868 2881 7871
rect 2056 7840 2881 7868
rect 566 7800 572 7812
rect 527 7772 572 7800
rect 566 7760 572 7772
rect 624 7760 630 7812
rect 1854 7800 1860 7812
rect 1794 7772 1860 7800
rect 1854 7760 1860 7772
rect 1912 7760 1918 7812
rect 2056 7744 2084 7840
rect 2869 7837 2881 7840
rect 2915 7868 2927 7871
rect 3237 7871 3295 7877
rect 3237 7868 3249 7871
rect 2915 7840 3249 7868
rect 2915 7837 2927 7840
rect 2869 7831 2927 7837
rect 3237 7837 3249 7840
rect 3283 7837 3295 7871
rect 3237 7831 3295 7837
rect 3421 7871 3479 7877
rect 3421 7837 3433 7871
rect 3467 7868 3479 7871
rect 3510 7868 3516 7880
rect 3467 7840 3516 7868
rect 3467 7837 3479 7840
rect 3421 7831 3479 7837
rect 3510 7828 3516 7840
rect 3568 7828 3574 7880
rect 3602 7828 3608 7880
rect 3660 7868 3666 7880
rect 4062 7868 4068 7880
rect 3660 7840 3705 7868
rect 4023 7840 4068 7868
rect 3660 7828 3666 7840
rect 4062 7828 4068 7840
rect 4120 7828 4126 7880
rect 4246 7828 4252 7880
rect 4304 7868 4310 7880
rect 4724 7877 4752 7908
rect 4893 7905 4905 7939
rect 4939 7936 4951 7939
rect 5077 7939 5135 7945
rect 5077 7936 5089 7939
rect 4939 7908 5089 7936
rect 4939 7905 4951 7908
rect 4893 7899 4951 7905
rect 5077 7905 5089 7908
rect 5123 7936 5135 7939
rect 5718 7936 5724 7948
rect 5123 7908 5724 7936
rect 5123 7905 5135 7908
rect 5077 7899 5135 7905
rect 5718 7896 5724 7908
rect 5776 7896 5782 7948
rect 9677 7939 9735 7945
rect 9677 7905 9689 7939
rect 9723 7936 9735 7939
rect 9858 7936 9864 7948
rect 9723 7908 9864 7936
rect 9723 7905 9735 7908
rect 9677 7899 9735 7905
rect 9858 7896 9864 7908
rect 9916 7896 9922 7948
rect 4433 7871 4491 7877
rect 4433 7868 4445 7871
rect 4304 7840 4445 7868
rect 4304 7828 4310 7840
rect 4433 7837 4445 7840
rect 4479 7837 4491 7871
rect 4433 7831 4491 7837
rect 4709 7871 4767 7877
rect 4709 7837 4721 7871
rect 4755 7837 4767 7871
rect 4709 7831 4767 7837
rect 4801 7871 4859 7877
rect 4801 7837 4813 7871
rect 4847 7837 4859 7871
rect 4801 7831 4859 7837
rect 4985 7871 5043 7877
rect 4985 7837 4997 7871
rect 5031 7868 5043 7871
rect 8018 7868 8024 7880
rect 5031 7840 6224 7868
rect 7931 7840 8024 7868
rect 5031 7837 5043 7840
rect 4985 7831 5043 7837
rect 2406 7760 2412 7812
rect 2464 7800 2470 7812
rect 2464 7772 4016 7800
rect 2464 7760 2470 7772
rect 2038 7732 2044 7744
rect 1999 7704 2044 7732
rect 2038 7692 2044 7704
rect 2096 7692 2102 7744
rect 2498 7692 2504 7744
rect 2556 7732 2562 7744
rect 2777 7735 2835 7741
rect 2777 7732 2789 7735
rect 2556 7704 2789 7732
rect 2556 7692 2562 7704
rect 2777 7701 2789 7704
rect 2823 7701 2835 7735
rect 3694 7732 3700 7744
rect 3655 7704 3700 7732
rect 2777 7695 2835 7701
rect 3694 7692 3700 7704
rect 3752 7692 3758 7744
rect 3878 7732 3884 7744
rect 3839 7704 3884 7732
rect 3878 7692 3884 7704
rect 3936 7692 3942 7744
rect 3988 7732 4016 7772
rect 4816 7732 4844 7831
rect 6196 7812 6224 7840
rect 8018 7828 8024 7840
rect 8076 7828 8082 7880
rect 9582 7828 9588 7880
rect 9640 7868 9646 7880
rect 9968 7877 9996 7976
rect 10873 7973 10885 8007
rect 10919 7973 10931 8007
rect 10873 7967 10931 7973
rect 10226 7936 10232 7948
rect 10187 7908 10232 7936
rect 10226 7896 10232 7908
rect 10284 7896 10290 7948
rect 10689 7939 10747 7945
rect 10689 7905 10701 7939
rect 10735 7905 10747 7939
rect 10689 7899 10747 7905
rect 10781 7939 10839 7945
rect 10781 7905 10793 7939
rect 10827 7936 10839 7939
rect 10890 7936 10918 7967
rect 11422 7964 11428 8016
rect 11480 8004 11486 8016
rect 13280 8013 13308 8044
rect 14366 8032 14372 8044
rect 14424 8032 14430 8084
rect 14550 8032 14556 8084
rect 14608 8072 14614 8084
rect 15013 8075 15071 8081
rect 15013 8072 15025 8075
rect 14608 8044 15025 8072
rect 14608 8032 14614 8044
rect 15013 8041 15025 8044
rect 15059 8041 15071 8075
rect 15013 8035 15071 8041
rect 12713 8007 12771 8013
rect 11480 7976 11525 8004
rect 11480 7964 11486 7976
rect 12713 7973 12725 8007
rect 12759 7973 12771 8007
rect 12713 7967 12771 7973
rect 13265 8007 13323 8013
rect 13265 7973 13277 8007
rect 13311 7973 13323 8007
rect 13265 7967 13323 7973
rect 10827 7908 10918 7936
rect 10827 7905 10839 7908
rect 10781 7899 10839 7905
rect 9953 7871 10011 7877
rect 9953 7868 9965 7871
rect 9640 7840 9965 7868
rect 9640 7828 9646 7840
rect 9953 7837 9965 7840
rect 9999 7837 10011 7871
rect 10502 7868 10508 7880
rect 10463 7840 10508 7868
rect 9953 7831 10011 7837
rect 10502 7828 10508 7840
rect 10560 7828 10566 7880
rect 5810 7800 5816 7812
rect 5771 7772 5816 7800
rect 5810 7760 5816 7772
rect 5868 7760 5874 7812
rect 6178 7800 6184 7812
rect 6139 7772 6184 7800
rect 6178 7760 6184 7772
rect 6236 7760 6242 7812
rect 6365 7803 6423 7809
rect 6365 7769 6377 7803
rect 6411 7800 6423 7803
rect 6546 7800 6552 7812
rect 6411 7772 6552 7800
rect 6411 7769 6423 7772
rect 6365 7763 6423 7769
rect 6546 7760 6552 7772
rect 6604 7760 6610 7812
rect 5902 7732 5908 7744
rect 3988 7704 4844 7732
rect 5815 7704 5908 7732
rect 5902 7692 5908 7704
rect 5960 7732 5966 7744
rect 6730 7732 6736 7744
rect 5960 7704 6736 7732
rect 5960 7692 5966 7704
rect 6730 7692 6736 7704
rect 6788 7692 6794 7744
rect 8036 7732 8064 7828
rect 9030 7760 9036 7812
rect 9088 7800 9094 7812
rect 9432 7803 9490 7809
rect 9432 7800 9444 7803
rect 9088 7772 9444 7800
rect 9088 7760 9094 7772
rect 9432 7769 9444 7772
rect 9478 7800 9490 7803
rect 10134 7800 10140 7812
rect 9478 7772 10140 7800
rect 9478 7769 9490 7772
rect 9432 7763 9490 7769
rect 10134 7760 10140 7772
rect 10192 7760 10198 7812
rect 10704 7800 10732 7899
rect 11238 7896 11244 7948
rect 11296 7936 11302 7948
rect 12253 7939 12311 7945
rect 12253 7936 12265 7939
rect 11296 7908 11341 7936
rect 11440 7908 12265 7936
rect 11296 7896 11302 7908
rect 10870 7868 10876 7880
rect 10831 7840 10876 7868
rect 10870 7828 10876 7840
rect 10928 7828 10934 7880
rect 10962 7828 10968 7880
rect 11020 7868 11026 7880
rect 11020 7840 11065 7868
rect 11020 7828 11026 7840
rect 11146 7828 11152 7880
rect 11204 7868 11210 7880
rect 11204 7840 11249 7868
rect 11204 7828 11210 7840
rect 11241 7803 11299 7809
rect 11241 7800 11253 7803
rect 10704 7772 11253 7800
rect 11241 7769 11253 7772
rect 11287 7769 11299 7803
rect 11241 7763 11299 7769
rect 11440 7732 11468 7908
rect 12253 7905 12265 7908
rect 12299 7905 12311 7939
rect 12728 7936 12756 7967
rect 13280 7936 13308 7967
rect 15838 7936 15844 7948
rect 12728 7908 13216 7936
rect 13280 7908 15844 7936
rect 12253 7899 12311 7905
rect 11609 7871 11667 7877
rect 11516 7849 11574 7855
rect 11516 7815 11528 7849
rect 11562 7815 11574 7849
rect 11609 7837 11621 7871
rect 11655 7868 11667 7871
rect 11790 7868 11796 7880
rect 11655 7840 11796 7868
rect 11655 7837 11667 7840
rect 11609 7831 11667 7837
rect 11790 7828 11796 7840
rect 11848 7828 11854 7880
rect 12342 7868 12348 7880
rect 12303 7840 12348 7868
rect 12342 7828 12348 7840
rect 12400 7828 12406 7880
rect 12986 7868 12992 7880
rect 12947 7840 12992 7868
rect 12986 7828 12992 7840
rect 13044 7828 13050 7880
rect 13188 7877 13216 7908
rect 15838 7896 15844 7908
rect 15896 7936 15902 7948
rect 15933 7939 15991 7945
rect 15933 7936 15945 7939
rect 15896 7908 15945 7936
rect 15896 7896 15902 7908
rect 15933 7905 15945 7908
rect 15979 7905 15991 7939
rect 15933 7899 15991 7905
rect 13173 7871 13231 7877
rect 13173 7837 13185 7871
rect 13219 7837 13231 7871
rect 13814 7868 13820 7880
rect 13775 7840 13820 7868
rect 13173 7831 13231 7837
rect 13814 7828 13820 7840
rect 13872 7828 13878 7880
rect 14001 7871 14059 7877
rect 14001 7837 14013 7871
rect 14047 7837 14059 7871
rect 14001 7831 14059 7837
rect 14599 7871 14657 7877
rect 14599 7837 14611 7871
rect 14645 7868 14657 7871
rect 14734 7868 14740 7880
rect 14645 7840 14740 7868
rect 14645 7837 14657 7840
rect 14599 7831 14657 7837
rect 11516 7812 11574 7815
rect 11514 7760 11520 7812
rect 11572 7760 11578 7812
rect 11698 7800 11704 7812
rect 11659 7772 11704 7800
rect 11698 7760 11704 7772
rect 11756 7760 11762 7812
rect 11882 7800 11888 7812
rect 11843 7772 11888 7800
rect 11882 7760 11888 7772
rect 11940 7760 11946 7812
rect 14016 7800 14044 7831
rect 14734 7828 14740 7840
rect 14792 7828 14798 7880
rect 14829 7871 14887 7877
rect 14829 7837 14841 7871
rect 14875 7837 14887 7871
rect 14829 7831 14887 7837
rect 14844 7800 14872 7831
rect 14918 7828 14924 7880
rect 14976 7868 14982 7880
rect 15194 7868 15200 7880
rect 14976 7840 15021 7868
rect 15155 7840 15200 7868
rect 14976 7828 14982 7840
rect 15194 7828 15200 7840
rect 15252 7828 15258 7880
rect 15473 7871 15531 7877
rect 15473 7837 15485 7871
rect 15519 7837 15531 7871
rect 15473 7831 15531 7837
rect 15105 7803 15163 7809
rect 15105 7800 15117 7803
rect 14016 7772 15117 7800
rect 15105 7769 15117 7772
rect 15151 7800 15163 7803
rect 15381 7803 15439 7809
rect 15381 7800 15393 7803
rect 15151 7772 15393 7800
rect 15151 7769 15163 7772
rect 15105 7763 15163 7769
rect 15381 7769 15393 7772
rect 15427 7769 15439 7803
rect 15381 7763 15439 7769
rect 14734 7732 14740 7744
rect 8036 7704 11468 7732
rect 14695 7704 14740 7732
rect 14734 7692 14740 7704
rect 14792 7692 14798 7744
rect 14918 7692 14924 7744
rect 14976 7732 14982 7744
rect 15488 7732 15516 7831
rect 15562 7760 15568 7812
rect 15620 7800 15626 7812
rect 16209 7803 16267 7809
rect 16209 7800 16221 7803
rect 15620 7772 16221 7800
rect 15620 7760 15626 7772
rect 16209 7769 16221 7772
rect 16255 7769 16267 7803
rect 16209 7763 16267 7769
rect 16298 7760 16304 7812
rect 16356 7800 16362 7812
rect 16356 7772 16698 7800
rect 16356 7760 16362 7772
rect 17586 7760 17592 7812
rect 17644 7800 17650 7812
rect 17957 7803 18015 7809
rect 17957 7800 17969 7803
rect 17644 7772 17969 7800
rect 17644 7760 17650 7772
rect 17957 7769 17969 7772
rect 18003 7769 18015 7803
rect 17957 7763 18015 7769
rect 17604 7732 17632 7760
rect 14976 7704 17632 7732
rect 14976 7692 14982 7704
rect 0 7642 18860 7664
rect 0 7590 4660 7642
rect 4712 7590 4724 7642
rect 4776 7590 4788 7642
rect 4840 7590 4852 7642
rect 4904 7590 4916 7642
rect 4968 7590 7760 7642
rect 7812 7590 7824 7642
rect 7876 7590 7888 7642
rect 7940 7590 7952 7642
rect 8004 7590 8016 7642
rect 8068 7590 10860 7642
rect 10912 7590 10924 7642
rect 10976 7590 10988 7642
rect 11040 7590 11052 7642
rect 11104 7590 11116 7642
rect 11168 7590 13960 7642
rect 14012 7590 14024 7642
rect 14076 7590 14088 7642
rect 14140 7590 14152 7642
rect 14204 7590 14216 7642
rect 14268 7590 17060 7642
rect 17112 7590 17124 7642
rect 17176 7590 17188 7642
rect 17240 7590 17252 7642
rect 17304 7590 17316 7642
rect 17368 7590 18860 7642
rect 0 7568 18860 7590
rect 566 7488 572 7540
rect 624 7528 630 7540
rect 1673 7531 1731 7537
rect 1673 7528 1685 7531
rect 624 7500 1685 7528
rect 624 7488 630 7500
rect 1673 7497 1685 7500
rect 1719 7497 1731 7531
rect 1946 7528 1952 7540
rect 1673 7491 1731 7497
rect 1780 7500 1952 7528
rect 1397 7395 1455 7401
rect 1397 7361 1409 7395
rect 1443 7392 1455 7395
rect 1780 7392 1808 7500
rect 1946 7488 1952 7500
rect 2004 7528 2010 7540
rect 2961 7531 3019 7537
rect 2961 7528 2973 7531
rect 2004 7500 2973 7528
rect 2004 7488 2010 7500
rect 2961 7497 2973 7500
rect 3007 7497 3019 7531
rect 2961 7491 3019 7497
rect 3142 7488 3148 7540
rect 3200 7528 3206 7540
rect 3694 7528 3700 7540
rect 3200 7500 3700 7528
rect 3200 7488 3206 7500
rect 3694 7488 3700 7500
rect 3752 7528 3758 7540
rect 5810 7528 5816 7540
rect 3752 7500 5816 7528
rect 3752 7488 3758 7500
rect 1857 7463 1915 7469
rect 1857 7429 1869 7463
rect 1903 7460 1915 7463
rect 2590 7460 2596 7472
rect 1903 7432 2596 7460
rect 1903 7429 1915 7432
rect 1857 7423 1915 7429
rect 2590 7420 2596 7432
rect 2648 7420 2654 7472
rect 3878 7460 3884 7472
rect 2792 7432 3884 7460
rect 2792 7404 2820 7432
rect 3878 7420 3884 7432
rect 3936 7420 3942 7472
rect 1443 7364 1808 7392
rect 1949 7395 2007 7401
rect 1443 7361 1455 7364
rect 1397 7355 1455 7361
rect 1949 7361 1961 7395
rect 1995 7392 2007 7395
rect 2038 7392 2044 7404
rect 1995 7364 2044 7392
rect 1995 7361 2007 7364
rect 1949 7355 2007 7361
rect 2038 7352 2044 7364
rect 2096 7352 2102 7404
rect 2317 7395 2375 7401
rect 2317 7361 2329 7395
rect 2363 7361 2375 7395
rect 2498 7392 2504 7404
rect 2459 7364 2504 7392
rect 2317 7355 2375 7361
rect 2332 7268 2360 7355
rect 2498 7352 2504 7364
rect 2556 7352 2562 7404
rect 2774 7352 2780 7404
rect 2832 7392 2838 7404
rect 3142 7392 3148 7404
rect 2832 7364 2925 7392
rect 3103 7364 3148 7392
rect 2832 7352 2838 7364
rect 3142 7352 3148 7364
rect 3200 7352 3206 7404
rect 3237 7395 3295 7401
rect 3237 7361 3249 7395
rect 3283 7361 3295 7395
rect 3237 7355 3295 7361
rect 2406 7284 2412 7336
rect 2464 7324 2470 7336
rect 3252 7324 3280 7355
rect 3326 7352 3332 7404
rect 3384 7392 3390 7404
rect 3384 7364 3429 7392
rect 3384 7352 3390 7364
rect 3510 7352 3516 7404
rect 3568 7392 3574 7404
rect 3697 7395 3755 7401
rect 3697 7392 3709 7395
rect 3568 7364 3709 7392
rect 3568 7352 3574 7364
rect 3697 7361 3709 7364
rect 3743 7361 3755 7395
rect 3697 7355 3755 7361
rect 4801 7395 4859 7401
rect 4801 7361 4813 7395
rect 4847 7392 4859 7395
rect 4908 7392 4936 7500
rect 5810 7488 5816 7500
rect 5868 7488 5874 7540
rect 5902 7488 5908 7540
rect 5960 7528 5966 7540
rect 6086 7528 6092 7540
rect 5960 7500 6092 7528
rect 5960 7488 5966 7500
rect 6086 7488 6092 7500
rect 6144 7488 6150 7540
rect 9582 7528 9588 7540
rect 6656 7500 9588 7528
rect 6178 7460 6184 7472
rect 5000 7432 6184 7460
rect 5000 7401 5028 7432
rect 6178 7420 6184 7432
rect 6236 7460 6242 7472
rect 6457 7463 6515 7469
rect 6457 7460 6469 7463
rect 6236 7432 6469 7460
rect 6236 7420 6242 7432
rect 6457 7429 6469 7432
rect 6503 7429 6515 7463
rect 6457 7423 6515 7429
rect 4847 7364 4936 7392
rect 4985 7395 5043 7401
rect 4847 7361 4859 7364
rect 4801 7355 4859 7361
rect 4985 7361 4997 7395
rect 5031 7361 5043 7395
rect 5258 7392 5264 7404
rect 5219 7364 5264 7392
rect 4985 7355 5043 7361
rect 5258 7352 5264 7364
rect 5316 7352 5322 7404
rect 5718 7392 5724 7404
rect 5679 7364 5724 7392
rect 5718 7352 5724 7364
rect 5776 7352 5782 7404
rect 5902 7392 5908 7404
rect 5863 7364 5908 7392
rect 5902 7352 5908 7364
rect 5960 7352 5966 7404
rect 6365 7395 6423 7401
rect 6365 7392 6377 7395
rect 6288 7364 6377 7392
rect 5074 7324 5080 7336
rect 2464 7296 2509 7324
rect 3252 7296 4108 7324
rect 4987 7296 5080 7324
rect 2464 7284 2470 7296
rect 4080 7268 4108 7296
rect 5074 7284 5080 7296
rect 5132 7324 5138 7336
rect 5997 7327 6055 7333
rect 5997 7324 6009 7327
rect 5132 7296 6009 7324
rect 5132 7284 5138 7296
rect 5997 7293 6009 7296
rect 6043 7324 6055 7327
rect 6086 7324 6092 7336
rect 6043 7296 6092 7324
rect 6043 7293 6055 7296
rect 5997 7287 6055 7293
rect 6086 7284 6092 7296
rect 6144 7284 6150 7336
rect 2314 7256 2320 7268
rect 2227 7228 2320 7256
rect 2314 7216 2320 7228
rect 2372 7256 2378 7268
rect 2372 7228 3188 7256
rect 2372 7216 2378 7228
rect 1489 7191 1547 7197
rect 1489 7157 1501 7191
rect 1535 7188 1547 7191
rect 2406 7188 2412 7200
rect 1535 7160 2412 7188
rect 1535 7157 1547 7160
rect 1489 7151 1547 7157
rect 2406 7148 2412 7160
rect 2464 7148 2470 7200
rect 2682 7188 2688 7200
rect 2643 7160 2688 7188
rect 2682 7148 2688 7160
rect 2740 7148 2746 7200
rect 3160 7188 3188 7228
rect 4062 7216 4068 7268
rect 4120 7256 4126 7268
rect 5258 7256 5264 7268
rect 4120 7228 5264 7256
rect 4120 7216 4126 7228
rect 5258 7216 5264 7228
rect 5316 7216 5322 7268
rect 3605 7191 3663 7197
rect 3605 7188 3617 7191
rect 3160 7160 3617 7188
rect 3605 7157 3617 7160
rect 3651 7157 3663 7191
rect 3605 7151 3663 7157
rect 4246 7148 4252 7200
rect 4304 7188 4310 7200
rect 6288 7188 6316 7364
rect 6365 7361 6377 7364
rect 6411 7392 6423 7395
rect 6656 7392 6684 7500
rect 9582 7488 9588 7500
rect 9640 7488 9646 7540
rect 9953 7531 10011 7537
rect 9953 7497 9965 7531
rect 9999 7528 10011 7531
rect 10410 7528 10416 7540
rect 9999 7500 10416 7528
rect 9999 7497 10011 7500
rect 9953 7491 10011 7497
rect 10410 7488 10416 7500
rect 10468 7488 10474 7540
rect 11422 7528 11428 7540
rect 10520 7500 11428 7528
rect 6748 7432 9076 7460
rect 6748 7401 6776 7432
rect 9048 7404 9076 7432
rect 6411 7364 6684 7392
rect 6733 7395 6791 7401
rect 6411 7361 6423 7364
rect 6365 7355 6423 7361
rect 6733 7361 6745 7395
rect 6779 7361 6791 7395
rect 6733 7355 6791 7361
rect 6638 7284 6644 7336
rect 6696 7324 6702 7336
rect 6748 7324 6776 7355
rect 6914 7352 6920 7404
rect 6972 7392 6978 7404
rect 7837 7395 7895 7401
rect 7837 7392 7849 7395
rect 6972 7364 7849 7392
rect 6972 7352 6978 7364
rect 7837 7361 7849 7364
rect 7883 7361 7895 7395
rect 8938 7392 8944 7404
rect 8899 7364 8944 7392
rect 7837 7355 7895 7361
rect 8938 7352 8944 7364
rect 8996 7352 9002 7404
rect 9030 7352 9036 7404
rect 9088 7392 9094 7404
rect 9088 7364 9133 7392
rect 9088 7352 9094 7364
rect 9214 7352 9220 7404
rect 9272 7392 9278 7404
rect 9585 7395 9643 7401
rect 9585 7392 9597 7395
rect 9272 7364 9597 7392
rect 9272 7352 9278 7364
rect 9585 7361 9597 7364
rect 9631 7361 9643 7395
rect 9585 7355 9643 7361
rect 9677 7395 9735 7401
rect 9677 7361 9689 7395
rect 9723 7361 9735 7395
rect 9677 7355 9735 7361
rect 9769 7395 9827 7401
rect 9769 7361 9781 7395
rect 9815 7392 9827 7395
rect 10410 7392 10416 7404
rect 9815 7364 10416 7392
rect 9815 7361 9827 7364
rect 9769 7355 9827 7361
rect 6696 7296 6776 7324
rect 6696 7284 6702 7296
rect 6822 7284 6828 7336
rect 6880 7324 6886 7336
rect 7929 7327 7987 7333
rect 6880 7296 6925 7324
rect 6880 7284 6886 7296
rect 7929 7293 7941 7327
rect 7975 7324 7987 7327
rect 8110 7324 8116 7336
rect 7975 7296 8116 7324
rect 7975 7293 7987 7296
rect 7929 7287 7987 7293
rect 8110 7284 8116 7296
rect 8168 7284 8174 7336
rect 9692 7324 9720 7355
rect 10410 7352 10416 7364
rect 10468 7352 10474 7404
rect 10520 7324 10548 7500
rect 11422 7488 11428 7500
rect 11480 7488 11486 7540
rect 15562 7528 15568 7540
rect 15523 7500 15568 7528
rect 15562 7488 15568 7500
rect 15620 7488 15626 7540
rect 17773 7531 17831 7537
rect 17773 7497 17785 7531
rect 17819 7528 17831 7531
rect 17954 7528 17960 7540
rect 17819 7500 17960 7528
rect 17819 7497 17831 7500
rect 17773 7491 17831 7497
rect 17954 7488 17960 7500
rect 18012 7488 18018 7540
rect 11974 7420 11980 7472
rect 12032 7420 12038 7472
rect 16298 7420 16304 7472
rect 16356 7420 16362 7472
rect 17037 7463 17095 7469
rect 17037 7429 17049 7463
rect 17083 7460 17095 7463
rect 18322 7460 18328 7472
rect 17083 7432 18328 7460
rect 17083 7429 17095 7432
rect 17037 7423 17095 7429
rect 18322 7420 18328 7432
rect 18380 7420 18386 7472
rect 10597 7395 10655 7401
rect 10597 7361 10609 7395
rect 10643 7392 10655 7395
rect 10643 7364 11100 7392
rect 10643 7361 10655 7364
rect 10597 7355 10655 7361
rect 9692 7296 9812 7324
rect 9784 7268 9812 7296
rect 10336 7296 10548 7324
rect 8205 7259 8263 7265
rect 8205 7225 8217 7259
rect 8251 7256 8263 7259
rect 8386 7256 8392 7268
rect 8251 7228 8392 7256
rect 8251 7225 8263 7228
rect 8205 7219 8263 7225
rect 8386 7216 8392 7228
rect 8444 7216 8450 7268
rect 9766 7216 9772 7268
rect 9824 7216 9830 7268
rect 4304 7160 6316 7188
rect 9217 7191 9275 7197
rect 4304 7148 4310 7160
rect 9217 7157 9229 7191
rect 9263 7188 9275 7191
rect 10336 7188 10364 7296
rect 10778 7284 10784 7336
rect 10836 7324 10842 7336
rect 10965 7327 11023 7333
rect 10965 7324 10977 7327
rect 10836 7296 10977 7324
rect 10836 7284 10842 7296
rect 10965 7293 10977 7296
rect 11011 7293 11023 7327
rect 11072 7324 11100 7364
rect 12342 7352 12348 7404
rect 12400 7401 12406 7404
rect 12400 7395 12449 7401
rect 12400 7361 12403 7395
rect 12437 7392 12449 7395
rect 12529 7395 12587 7401
rect 12529 7392 12541 7395
rect 12437 7364 12541 7392
rect 12437 7361 12449 7364
rect 12400 7355 12449 7361
rect 12529 7361 12541 7364
rect 12575 7361 12587 7395
rect 12529 7355 12587 7361
rect 12400 7352 12406 7355
rect 14734 7352 14740 7404
rect 14792 7392 14798 7404
rect 15105 7395 15163 7401
rect 15105 7392 15117 7395
rect 14792 7364 15117 7392
rect 14792 7352 14798 7364
rect 15105 7361 15117 7364
rect 15151 7392 15163 7395
rect 15194 7392 15200 7404
rect 15151 7364 15200 7392
rect 15151 7361 15163 7364
rect 15105 7355 15163 7361
rect 15194 7352 15200 7364
rect 15252 7352 15258 7404
rect 17313 7395 17371 7401
rect 17313 7361 17325 7395
rect 17359 7392 17371 7395
rect 17494 7392 17500 7404
rect 17359 7364 17500 7392
rect 17359 7361 17371 7364
rect 17313 7355 17371 7361
rect 17494 7352 17500 7364
rect 17552 7352 17558 7404
rect 11330 7324 11336 7336
rect 11072 7296 11336 7324
rect 10965 7287 11023 7293
rect 11330 7284 11336 7296
rect 11388 7284 11394 7336
rect 17862 7324 17868 7336
rect 17823 7296 17868 7324
rect 17862 7284 17868 7296
rect 17920 7284 17926 7336
rect 17957 7327 18015 7333
rect 17957 7293 17969 7327
rect 18003 7293 18015 7327
rect 17957 7287 18015 7293
rect 17972 7256 18000 7287
rect 17236 7228 18000 7256
rect 9263 7160 10364 7188
rect 9263 7157 9275 7160
rect 9217 7151 9275 7157
rect 10410 7148 10416 7200
rect 10468 7188 10474 7200
rect 12621 7191 12679 7197
rect 12621 7188 12633 7191
rect 10468 7160 12633 7188
rect 10468 7148 10474 7160
rect 12621 7157 12633 7160
rect 12667 7157 12679 7191
rect 15010 7188 15016 7200
rect 14923 7160 15016 7188
rect 12621 7151 12679 7157
rect 15010 7148 15016 7160
rect 15068 7188 15074 7200
rect 17236 7188 17264 7228
rect 17402 7188 17408 7200
rect 15068 7160 17264 7188
rect 17363 7160 17408 7188
rect 15068 7148 15074 7160
rect 17402 7148 17408 7160
rect 17460 7148 17466 7200
rect 0 7098 18860 7120
rect 0 7046 3110 7098
rect 3162 7046 3174 7098
rect 3226 7046 3238 7098
rect 3290 7046 3302 7098
rect 3354 7046 3366 7098
rect 3418 7046 6210 7098
rect 6262 7046 6274 7098
rect 6326 7046 6338 7098
rect 6390 7046 6402 7098
rect 6454 7046 6466 7098
rect 6518 7046 9310 7098
rect 9362 7046 9374 7098
rect 9426 7046 9438 7098
rect 9490 7046 9502 7098
rect 9554 7046 9566 7098
rect 9618 7046 12410 7098
rect 12462 7046 12474 7098
rect 12526 7046 12538 7098
rect 12590 7046 12602 7098
rect 12654 7046 12666 7098
rect 12718 7046 15510 7098
rect 15562 7046 15574 7098
rect 15626 7046 15638 7098
rect 15690 7046 15702 7098
rect 15754 7046 15766 7098
rect 15818 7046 18860 7098
rect 0 7024 18860 7046
rect 5626 6944 5632 6996
rect 5684 6984 5690 6996
rect 6638 6984 6644 6996
rect 5684 6956 6644 6984
rect 5684 6944 5690 6956
rect 6638 6944 6644 6956
rect 6696 6944 6702 6996
rect 10134 6984 10140 6996
rect 10095 6956 10140 6984
rect 10134 6944 10140 6956
rect 10192 6944 10198 6996
rect 10410 6984 10416 6996
rect 10371 6956 10416 6984
rect 10410 6944 10416 6956
rect 10468 6944 10474 6996
rect 12986 6984 12992 6996
rect 10612 6956 12992 6984
rect 2409 6919 2467 6925
rect 2409 6885 2421 6919
rect 2455 6916 2467 6919
rect 2774 6916 2780 6928
rect 2455 6888 2780 6916
rect 2455 6885 2467 6888
rect 2409 6879 2467 6885
rect 2774 6876 2780 6888
rect 2832 6876 2838 6928
rect 3234 6876 3240 6928
rect 3292 6916 3298 6928
rect 3602 6916 3608 6928
rect 3292 6888 3608 6916
rect 3292 6876 3298 6888
rect 3602 6876 3608 6888
rect 3660 6876 3666 6928
rect 5902 6876 5908 6928
rect 5960 6916 5966 6928
rect 9401 6919 9459 6925
rect 5960 6888 7328 6916
rect 5960 6876 5966 6888
rect 1946 6848 1952 6860
rect 1907 6820 1952 6848
rect 1946 6808 1952 6820
rect 2004 6808 2010 6860
rect 2958 6848 2964 6860
rect 2871 6820 2964 6848
rect 2958 6808 2964 6820
rect 3016 6848 3022 6860
rect 3016 6820 3372 6848
rect 3016 6808 3022 6820
rect 1489 6783 1547 6789
rect 1489 6749 1501 6783
rect 1535 6749 1547 6783
rect 1489 6743 1547 6749
rect 1581 6783 1639 6789
rect 1581 6749 1593 6783
rect 1627 6780 1639 6783
rect 2682 6780 2688 6792
rect 1627 6752 2688 6780
rect 1627 6749 1639 6752
rect 1581 6743 1639 6749
rect 1504 6712 1532 6743
rect 2682 6740 2688 6752
rect 2740 6780 2746 6792
rect 2777 6783 2835 6789
rect 2777 6780 2789 6783
rect 2740 6752 2789 6780
rect 2740 6740 2746 6752
rect 2777 6749 2789 6752
rect 2823 6749 2835 6783
rect 2777 6743 2835 6749
rect 2038 6712 2044 6724
rect 1504 6684 2044 6712
rect 2038 6672 2044 6684
rect 2096 6712 2102 6724
rect 2976 6712 3004 6808
rect 3053 6783 3111 6789
rect 3053 6749 3065 6783
rect 3099 6749 3111 6783
rect 3234 6780 3240 6792
rect 3195 6752 3240 6780
rect 3053 6743 3111 6749
rect 2096 6684 3004 6712
rect 3068 6712 3096 6743
rect 3234 6740 3240 6752
rect 3292 6740 3298 6792
rect 3344 6789 3372 6820
rect 6086 6808 6092 6860
rect 6144 6848 6150 6860
rect 6365 6851 6423 6857
rect 6365 6848 6377 6851
rect 6144 6820 6377 6848
rect 6144 6808 6150 6820
rect 6365 6817 6377 6820
rect 6411 6848 6423 6851
rect 7300 6848 7328 6888
rect 7760 6888 8800 6916
rect 7561 6851 7619 6857
rect 7561 6848 7573 6851
rect 6411 6820 7236 6848
rect 7300 6820 7573 6848
rect 6411 6817 6423 6820
rect 6365 6811 6423 6817
rect 3329 6783 3387 6789
rect 3329 6749 3341 6783
rect 3375 6749 3387 6783
rect 3510 6780 3516 6792
rect 3471 6752 3516 6780
rect 3329 6743 3387 6749
rect 3510 6740 3516 6752
rect 3568 6740 3574 6792
rect 4062 6780 4068 6792
rect 4023 6752 4068 6780
rect 4062 6740 4068 6752
rect 4120 6740 4126 6792
rect 6457 6783 6515 6789
rect 6457 6749 6469 6783
rect 6503 6780 6515 6783
rect 7208 6780 7236 6820
rect 7561 6817 7573 6820
rect 7607 6848 7619 6851
rect 7760 6848 7788 6888
rect 7607 6820 7788 6848
rect 7837 6851 7895 6857
rect 7607 6817 7619 6820
rect 7561 6811 7619 6817
rect 7837 6817 7849 6851
rect 7883 6848 7895 6851
rect 8018 6848 8024 6860
rect 7883 6820 8024 6848
rect 7883 6817 7895 6820
rect 7837 6811 7895 6817
rect 8018 6808 8024 6820
rect 8076 6848 8082 6860
rect 8481 6851 8539 6857
rect 8481 6848 8493 6851
rect 8076 6820 8493 6848
rect 8076 6808 8082 6820
rect 8481 6817 8493 6820
rect 8527 6817 8539 6851
rect 8662 6848 8668 6860
rect 8623 6820 8668 6848
rect 8481 6811 8539 6817
rect 8662 6808 8668 6820
rect 8720 6808 8726 6860
rect 8772 6848 8800 6888
rect 9401 6885 9413 6919
rect 9447 6916 9459 6919
rect 10502 6916 10508 6928
rect 9447 6888 10508 6916
rect 9447 6885 9459 6888
rect 9401 6879 9459 6885
rect 10502 6876 10508 6888
rect 10560 6876 10566 6928
rect 8772 6820 9628 6848
rect 8386 6780 8392 6792
rect 6503 6752 6960 6780
rect 7208 6752 8156 6780
rect 8347 6752 8392 6780
rect 6503 6749 6515 6752
rect 6457 6743 6515 6749
rect 3421 6715 3479 6721
rect 3421 6712 3433 6715
rect 3068 6684 3433 6712
rect 2096 6672 2102 6684
rect 3421 6681 3433 6684
rect 3467 6681 3479 6715
rect 4338 6712 4344 6724
rect 4299 6684 4344 6712
rect 3421 6675 3479 6681
rect 4338 6672 4344 6684
rect 4396 6672 4402 6724
rect 4430 6672 4436 6724
rect 4488 6712 4494 6724
rect 4488 6684 4830 6712
rect 4488 6672 4494 6684
rect 566 6604 572 6656
rect 624 6644 630 6656
rect 1305 6647 1363 6653
rect 1305 6644 1317 6647
rect 624 6616 1317 6644
rect 624 6604 630 6616
rect 1305 6613 1317 6616
rect 1351 6613 1363 6647
rect 1305 6607 1363 6613
rect 2406 6604 2412 6656
rect 2464 6644 2470 6656
rect 2501 6647 2559 6653
rect 2501 6644 2513 6647
rect 2464 6616 2513 6644
rect 2464 6604 2470 6616
rect 2501 6613 2513 6616
rect 2547 6613 2559 6647
rect 2501 6607 2559 6613
rect 2590 6604 2596 6656
rect 2648 6644 2654 6656
rect 2961 6647 3019 6653
rect 2961 6644 2973 6647
rect 2648 6616 2973 6644
rect 2648 6604 2654 6616
rect 2961 6613 2973 6616
rect 3007 6613 3019 6647
rect 2961 6607 3019 6613
rect 5813 6647 5871 6653
rect 5813 6613 5825 6647
rect 5859 6644 5871 6647
rect 5902 6644 5908 6656
rect 5859 6616 5908 6644
rect 5859 6613 5871 6616
rect 5813 6607 5871 6613
rect 5902 6604 5908 6616
rect 5960 6604 5966 6656
rect 6086 6604 6092 6656
rect 6144 6644 6150 6656
rect 6181 6647 6239 6653
rect 6181 6644 6193 6647
rect 6144 6616 6193 6644
rect 6144 6604 6150 6616
rect 6181 6613 6193 6616
rect 6227 6613 6239 6647
rect 6822 6644 6828 6656
rect 6783 6616 6828 6644
rect 6181 6607 6239 6613
rect 6822 6604 6828 6616
rect 6880 6604 6886 6656
rect 6932 6653 6960 6752
rect 7285 6715 7343 6721
rect 7285 6681 7297 6715
rect 7331 6712 7343 6715
rect 8128 6712 8156 6752
rect 8386 6740 8392 6752
rect 8444 6740 8450 6792
rect 8570 6740 8576 6792
rect 8628 6780 8634 6792
rect 9214 6780 9220 6792
rect 8628 6752 9220 6780
rect 8628 6740 8634 6752
rect 9214 6740 9220 6752
rect 9272 6780 9278 6792
rect 9493 6783 9551 6789
rect 9493 6780 9505 6783
rect 9272 6752 9505 6780
rect 9272 6740 9278 6752
rect 9493 6749 9505 6752
rect 9539 6749 9551 6783
rect 9600 6780 9628 6820
rect 9766 6808 9772 6860
rect 9824 6848 9830 6860
rect 10612 6848 10640 6956
rect 12986 6944 12992 6956
rect 13044 6944 13050 6996
rect 15194 6984 15200 6996
rect 15155 6956 15200 6984
rect 15194 6944 15200 6956
rect 15252 6944 15258 6996
rect 17773 6987 17831 6993
rect 17773 6953 17785 6987
rect 17819 6984 17831 6987
rect 17862 6984 17868 6996
rect 17819 6956 17868 6984
rect 17819 6953 17831 6956
rect 17773 6947 17831 6953
rect 17862 6944 17868 6956
rect 17920 6944 17926 6996
rect 18322 6984 18328 6996
rect 18283 6956 18328 6984
rect 18322 6944 18328 6956
rect 18380 6944 18386 6996
rect 11333 6851 11391 6857
rect 11333 6848 11345 6851
rect 9824 6820 10640 6848
rect 10888 6820 11345 6848
rect 9824 6808 9830 6820
rect 9858 6780 9864 6792
rect 9600 6752 9864 6780
rect 9493 6743 9551 6749
rect 9401 6715 9459 6721
rect 9401 6712 9413 6715
rect 7331 6684 8064 6712
rect 8128 6684 9413 6712
rect 7331 6681 7343 6684
rect 7285 6675 7343 6681
rect 8036 6653 8064 6684
rect 9401 6681 9413 6684
rect 9447 6681 9459 6715
rect 9508 6712 9536 6743
rect 9858 6740 9864 6752
rect 9916 6740 9922 6792
rect 9968 6789 9996 6820
rect 10244 6792 10272 6820
rect 9953 6783 10011 6789
rect 9953 6749 9965 6783
rect 9999 6749 10011 6783
rect 9953 6743 10011 6749
rect 10137 6783 10195 6789
rect 10137 6749 10149 6783
rect 10183 6749 10195 6783
rect 10137 6743 10195 6749
rect 10152 6712 10180 6743
rect 10226 6740 10232 6792
rect 10284 6740 10290 6792
rect 10318 6740 10324 6792
rect 10376 6780 10382 6792
rect 10888 6780 10916 6820
rect 11333 6817 11345 6820
rect 11379 6817 11391 6851
rect 11882 6848 11888 6860
rect 11333 6811 11391 6817
rect 11440 6820 11888 6848
rect 10376 6752 10916 6780
rect 11149 6783 11207 6789
rect 10376 6740 10382 6752
rect 11149 6749 11161 6783
rect 11195 6780 11207 6783
rect 11238 6780 11244 6792
rect 11195 6752 11244 6780
rect 11195 6749 11207 6752
rect 11149 6743 11207 6749
rect 11238 6740 11244 6752
rect 11296 6740 11302 6792
rect 11440 6780 11468 6820
rect 11882 6808 11888 6820
rect 11940 6848 11946 6860
rect 13909 6851 13967 6857
rect 13909 6848 13921 6851
rect 11940 6820 13921 6848
rect 11940 6808 11946 6820
rect 13909 6817 13921 6820
rect 13955 6848 13967 6851
rect 14826 6848 14832 6860
rect 13955 6820 14832 6848
rect 13955 6817 13967 6820
rect 13909 6811 13967 6817
rect 14826 6808 14832 6820
rect 14884 6808 14890 6860
rect 15010 6848 15016 6860
rect 14971 6820 15016 6848
rect 15010 6808 15016 6820
rect 15068 6808 15074 6860
rect 15562 6848 15568 6860
rect 15475 6820 15568 6848
rect 15562 6808 15568 6820
rect 15620 6848 15626 6860
rect 17313 6851 17371 6857
rect 15620 6820 16344 6848
rect 15620 6808 15626 6820
rect 11348 6752 11468 6780
rect 9508 6684 10180 6712
rect 9401 6675 9459 6681
rect 10686 6672 10692 6724
rect 10744 6712 10750 6724
rect 11348 6712 11376 6752
rect 11514 6740 11520 6792
rect 11572 6780 11578 6792
rect 11609 6783 11667 6789
rect 11609 6780 11621 6783
rect 11572 6752 11621 6780
rect 11572 6740 11578 6752
rect 11609 6749 11621 6752
rect 11655 6749 11667 6783
rect 11609 6743 11667 6749
rect 13538 6740 13544 6792
rect 13596 6780 13602 6792
rect 14737 6783 14795 6789
rect 14737 6780 14749 6783
rect 13596 6752 14749 6780
rect 13596 6740 13602 6752
rect 14737 6749 14749 6752
rect 14783 6749 14795 6783
rect 14737 6743 14795 6749
rect 15194 6740 15200 6792
rect 15252 6780 15258 6792
rect 15381 6783 15439 6789
rect 15381 6780 15393 6783
rect 15252 6752 15393 6780
rect 15252 6740 15258 6752
rect 15381 6749 15393 6752
rect 15427 6749 15439 6783
rect 15381 6743 15439 6749
rect 15470 6740 15476 6792
rect 15528 6780 15534 6792
rect 15528 6752 15573 6780
rect 15528 6740 15534 6752
rect 10744 6684 11376 6712
rect 10744 6672 10750 6684
rect 6917 6647 6975 6653
rect 6917 6613 6929 6647
rect 6963 6613 6975 6647
rect 6917 6607 6975 6613
rect 7377 6647 7435 6653
rect 7377 6613 7389 6647
rect 7423 6644 7435 6647
rect 7837 6647 7895 6653
rect 7837 6644 7849 6647
rect 7423 6616 7849 6644
rect 7423 6613 7435 6616
rect 7377 6607 7435 6613
rect 7837 6613 7849 6616
rect 7883 6613 7895 6647
rect 7837 6607 7895 6613
rect 8021 6647 8079 6653
rect 8021 6613 8033 6647
rect 8067 6613 8079 6647
rect 9582 6644 9588 6656
rect 9543 6616 9588 6644
rect 8021 6607 8079 6613
rect 9582 6604 9588 6616
rect 9640 6604 9646 6656
rect 10778 6644 10784 6656
rect 10739 6616 10784 6644
rect 10778 6604 10784 6616
rect 10836 6604 10842 6656
rect 11241 6647 11299 6653
rect 11241 6613 11253 6647
rect 11287 6644 11299 6647
rect 11348 6644 11376 6684
rect 13633 6715 13691 6721
rect 13633 6681 13645 6715
rect 13679 6712 13691 6715
rect 16316 6712 16344 6820
rect 17313 6817 17325 6851
rect 17359 6848 17371 6851
rect 17586 6848 17592 6860
rect 17359 6820 17592 6848
rect 17359 6817 17371 6820
rect 17313 6811 17371 6817
rect 17586 6808 17592 6820
rect 17644 6808 17650 6860
rect 17129 6783 17187 6789
rect 17129 6749 17141 6783
rect 17175 6780 17187 6783
rect 17402 6780 17408 6792
rect 17175 6752 17408 6780
rect 17175 6749 17187 6752
rect 17129 6743 17187 6749
rect 17402 6740 17408 6752
rect 17460 6740 17466 6792
rect 17770 6780 17776 6792
rect 17731 6752 17776 6780
rect 17770 6740 17776 6752
rect 17828 6740 17834 6792
rect 18506 6780 18512 6792
rect 18467 6752 18512 6780
rect 18506 6740 18512 6752
rect 18564 6740 18570 6792
rect 17221 6715 17279 6721
rect 17221 6712 17233 6715
rect 13679 6684 14412 6712
rect 16316 6684 17233 6712
rect 13679 6681 13691 6684
rect 13633 6675 13691 6681
rect 11287 6616 11376 6644
rect 11287 6613 11299 6616
rect 11241 6607 11299 6613
rect 11514 6604 11520 6656
rect 11572 6644 11578 6656
rect 11793 6647 11851 6653
rect 11793 6644 11805 6647
rect 11572 6616 11805 6644
rect 11572 6604 11578 6616
rect 11793 6613 11805 6616
rect 11839 6613 11851 6647
rect 11793 6607 11851 6613
rect 13170 6604 13176 6656
rect 13228 6644 13234 6656
rect 13265 6647 13323 6653
rect 13265 6644 13277 6647
rect 13228 6616 13277 6644
rect 13228 6604 13234 6616
rect 13265 6613 13277 6616
rect 13311 6613 13323 6647
rect 13265 6607 13323 6613
rect 13725 6647 13783 6653
rect 13725 6613 13737 6647
rect 13771 6644 13783 6647
rect 13814 6644 13820 6656
rect 13771 6616 13820 6644
rect 13771 6613 13783 6616
rect 13725 6607 13783 6613
rect 13814 6604 13820 6616
rect 13872 6604 13878 6656
rect 14384 6653 14412 6684
rect 17221 6681 17233 6684
rect 17267 6712 17279 6715
rect 17788 6712 17816 6740
rect 17267 6684 17816 6712
rect 17267 6681 17279 6684
rect 17221 6675 17279 6681
rect 14369 6647 14427 6653
rect 14369 6613 14381 6647
rect 14415 6613 14427 6647
rect 14369 6607 14427 6613
rect 14826 6604 14832 6656
rect 14884 6644 14890 6656
rect 14884 6616 14929 6644
rect 14884 6604 14890 6616
rect 16390 6604 16396 6656
rect 16448 6644 16454 6656
rect 16761 6647 16819 6653
rect 16761 6644 16773 6647
rect 16448 6616 16773 6644
rect 16448 6604 16454 6616
rect 16761 6613 16773 6616
rect 16807 6613 16819 6647
rect 16761 6607 16819 6613
rect 0 6554 18860 6576
rect 0 6502 4660 6554
rect 4712 6502 4724 6554
rect 4776 6502 4788 6554
rect 4840 6502 4852 6554
rect 4904 6502 4916 6554
rect 4968 6502 7760 6554
rect 7812 6502 7824 6554
rect 7876 6502 7888 6554
rect 7940 6502 7952 6554
rect 8004 6502 8016 6554
rect 8068 6502 10860 6554
rect 10912 6502 10924 6554
rect 10976 6502 10988 6554
rect 11040 6502 11052 6554
rect 11104 6502 11116 6554
rect 11168 6502 13960 6554
rect 14012 6502 14024 6554
rect 14076 6502 14088 6554
rect 14140 6502 14152 6554
rect 14204 6502 14216 6554
rect 14268 6502 17060 6554
rect 17112 6502 17124 6554
rect 17176 6502 17188 6554
rect 17240 6502 17252 6554
rect 17304 6502 17316 6554
rect 17368 6502 18860 6554
rect 0 6480 18860 6502
rect 2038 6440 2044 6452
rect 1999 6412 2044 6440
rect 2038 6400 2044 6412
rect 2096 6400 2102 6452
rect 4338 6400 4344 6452
rect 4396 6440 4402 6452
rect 4433 6443 4491 6449
rect 4433 6440 4445 6443
rect 4396 6412 4445 6440
rect 4396 6400 4402 6412
rect 4433 6409 4445 6412
rect 4479 6409 4491 6443
rect 4433 6403 4491 6409
rect 5077 6443 5135 6449
rect 5077 6409 5089 6443
rect 5123 6440 5135 6443
rect 6181 6443 6239 6449
rect 6181 6440 6193 6443
rect 5123 6412 6193 6440
rect 5123 6409 5135 6412
rect 5077 6403 5135 6409
rect 6181 6409 6193 6412
rect 6227 6409 6239 6443
rect 6822 6440 6828 6452
rect 6783 6412 6828 6440
rect 6181 6403 6239 6409
rect 6822 6400 6828 6412
rect 6880 6400 6886 6452
rect 8021 6443 8079 6449
rect 8021 6440 8033 6443
rect 6932 6412 8033 6440
rect 566 6372 572 6384
rect 527 6344 572 6372
rect 566 6332 572 6344
rect 624 6332 630 6384
rect 5629 6375 5687 6381
rect 5629 6341 5641 6375
rect 5675 6372 5687 6375
rect 6932 6372 6960 6412
rect 8021 6409 8033 6412
rect 8067 6409 8079 6443
rect 8021 6403 8079 6409
rect 8481 6443 8539 6449
rect 8481 6409 8493 6443
rect 8527 6440 8539 6443
rect 9030 6440 9036 6452
rect 8527 6412 9036 6440
rect 8527 6409 8539 6412
rect 8481 6403 8539 6409
rect 9030 6400 9036 6412
rect 9088 6400 9094 6452
rect 10229 6443 10287 6449
rect 10229 6409 10241 6443
rect 10275 6440 10287 6443
rect 10413 6443 10471 6449
rect 10413 6440 10425 6443
rect 10275 6412 10425 6440
rect 10275 6409 10287 6412
rect 10229 6403 10287 6409
rect 10413 6409 10425 6412
rect 10459 6409 10471 6443
rect 11149 6443 11207 6449
rect 10413 6403 10471 6409
rect 10695 6412 11008 6440
rect 8662 6372 8668 6384
rect 5675 6344 6960 6372
rect 8575 6344 8668 6372
rect 5675 6341 5687 6344
rect 5629 6335 5687 6341
rect 8662 6332 8668 6344
rect 8720 6372 8726 6384
rect 9582 6372 9588 6384
rect 8720 6344 9588 6372
rect 8720 6332 8726 6344
rect 9582 6332 9588 6344
rect 9640 6372 9646 6384
rect 10695 6372 10723 6412
rect 9640 6344 10723 6372
rect 9640 6332 9646 6344
rect 2314 6304 2320 6316
rect 290 6236 296 6248
rect 251 6208 296 6236
rect 290 6196 296 6208
rect 348 6196 354 6248
rect 1688 6168 1716 6290
rect 2275 6276 2320 6304
rect 2314 6264 2320 6276
rect 2372 6264 2378 6316
rect 2406 6264 2412 6316
rect 2464 6304 2470 6316
rect 4617 6307 4675 6313
rect 2464 6276 2509 6304
rect 2464 6264 2470 6276
rect 4617 6273 4629 6307
rect 4663 6304 4675 6307
rect 5074 6304 5080 6316
rect 4663 6276 5080 6304
rect 4663 6273 4675 6276
rect 4617 6267 4675 6273
rect 5074 6264 5080 6276
rect 5132 6264 5138 6316
rect 5718 6304 5724 6316
rect 5679 6276 5724 6304
rect 5718 6264 5724 6276
rect 5776 6264 5782 6316
rect 5902 6264 5908 6316
rect 5960 6304 5966 6316
rect 6089 6307 6147 6313
rect 6089 6304 6101 6307
rect 5960 6276 6101 6304
rect 5960 6264 5966 6276
rect 6089 6273 6101 6276
rect 6135 6273 6147 6307
rect 6270 6304 6276 6316
rect 6231 6276 6276 6304
rect 6089 6267 6147 6273
rect 2590 6236 2596 6248
rect 2551 6208 2596 6236
rect 2590 6196 2596 6208
rect 2648 6196 2654 6248
rect 4709 6239 4767 6245
rect 4709 6205 4721 6239
rect 4755 6205 4767 6239
rect 5810 6236 5816 6248
rect 5771 6208 5816 6236
rect 4709 6199 4767 6205
rect 1854 6168 1860 6180
rect 1688 6140 1860 6168
rect 1854 6128 1860 6140
rect 1912 6168 1918 6180
rect 2406 6168 2412 6180
rect 1912 6140 2412 6168
rect 1912 6128 1918 6140
rect 2406 6128 2412 6140
rect 2464 6168 2470 6180
rect 4430 6168 4436 6180
rect 2464 6140 4436 6168
rect 2464 6128 2470 6140
rect 4430 6128 4436 6140
rect 4488 6128 4494 6180
rect 4724 6168 4752 6199
rect 5810 6196 5816 6208
rect 5868 6196 5874 6248
rect 6104 6236 6132 6267
rect 6270 6264 6276 6276
rect 6328 6264 6334 6316
rect 6365 6307 6423 6313
rect 6365 6273 6377 6307
rect 6411 6304 6423 6307
rect 6546 6304 6552 6316
rect 6411 6276 6552 6304
rect 6411 6273 6423 6276
rect 6365 6267 6423 6273
rect 6546 6264 6552 6276
rect 6604 6304 6610 6316
rect 6641 6307 6699 6313
rect 6641 6304 6653 6307
rect 6604 6276 6653 6304
rect 6604 6264 6610 6276
rect 6641 6273 6653 6276
rect 6687 6273 6699 6307
rect 6641 6267 6699 6273
rect 6730 6264 6736 6316
rect 6788 6304 6794 6316
rect 6914 6304 6920 6316
rect 6788 6276 6833 6304
rect 6875 6276 6920 6304
rect 6788 6264 6794 6276
rect 6914 6264 6920 6276
rect 6972 6264 6978 6316
rect 8386 6304 8392 6316
rect 8347 6276 8392 6304
rect 8386 6264 8392 6276
rect 8444 6264 8450 6316
rect 7466 6236 7472 6248
rect 6104 6208 7472 6236
rect 7466 6196 7472 6208
rect 7524 6196 7530 6248
rect 8680 6245 8708 6332
rect 9950 6304 9956 6316
rect 9911 6276 9956 6304
rect 9950 6264 9956 6276
rect 10008 6264 10014 6316
rect 10137 6307 10195 6313
rect 10137 6304 10149 6307
rect 10060 6276 10149 6304
rect 8665 6239 8723 6245
rect 8665 6205 8677 6239
rect 8711 6205 8723 6239
rect 9766 6236 9772 6248
rect 8665 6199 8723 6205
rect 8772 6208 9772 6236
rect 5261 6171 5319 6177
rect 5261 6168 5273 6171
rect 4724 6140 5273 6168
rect 5261 6137 5273 6140
rect 5307 6137 5319 6171
rect 5261 6131 5319 6137
rect 6270 6128 6276 6180
rect 6328 6168 6334 6180
rect 6549 6171 6607 6177
rect 6328 6140 6408 6168
rect 6328 6128 6334 6140
rect 2501 6103 2559 6109
rect 2501 6069 2513 6103
rect 2547 6100 2559 6103
rect 2958 6100 2964 6112
rect 2547 6072 2964 6100
rect 2547 6069 2559 6072
rect 2501 6063 2559 6069
rect 2958 6060 2964 6072
rect 3016 6060 3022 6112
rect 6380 6100 6408 6140
rect 6549 6137 6561 6171
rect 6595 6168 6607 6171
rect 8772 6168 8800 6208
rect 9766 6196 9772 6208
rect 9824 6196 9830 6248
rect 6595 6140 8800 6168
rect 6595 6137 6607 6140
rect 6549 6131 6607 6137
rect 6730 6100 6736 6112
rect 6380 6072 6736 6100
rect 6730 6060 6736 6072
rect 6788 6100 6794 6112
rect 10060 6100 10088 6276
rect 10137 6273 10149 6276
rect 10183 6273 10195 6307
rect 10137 6267 10195 6273
rect 10226 6264 10232 6316
rect 10284 6304 10290 6316
rect 10778 6304 10784 6316
rect 10284 6276 10329 6304
rect 10739 6276 10784 6304
rect 10284 6264 10290 6276
rect 10778 6264 10784 6276
rect 10836 6264 10842 6316
rect 10980 6304 11008 6412
rect 11149 6409 11161 6443
rect 11195 6440 11207 6443
rect 11238 6440 11244 6452
rect 11195 6412 11244 6440
rect 11195 6409 11207 6412
rect 11149 6403 11207 6409
rect 11238 6400 11244 6412
rect 11296 6400 11302 6452
rect 11514 6440 11520 6452
rect 11475 6412 11520 6440
rect 11514 6400 11520 6412
rect 11572 6400 11578 6452
rect 11609 6443 11667 6449
rect 11609 6409 11621 6443
rect 11655 6440 11667 6443
rect 11882 6440 11888 6452
rect 11655 6412 11888 6440
rect 11655 6409 11667 6412
rect 11609 6403 11667 6409
rect 11882 6400 11888 6412
rect 11940 6400 11946 6452
rect 13814 6400 13820 6452
rect 13872 6440 13878 6452
rect 14001 6443 14059 6449
rect 14001 6440 14013 6443
rect 13872 6412 14013 6440
rect 13872 6400 13878 6412
rect 14001 6409 14013 6412
rect 14047 6440 14059 6443
rect 14645 6443 14703 6449
rect 14047 6412 14320 6440
rect 14047 6409 14059 6412
rect 14001 6403 14059 6409
rect 11330 6332 11336 6384
rect 11388 6372 11394 6384
rect 11790 6372 11796 6384
rect 11388 6344 11796 6372
rect 11388 6332 11394 6344
rect 11790 6332 11796 6344
rect 11848 6372 11854 6384
rect 14292 6372 14320 6412
rect 14645 6409 14657 6443
rect 14691 6440 14703 6443
rect 14826 6440 14832 6452
rect 14691 6412 14832 6440
rect 14691 6409 14703 6412
rect 14645 6403 14703 6409
rect 14826 6400 14832 6412
rect 14884 6400 14890 6452
rect 16577 6443 16635 6449
rect 16577 6409 16589 6443
rect 16623 6440 16635 6443
rect 16623 6412 16804 6440
rect 16623 6409 16635 6412
rect 16577 6403 16635 6409
rect 15013 6375 15071 6381
rect 15013 6372 15025 6375
rect 11848 6344 12296 6372
rect 11848 6332 11854 6344
rect 12268 6313 12296 6344
rect 14292 6344 15025 6372
rect 12253 6307 12311 6313
rect 10980 6276 11744 6304
rect 10502 6196 10508 6248
rect 10560 6236 10566 6248
rect 11716 6245 11744 6276
rect 12253 6273 12265 6307
rect 12299 6273 12311 6307
rect 13814 6304 13820 6316
rect 13662 6276 13820 6304
rect 12253 6267 12311 6273
rect 13814 6264 13820 6276
rect 13872 6264 13878 6316
rect 14292 6313 14320 6344
rect 15013 6341 15025 6344
rect 15059 6372 15071 6375
rect 15470 6372 15476 6384
rect 15059 6344 15476 6372
rect 15059 6341 15071 6344
rect 15013 6335 15071 6341
rect 15470 6332 15476 6344
rect 15528 6332 15534 6384
rect 14277 6307 14335 6313
rect 14277 6273 14289 6307
rect 14323 6273 14335 6307
rect 14277 6267 14335 6273
rect 14737 6307 14795 6313
rect 14737 6273 14749 6307
rect 14783 6304 14795 6307
rect 15562 6304 15568 6316
rect 14783 6276 15568 6304
rect 14783 6273 14795 6276
rect 14737 6267 14795 6273
rect 10873 6239 10931 6245
rect 10873 6236 10885 6239
rect 10560 6208 10885 6236
rect 10560 6196 10566 6208
rect 10873 6205 10885 6208
rect 10919 6205 10931 6239
rect 10873 6199 10931 6205
rect 11701 6239 11759 6245
rect 11701 6205 11713 6239
rect 11747 6205 11759 6239
rect 11701 6199 11759 6205
rect 12529 6239 12587 6245
rect 12529 6205 12541 6239
rect 12575 6236 12587 6239
rect 12986 6236 12992 6248
rect 12575 6208 12992 6236
rect 12575 6205 12587 6208
rect 12529 6199 12587 6205
rect 12986 6196 12992 6208
rect 13044 6196 13050 6248
rect 14369 6239 14427 6245
rect 14369 6205 14381 6239
rect 14415 6236 14427 6239
rect 14752 6236 14780 6267
rect 15562 6264 15568 6276
rect 15620 6264 15626 6316
rect 16390 6304 16396 6316
rect 16351 6276 16396 6304
rect 16390 6264 16396 6276
rect 16448 6264 16454 6316
rect 16776 6304 16804 6412
rect 17770 6400 17776 6452
rect 17828 6440 17834 6452
rect 18463 6443 18521 6449
rect 18463 6440 18475 6443
rect 17828 6412 18475 6440
rect 17828 6400 17834 6412
rect 18463 6409 18475 6412
rect 18509 6409 18521 6443
rect 18463 6403 18521 6409
rect 17402 6332 17408 6384
rect 17460 6332 17466 6384
rect 17037 6307 17095 6313
rect 17037 6304 17049 6307
rect 16776 6276 17049 6304
rect 17037 6273 17049 6276
rect 17083 6273 17095 6307
rect 17037 6267 17095 6273
rect 14415 6208 14780 6236
rect 14829 6239 14887 6245
rect 14415 6205 14427 6208
rect 14369 6199 14427 6205
rect 14829 6205 14841 6239
rect 14875 6236 14887 6239
rect 14918 6236 14924 6248
rect 14875 6208 14924 6236
rect 14875 6205 14887 6208
rect 14829 6199 14887 6205
rect 14918 6196 14924 6208
rect 14976 6196 14982 6248
rect 16666 6236 16672 6248
rect 16627 6208 16672 6236
rect 16666 6196 16672 6208
rect 16724 6196 16730 6248
rect 11606 6168 11612 6180
rect 10198 6140 11612 6168
rect 10198 6100 10226 6140
rect 11606 6128 11612 6140
rect 11664 6128 11670 6180
rect 6788 6072 10226 6100
rect 11057 6103 11115 6109
rect 6788 6060 6794 6072
rect 11057 6069 11069 6103
rect 11103 6100 11115 6103
rect 11514 6100 11520 6112
rect 11103 6072 11520 6100
rect 11103 6069 11115 6072
rect 11057 6063 11115 6069
rect 11514 6060 11520 6072
rect 11572 6060 11578 6112
rect 14918 6100 14924 6112
rect 14879 6072 14924 6100
rect 14918 6060 14924 6072
rect 14976 6060 14982 6112
rect 0 6010 18860 6032
rect 0 5958 3110 6010
rect 3162 5958 3174 6010
rect 3226 5958 3238 6010
rect 3290 5958 3302 6010
rect 3354 5958 3366 6010
rect 3418 5958 6210 6010
rect 6262 5958 6274 6010
rect 6326 5958 6338 6010
rect 6390 5958 6402 6010
rect 6454 5958 6466 6010
rect 6518 5958 9310 6010
rect 9362 5958 9374 6010
rect 9426 5958 9438 6010
rect 9490 5958 9502 6010
rect 9554 5958 9566 6010
rect 9618 5958 12410 6010
rect 12462 5958 12474 6010
rect 12526 5958 12538 6010
rect 12590 5958 12602 6010
rect 12654 5958 12666 6010
rect 12718 5958 15510 6010
rect 15562 5958 15574 6010
rect 15626 5958 15638 6010
rect 15690 5958 15702 6010
rect 15754 5958 15766 6010
rect 15818 5958 18860 6010
rect 0 5936 18860 5958
rect 3510 5856 3516 5908
rect 3568 5896 3574 5908
rect 4479 5899 4537 5905
rect 4479 5896 4491 5899
rect 3568 5868 4491 5896
rect 3568 5856 3574 5868
rect 4479 5865 4491 5868
rect 4525 5865 4537 5899
rect 4479 5859 4537 5865
rect 6914 5856 6920 5908
rect 6972 5896 6978 5908
rect 7607 5899 7665 5905
rect 7607 5896 7619 5899
rect 6972 5868 7619 5896
rect 6972 5856 6978 5868
rect 7607 5865 7619 5868
rect 7653 5865 7665 5899
rect 7607 5859 7665 5865
rect 8202 5856 8208 5908
rect 8260 5896 8266 5908
rect 9950 5896 9956 5908
rect 8260 5868 9956 5896
rect 8260 5856 8266 5868
rect 9950 5856 9956 5868
rect 10008 5896 10014 5908
rect 10045 5899 10103 5905
rect 10045 5896 10057 5899
rect 10008 5868 10057 5896
rect 10008 5856 10014 5868
rect 10045 5865 10057 5868
rect 10091 5865 10103 5899
rect 12986 5896 12992 5908
rect 12947 5868 12992 5896
rect 10045 5859 10103 5865
rect 12986 5856 12992 5868
rect 13044 5856 13050 5908
rect 15105 5899 15163 5905
rect 15105 5865 15117 5899
rect 15151 5896 15163 5899
rect 16681 5899 16739 5905
rect 16681 5896 16693 5899
rect 15151 5868 16693 5896
rect 15151 5865 15163 5868
rect 15105 5859 15163 5865
rect 16681 5865 16693 5868
rect 16727 5865 16739 5899
rect 16681 5859 16739 5865
rect 15378 5828 15384 5840
rect 12406 5800 15384 5828
rect 290 5720 296 5772
rect 348 5760 354 5772
rect 4062 5760 4068 5772
rect 348 5732 4068 5760
rect 348 5720 354 5732
rect 2332 5701 2360 5732
rect 4062 5720 4068 5732
rect 4120 5760 4126 5772
rect 5813 5763 5871 5769
rect 5813 5760 5825 5763
rect 4120 5732 5825 5760
rect 4120 5720 4126 5732
rect 5813 5729 5825 5732
rect 5859 5760 5871 5763
rect 5994 5760 6000 5772
rect 5859 5732 6000 5760
rect 5859 5729 5871 5732
rect 5813 5723 5871 5729
rect 5994 5720 6000 5732
rect 6052 5720 6058 5772
rect 6086 5720 6092 5772
rect 6144 5760 6150 5772
rect 6181 5763 6239 5769
rect 6181 5760 6193 5763
rect 6144 5732 6193 5760
rect 6144 5720 6150 5732
rect 6181 5729 6193 5732
rect 6227 5729 6239 5763
rect 12406 5760 12434 5800
rect 15378 5788 15384 5800
rect 15436 5788 15442 5840
rect 6181 5723 6239 5729
rect 9876 5732 12434 5760
rect 14829 5763 14887 5769
rect 2317 5695 2375 5701
rect 2317 5661 2329 5695
rect 2363 5661 2375 5695
rect 2317 5655 2375 5661
rect 2409 5695 2467 5701
rect 2409 5661 2421 5695
rect 2455 5692 2467 5695
rect 2685 5695 2743 5701
rect 2685 5692 2697 5695
rect 2455 5664 2697 5692
rect 2455 5661 2467 5664
rect 2409 5655 2467 5661
rect 2685 5661 2697 5664
rect 2731 5661 2743 5695
rect 2685 5655 2743 5661
rect 2958 5652 2964 5704
rect 3016 5692 3022 5704
rect 9876 5701 9904 5732
rect 14829 5729 14841 5763
rect 14875 5760 14887 5763
rect 14918 5760 14924 5772
rect 14875 5732 14924 5760
rect 14875 5729 14887 5732
rect 14829 5723 14887 5729
rect 14918 5720 14924 5732
rect 14976 5720 14982 5772
rect 15194 5760 15200 5772
rect 15155 5732 15200 5760
rect 15194 5720 15200 5732
rect 15252 5720 15258 5772
rect 16666 5720 16672 5772
rect 16724 5760 16730 5772
rect 16945 5763 17003 5769
rect 16945 5760 16957 5763
rect 16724 5732 16957 5760
rect 16724 5720 16730 5732
rect 16945 5729 16957 5732
rect 16991 5729 17003 5763
rect 16945 5723 17003 5729
rect 3053 5695 3111 5701
rect 3053 5692 3065 5695
rect 3016 5664 3065 5692
rect 3016 5652 3022 5664
rect 3053 5661 3065 5664
rect 3099 5661 3111 5695
rect 3053 5655 3111 5661
rect 9861 5695 9919 5701
rect 9861 5661 9873 5695
rect 9907 5661 9919 5695
rect 9861 5655 9919 5661
rect 11790 5652 11796 5704
rect 11848 5692 11854 5704
rect 13170 5692 13176 5704
rect 11848 5664 11893 5692
rect 13131 5664 13176 5692
rect 11848 5652 11854 5664
rect 13170 5652 13176 5664
rect 13228 5652 13234 5704
rect 14737 5695 14795 5701
rect 14737 5661 14749 5695
rect 14783 5692 14795 5695
rect 15212 5692 15240 5720
rect 18506 5692 18512 5704
rect 14783 5664 15240 5692
rect 18467 5664 18512 5692
rect 14783 5661 14795 5664
rect 14737 5655 14795 5661
rect 18506 5652 18512 5664
rect 18564 5652 18570 5704
rect 3786 5584 3792 5636
rect 3844 5584 3850 5636
rect 11514 5624 11520 5636
rect 2406 5516 2412 5568
rect 2464 5556 2470 5568
rect 3804 5556 3832 5584
rect 6564 5556 6592 5610
rect 8312 5596 9674 5624
rect 8312 5568 8340 5596
rect 8294 5556 8300 5568
rect 2464 5528 8300 5556
rect 2464 5516 2470 5528
rect 8294 5516 8300 5528
rect 8352 5516 8358 5568
rect 8573 5559 8631 5565
rect 8573 5525 8585 5559
rect 8619 5556 8631 5559
rect 8846 5556 8852 5568
rect 8619 5528 8852 5556
rect 8619 5525 8631 5528
rect 8573 5519 8631 5525
rect 8846 5516 8852 5528
rect 8904 5516 8910 5568
rect 9646 5556 9674 5596
rect 11072 5556 11100 5610
rect 11475 5596 11520 5624
rect 11514 5584 11520 5596
rect 11572 5584 11578 5636
rect 15102 5584 15108 5636
rect 15160 5624 15166 5636
rect 15160 5596 15502 5624
rect 15160 5584 15166 5596
rect 13814 5556 13820 5568
rect 9646 5528 13820 5556
rect 13814 5516 13820 5528
rect 13872 5516 13878 5568
rect 18230 5516 18236 5568
rect 18288 5556 18294 5568
rect 18325 5559 18383 5565
rect 18325 5556 18337 5559
rect 18288 5528 18337 5556
rect 18288 5516 18294 5528
rect 18325 5525 18337 5528
rect 18371 5525 18383 5559
rect 18325 5519 18383 5525
rect 0 5466 18860 5488
rect 0 5414 4660 5466
rect 4712 5414 4724 5466
rect 4776 5414 4788 5466
rect 4840 5414 4852 5466
rect 4904 5414 4916 5466
rect 4968 5414 7760 5466
rect 7812 5414 7824 5466
rect 7876 5414 7888 5466
rect 7940 5414 7952 5466
rect 8004 5414 8016 5466
rect 8068 5414 10860 5466
rect 10912 5414 10924 5466
rect 10976 5414 10988 5466
rect 11040 5414 11052 5466
rect 11104 5414 11116 5466
rect 11168 5414 13960 5466
rect 14012 5414 14024 5466
rect 14076 5414 14088 5466
rect 14140 5414 14152 5466
rect 14204 5414 14216 5466
rect 14268 5414 17060 5466
rect 17112 5414 17124 5466
rect 17176 5414 17188 5466
rect 17240 5414 17252 5466
rect 17304 5414 17316 5466
rect 17368 5414 18860 5466
rect 0 5392 18860 5414
rect 9309 5355 9367 5361
rect 9309 5352 9321 5355
rect 8772 5324 9321 5352
rect 7466 5244 7472 5296
rect 7524 5284 7530 5296
rect 7524 5256 8064 5284
rect 7524 5244 7530 5256
rect 5074 5176 5080 5228
rect 5132 5216 5138 5228
rect 5721 5219 5779 5225
rect 5721 5216 5733 5219
rect 5132 5188 5733 5216
rect 5132 5176 5138 5188
rect 5721 5185 5733 5188
rect 5767 5185 5779 5219
rect 5721 5179 5779 5185
rect 6914 5176 6920 5228
rect 6972 5216 6978 5228
rect 7561 5219 7619 5225
rect 7561 5216 7573 5219
rect 6972 5188 7573 5216
rect 6972 5176 6978 5188
rect 7561 5185 7573 5188
rect 7607 5185 7619 5219
rect 7561 5179 7619 5185
rect 7745 5219 7803 5225
rect 7745 5185 7757 5219
rect 7791 5216 7803 5219
rect 7834 5216 7840 5228
rect 7791 5188 7840 5216
rect 7791 5185 7803 5188
rect 7745 5179 7803 5185
rect 5813 5015 5871 5021
rect 5813 4981 5825 5015
rect 5859 5012 5871 5015
rect 6914 5012 6920 5024
rect 5859 4984 6920 5012
rect 5859 4981 5871 4984
rect 5813 4975 5871 4981
rect 6914 4972 6920 4984
rect 6972 4972 6978 5024
rect 7576 5012 7604 5179
rect 7834 5176 7840 5188
rect 7892 5176 7898 5228
rect 8036 5225 8064 5256
rect 8202 5244 8208 5296
rect 8260 5284 8266 5296
rect 8772 5293 8800 5324
rect 9309 5321 9321 5324
rect 9355 5321 9367 5355
rect 9309 5315 9367 5321
rect 10594 5312 10600 5364
rect 10652 5352 10658 5364
rect 10873 5355 10931 5361
rect 10873 5352 10885 5355
rect 10652 5324 10885 5352
rect 10652 5312 10658 5324
rect 10873 5321 10885 5324
rect 10919 5321 10931 5355
rect 17402 5352 17408 5364
rect 10873 5315 10931 5321
rect 17052 5324 17408 5352
rect 8573 5287 8631 5293
rect 8573 5284 8585 5287
rect 8260 5256 8585 5284
rect 8260 5244 8266 5256
rect 8573 5253 8585 5256
rect 8619 5253 8631 5287
rect 8573 5247 8631 5253
rect 8757 5287 8815 5293
rect 8757 5253 8769 5287
rect 8803 5253 8815 5287
rect 9033 5287 9091 5293
rect 9033 5284 9045 5287
rect 8757 5247 8815 5253
rect 8862 5256 9045 5284
rect 8862 5225 8890 5256
rect 9033 5253 9045 5256
rect 9079 5253 9091 5287
rect 9033 5247 9091 5253
rect 9122 5244 9128 5296
rect 9180 5284 9186 5296
rect 10781 5287 10839 5293
rect 10781 5284 10793 5287
rect 9180 5256 10793 5284
rect 9180 5244 9186 5256
rect 10781 5253 10793 5256
rect 10827 5253 10839 5287
rect 10781 5247 10839 5253
rect 13814 5244 13820 5296
rect 13872 5284 13878 5296
rect 15102 5284 15108 5296
rect 13872 5256 15108 5284
rect 13872 5244 13878 5256
rect 15102 5244 15108 5256
rect 15160 5244 15166 5296
rect 16298 5244 16304 5296
rect 16356 5284 16362 5296
rect 17052 5284 17080 5324
rect 17402 5312 17408 5324
rect 17460 5312 17466 5364
rect 16356 5270 17080 5284
rect 16356 5256 17066 5270
rect 16356 5244 16362 5256
rect 17954 5244 17960 5296
rect 18012 5284 18018 5296
rect 18012 5256 18552 5284
rect 18012 5244 18018 5256
rect 8021 5219 8079 5225
rect 8021 5185 8033 5219
rect 8067 5185 8079 5219
rect 8021 5179 8079 5185
rect 8847 5219 8905 5225
rect 8847 5185 8859 5219
rect 8893 5185 8905 5219
rect 9217 5219 9275 5225
rect 8847 5179 8905 5185
rect 8938 5166 8944 5218
rect 8996 5206 9002 5218
rect 8996 5178 9041 5206
rect 9217 5185 9229 5219
rect 9263 5185 9275 5219
rect 9766 5216 9772 5228
rect 9727 5188 9772 5216
rect 9217 5179 9275 5185
rect 8996 5166 9002 5178
rect 7653 5151 7711 5157
rect 7653 5117 7665 5151
rect 7699 5148 7711 5151
rect 7929 5151 7987 5157
rect 7929 5148 7941 5151
rect 7699 5120 7941 5148
rect 7699 5117 7711 5120
rect 7653 5111 7711 5117
rect 7929 5117 7941 5120
rect 7975 5117 7987 5151
rect 8386 5148 8392 5160
rect 8347 5120 8392 5148
rect 7929 5111 7987 5117
rect 8386 5108 8392 5120
rect 8444 5108 8450 5160
rect 9232 5148 9260 5179
rect 9766 5176 9772 5188
rect 9824 5176 9830 5228
rect 18524 5225 18552 5256
rect 12345 5219 12403 5225
rect 12345 5185 12357 5219
rect 12391 5185 12403 5219
rect 12345 5179 12403 5185
rect 18509 5219 18567 5225
rect 18509 5185 18521 5219
rect 18555 5185 18567 5219
rect 18509 5179 18567 5185
rect 12250 5148 12256 5160
rect 9232 5120 9444 5148
rect 12211 5120 12256 5148
rect 8478 5040 8484 5092
rect 8536 5080 8542 5092
rect 8665 5083 8723 5089
rect 8665 5080 8677 5083
rect 8536 5052 8677 5080
rect 8536 5040 8542 5052
rect 8665 5049 8677 5052
rect 8711 5049 8723 5083
rect 8665 5043 8723 5049
rect 9416 5012 9444 5120
rect 12250 5108 12256 5120
rect 12308 5108 12314 5160
rect 12360 5080 12388 5179
rect 12713 5151 12771 5157
rect 12713 5117 12725 5151
rect 12759 5148 12771 5151
rect 14277 5151 14335 5157
rect 14277 5148 14289 5151
rect 12759 5120 14289 5148
rect 12759 5117 12771 5120
rect 12713 5111 12771 5117
rect 14277 5117 14289 5120
rect 14323 5117 14335 5151
rect 14550 5148 14556 5160
rect 14511 5120 14556 5148
rect 14277 5111 14335 5117
rect 14550 5108 14556 5120
rect 14608 5108 14614 5160
rect 18230 5148 18236 5160
rect 18191 5120 18236 5148
rect 18230 5108 18236 5120
rect 18288 5108 18294 5160
rect 12802 5080 12808 5092
rect 12360 5052 12808 5080
rect 12802 5040 12808 5052
rect 12860 5040 12866 5092
rect 7576 4984 9444 5012
rect 9953 5015 10011 5021
rect 9953 4981 9965 5015
rect 9999 5012 10011 5015
rect 10042 5012 10048 5024
rect 9999 4984 10048 5012
rect 9999 4981 10011 4984
rect 9953 4975 10011 4981
rect 10042 4972 10048 4984
rect 10100 4972 10106 5024
rect 16761 5015 16819 5021
rect 16761 4981 16773 5015
rect 16807 5012 16819 5015
rect 17678 5012 17684 5024
rect 16807 4984 17684 5012
rect 16807 4981 16819 4984
rect 16761 4975 16819 4981
rect 17678 4972 17684 4984
rect 17736 4972 17742 5024
rect 0 4922 18860 4944
rect 0 4870 3110 4922
rect 3162 4870 3174 4922
rect 3226 4870 3238 4922
rect 3290 4870 3302 4922
rect 3354 4870 3366 4922
rect 3418 4870 6210 4922
rect 6262 4870 6274 4922
rect 6326 4870 6338 4922
rect 6390 4870 6402 4922
rect 6454 4870 6466 4922
rect 6518 4870 9310 4922
rect 9362 4870 9374 4922
rect 9426 4870 9438 4922
rect 9490 4870 9502 4922
rect 9554 4870 9566 4922
rect 9618 4870 12410 4922
rect 12462 4870 12474 4922
rect 12526 4870 12538 4922
rect 12590 4870 12602 4922
rect 12654 4870 12666 4922
rect 12718 4870 15510 4922
rect 15562 4870 15574 4922
rect 15626 4870 15638 4922
rect 15690 4870 15702 4922
rect 15754 4870 15766 4922
rect 15818 4870 18860 4922
rect 0 4848 18860 4870
rect 5074 4808 5080 4820
rect 5035 4780 5080 4808
rect 5074 4768 5080 4780
rect 5132 4768 5138 4820
rect 9858 4768 9864 4820
rect 9916 4768 9922 4820
rect 12250 4808 12256 4820
rect 12211 4780 12256 4808
rect 12250 4768 12256 4780
rect 12308 4768 12314 4820
rect 14093 4811 14151 4817
rect 14093 4777 14105 4811
rect 14139 4808 14151 4811
rect 14458 4808 14464 4820
rect 14139 4780 14464 4808
rect 14139 4777 14151 4780
rect 14093 4771 14151 4777
rect 14458 4768 14464 4780
rect 14516 4768 14522 4820
rect 9876 4740 9904 4768
rect 9692 4712 9904 4740
rect 8754 4672 8760 4684
rect 2332 4644 6868 4672
rect 2332 4616 2360 4644
rect 2314 4604 2320 4616
rect 2227 4576 2320 4604
rect 2314 4564 2320 4576
rect 2372 4564 2378 4616
rect 2409 4607 2467 4613
rect 2409 4573 2421 4607
rect 2455 4604 2467 4607
rect 2685 4607 2743 4613
rect 2685 4604 2697 4607
rect 2455 4576 2697 4604
rect 2455 4573 2467 4576
rect 2409 4567 2467 4573
rect 2685 4573 2697 4576
rect 2731 4573 2743 4607
rect 3050 4604 3056 4616
rect 3011 4576 3056 4604
rect 2685 4567 2743 4573
rect 3050 4564 3056 4576
rect 3108 4564 3114 4616
rect 4479 4607 4537 4613
rect 4479 4573 4491 4607
rect 4525 4604 4537 4607
rect 4801 4607 4859 4613
rect 4801 4604 4813 4607
rect 4525 4576 4813 4604
rect 4525 4573 4537 4576
rect 4479 4567 4537 4573
rect 4801 4573 4813 4576
rect 4847 4604 4859 4607
rect 4982 4604 4988 4616
rect 4847 4576 4988 4604
rect 4847 4573 4859 4576
rect 4801 4567 4859 4573
rect 4982 4564 4988 4576
rect 5040 4564 5046 4616
rect 6840 4613 6868 4644
rect 7208 4644 8760 4672
rect 7208 4613 7236 4644
rect 8754 4632 8760 4644
rect 8812 4632 8818 4684
rect 9692 4681 9720 4712
rect 9677 4675 9735 4681
rect 9677 4641 9689 4675
rect 9723 4641 9735 4675
rect 9677 4635 9735 4641
rect 9769 4675 9827 4681
rect 9769 4641 9781 4675
rect 9815 4672 9827 4675
rect 10594 4672 10600 4684
rect 9815 4644 10600 4672
rect 9815 4641 9827 4644
rect 9769 4635 9827 4641
rect 10594 4632 10600 4644
rect 10652 4632 10658 4684
rect 12066 4632 12072 4684
rect 12124 4672 12130 4684
rect 12124 4644 12468 4672
rect 12124 4632 12130 4644
rect 6825 4607 6883 4613
rect 6825 4573 6837 4607
rect 6871 4604 6883 4607
rect 7193 4607 7251 4613
rect 6871 4576 7052 4604
rect 6871 4573 6883 4576
rect 6825 4567 6883 4573
rect 7024 4545 7052 4576
rect 7193 4573 7205 4607
rect 7239 4573 7251 4607
rect 7193 4567 7251 4573
rect 7650 4564 7656 4616
rect 7708 4604 7714 4616
rect 7837 4607 7895 4613
rect 7837 4604 7849 4607
rect 7708 4576 7849 4604
rect 7708 4564 7714 4576
rect 7837 4573 7849 4576
rect 7883 4573 7895 4607
rect 8202 4604 8208 4616
rect 8163 4576 8208 4604
rect 7837 4567 7895 4573
rect 8202 4564 8208 4576
rect 8260 4564 8266 4616
rect 9030 4604 9036 4616
rect 8956 4576 9036 4604
rect 6549 4539 6607 4545
rect 4094 4522 5382 4536
rect 4080 4508 5382 4522
rect 2406 4428 2412 4480
rect 2464 4468 2470 4480
rect 4080 4468 4108 4508
rect 6549 4505 6561 4539
rect 6595 4505 6607 4539
rect 6549 4499 6607 4505
rect 7009 4539 7067 4545
rect 7009 4505 7021 4539
rect 7055 4536 7067 4539
rect 7374 4536 7380 4548
rect 7055 4508 7380 4536
rect 7055 4505 7067 4508
rect 7009 4499 7067 4505
rect 2464 4440 4108 4468
rect 4709 4471 4767 4477
rect 2464 4428 2470 4440
rect 4709 4437 4721 4471
rect 4755 4468 4767 4471
rect 5166 4468 5172 4480
rect 4755 4440 5172 4468
rect 4755 4437 4767 4440
rect 4709 4431 4767 4437
rect 5166 4428 5172 4440
rect 5224 4428 5230 4480
rect 5626 4428 5632 4480
rect 5684 4468 5690 4480
rect 6564 4468 6592 4499
rect 7374 4496 7380 4508
rect 7432 4536 7438 4548
rect 7668 4536 7696 4564
rect 7432 4508 7696 4536
rect 7432 4496 7438 4508
rect 5684 4440 6592 4468
rect 7668 4468 7696 4508
rect 8478 4496 8484 4548
rect 8536 4536 8542 4548
rect 8536 4530 8602 4536
rect 8956 4530 8984 4576
rect 9030 4564 9036 4576
rect 9088 4604 9094 4616
rect 12440 4613 12468 4644
rect 14550 4632 14556 4684
rect 14608 4672 14614 4684
rect 15841 4675 15899 4681
rect 15841 4672 15853 4675
rect 14608 4644 15853 4672
rect 14608 4632 14614 4644
rect 15841 4641 15853 4644
rect 15887 4641 15899 4675
rect 17678 4672 17684 4684
rect 17639 4644 17684 4672
rect 15841 4635 15899 4641
rect 17678 4632 17684 4644
rect 17736 4632 17742 4684
rect 12345 4607 12403 4613
rect 9088 4592 9674 4604
rect 9088 4576 9634 4592
rect 9088 4564 9094 4576
rect 9628 4540 9634 4576
rect 9686 4540 9692 4592
rect 12345 4573 12357 4607
rect 12391 4573 12403 4607
rect 12345 4567 12403 4573
rect 12431 4607 12489 4613
rect 12431 4573 12443 4607
rect 12477 4573 12489 4607
rect 12431 4567 12489 4573
rect 12535 4607 12593 4613
rect 12535 4573 12547 4607
rect 12581 4573 12593 4607
rect 12535 4567 12593 4573
rect 12713 4607 12771 4613
rect 12713 4573 12725 4607
rect 12759 4604 12771 4607
rect 12802 4604 12808 4616
rect 12759 4576 12808 4604
rect 12759 4573 12771 4576
rect 12713 4567 12771 4573
rect 10042 4536 10048 4548
rect 8536 4508 8984 4530
rect 10003 4508 10048 4536
rect 8536 4496 8542 4508
rect 8588 4502 8984 4508
rect 10042 4496 10048 4508
rect 10100 4496 10106 4548
rect 11330 4536 11336 4548
rect 11270 4508 11336 4536
rect 11330 4496 11336 4508
rect 11388 4496 11394 4548
rect 11422 4496 11428 4548
rect 11480 4536 11486 4548
rect 12161 4539 12219 4545
rect 12161 4536 12173 4539
rect 11480 4508 12173 4536
rect 11480 4496 11486 4508
rect 12161 4505 12173 4508
rect 12207 4536 12219 4539
rect 12250 4536 12256 4548
rect 12207 4508 12256 4536
rect 12207 4505 12219 4508
rect 12161 4499 12219 4505
rect 12250 4496 12256 4508
rect 12308 4496 12314 4548
rect 12360 4536 12388 4567
rect 12550 4536 12578 4567
rect 12802 4564 12808 4576
rect 12860 4564 12866 4616
rect 17954 4564 17960 4616
rect 18012 4604 18018 4616
rect 18506 4604 18512 4616
rect 18012 4576 18057 4604
rect 18467 4576 18512 4604
rect 18012 4564 18018 4576
rect 18506 4564 18512 4576
rect 18564 4564 18570 4616
rect 12360 4508 12578 4536
rect 9122 4468 9128 4480
rect 7668 4440 9128 4468
rect 5684 4428 5690 4440
rect 9122 4428 9128 4440
rect 9180 4428 9186 4480
rect 11514 4468 11520 4480
rect 11475 4440 11520 4468
rect 11514 4428 11520 4440
rect 11572 4468 11578 4480
rect 12360 4468 12388 4508
rect 15102 4496 15108 4548
rect 15160 4496 15166 4548
rect 15565 4539 15623 4545
rect 15565 4505 15577 4539
rect 15611 4505 15623 4539
rect 15930 4536 15936 4548
rect 15891 4508 15936 4536
rect 15565 4499 15623 4505
rect 12618 4468 12624 4480
rect 11572 4440 12388 4468
rect 12579 4440 12624 4468
rect 11572 4428 11578 4440
rect 12618 4428 12624 4440
rect 12676 4428 12682 4480
rect 15580 4468 15608 4499
rect 15930 4496 15936 4508
rect 15988 4496 15994 4548
rect 16298 4496 16304 4548
rect 16356 4536 16362 4548
rect 18230 4536 18236 4548
rect 16356 4508 16514 4536
rect 17328 4508 18236 4536
rect 16356 4496 16362 4508
rect 17328 4468 17356 4508
rect 18230 4496 18236 4508
rect 18288 4496 18294 4548
rect 15580 4440 17356 4468
rect 17402 4428 17408 4480
rect 17460 4468 17466 4480
rect 18325 4471 18383 4477
rect 18325 4468 18337 4471
rect 17460 4440 18337 4468
rect 17460 4428 17466 4440
rect 18325 4437 18337 4440
rect 18371 4437 18383 4471
rect 18325 4431 18383 4437
rect 0 4378 18860 4400
rect 0 4326 4660 4378
rect 4712 4326 4724 4378
rect 4776 4326 4788 4378
rect 4840 4326 4852 4378
rect 4904 4326 4916 4378
rect 4968 4326 7760 4378
rect 7812 4326 7824 4378
rect 7876 4326 7888 4378
rect 7940 4326 7952 4378
rect 8004 4326 8016 4378
rect 8068 4326 10860 4378
rect 10912 4326 10924 4378
rect 10976 4326 10988 4378
rect 11040 4326 11052 4378
rect 11104 4326 11116 4378
rect 11168 4326 13960 4378
rect 14012 4326 14024 4378
rect 14076 4326 14088 4378
rect 14140 4326 14152 4378
rect 14204 4326 14216 4378
rect 14268 4326 17060 4378
rect 17112 4326 17124 4378
rect 17176 4326 17188 4378
rect 17240 4326 17252 4378
rect 17304 4326 17316 4378
rect 17368 4326 18860 4378
rect 0 4304 18860 4326
rect 3050 4224 3056 4276
rect 3108 4264 3114 4276
rect 3237 4267 3295 4273
rect 3237 4264 3249 4267
rect 3108 4236 3249 4264
rect 3108 4224 3114 4236
rect 3237 4233 3249 4236
rect 3283 4233 3295 4267
rect 3237 4227 3295 4233
rect 8021 4267 8079 4273
rect 8021 4233 8033 4267
rect 8067 4264 8079 4267
rect 8202 4264 8208 4276
rect 8067 4236 8208 4264
rect 8067 4233 8079 4236
rect 8021 4227 8079 4233
rect 8202 4224 8208 4236
rect 8260 4224 8266 4276
rect 8757 4267 8815 4273
rect 8757 4233 8769 4267
rect 8803 4264 8815 4267
rect 9217 4267 9275 4273
rect 9217 4264 9229 4267
rect 8803 4236 9229 4264
rect 8803 4233 8815 4236
rect 8757 4227 8815 4233
rect 9217 4233 9229 4236
rect 9263 4233 9275 4267
rect 9217 4227 9275 4233
rect 9766 4224 9772 4276
rect 9824 4264 9830 4276
rect 10413 4267 10471 4273
rect 10413 4264 10425 4267
rect 9824 4236 10425 4264
rect 9824 4224 9830 4236
rect 10413 4233 10425 4236
rect 10459 4233 10471 4267
rect 10413 4227 10471 4233
rect 10781 4267 10839 4273
rect 10781 4233 10793 4267
rect 10827 4264 10839 4267
rect 11241 4267 11299 4273
rect 11241 4264 11253 4267
rect 10827 4236 11253 4264
rect 10827 4233 10839 4236
rect 10781 4227 10839 4233
rect 11241 4233 11253 4236
rect 11287 4233 11299 4267
rect 15930 4264 15936 4276
rect 11241 4227 11299 4233
rect 11624 4236 15936 4264
rect 11624 4208 11652 4236
rect 15930 4224 15936 4236
rect 15988 4264 15994 4276
rect 15988 4236 16344 4264
rect 15988 4224 15994 4236
rect 4982 4196 4988 4208
rect 4895 4168 4988 4196
rect 4908 4137 4936 4168
rect 4982 4156 4988 4168
rect 5040 4196 5046 4208
rect 5442 4196 5448 4208
rect 5040 4168 5448 4196
rect 5040 4156 5046 4168
rect 5442 4156 5448 4168
rect 5500 4156 5506 4208
rect 8938 4156 8944 4208
rect 8996 4196 9002 4208
rect 9585 4199 9643 4205
rect 9585 4196 9597 4199
rect 8996 4168 9597 4196
rect 8996 4156 9002 4168
rect 9585 4165 9597 4168
rect 9631 4165 9643 4199
rect 11606 4196 11612 4208
rect 11567 4168 11612 4196
rect 9585 4159 9643 4165
rect 11606 4156 11612 4168
rect 11664 4156 11670 4208
rect 16316 4205 16344 4236
rect 16301 4199 16359 4205
rect 12084 4168 12572 4196
rect 12084 4140 12112 4168
rect 3513 4131 3571 4137
rect 3513 4097 3525 4131
rect 3559 4097 3571 4131
rect 3513 4091 3571 4097
rect 4893 4131 4951 4137
rect 4893 4097 4905 4131
rect 4939 4097 4951 4131
rect 5074 4128 5080 4140
rect 5035 4100 5080 4128
rect 4893 4091 4951 4097
rect 3237 4063 3295 4069
rect 3237 4029 3249 4063
rect 3283 4029 3295 4063
rect 3528 4060 3556 4091
rect 5074 4088 5080 4100
rect 5132 4088 5138 4140
rect 5166 4088 5172 4140
rect 5224 4128 5230 4140
rect 6733 4131 6791 4137
rect 6733 4128 6745 4131
rect 5224 4100 6745 4128
rect 5224 4088 5230 4100
rect 6733 4097 6745 4100
rect 6779 4097 6791 4131
rect 6914 4128 6920 4140
rect 6875 4100 6920 4128
rect 6733 4091 6791 4097
rect 6914 4088 6920 4100
rect 6972 4088 6978 4140
rect 7193 4131 7251 4137
rect 7193 4097 7205 4131
rect 7239 4097 7251 4131
rect 7466 4128 7472 4140
rect 7427 4100 7472 4128
rect 7193 4091 7251 4097
rect 5184 4060 5212 4088
rect 3528 4032 5212 4060
rect 6365 4063 6423 4069
rect 3237 4023 3295 4029
rect 6365 4029 6377 4063
rect 6411 4060 6423 4063
rect 6546 4060 6552 4072
rect 6411 4032 6552 4060
rect 6411 4029 6423 4032
rect 6365 4023 6423 4029
rect 3252 3992 3280 4023
rect 6546 4020 6552 4032
rect 6604 4020 6610 4072
rect 6638 4020 6644 4072
rect 6696 4060 6702 4072
rect 7098 4060 7104 4072
rect 6696 4032 6741 4060
rect 7059 4032 7104 4060
rect 6696 4020 6702 4032
rect 7098 4020 7104 4032
rect 7156 4020 7162 4072
rect 3970 3992 3976 4004
rect 3252 3964 3976 3992
rect 3970 3952 3976 3964
rect 4028 3952 4034 4004
rect 4522 3952 4528 4004
rect 4580 3992 4586 4004
rect 5902 3992 5908 4004
rect 4580 3964 5908 3992
rect 4580 3952 4586 3964
rect 5902 3952 5908 3964
rect 5960 3952 5966 4004
rect 7208 3992 7236 4091
rect 7466 4088 7472 4100
rect 7524 4088 7530 4140
rect 7837 4131 7895 4137
rect 7837 4097 7849 4131
rect 7883 4128 7895 4131
rect 8849 4131 8907 4137
rect 7883 4100 8432 4128
rect 7883 4097 7895 4100
rect 7837 4091 7895 4097
rect 8404 4001 8432 4100
rect 8849 4097 8861 4131
rect 8895 4128 8907 4131
rect 9766 4128 9772 4140
rect 8895 4100 9772 4128
rect 8895 4097 8907 4100
rect 8849 4091 8907 4097
rect 9766 4088 9772 4100
rect 9824 4088 9830 4140
rect 10778 4128 10784 4140
rect 9876 4100 10784 4128
rect 8754 4020 8760 4072
rect 8812 4060 8818 4072
rect 8941 4063 8999 4069
rect 8941 4060 8953 4063
rect 8812 4032 8953 4060
rect 8812 4020 8818 4032
rect 8941 4029 8953 4032
rect 8987 4029 8999 4063
rect 9674 4060 9680 4072
rect 9635 4032 9680 4060
rect 8941 4023 8999 4029
rect 6840 3964 7236 3992
rect 8389 3995 8447 4001
rect 6840 3936 6868 3964
rect 8389 3961 8401 3995
rect 8435 3961 8447 3995
rect 8389 3955 8447 3961
rect 3421 3927 3479 3933
rect 3421 3893 3433 3927
rect 3467 3924 3479 3927
rect 3510 3924 3516 3936
rect 3467 3896 3516 3924
rect 3467 3893 3479 3896
rect 3421 3887 3479 3893
rect 3510 3884 3516 3896
rect 3568 3884 3574 3936
rect 4893 3927 4951 3933
rect 4893 3893 4905 3927
rect 4939 3924 4951 3927
rect 5534 3924 5540 3936
rect 4939 3896 5540 3924
rect 4939 3893 4951 3896
rect 4893 3887 4951 3893
rect 5534 3884 5540 3896
rect 5592 3884 5598 3936
rect 6822 3924 6828 3936
rect 6783 3896 6828 3924
rect 6822 3884 6828 3896
rect 6880 3884 6886 3936
rect 8956 3924 8984 4023
rect 9674 4020 9680 4032
rect 9732 4020 9738 4072
rect 9876 4069 9904 4100
rect 10778 4088 10784 4100
rect 10836 4088 10842 4140
rect 10870 4088 10876 4140
rect 10928 4128 10934 4140
rect 11514 4128 11520 4140
rect 10928 4100 11520 4128
rect 10928 4088 10934 4100
rect 11514 4088 11520 4100
rect 11572 4088 11578 4140
rect 12066 4128 12072 4140
rect 12027 4100 12072 4128
rect 12066 4088 12072 4100
rect 12124 4088 12130 4140
rect 12253 4131 12311 4137
rect 12253 4097 12265 4131
rect 12299 4097 12311 4131
rect 12253 4091 12311 4097
rect 9861 4063 9919 4069
rect 9861 4029 9873 4063
rect 9907 4029 9919 4063
rect 10965 4063 11023 4069
rect 10965 4060 10977 4063
rect 9861 4023 9919 4029
rect 10428 4032 10977 4060
rect 10428 3924 10456 4032
rect 10965 4029 10977 4032
rect 11011 4060 11023 4063
rect 11422 4060 11428 4072
rect 11011 4032 11428 4060
rect 11011 4029 11023 4032
rect 10965 4023 11023 4029
rect 11422 4020 11428 4032
rect 11480 4020 11486 4072
rect 11698 4060 11704 4072
rect 11659 4032 11704 4060
rect 11698 4020 11704 4032
rect 11756 4020 11762 4072
rect 11793 4063 11851 4069
rect 11793 4029 11805 4063
rect 11839 4029 11851 4063
rect 11793 4023 11851 4029
rect 10778 3952 10784 4004
rect 10836 3992 10842 4004
rect 11808 3992 11836 4023
rect 12161 3995 12219 4001
rect 12161 3992 12173 3995
rect 10836 3964 12173 3992
rect 10836 3952 10842 3964
rect 12161 3961 12173 3964
rect 12207 3961 12219 3995
rect 12268 3992 12296 4091
rect 12342 4088 12348 4140
rect 12400 4128 12406 4140
rect 12544 4137 12572 4168
rect 16301 4165 16313 4199
rect 16347 4165 16359 4199
rect 16301 4159 16359 4165
rect 12618 4137 12624 4140
rect 12437 4131 12495 4137
rect 12437 4128 12449 4131
rect 12400 4100 12449 4128
rect 12400 4088 12406 4100
rect 12437 4097 12449 4100
rect 12483 4097 12495 4131
rect 12437 4091 12495 4097
rect 12529 4131 12587 4137
rect 12529 4097 12541 4131
rect 12575 4097 12587 4131
rect 12529 4091 12587 4097
rect 12617 4091 12624 4137
rect 12676 4128 12682 4140
rect 13354 4128 13360 4140
rect 12676 4100 12717 4128
rect 13315 4100 13360 4128
rect 12618 4088 12624 4091
rect 12676 4088 12682 4100
rect 13354 4088 13360 4100
rect 13412 4088 13418 4140
rect 14369 4131 14427 4137
rect 14369 4097 14381 4131
rect 14415 4097 14427 4131
rect 14369 4091 14427 4097
rect 14553 4131 14611 4137
rect 14553 4097 14565 4131
rect 14599 4128 14611 4131
rect 15194 4128 15200 4140
rect 14599 4100 15200 4128
rect 14599 4097 14611 4100
rect 14553 4091 14611 4097
rect 12805 4063 12863 4069
rect 12805 4029 12817 4063
rect 12851 4060 12863 4063
rect 13265 4063 13323 4069
rect 13265 4060 13277 4063
rect 12851 4032 13277 4060
rect 12851 4029 12863 4032
rect 12805 4023 12863 4029
rect 13265 4029 13277 4032
rect 13311 4029 13323 4063
rect 14384 4060 14412 4091
rect 15194 4088 15200 4100
rect 15252 4128 15258 4140
rect 16117 4131 16175 4137
rect 16117 4128 16129 4131
rect 15252 4100 16129 4128
rect 15252 4088 15258 4100
rect 16117 4097 16129 4100
rect 16163 4097 16175 4131
rect 18138 4128 18144 4140
rect 16117 4091 16175 4097
rect 17788 4100 18144 4128
rect 17788 4060 17816 4100
rect 18138 4088 18144 4100
rect 18196 4088 18202 4140
rect 14384 4032 17816 4060
rect 17865 4063 17923 4069
rect 13265 4023 13323 4029
rect 17865 4029 17877 4063
rect 17911 4029 17923 4063
rect 17865 4023 17923 4029
rect 12618 3992 12624 4004
rect 12268 3964 12624 3992
rect 12161 3955 12219 3961
rect 12618 3952 12624 3964
rect 12676 3952 12682 4004
rect 17586 3992 17592 4004
rect 12820 3964 17592 3992
rect 12820 3936 12848 3964
rect 17586 3952 17592 3964
rect 17644 3992 17650 4004
rect 17880 3992 17908 4023
rect 18322 4020 18328 4072
rect 18380 4060 18386 4072
rect 18509 4063 18567 4069
rect 18509 4060 18521 4063
rect 18380 4032 18521 4060
rect 18380 4020 18386 4032
rect 18509 4029 18521 4032
rect 18555 4029 18567 4063
rect 18509 4023 18567 4029
rect 17644 3964 17908 3992
rect 17644 3952 17650 3964
rect 8956 3896 10456 3924
rect 12802 3884 12808 3936
rect 12860 3884 12866 3936
rect 13633 3927 13691 3933
rect 13633 3893 13645 3927
rect 13679 3924 13691 3927
rect 14182 3924 14188 3936
rect 13679 3896 14188 3924
rect 13679 3893 13691 3896
rect 13633 3887 13691 3893
rect 14182 3884 14188 3896
rect 14240 3884 14246 3936
rect 14369 3927 14427 3933
rect 14369 3893 14381 3927
rect 14415 3924 14427 3927
rect 14642 3924 14648 3936
rect 14415 3896 14648 3924
rect 14415 3893 14427 3896
rect 14369 3887 14427 3893
rect 14642 3884 14648 3896
rect 14700 3884 14706 3936
rect 16942 3884 16948 3936
rect 17000 3924 17006 3936
rect 17405 3927 17463 3933
rect 17405 3924 17417 3927
rect 17000 3896 17417 3924
rect 17000 3884 17006 3896
rect 17405 3893 17417 3896
rect 17451 3893 17463 3927
rect 18046 3924 18052 3936
rect 18007 3896 18052 3924
rect 17405 3887 17463 3893
rect 18046 3884 18052 3896
rect 18104 3884 18110 3936
rect 0 3834 18860 3856
rect 0 3782 3110 3834
rect 3162 3782 3174 3834
rect 3226 3782 3238 3834
rect 3290 3782 3302 3834
rect 3354 3782 3366 3834
rect 3418 3782 6210 3834
rect 6262 3782 6274 3834
rect 6326 3782 6338 3834
rect 6390 3782 6402 3834
rect 6454 3782 6466 3834
rect 6518 3782 9310 3834
rect 9362 3782 9374 3834
rect 9426 3782 9438 3834
rect 9490 3782 9502 3834
rect 9554 3782 9566 3834
rect 9618 3782 12410 3834
rect 12462 3782 12474 3834
rect 12526 3782 12538 3834
rect 12590 3782 12602 3834
rect 12654 3782 12666 3834
rect 12718 3782 15510 3834
rect 15562 3782 15574 3834
rect 15626 3782 15638 3834
rect 15690 3782 15702 3834
rect 15754 3782 15766 3834
rect 15818 3782 18860 3834
rect 0 3760 18860 3782
rect 4157 3723 4215 3729
rect 4157 3720 4169 3723
rect 3712 3692 4169 3720
rect 750 3584 756 3596
rect 663 3556 756 3584
rect 750 3544 756 3556
rect 808 3584 814 3596
rect 2314 3584 2320 3596
rect 808 3556 2320 3584
rect 808 3544 814 3556
rect 2314 3544 2320 3556
rect 2372 3544 2378 3596
rect 2501 3587 2559 3593
rect 2501 3553 2513 3587
rect 2547 3584 2559 3587
rect 3329 3587 3387 3593
rect 2547 3556 2774 3584
rect 2547 3553 2559 3556
rect 2501 3547 2559 3553
rect 2406 3516 2412 3528
rect 2162 3488 2412 3516
rect 2406 3476 2412 3488
rect 2464 3476 2470 3528
rect 2746 3516 2774 3556
rect 3329 3553 3341 3587
rect 3375 3584 3387 3587
rect 3712 3584 3740 3692
rect 4157 3689 4169 3692
rect 4203 3720 4215 3723
rect 5350 3720 5356 3732
rect 4203 3692 5356 3720
rect 4203 3689 4215 3692
rect 4157 3683 4215 3689
rect 5350 3680 5356 3692
rect 5408 3680 5414 3732
rect 5626 3720 5632 3732
rect 5587 3692 5632 3720
rect 5626 3680 5632 3692
rect 5684 3680 5690 3732
rect 5721 3723 5779 3729
rect 5721 3689 5733 3723
rect 5767 3720 5779 3723
rect 6822 3720 6828 3732
rect 5767 3692 6828 3720
rect 5767 3689 5779 3692
rect 5721 3683 5779 3689
rect 6822 3680 6828 3692
rect 6880 3680 6886 3732
rect 7466 3680 7472 3732
rect 7524 3720 7530 3732
rect 7929 3723 7987 3729
rect 7929 3720 7941 3723
rect 7524 3692 7941 3720
rect 7524 3680 7530 3692
rect 7929 3689 7941 3692
rect 7975 3689 7987 3723
rect 7929 3683 7987 3689
rect 9585 3723 9643 3729
rect 9585 3689 9597 3723
rect 9631 3720 9643 3723
rect 9674 3720 9680 3732
rect 9631 3692 9680 3720
rect 9631 3689 9643 3692
rect 9585 3683 9643 3689
rect 9674 3680 9680 3692
rect 9732 3680 9738 3732
rect 10873 3723 10931 3729
rect 10873 3689 10885 3723
rect 10919 3720 10931 3723
rect 11698 3720 11704 3732
rect 10919 3692 11704 3720
rect 10919 3689 10931 3692
rect 10873 3683 10931 3689
rect 11698 3680 11704 3692
rect 11756 3680 11762 3732
rect 12802 3720 12808 3732
rect 12406 3692 12808 3720
rect 3878 3652 3884 3664
rect 3839 3624 3884 3652
rect 3878 3612 3884 3624
rect 3936 3612 3942 3664
rect 4062 3612 4068 3664
rect 4120 3652 4126 3664
rect 5905 3655 5963 3661
rect 5905 3652 5917 3655
rect 4120 3624 5917 3652
rect 4120 3612 4126 3624
rect 5905 3621 5917 3624
rect 5951 3621 5963 3655
rect 5905 3615 5963 3621
rect 6273 3655 6331 3661
rect 6273 3621 6285 3655
rect 6319 3621 6331 3655
rect 6273 3615 6331 3621
rect 6288 3584 6316 3615
rect 6362 3612 6368 3664
rect 6420 3652 6426 3664
rect 6638 3652 6644 3664
rect 6420 3624 6644 3652
rect 6420 3612 6426 3624
rect 6638 3612 6644 3624
rect 6696 3652 6702 3664
rect 8573 3655 8631 3661
rect 8573 3652 8585 3655
rect 6696 3624 8585 3652
rect 6696 3612 6702 3624
rect 8573 3621 8585 3624
rect 8619 3621 8631 3655
rect 12406 3652 12434 3692
rect 12802 3680 12808 3692
rect 12860 3680 12866 3732
rect 12894 3680 12900 3732
rect 12952 3720 12958 3732
rect 12952 3692 15884 3720
rect 12952 3680 12958 3692
rect 8573 3615 8631 3621
rect 9048 3624 12434 3652
rect 3375 3556 3740 3584
rect 4448 3556 6316 3584
rect 6917 3587 6975 3593
rect 3375 3553 3387 3556
rect 3329 3547 3387 3553
rect 2866 3516 2872 3528
rect 2746 3488 2872 3516
rect 2866 3476 2872 3488
rect 2924 3476 2930 3528
rect 2961 3519 3019 3525
rect 2961 3485 2973 3519
rect 3007 3516 3019 3519
rect 3602 3516 3608 3528
rect 3007 3488 3608 3516
rect 3007 3485 3019 3488
rect 2961 3479 3019 3485
rect 3602 3476 3608 3488
rect 3660 3476 3666 3528
rect 3878 3516 3884 3528
rect 3839 3488 3884 3516
rect 3878 3476 3884 3488
rect 3936 3476 3942 3528
rect 4065 3519 4123 3525
rect 4065 3485 4077 3519
rect 4111 3516 4123 3519
rect 4154 3516 4160 3528
rect 4111 3488 4160 3516
rect 4111 3485 4123 3488
rect 4065 3479 4123 3485
rect 4154 3476 4160 3488
rect 4212 3476 4218 3528
rect 4338 3516 4344 3528
rect 4299 3488 4344 3516
rect 4338 3476 4344 3488
rect 4396 3476 4402 3528
rect 4448 3525 4476 3556
rect 4433 3519 4491 3525
rect 4433 3485 4445 3519
rect 4479 3485 4491 3519
rect 4433 3479 4491 3485
rect 4522 3476 4528 3528
rect 4580 3516 4586 3528
rect 5000 3525 5028 3556
rect 6917 3553 6929 3587
rect 6963 3584 6975 3587
rect 7098 3584 7104 3596
rect 6963 3556 7104 3584
rect 6963 3553 6975 3556
rect 6917 3547 6975 3553
rect 7098 3544 7104 3556
rect 7156 3544 7162 3596
rect 9048 3593 9076 3624
rect 15856 3596 15884 3692
rect 18138 3652 18144 3664
rect 18099 3624 18144 3652
rect 18138 3612 18144 3624
rect 18196 3612 18202 3664
rect 9033 3587 9091 3593
rect 9033 3584 9045 3587
rect 8220 3556 9045 3584
rect 4985 3519 5043 3525
rect 4580 3488 4625 3516
rect 4580 3476 4586 3488
rect 4985 3485 4997 3519
rect 5031 3485 5043 3519
rect 4985 3479 5043 3485
rect 5074 3476 5080 3528
rect 5132 3516 5138 3528
rect 5261 3519 5319 3525
rect 5261 3516 5273 3519
rect 5132 3488 5273 3516
rect 5132 3476 5138 3488
rect 5261 3485 5273 3488
rect 5307 3485 5319 3519
rect 5261 3479 5319 3485
rect 5350 3476 5356 3528
rect 5408 3516 5414 3528
rect 5813 3519 5871 3525
rect 5813 3516 5825 3519
rect 5408 3488 5825 3516
rect 5408 3476 5414 3488
rect 5813 3485 5825 3488
rect 5859 3485 5871 3519
rect 5813 3479 5871 3485
rect 5902 3476 5908 3528
rect 5960 3516 5966 3528
rect 6089 3519 6147 3525
rect 5960 3488 6005 3516
rect 5960 3476 5966 3488
rect 6089 3485 6101 3519
rect 6135 3485 6147 3519
rect 6089 3479 6147 3485
rect 1029 3451 1087 3457
rect 1029 3417 1041 3451
rect 1075 3417 1087 3451
rect 2685 3451 2743 3457
rect 2685 3448 2697 3451
rect 1029 3411 1087 3417
rect 2332 3420 2697 3448
rect 1044 3380 1072 3411
rect 2332 3380 2360 3420
rect 2685 3417 2697 3420
rect 2731 3417 2743 3451
rect 2685 3411 2743 3417
rect 3970 3408 3976 3460
rect 4028 3448 4034 3460
rect 4028 3420 5396 3448
rect 4028 3408 4034 3420
rect 1044 3352 2360 3380
rect 3878 3340 3884 3392
rect 3936 3380 3942 3392
rect 5368 3389 5396 3420
rect 5442 3408 5448 3460
rect 5500 3448 5506 3460
rect 6104 3448 6132 3479
rect 7282 3476 7288 3528
rect 7340 3516 7346 3528
rect 8220 3525 8248 3556
rect 9033 3553 9045 3556
rect 9079 3553 9091 3587
rect 9033 3547 9091 3553
rect 10505 3587 10563 3593
rect 10505 3553 10517 3587
rect 10551 3553 10563 3587
rect 10870 3584 10876 3596
rect 10505 3547 10563 3553
rect 10612 3556 10876 3584
rect 8021 3519 8079 3525
rect 8021 3516 8033 3519
rect 7340 3488 8033 3516
rect 7340 3476 7346 3488
rect 8021 3485 8033 3488
rect 8067 3485 8079 3519
rect 8021 3479 8079 3485
rect 8205 3519 8263 3525
rect 8205 3485 8217 3519
rect 8251 3485 8263 3519
rect 8205 3479 8263 3485
rect 9122 3476 9128 3528
rect 9180 3516 9186 3528
rect 9766 3516 9772 3528
rect 9180 3488 9225 3516
rect 9679 3488 9772 3516
rect 9180 3476 9186 3488
rect 9766 3476 9772 3488
rect 9824 3516 9830 3528
rect 10520 3516 10548 3547
rect 10612 3525 10640 3556
rect 10870 3544 10876 3556
rect 10928 3544 10934 3596
rect 13817 3587 13875 3593
rect 13817 3553 13829 3587
rect 13863 3584 13875 3587
rect 14550 3584 14556 3596
rect 13863 3556 14556 3584
rect 13863 3553 13875 3556
rect 13817 3547 13875 3553
rect 9824 3488 10548 3516
rect 9824 3476 9830 3488
rect 7837 3451 7895 3457
rect 7837 3448 7849 3451
rect 5500 3420 6132 3448
rect 6472 3420 7849 3448
rect 5500 3408 5506 3420
rect 4801 3383 4859 3389
rect 4801 3380 4813 3383
rect 3936 3352 4813 3380
rect 3936 3340 3942 3352
rect 4801 3349 4813 3352
rect 4847 3349 4859 3383
rect 4801 3343 4859 3349
rect 5353 3383 5411 3389
rect 5353 3349 5365 3383
rect 5399 3349 5411 3383
rect 5353 3343 5411 3349
rect 5626 3340 5632 3392
rect 5684 3380 5690 3392
rect 6472 3380 6500 3420
rect 7837 3417 7849 3420
rect 7883 3448 7895 3451
rect 8754 3448 8760 3460
rect 7883 3420 8760 3448
rect 7883 3417 7895 3420
rect 7837 3411 7895 3417
rect 8754 3408 8760 3420
rect 8812 3408 8818 3460
rect 10520 3448 10548 3488
rect 10597 3519 10655 3525
rect 10597 3485 10609 3519
rect 10643 3485 10655 3519
rect 10597 3479 10655 3485
rect 10686 3476 10692 3528
rect 10744 3516 10750 3528
rect 13078 3516 13084 3528
rect 10744 3488 13084 3516
rect 10744 3476 10750 3488
rect 13078 3476 13084 3488
rect 13136 3516 13142 3528
rect 13832 3516 13860 3547
rect 14550 3544 14556 3556
rect 14608 3544 14614 3596
rect 15838 3584 15844 3596
rect 15751 3556 15844 3584
rect 15838 3544 15844 3556
rect 15896 3544 15902 3596
rect 17586 3584 17592 3596
rect 17547 3556 17592 3584
rect 17586 3544 17592 3556
rect 17644 3544 17650 3596
rect 14182 3516 14188 3528
rect 13136 3488 13860 3516
rect 14143 3488 14188 3516
rect 13136 3476 13142 3488
rect 14182 3476 14188 3488
rect 14240 3476 14246 3528
rect 15102 3476 15108 3528
rect 15160 3516 15166 3528
rect 16206 3516 16212 3528
rect 15160 3488 15240 3516
rect 16167 3488 16212 3516
rect 15160 3476 15166 3488
rect 12066 3448 12072 3460
rect 10520 3420 12072 3448
rect 12066 3408 12072 3420
rect 12124 3408 12130 3460
rect 12250 3408 12256 3460
rect 12308 3448 12314 3460
rect 13814 3448 13820 3460
rect 12308 3420 13820 3448
rect 12308 3408 12314 3420
rect 13814 3408 13820 3420
rect 13872 3408 13878 3460
rect 15212 3448 15240 3488
rect 16206 3476 16212 3488
rect 16264 3476 16270 3528
rect 18322 3516 18328 3528
rect 18283 3488 18328 3516
rect 18322 3476 18328 3488
rect 18380 3476 18386 3528
rect 15212 3434 15792 3448
rect 15226 3420 15792 3434
rect 6638 3380 6644 3392
rect 5684 3352 6500 3380
rect 6599 3352 6644 3380
rect 5684 3340 5690 3352
rect 6638 3340 6644 3352
rect 6696 3340 6702 3392
rect 6730 3340 6736 3392
rect 6788 3380 6794 3392
rect 6788 3352 6833 3380
rect 6788 3340 6794 3352
rect 7098 3340 7104 3392
rect 7156 3380 7162 3392
rect 7561 3383 7619 3389
rect 7561 3380 7573 3383
rect 7156 3352 7573 3380
rect 7156 3340 7162 3352
rect 7561 3349 7573 3352
rect 7607 3349 7619 3383
rect 7561 3343 7619 3349
rect 8662 3340 8668 3392
rect 8720 3380 8726 3392
rect 9217 3383 9275 3389
rect 9217 3380 9229 3383
rect 8720 3352 9229 3380
rect 8720 3340 8726 3352
rect 9217 3349 9229 3352
rect 9263 3349 9275 3383
rect 9217 3343 9275 3349
rect 13354 3340 13360 3392
rect 13412 3380 13418 3392
rect 15611 3383 15669 3389
rect 15611 3380 15623 3383
rect 13412 3352 15623 3380
rect 13412 3340 13418 3352
rect 15611 3349 15623 3352
rect 15657 3349 15669 3383
rect 15764 3380 15792 3420
rect 16298 3380 16304 3392
rect 15764 3352 16304 3380
rect 15611 3343 15669 3349
rect 16298 3340 16304 3352
rect 16356 3380 16362 3392
rect 16592 3380 16620 3434
rect 16356 3352 16620 3380
rect 16356 3340 16362 3352
rect 0 3290 18860 3312
rect 0 3238 4660 3290
rect 4712 3238 4724 3290
rect 4776 3238 4788 3290
rect 4840 3238 4852 3290
rect 4904 3238 4916 3290
rect 4968 3238 7760 3290
rect 7812 3238 7824 3290
rect 7876 3238 7888 3290
rect 7940 3238 7952 3290
rect 8004 3238 8016 3290
rect 8068 3238 10860 3290
rect 10912 3238 10924 3290
rect 10976 3238 10988 3290
rect 11040 3238 11052 3290
rect 11104 3238 11116 3290
rect 11168 3238 13960 3290
rect 14012 3238 14024 3290
rect 14076 3238 14088 3290
rect 14140 3238 14152 3290
rect 14204 3238 14216 3290
rect 14268 3238 17060 3290
rect 17112 3238 17124 3290
rect 17176 3238 17188 3290
rect 17240 3238 17252 3290
rect 17304 3238 17316 3290
rect 17368 3238 18860 3290
rect 0 3216 18860 3238
rect 3421 3179 3479 3185
rect 3421 3145 3433 3179
rect 3467 3176 3479 3179
rect 3510 3176 3516 3188
rect 3467 3148 3516 3176
rect 3467 3145 3479 3148
rect 3421 3139 3479 3145
rect 3510 3136 3516 3148
rect 3568 3136 3574 3188
rect 3602 3136 3608 3188
rect 3660 3176 3666 3188
rect 4430 3176 4436 3188
rect 3660 3148 3705 3176
rect 3804 3148 4436 3176
rect 3660 3136 3666 3148
rect 2866 3068 2872 3120
rect 2924 3108 2930 3120
rect 2961 3111 3019 3117
rect 2961 3108 2973 3111
rect 2924 3080 2973 3108
rect 2924 3068 2930 3080
rect 2961 3077 2973 3080
rect 3007 3108 3019 3111
rect 3804 3108 3832 3148
rect 4430 3136 4436 3148
rect 4488 3136 4494 3188
rect 5537 3179 5595 3185
rect 5537 3145 5549 3179
rect 5583 3145 5595 3179
rect 14550 3176 14556 3188
rect 5537 3139 5595 3145
rect 8312 3148 12434 3176
rect 14511 3148 14556 3176
rect 3007 3080 3832 3108
rect 5552 3108 5580 3139
rect 8312 3120 8340 3148
rect 5810 3108 5816 3120
rect 5552 3080 5816 3108
rect 3007 3077 3019 3080
rect 2961 3071 3019 3077
rect 5810 3068 5816 3080
rect 5868 3108 5874 3120
rect 6362 3108 6368 3120
rect 5868 3080 6040 3108
rect 5868 3068 5874 3080
rect 3697 3043 3755 3049
rect 3697 3009 3709 3043
rect 3743 3040 3755 3043
rect 3878 3040 3884 3052
rect 3743 3012 3884 3040
rect 3743 3009 3755 3012
rect 3697 3003 3755 3009
rect 3329 2907 3387 2913
rect 3329 2873 3341 2907
rect 3375 2904 3387 2907
rect 3712 2904 3740 3003
rect 3878 3000 3884 3012
rect 3936 3000 3942 3052
rect 4154 3000 4160 3052
rect 4212 3040 4218 3052
rect 4522 3040 4528 3052
rect 4212 3012 4528 3040
rect 4212 3000 4218 3012
rect 4522 3000 4528 3012
rect 4580 3040 4586 3052
rect 4798 3040 4804 3052
rect 4580 3012 4804 3040
rect 4580 3000 4586 3012
rect 4798 3000 4804 3012
rect 4856 3000 4862 3052
rect 5534 3040 5540 3052
rect 5495 3012 5540 3040
rect 5534 3000 5540 3012
rect 5592 3000 5598 3052
rect 5902 3040 5908 3052
rect 5863 3012 5908 3040
rect 5902 3000 5908 3012
rect 5960 3000 5966 3052
rect 6012 3049 6040 3080
rect 6104 3080 6368 3108
rect 5997 3043 6055 3049
rect 5997 3009 6009 3043
rect 6043 3009 6055 3043
rect 5997 3003 6055 3009
rect 4338 2932 4344 2984
rect 4396 2972 4402 2984
rect 4893 2975 4951 2981
rect 4893 2972 4905 2975
rect 4396 2944 4905 2972
rect 4396 2932 4402 2944
rect 4893 2941 4905 2944
rect 4939 2972 4951 2975
rect 5353 2975 5411 2981
rect 5353 2972 5365 2975
rect 4939 2944 5365 2972
rect 4939 2941 4951 2944
rect 4893 2935 4951 2941
rect 5353 2941 5365 2944
rect 5399 2941 5411 2975
rect 5626 2972 5632 2984
rect 5587 2944 5632 2972
rect 5353 2935 5411 2941
rect 5626 2932 5632 2944
rect 5684 2932 5690 2984
rect 5813 2975 5871 2981
rect 5813 2941 5825 2975
rect 5859 2972 5871 2975
rect 6104 2972 6132 3080
rect 6362 3068 6368 3080
rect 6420 3068 6426 3120
rect 7466 3108 7472 3120
rect 7392 3080 7472 3108
rect 6181 3043 6239 3049
rect 6181 3009 6193 3043
rect 6227 3040 6239 3043
rect 7101 3043 7159 3049
rect 7101 3040 7113 3043
rect 6227 3012 7113 3040
rect 6227 3009 6239 3012
rect 6181 3003 6239 3009
rect 7101 3009 7113 3012
rect 7147 3040 7159 3043
rect 7190 3040 7196 3052
rect 7147 3012 7196 3040
rect 7147 3009 7159 3012
rect 7101 3003 7159 3009
rect 5859 2944 6132 2972
rect 5859 2941 5871 2944
rect 5813 2935 5871 2941
rect 3375 2876 3740 2904
rect 3375 2873 3387 2876
rect 3329 2867 3387 2873
rect 4430 2864 4436 2916
rect 4488 2904 4494 2916
rect 6089 2907 6147 2913
rect 6089 2904 6101 2907
rect 4488 2876 6101 2904
rect 4488 2864 4494 2876
rect 6089 2873 6101 2876
rect 6135 2873 6147 2907
rect 6089 2867 6147 2873
rect 5353 2839 5411 2845
rect 5353 2805 5365 2839
rect 5399 2836 5411 2839
rect 6196 2836 6224 3003
rect 7190 3000 7196 3012
rect 7248 3000 7254 3052
rect 7392 3049 7420 3080
rect 7466 3068 7472 3080
rect 7524 3108 7530 3120
rect 8113 3111 8171 3117
rect 8113 3108 8125 3111
rect 7524 3080 8125 3108
rect 7524 3068 7530 3080
rect 8113 3077 8125 3080
rect 8159 3077 8171 3111
rect 8113 3071 8171 3077
rect 8294 3068 8300 3120
rect 8352 3108 8358 3120
rect 8352 3080 8445 3108
rect 8352 3068 8358 3080
rect 9122 3068 9128 3120
rect 9180 3068 9186 3120
rect 11330 3068 11336 3120
rect 11388 3068 11394 3120
rect 7377 3043 7435 3049
rect 7377 3009 7389 3043
rect 7423 3009 7435 3043
rect 7558 3040 7564 3052
rect 7519 3012 7564 3040
rect 7377 3003 7435 3009
rect 7558 3000 7564 3012
rect 7616 3000 7622 3052
rect 7650 3000 7656 3052
rect 7708 3040 7714 3052
rect 7834 3040 7840 3052
rect 7708 3012 7753 3040
rect 7795 3012 7840 3040
rect 7708 3000 7714 3012
rect 7834 3000 7840 3012
rect 7892 3000 7898 3052
rect 8389 3043 8447 3049
rect 8389 3009 8401 3043
rect 8435 3040 8447 3043
rect 8662 3040 8668 3052
rect 8435 3012 8668 3040
rect 8435 3009 8447 3012
rect 8389 3003 8447 3009
rect 8662 3000 8668 3012
rect 8720 3000 8726 3052
rect 12406 3040 12434 3148
rect 14550 3136 14556 3148
rect 14608 3176 14614 3188
rect 15378 3176 15384 3188
rect 14608 3148 15384 3176
rect 14608 3136 14614 3148
rect 15378 3136 15384 3148
rect 15436 3136 15442 3188
rect 15979 3179 16037 3185
rect 15979 3145 15991 3179
rect 16025 3176 16037 3179
rect 16206 3176 16212 3188
rect 16025 3148 16212 3176
rect 16025 3145 16037 3148
rect 15979 3139 16037 3145
rect 16206 3136 16212 3148
rect 16264 3136 16270 3188
rect 18322 3176 18328 3188
rect 18283 3148 18328 3176
rect 18322 3136 18328 3148
rect 18380 3136 18386 3188
rect 12894 3108 12900 3120
rect 12855 3080 12900 3108
rect 12894 3068 12900 3080
rect 12952 3068 12958 3120
rect 13354 3068 13360 3120
rect 13412 3108 13418 3120
rect 14461 3111 14519 3117
rect 14461 3108 14473 3111
rect 13412 3080 14473 3108
rect 13412 3068 13418 3080
rect 14461 3077 14473 3080
rect 14507 3077 14519 3111
rect 14461 3071 14519 3077
rect 16390 3068 16396 3120
rect 16448 3068 16454 3120
rect 12529 3043 12587 3049
rect 12529 3040 12541 3043
rect 12406 3012 12541 3040
rect 12529 3009 12541 3012
rect 12575 3009 12587 3043
rect 12802 3040 12808 3052
rect 12763 3012 12808 3040
rect 12529 3003 12587 3009
rect 8757 2975 8815 2981
rect 8757 2972 8769 2975
rect 7760 2944 8769 2972
rect 7760 2913 7788 2944
rect 8757 2941 8769 2944
rect 8803 2941 8815 2975
rect 8757 2935 8815 2941
rect 10413 2975 10471 2981
rect 10413 2941 10425 2975
rect 10459 2972 10471 2975
rect 10594 2972 10600 2984
rect 10459 2944 10600 2972
rect 10459 2941 10471 2944
rect 10413 2935 10471 2941
rect 10594 2932 10600 2944
rect 10652 2932 10658 2984
rect 10781 2975 10839 2981
rect 10781 2941 10793 2975
rect 10827 2972 10839 2975
rect 12250 2972 12256 2984
rect 10827 2944 12256 2972
rect 10827 2941 10839 2944
rect 10781 2935 10839 2941
rect 12250 2932 12256 2944
rect 12308 2932 12314 2984
rect 12544 2972 12572 3003
rect 12802 3000 12808 3012
rect 12860 3000 12866 3052
rect 13173 3043 13231 3049
rect 13173 3009 13185 3043
rect 13219 3040 13231 3043
rect 13219 3012 13584 3040
rect 13219 3009 13231 3012
rect 13173 3003 13231 3009
rect 12894 2972 12900 2984
rect 12544 2944 12900 2972
rect 12894 2932 12900 2944
rect 12952 2932 12958 2984
rect 13556 2913 13584 3012
rect 13814 3000 13820 3052
rect 13872 3040 13878 3052
rect 14001 3043 14059 3049
rect 14001 3040 14013 3043
rect 13872 3012 14013 3040
rect 13872 3000 13878 3012
rect 14001 3009 14013 3012
rect 14047 3009 14059 3043
rect 17773 3043 17831 3049
rect 17773 3040 17785 3043
rect 14001 3003 14059 3009
rect 17328 3012 17785 3040
rect 14642 2972 14648 2984
rect 14603 2944 14648 2972
rect 14642 2932 14648 2944
rect 14700 2932 14706 2984
rect 15838 2932 15844 2984
rect 15896 2972 15902 2984
rect 17328 2972 17356 3012
rect 17773 3009 17785 3012
rect 17819 3040 17831 3043
rect 17954 3040 17960 3052
rect 17819 3012 17960 3040
rect 17819 3009 17831 3012
rect 17773 3003 17831 3009
rect 17954 3000 17960 3012
rect 18012 3000 18018 3052
rect 15896 2944 17356 2972
rect 15896 2932 15902 2944
rect 17402 2932 17408 2984
rect 17460 2972 17466 2984
rect 17460 2944 17505 2972
rect 17460 2932 17466 2944
rect 17586 2932 17592 2984
rect 17644 2972 17650 2984
rect 17865 2975 17923 2981
rect 17865 2972 17877 2975
rect 17644 2944 17877 2972
rect 17644 2932 17650 2944
rect 17865 2941 17877 2944
rect 17911 2941 17923 2975
rect 17865 2935 17923 2941
rect 7745 2907 7803 2913
rect 7745 2873 7757 2907
rect 7791 2873 7803 2907
rect 7745 2867 7803 2873
rect 13541 2907 13599 2913
rect 13541 2873 13553 2907
rect 13587 2873 13599 2907
rect 13541 2867 13599 2873
rect 13725 2907 13783 2913
rect 13725 2873 13737 2907
rect 13771 2904 13783 2907
rect 14093 2907 14151 2913
rect 14093 2904 14105 2907
rect 13771 2876 14105 2904
rect 13771 2873 13783 2876
rect 13725 2867 13783 2873
rect 14093 2873 14105 2876
rect 14139 2873 14151 2907
rect 14093 2867 14151 2873
rect 5399 2808 6224 2836
rect 5399 2805 5411 2808
rect 5353 2799 5411 2805
rect 6638 2796 6644 2848
rect 6696 2836 6702 2848
rect 7193 2839 7251 2845
rect 7193 2836 7205 2839
rect 6696 2808 7205 2836
rect 6696 2796 6702 2808
rect 7193 2805 7205 2808
rect 7239 2836 7251 2839
rect 8754 2836 8760 2848
rect 7239 2808 8760 2836
rect 7239 2805 7251 2808
rect 7193 2799 7251 2805
rect 8754 2796 8760 2808
rect 8812 2796 8818 2848
rect 10226 2845 10232 2848
rect 10183 2839 10232 2845
rect 10183 2805 10195 2839
rect 10229 2805 10232 2839
rect 10183 2799 10232 2805
rect 10226 2796 10232 2799
rect 10284 2796 10290 2848
rect 11790 2796 11796 2848
rect 11848 2836 11854 2848
rect 12207 2839 12265 2845
rect 12207 2836 12219 2839
rect 11848 2808 12219 2836
rect 11848 2796 11854 2808
rect 12207 2805 12219 2808
rect 12253 2805 12265 2839
rect 12207 2799 12265 2805
rect 0 2746 18860 2768
rect 0 2694 3110 2746
rect 3162 2694 3174 2746
rect 3226 2694 3238 2746
rect 3290 2694 3302 2746
rect 3354 2694 3366 2746
rect 3418 2694 6210 2746
rect 6262 2694 6274 2746
rect 6326 2694 6338 2746
rect 6390 2694 6402 2746
rect 6454 2694 6466 2746
rect 6518 2694 9310 2746
rect 9362 2694 9374 2746
rect 9426 2694 9438 2746
rect 9490 2694 9502 2746
rect 9554 2694 9566 2746
rect 9618 2694 12410 2746
rect 12462 2694 12474 2746
rect 12526 2694 12538 2746
rect 12590 2694 12602 2746
rect 12654 2694 12666 2746
rect 12718 2694 15510 2746
rect 15562 2694 15574 2746
rect 15626 2694 15638 2746
rect 15690 2694 15702 2746
rect 15754 2694 15766 2746
rect 15818 2694 18860 2746
rect 0 2672 18860 2694
rect 6825 2635 6883 2641
rect 6825 2601 6837 2635
rect 6871 2632 6883 2635
rect 7558 2632 7564 2644
rect 6871 2604 7564 2632
rect 6871 2601 6883 2604
rect 6825 2595 6883 2601
rect 7558 2592 7564 2604
rect 7616 2592 7622 2644
rect 12250 2632 12256 2644
rect 12211 2604 12256 2632
rect 12250 2592 12256 2604
rect 12308 2592 12314 2644
rect 3145 2567 3203 2573
rect 3145 2564 3157 2567
rect 2056 2536 3157 2564
rect 750 2496 756 2508
rect 711 2468 756 2496
rect 750 2456 756 2468
rect 808 2456 814 2508
rect 1029 2499 1087 2505
rect 1029 2465 1041 2499
rect 1075 2496 1087 2499
rect 2056 2496 2084 2536
rect 3145 2533 3157 2536
rect 3191 2533 3203 2567
rect 3145 2527 3203 2533
rect 3237 2567 3295 2573
rect 3237 2533 3249 2567
rect 3283 2564 3295 2567
rect 3878 2564 3884 2576
rect 3283 2536 3884 2564
rect 3283 2533 3295 2536
rect 3237 2527 3295 2533
rect 3878 2524 3884 2536
rect 3936 2564 3942 2576
rect 5626 2564 5632 2576
rect 3936 2536 4200 2564
rect 3936 2524 3942 2536
rect 1075 2468 2084 2496
rect 3053 2499 3111 2505
rect 1075 2465 1087 2468
rect 1029 2459 1087 2465
rect 3053 2465 3065 2499
rect 3099 2496 3111 2499
rect 3694 2496 3700 2508
rect 3099 2468 3700 2496
rect 3099 2465 3111 2468
rect 3053 2459 3111 2465
rect 3694 2456 3700 2468
rect 3752 2456 3758 2508
rect 4172 2505 4200 2536
rect 5000 2536 5632 2564
rect 5000 2505 5028 2536
rect 5626 2524 5632 2536
rect 5684 2524 5690 2576
rect 5813 2567 5871 2573
rect 5813 2533 5825 2567
rect 5859 2564 5871 2567
rect 7650 2564 7656 2576
rect 5859 2536 7656 2564
rect 5859 2533 5871 2536
rect 5813 2527 5871 2533
rect 7650 2524 7656 2536
rect 7708 2524 7714 2576
rect 12161 2567 12219 2573
rect 12161 2533 12173 2567
rect 12207 2564 12219 2567
rect 12802 2564 12808 2576
rect 12207 2536 12808 2564
rect 12207 2533 12219 2536
rect 12161 2527 12219 2533
rect 12802 2524 12808 2536
rect 12860 2524 12866 2576
rect 16482 2564 16488 2576
rect 15396 2536 16488 2564
rect 15396 2508 15424 2536
rect 16482 2524 16488 2536
rect 16540 2524 16546 2576
rect 4157 2499 4215 2505
rect 4157 2465 4169 2499
rect 4203 2465 4215 2499
rect 4157 2459 4215 2465
rect 4985 2499 5043 2505
rect 4985 2465 4997 2499
rect 5031 2465 5043 2499
rect 4985 2459 5043 2465
rect 5169 2499 5227 2505
rect 5169 2465 5181 2499
rect 5215 2496 5227 2499
rect 5258 2496 5264 2508
rect 5215 2468 5264 2496
rect 5215 2465 5227 2468
rect 5169 2459 5227 2465
rect 5258 2456 5264 2468
rect 5316 2456 5322 2508
rect 5718 2496 5724 2508
rect 5644 2468 5724 2496
rect 3329 2431 3387 2437
rect 3329 2397 3341 2431
rect 3375 2397 3387 2431
rect 4430 2428 4436 2440
rect 4391 2400 4436 2428
rect 3329 2391 3387 2397
rect 2406 2360 2412 2372
rect 2254 2332 2412 2360
rect 2406 2320 2412 2332
rect 2464 2360 2470 2372
rect 2682 2360 2688 2372
rect 2464 2332 2688 2360
rect 2464 2320 2470 2332
rect 2682 2320 2688 2332
rect 2740 2320 2746 2372
rect 3344 2360 3372 2391
rect 4430 2388 4436 2400
rect 4488 2388 4494 2440
rect 5644 2437 5672 2468
rect 5718 2456 5724 2468
rect 5776 2456 5782 2508
rect 10137 2499 10195 2505
rect 10137 2496 10149 2499
rect 6748 2468 10149 2496
rect 5629 2431 5687 2437
rect 5629 2397 5641 2431
rect 5675 2397 5687 2431
rect 5810 2428 5816 2440
rect 5771 2400 5816 2428
rect 5629 2391 5687 2397
rect 5810 2388 5816 2400
rect 5868 2388 5874 2440
rect 6748 2437 6776 2468
rect 10137 2465 10149 2468
rect 10183 2465 10195 2499
rect 10137 2459 10195 2465
rect 11701 2499 11759 2505
rect 11701 2465 11713 2499
rect 11747 2465 11759 2499
rect 15378 2496 15384 2508
rect 11701 2459 11759 2465
rect 11808 2468 12434 2496
rect 15339 2468 15384 2496
rect 6089 2431 6147 2437
rect 6089 2397 6101 2431
rect 6135 2428 6147 2431
rect 6733 2431 6791 2437
rect 6733 2428 6745 2431
rect 6135 2400 6745 2428
rect 6135 2397 6147 2400
rect 6089 2391 6147 2397
rect 6733 2397 6745 2400
rect 6779 2397 6791 2431
rect 6733 2391 6791 2397
rect 6825 2431 6883 2437
rect 6825 2397 6837 2431
rect 6871 2428 6883 2431
rect 7098 2428 7104 2440
rect 6871 2400 7104 2428
rect 6871 2397 6883 2400
rect 6825 2391 6883 2397
rect 7098 2388 7104 2400
rect 7156 2388 7162 2440
rect 7190 2388 7196 2440
rect 7248 2428 7254 2440
rect 7469 2431 7527 2437
rect 7469 2428 7481 2431
rect 7248 2400 7481 2428
rect 7248 2388 7254 2400
rect 7469 2397 7481 2400
rect 7515 2397 7527 2431
rect 7469 2391 7527 2397
rect 8294 2388 8300 2440
rect 8352 2428 8358 2440
rect 8570 2428 8576 2440
rect 8352 2400 8576 2428
rect 8352 2388 8358 2400
rect 8570 2388 8576 2400
rect 8628 2388 8634 2440
rect 8662 2388 8668 2440
rect 8720 2428 8726 2440
rect 10226 2428 10232 2440
rect 8720 2400 8765 2428
rect 10139 2400 10232 2428
rect 8720 2388 8726 2400
rect 10226 2388 10232 2400
rect 10284 2428 10290 2440
rect 11716 2428 11744 2459
rect 11808 2440 11836 2468
rect 10284 2400 11744 2428
rect 10284 2388 10290 2400
rect 11790 2388 11796 2440
rect 11848 2428 11854 2440
rect 12250 2428 12256 2440
rect 11848 2400 11893 2428
rect 12211 2400 12256 2428
rect 11848 2388 11854 2400
rect 12250 2388 12256 2400
rect 12308 2388 12314 2440
rect 12406 2428 12434 2468
rect 15378 2456 15384 2468
rect 15436 2456 15442 2508
rect 15746 2456 15752 2508
rect 15804 2496 15810 2508
rect 17954 2496 17960 2508
rect 15804 2468 15849 2496
rect 17915 2468 17960 2496
rect 15804 2456 15810 2468
rect 17954 2456 17960 2468
rect 18012 2456 18018 2508
rect 12621 2431 12679 2437
rect 12621 2428 12633 2431
rect 12406 2400 12633 2428
rect 12621 2397 12633 2400
rect 12667 2397 12679 2431
rect 12621 2391 12679 2397
rect 14550 2388 14556 2440
rect 14608 2428 14614 2440
rect 15473 2431 15531 2437
rect 15473 2428 15485 2431
rect 14608 2400 15485 2428
rect 14608 2388 14614 2400
rect 15473 2397 15485 2400
rect 15519 2397 15531 2431
rect 15473 2391 15531 2397
rect 15562 2388 15568 2440
rect 15620 2428 15626 2440
rect 18506 2428 18512 2440
rect 15620 2400 15665 2428
rect 18467 2400 18512 2428
rect 15620 2388 15626 2400
rect 18506 2388 18512 2400
rect 18564 2388 18570 2440
rect 3510 2360 3516 2372
rect 3344 2332 3516 2360
rect 3510 2320 3516 2332
rect 3568 2360 3574 2372
rect 4893 2363 4951 2369
rect 4893 2360 4905 2363
rect 3568 2332 4905 2360
rect 3568 2320 3574 2332
rect 4893 2329 4905 2332
rect 4939 2329 4951 2363
rect 4893 2323 4951 2329
rect 5258 2320 5264 2372
rect 5316 2360 5322 2372
rect 6549 2363 6607 2369
rect 6549 2360 6561 2363
rect 5316 2332 6561 2360
rect 5316 2320 5322 2332
rect 6549 2329 6561 2332
rect 6595 2329 6607 2363
rect 6549 2323 6607 2329
rect 7834 2320 7840 2372
rect 7892 2320 7898 2372
rect 8849 2363 8907 2369
rect 8849 2360 8861 2363
rect 8680 2332 8861 2360
rect 2501 2295 2559 2301
rect 2501 2261 2513 2295
rect 2547 2292 2559 2295
rect 2958 2292 2964 2304
rect 2547 2264 2964 2292
rect 2547 2261 2559 2264
rect 2501 2255 2559 2261
rect 2958 2252 2964 2264
rect 3016 2292 3022 2304
rect 3602 2292 3608 2304
rect 3016 2264 3608 2292
rect 3016 2252 3022 2264
rect 3602 2252 3608 2264
rect 3660 2292 3666 2304
rect 4062 2292 4068 2304
rect 3660 2264 4068 2292
rect 3660 2252 3666 2264
rect 4062 2252 4068 2264
rect 4120 2252 4126 2304
rect 4338 2252 4344 2304
rect 4396 2292 4402 2304
rect 4525 2295 4583 2301
rect 4525 2292 4537 2295
rect 4396 2264 4537 2292
rect 4396 2252 4402 2264
rect 4525 2261 4537 2264
rect 4571 2261 4583 2295
rect 4525 2255 4583 2261
rect 7561 2295 7619 2301
rect 7561 2261 7573 2295
rect 7607 2292 7619 2295
rect 7852 2292 7880 2320
rect 8202 2292 8208 2304
rect 7607 2264 8208 2292
rect 7607 2261 7619 2264
rect 7561 2255 7619 2261
rect 8202 2252 8208 2264
rect 8260 2292 8266 2304
rect 8680 2292 8708 2332
rect 8849 2329 8861 2332
rect 8895 2360 8907 2363
rect 12158 2360 12164 2372
rect 8895 2332 12164 2360
rect 8895 2329 8907 2332
rect 8849 2323 8907 2329
rect 12158 2320 12164 2332
rect 12216 2360 12222 2372
rect 12345 2363 12403 2369
rect 12345 2360 12357 2363
rect 12216 2332 12357 2360
rect 12216 2320 12222 2332
rect 12345 2329 12357 2332
rect 12391 2329 12403 2363
rect 12345 2323 12403 2329
rect 12529 2363 12587 2369
rect 12529 2329 12541 2363
rect 12575 2360 12587 2363
rect 13170 2360 13176 2372
rect 12575 2332 13176 2360
rect 12575 2329 12587 2332
rect 12529 2323 12587 2329
rect 13170 2320 13176 2332
rect 13228 2320 13234 2372
rect 15194 2369 15200 2372
rect 15136 2363 15200 2369
rect 15136 2329 15148 2363
rect 15182 2329 15200 2363
rect 15136 2323 15200 2329
rect 15194 2320 15200 2323
rect 15252 2320 15258 2372
rect 15378 2320 15384 2372
rect 15436 2360 15442 2372
rect 15933 2363 15991 2369
rect 15933 2360 15945 2363
rect 15436 2332 15945 2360
rect 15436 2320 15442 2332
rect 15933 2329 15945 2332
rect 15979 2360 15991 2363
rect 16298 2360 16304 2372
rect 15979 2332 16304 2360
rect 15979 2329 15991 2332
rect 15933 2323 15991 2329
rect 16298 2320 16304 2332
rect 16356 2320 16362 2372
rect 16390 2320 16396 2372
rect 16448 2360 16454 2372
rect 16448 2332 16514 2360
rect 16448 2320 16454 2332
rect 17402 2320 17408 2372
rect 17460 2360 17466 2372
rect 17681 2363 17739 2369
rect 17681 2360 17693 2363
rect 17460 2332 17693 2360
rect 17460 2320 17466 2332
rect 17681 2329 17693 2332
rect 17727 2329 17739 2363
rect 17681 2323 17739 2329
rect 8260 2264 8708 2292
rect 8757 2295 8815 2301
rect 8260 2252 8266 2264
rect 8757 2261 8769 2295
rect 8803 2292 8815 2295
rect 9122 2292 9128 2304
rect 8803 2264 9128 2292
rect 8803 2261 8815 2264
rect 8757 2255 8815 2261
rect 9122 2252 9128 2264
rect 9180 2252 9186 2304
rect 12710 2292 12716 2304
rect 12671 2264 12716 2292
rect 12710 2252 12716 2264
rect 12768 2252 12774 2304
rect 14001 2295 14059 2301
rect 14001 2261 14013 2295
rect 14047 2292 14059 2295
rect 14366 2292 14372 2304
rect 14047 2264 14372 2292
rect 14047 2261 14059 2264
rect 14001 2255 14059 2261
rect 14366 2252 14372 2264
rect 14424 2252 14430 2304
rect 15746 2292 15752 2304
rect 15707 2264 15752 2292
rect 15746 2252 15752 2264
rect 15804 2252 15810 2304
rect 16022 2252 16028 2304
rect 16080 2292 16086 2304
rect 18325 2295 18383 2301
rect 18325 2292 18337 2295
rect 16080 2264 18337 2292
rect 16080 2252 16086 2264
rect 18325 2261 18337 2264
rect 18371 2261 18383 2295
rect 18325 2255 18383 2261
rect 0 2202 18860 2224
rect 0 2150 4660 2202
rect 4712 2150 4724 2202
rect 4776 2150 4788 2202
rect 4840 2150 4852 2202
rect 4904 2150 4916 2202
rect 4968 2150 7760 2202
rect 7812 2150 7824 2202
rect 7876 2150 7888 2202
rect 7940 2150 7952 2202
rect 8004 2150 8016 2202
rect 8068 2150 10860 2202
rect 10912 2150 10924 2202
rect 10976 2150 10988 2202
rect 11040 2150 11052 2202
rect 11104 2150 11116 2202
rect 11168 2150 13960 2202
rect 14012 2150 14024 2202
rect 14076 2150 14088 2202
rect 14140 2150 14152 2202
rect 14204 2150 14216 2202
rect 14268 2150 17060 2202
rect 17112 2150 17124 2202
rect 17176 2150 17188 2202
rect 17240 2150 17252 2202
rect 17304 2150 17316 2202
rect 17368 2150 18860 2202
rect 0 2128 18860 2150
rect 3510 2088 3516 2100
rect 3471 2060 3516 2088
rect 3510 2048 3516 2060
rect 3568 2048 3574 2100
rect 3694 2088 3700 2100
rect 3655 2060 3700 2088
rect 3694 2048 3700 2060
rect 3752 2048 3758 2100
rect 4338 2088 4344 2100
rect 4299 2060 4344 2088
rect 4338 2048 4344 2060
rect 4396 2048 4402 2100
rect 5902 2048 5908 2100
rect 5960 2088 5966 2100
rect 6457 2091 6515 2097
rect 6457 2088 6469 2091
rect 5960 2060 6469 2088
rect 5960 2048 5966 2060
rect 6457 2057 6469 2060
rect 6503 2088 6515 2091
rect 7282 2088 7288 2100
rect 6503 2060 7288 2088
rect 6503 2057 6515 2060
rect 6457 2051 6515 2057
rect 7282 2048 7288 2060
rect 7340 2048 7346 2100
rect 8662 2048 8668 2100
rect 8720 2088 8726 2100
rect 9125 2091 9183 2097
rect 9125 2088 9137 2091
rect 8720 2060 9137 2088
rect 8720 2048 8726 2060
rect 9125 2057 9137 2060
rect 9171 2057 9183 2091
rect 9125 2051 9183 2057
rect 9861 2091 9919 2097
rect 9861 2057 9873 2091
rect 9907 2088 9919 2091
rect 10505 2091 10563 2097
rect 10505 2088 10517 2091
rect 9907 2060 10517 2088
rect 9907 2057 9919 2060
rect 9861 2051 9919 2057
rect 10505 2057 10517 2060
rect 10551 2057 10563 2091
rect 10505 2051 10563 2057
rect 10965 2091 11023 2097
rect 10965 2057 10977 2091
rect 11011 2088 11023 2091
rect 11606 2088 11612 2100
rect 11011 2060 11612 2088
rect 11011 2057 11023 2060
rect 10965 2051 11023 2057
rect 4430 2020 4436 2032
rect 3712 1992 4436 2020
rect 3602 1952 3608 1964
rect 3563 1924 3608 1952
rect 3602 1912 3608 1924
rect 3660 1912 3666 1964
rect 3712 1961 3740 1992
rect 4430 1980 4436 1992
rect 4488 1980 4494 2032
rect 5258 1980 5264 2032
rect 5316 2020 5322 2032
rect 9030 2020 9036 2032
rect 5316 1992 6592 2020
rect 8878 1992 9036 2020
rect 5316 1980 5322 1992
rect 3697 1955 3755 1961
rect 3697 1921 3709 1955
rect 3743 1921 3755 1955
rect 3697 1915 3755 1921
rect 3881 1955 3939 1961
rect 3881 1921 3893 1955
rect 3927 1952 3939 1955
rect 3927 1924 4016 1952
rect 3927 1921 3939 1924
rect 3881 1915 3939 1921
rect 3988 1825 4016 1924
rect 5166 1912 5172 1964
rect 5224 1952 5230 1964
rect 5445 1955 5503 1961
rect 5445 1952 5457 1955
rect 5224 1924 5457 1952
rect 5224 1912 5230 1924
rect 5445 1921 5457 1924
rect 5491 1921 5503 1955
rect 6365 1955 6423 1961
rect 6365 1952 6377 1955
rect 5445 1915 5503 1921
rect 5828 1924 6377 1952
rect 4433 1887 4491 1893
rect 4433 1853 4445 1887
rect 4479 1853 4491 1887
rect 4433 1847 4491 1853
rect 3973 1819 4031 1825
rect 3973 1785 3985 1819
rect 4019 1785 4031 1819
rect 4448 1816 4476 1847
rect 4522 1844 4528 1896
rect 4580 1884 4586 1896
rect 5534 1884 5540 1896
rect 4580 1856 4625 1884
rect 5495 1856 5540 1884
rect 4580 1844 4586 1856
rect 5534 1844 5540 1856
rect 5592 1844 5598 1896
rect 5828 1893 5856 1924
rect 6365 1921 6377 1924
rect 6411 1921 6423 1955
rect 6365 1915 6423 1921
rect 6564 1893 6592 1992
rect 9030 1980 9036 1992
rect 9088 1980 9094 2032
rect 10980 2020 11008 2051
rect 11606 2048 11612 2060
rect 11664 2048 11670 2100
rect 12250 2088 12256 2100
rect 12211 2060 12256 2088
rect 12250 2048 12256 2060
rect 12308 2048 12314 2100
rect 12710 2088 12716 2100
rect 12406 2060 12716 2088
rect 9140 1992 11008 2020
rect 7374 1952 7380 1964
rect 7335 1924 7380 1952
rect 7374 1912 7380 1924
rect 7432 1912 7438 1964
rect 5813 1887 5871 1893
rect 5813 1853 5825 1887
rect 5859 1853 5871 1887
rect 5813 1847 5871 1853
rect 6549 1887 6607 1893
rect 6549 1853 6561 1887
rect 6595 1853 6607 1887
rect 7650 1884 7656 1896
rect 7611 1856 7656 1884
rect 6549 1847 6607 1853
rect 7650 1844 7656 1856
rect 7708 1844 7714 1896
rect 5626 1816 5632 1828
rect 4448 1788 5632 1816
rect 3973 1779 4031 1785
rect 5626 1776 5632 1788
rect 5684 1776 5690 1828
rect 5994 1748 6000 1760
rect 5955 1720 6000 1748
rect 5994 1708 6000 1720
rect 6052 1708 6058 1760
rect 7282 1708 7288 1760
rect 7340 1748 7346 1760
rect 9140 1748 9168 1992
rect 10870 1952 10876 1964
rect 10831 1924 10876 1952
rect 10870 1912 10876 1924
rect 10928 1912 10934 1964
rect 12406 1961 12434 2060
rect 12710 2048 12716 2060
rect 12768 2088 12774 2100
rect 13081 2091 13139 2097
rect 12768 2060 13032 2088
rect 12768 2048 12774 2060
rect 13004 2020 13032 2060
rect 13081 2057 13093 2091
rect 13127 2088 13139 2091
rect 13170 2088 13176 2100
rect 13127 2060 13176 2088
rect 13127 2057 13139 2060
rect 13081 2051 13139 2057
rect 13170 2048 13176 2060
rect 13228 2048 13234 2100
rect 14277 2091 14335 2097
rect 14277 2057 14289 2091
rect 14323 2088 14335 2091
rect 14550 2088 14556 2100
rect 14323 2060 14556 2088
rect 14323 2057 14335 2060
rect 14277 2051 14335 2057
rect 14550 2048 14556 2060
rect 14608 2048 14614 2100
rect 14829 2091 14887 2097
rect 14829 2057 14841 2091
rect 14875 2088 14887 2091
rect 15562 2088 15568 2100
rect 14875 2060 15568 2088
rect 14875 2057 14887 2060
rect 14829 2051 14887 2057
rect 15562 2048 15568 2060
rect 15620 2048 15626 2100
rect 17402 2088 17408 2100
rect 17363 2060 17408 2088
rect 17402 2048 17408 2060
rect 17460 2048 17466 2100
rect 13004 1992 13308 2020
rect 12406 1955 12483 1961
rect 12406 1924 12437 1955
rect 12425 1921 12437 1924
rect 12471 1921 12483 1955
rect 12425 1915 12483 1921
rect 12529 1955 12587 1961
rect 12529 1921 12541 1955
rect 12575 1921 12587 1955
rect 12529 1915 12587 1921
rect 12621 1955 12679 1961
rect 12621 1921 12633 1955
rect 12667 1950 12679 1955
rect 12805 1955 12863 1961
rect 12667 1922 12756 1950
rect 12667 1921 12679 1922
rect 12621 1915 12679 1921
rect 9953 1887 10011 1893
rect 9953 1853 9965 1887
rect 9999 1853 10011 1887
rect 9953 1847 10011 1853
rect 10137 1887 10195 1893
rect 10137 1853 10149 1887
rect 10183 1884 10195 1887
rect 10318 1884 10324 1896
rect 10183 1856 10324 1884
rect 10183 1853 10195 1856
rect 10137 1847 10195 1853
rect 7340 1720 9168 1748
rect 7340 1708 7346 1720
rect 9214 1708 9220 1760
rect 9272 1748 9278 1760
rect 9493 1751 9551 1757
rect 9493 1748 9505 1751
rect 9272 1720 9505 1748
rect 9272 1708 9278 1720
rect 9493 1717 9505 1720
rect 9539 1717 9551 1751
rect 9968 1748 9996 1847
rect 10318 1844 10324 1856
rect 10376 1844 10382 1896
rect 11149 1887 11207 1893
rect 11149 1853 11161 1887
rect 11195 1884 11207 1887
rect 11330 1884 11336 1896
rect 11195 1856 11336 1884
rect 11195 1853 11207 1856
rect 11149 1847 11207 1853
rect 11330 1844 11336 1856
rect 11388 1844 11394 1896
rect 12544 1816 12572 1915
rect 12728 1884 12756 1922
rect 12805 1921 12817 1955
rect 12851 1952 12863 1955
rect 12894 1952 12900 1964
rect 12851 1924 12900 1952
rect 12851 1921 12863 1924
rect 12805 1915 12863 1921
rect 12894 1912 12900 1924
rect 12952 1912 12958 1964
rect 12986 1912 12992 1964
rect 13044 1952 13050 1964
rect 13280 1961 13308 1992
rect 13814 1980 13820 2032
rect 13872 2020 13878 2032
rect 15378 2020 15384 2032
rect 13872 1992 15384 2020
rect 13872 1980 13878 1992
rect 13265 1955 13323 1961
rect 13044 1924 13089 1952
rect 13044 1912 13050 1924
rect 13265 1921 13277 1955
rect 13311 1921 13323 1955
rect 13265 1915 13323 1921
rect 14093 1955 14151 1961
rect 14093 1921 14105 1955
rect 14139 1952 14151 1955
rect 14185 1955 14243 1961
rect 14185 1952 14197 1955
rect 14139 1924 14197 1952
rect 14139 1921 14151 1924
rect 14093 1915 14151 1921
rect 14185 1921 14197 1924
rect 14231 1921 14243 1955
rect 14366 1952 14372 1964
rect 14327 1924 14372 1952
rect 14185 1915 14243 1921
rect 13004 1884 13032 1912
rect 12728 1856 13032 1884
rect 14200 1884 14228 1915
rect 14366 1912 14372 1924
rect 14424 1952 14430 1964
rect 15120 1961 15148 1992
rect 15378 1980 15384 1992
rect 15436 1980 15442 2032
rect 15838 2020 15844 2032
rect 15672 1992 15844 2020
rect 15672 1961 15700 1992
rect 15838 1980 15844 1992
rect 15896 1980 15902 2032
rect 15933 2023 15991 2029
rect 15933 1989 15945 2023
rect 15979 2020 15991 2023
rect 16022 2020 16028 2032
rect 15979 1992 16028 2020
rect 15979 1989 15991 1992
rect 15933 1983 15991 1989
rect 16022 1980 16028 1992
rect 16080 1980 16086 2032
rect 16390 1980 16396 2032
rect 16448 1980 16454 2032
rect 14645 1955 14703 1961
rect 14645 1952 14657 1955
rect 14424 1924 14657 1952
rect 14424 1912 14430 1924
rect 14645 1921 14657 1924
rect 14691 1921 14703 1955
rect 14645 1915 14703 1921
rect 15105 1955 15163 1961
rect 15105 1921 15117 1955
rect 15151 1921 15163 1955
rect 15105 1915 15163 1921
rect 15657 1955 15715 1961
rect 15657 1921 15669 1955
rect 15703 1921 15715 1955
rect 15657 1915 15715 1921
rect 14461 1887 14519 1893
rect 14461 1884 14473 1887
rect 14200 1856 14473 1884
rect 14461 1853 14473 1856
rect 14507 1884 14519 1887
rect 15194 1884 15200 1896
rect 14507 1856 15200 1884
rect 14507 1853 14519 1856
rect 14461 1847 14519 1853
rect 15194 1844 15200 1856
rect 15252 1884 15258 1896
rect 15381 1887 15439 1893
rect 15381 1884 15393 1887
rect 15252 1856 15393 1884
rect 15252 1844 15258 1856
rect 15381 1853 15393 1856
rect 15427 1853 15439 1887
rect 15381 1847 15439 1853
rect 14921 1819 14979 1825
rect 14921 1816 14933 1819
rect 12544 1788 14933 1816
rect 14921 1785 14933 1788
rect 14967 1816 14979 1819
rect 15654 1816 15660 1828
rect 14967 1788 15660 1816
rect 14967 1785 14979 1788
rect 14921 1779 14979 1785
rect 15654 1776 15660 1788
rect 15712 1776 15718 1828
rect 14093 1751 14151 1757
rect 14093 1748 14105 1751
rect 9968 1720 14105 1748
rect 9493 1711 9551 1717
rect 14093 1717 14105 1720
rect 14139 1717 14151 1751
rect 14093 1711 14151 1717
rect 15289 1751 15347 1757
rect 15289 1717 15301 1751
rect 15335 1748 15347 1751
rect 16942 1748 16948 1760
rect 15335 1720 16948 1748
rect 15335 1717 15347 1720
rect 15289 1711 15347 1717
rect 16942 1708 16948 1720
rect 17000 1708 17006 1760
rect 0 1658 18860 1680
rect 0 1606 3110 1658
rect 3162 1606 3174 1658
rect 3226 1606 3238 1658
rect 3290 1606 3302 1658
rect 3354 1606 3366 1658
rect 3418 1606 6210 1658
rect 6262 1606 6274 1658
rect 6326 1606 6338 1658
rect 6390 1606 6402 1658
rect 6454 1606 6466 1658
rect 6518 1606 9310 1658
rect 9362 1606 9374 1658
rect 9426 1606 9438 1658
rect 9490 1606 9502 1658
rect 9554 1606 9566 1658
rect 9618 1606 12410 1658
rect 12462 1606 12474 1658
rect 12526 1606 12538 1658
rect 12590 1606 12602 1658
rect 12654 1606 12666 1658
rect 12718 1606 15510 1658
rect 15562 1606 15574 1658
rect 15626 1606 15638 1658
rect 15690 1606 15702 1658
rect 15754 1606 15766 1658
rect 15818 1606 18860 1658
rect 0 1584 18860 1606
rect 2961 1547 3019 1553
rect 2961 1513 2973 1547
rect 3007 1544 3019 1547
rect 3878 1544 3884 1556
rect 3007 1516 3884 1544
rect 3007 1513 3019 1516
rect 2961 1507 3019 1513
rect 3878 1504 3884 1516
rect 3936 1504 3942 1556
rect 5534 1544 5540 1556
rect 5495 1516 5540 1544
rect 5534 1504 5540 1516
rect 5592 1504 5598 1556
rect 10597 1547 10655 1553
rect 10597 1513 10609 1547
rect 10643 1544 10655 1547
rect 10870 1544 10876 1556
rect 10643 1516 10876 1544
rect 10643 1513 10655 1516
rect 10597 1507 10655 1513
rect 10870 1504 10876 1516
rect 10928 1504 10934 1556
rect 2869 1479 2927 1485
rect 2869 1476 2881 1479
rect 2056 1448 2881 1476
rect 750 1408 756 1420
rect 711 1380 756 1408
rect 750 1368 756 1380
rect 808 1368 814 1420
rect 1029 1411 1087 1417
rect 1029 1377 1041 1411
rect 1075 1408 1087 1411
rect 2056 1408 2084 1448
rect 2869 1445 2881 1448
rect 2915 1445 2927 1479
rect 2869 1439 2927 1445
rect 3513 1479 3571 1485
rect 3513 1445 3525 1479
rect 3559 1476 3571 1479
rect 5718 1476 5724 1488
rect 3559 1448 5724 1476
rect 3559 1445 3571 1448
rect 3513 1439 3571 1445
rect 5718 1436 5724 1448
rect 5776 1436 5782 1488
rect 8662 1436 8668 1488
rect 8720 1476 8726 1488
rect 8720 1448 9628 1476
rect 8720 1436 8726 1448
rect 1075 1380 2084 1408
rect 2777 1411 2835 1417
rect 1075 1377 1087 1380
rect 1029 1371 1087 1377
rect 2777 1377 2789 1411
rect 2823 1408 2835 1411
rect 3973 1411 4031 1417
rect 3973 1408 3985 1411
rect 2823 1380 3985 1408
rect 2823 1377 2835 1380
rect 2777 1371 2835 1377
rect 3973 1377 3985 1380
rect 4019 1377 4031 1411
rect 3973 1371 4031 1377
rect 5000 1380 5304 1408
rect 3053 1343 3111 1349
rect 3053 1309 3065 1343
rect 3099 1340 3111 1343
rect 3513 1343 3571 1349
rect 3513 1340 3525 1343
rect 3099 1312 3525 1340
rect 3099 1309 3111 1312
rect 3053 1303 3111 1309
rect 3513 1309 3525 1312
rect 3559 1340 3571 1343
rect 3697 1343 3755 1349
rect 3697 1340 3709 1343
rect 3559 1312 3709 1340
rect 3559 1309 3571 1312
rect 3513 1303 3571 1309
rect 3697 1309 3709 1312
rect 3743 1309 3755 1343
rect 3697 1303 3755 1309
rect 3789 1343 3847 1349
rect 3789 1309 3801 1343
rect 3835 1309 3847 1343
rect 3789 1303 3847 1309
rect 2682 1272 2688 1284
rect 2254 1244 2688 1272
rect 2682 1232 2688 1244
rect 2740 1232 2746 1284
rect 2958 1232 2964 1284
rect 3016 1272 3022 1284
rect 3237 1275 3295 1281
rect 3237 1272 3249 1275
rect 3016 1244 3249 1272
rect 3016 1232 3022 1244
rect 3237 1241 3249 1244
rect 3283 1241 3295 1275
rect 3418 1272 3424 1284
rect 3379 1244 3424 1272
rect 3237 1235 3295 1241
rect 3418 1232 3424 1244
rect 3476 1232 3482 1284
rect 2501 1207 2559 1213
rect 2501 1173 2513 1207
rect 2547 1204 2559 1207
rect 3804 1204 3832 1303
rect 3878 1300 3884 1352
rect 3936 1340 3942 1352
rect 4065 1343 4123 1349
rect 3936 1312 3981 1340
rect 3936 1300 3942 1312
rect 4065 1309 4077 1343
rect 4111 1309 4123 1343
rect 4065 1303 4123 1309
rect 4080 1272 4108 1303
rect 4154 1300 4160 1352
rect 4212 1340 4218 1352
rect 5000 1349 5028 1380
rect 4433 1343 4491 1349
rect 4433 1340 4445 1343
rect 4212 1312 4445 1340
rect 4212 1300 4218 1312
rect 4433 1309 4445 1312
rect 4479 1309 4491 1343
rect 4433 1303 4491 1309
rect 4985 1343 5043 1349
rect 4985 1309 4997 1343
rect 5031 1309 5043 1343
rect 4985 1303 5043 1309
rect 5074 1300 5080 1352
rect 5132 1342 5138 1352
rect 5169 1343 5227 1349
rect 5169 1342 5181 1343
rect 5132 1314 5181 1342
rect 5132 1300 5138 1314
rect 5169 1309 5181 1314
rect 5215 1309 5227 1343
rect 5276 1340 5304 1380
rect 5902 1368 5908 1420
rect 5960 1408 5966 1420
rect 6089 1411 6147 1417
rect 6089 1408 6101 1411
rect 5960 1380 6101 1408
rect 5960 1368 5966 1380
rect 6089 1377 6101 1380
rect 6135 1377 6147 1411
rect 6089 1371 6147 1377
rect 6273 1411 6331 1417
rect 6273 1377 6285 1411
rect 6319 1377 6331 1411
rect 6273 1371 6331 1377
rect 8757 1411 8815 1417
rect 8757 1377 8769 1411
rect 8803 1408 8815 1411
rect 9214 1408 9220 1420
rect 8803 1380 9220 1408
rect 8803 1377 8815 1380
rect 8757 1371 8815 1377
rect 5350 1340 5356 1352
rect 5276 1312 5356 1340
rect 5169 1303 5227 1309
rect 5350 1300 5356 1312
rect 5408 1300 5414 1352
rect 5534 1340 5540 1352
rect 5495 1312 5540 1340
rect 5534 1300 5540 1312
rect 5592 1300 5598 1352
rect 5994 1340 6000 1352
rect 5955 1312 6000 1340
rect 5994 1300 6000 1312
rect 6052 1300 6058 1352
rect 6288 1272 6316 1371
rect 9214 1368 9220 1380
rect 9272 1368 9278 1420
rect 6457 1343 6515 1349
rect 6457 1309 6469 1343
rect 6503 1340 6515 1343
rect 6546 1340 6552 1352
rect 6503 1312 6552 1340
rect 6503 1309 6515 1312
rect 6457 1303 6515 1309
rect 6546 1300 6552 1312
rect 6604 1300 6610 1352
rect 7650 1300 7656 1352
rect 7708 1340 7714 1352
rect 8481 1343 8539 1349
rect 8481 1340 8493 1343
rect 7708 1312 8493 1340
rect 7708 1300 7714 1312
rect 8481 1309 8493 1312
rect 8527 1309 8539 1343
rect 8662 1340 8668 1352
rect 8623 1312 8668 1340
rect 8481 1303 8539 1309
rect 8662 1300 8668 1312
rect 8720 1300 8726 1352
rect 9122 1340 9128 1352
rect 9083 1312 9128 1340
rect 9122 1300 9128 1312
rect 9180 1300 9186 1352
rect 9600 1340 9628 1448
rect 10134 1408 10140 1420
rect 10095 1380 10140 1408
rect 10134 1368 10140 1380
rect 10192 1368 10198 1420
rect 11072 1380 11284 1408
rect 10229 1343 10287 1349
rect 10229 1340 10241 1343
rect 9600 1312 10241 1340
rect 10229 1309 10241 1312
rect 10275 1340 10287 1343
rect 11072 1340 11100 1380
rect 11256 1349 11284 1380
rect 11330 1368 11336 1420
rect 11388 1408 11394 1420
rect 14093 1411 14151 1417
rect 14093 1408 14105 1411
rect 11388 1380 14105 1408
rect 11388 1368 11394 1380
rect 12636 1349 12664 1380
rect 14093 1377 14105 1380
rect 14139 1377 14151 1411
rect 16482 1408 16488 1420
rect 16443 1380 16488 1408
rect 14093 1371 14151 1377
rect 16482 1368 16488 1380
rect 16540 1408 16546 1420
rect 16577 1411 16635 1417
rect 16577 1408 16589 1411
rect 16540 1380 16589 1408
rect 16540 1368 16546 1380
rect 16577 1377 16589 1380
rect 16623 1377 16635 1411
rect 16577 1371 16635 1377
rect 10275 1312 11100 1340
rect 11149 1343 11207 1349
rect 10275 1309 10287 1312
rect 10229 1303 10287 1309
rect 11149 1309 11161 1343
rect 11195 1309 11207 1343
rect 11149 1303 11207 1309
rect 11241 1343 11299 1349
rect 11241 1309 11253 1343
rect 11287 1309 11299 1343
rect 11241 1303 11299 1309
rect 12621 1343 12679 1349
rect 12621 1309 12633 1343
rect 12667 1309 12679 1343
rect 12621 1303 12679 1309
rect 12713 1343 12771 1349
rect 12713 1309 12725 1343
rect 12759 1340 12771 1343
rect 12986 1340 12992 1352
rect 12759 1312 12992 1340
rect 12759 1309 12771 1312
rect 12713 1303 12771 1309
rect 6638 1272 6644 1284
rect 4080 1244 5672 1272
rect 6288 1244 6644 1272
rect 5074 1204 5080 1216
rect 2547 1176 5080 1204
rect 2547 1173 2559 1176
rect 2501 1167 2559 1173
rect 5074 1164 5080 1176
rect 5132 1164 5138 1216
rect 5169 1207 5227 1213
rect 5169 1173 5181 1207
rect 5215 1204 5227 1207
rect 5258 1204 5264 1216
rect 5215 1176 5264 1204
rect 5215 1173 5227 1176
rect 5169 1167 5227 1173
rect 5258 1164 5264 1176
rect 5316 1164 5322 1216
rect 5644 1213 5672 1244
rect 6638 1232 6644 1244
rect 6696 1272 6702 1284
rect 10318 1272 10324 1284
rect 6696 1244 10324 1272
rect 6696 1232 6702 1244
rect 10318 1232 10324 1244
rect 10376 1232 10382 1284
rect 10778 1232 10784 1284
rect 10836 1272 10842 1284
rect 10873 1275 10931 1281
rect 10873 1272 10885 1275
rect 10836 1244 10885 1272
rect 10836 1232 10842 1244
rect 10873 1241 10885 1244
rect 10919 1241 10931 1275
rect 11054 1272 11060 1284
rect 11015 1244 11060 1272
rect 10873 1235 10931 1241
rect 11054 1232 11060 1244
rect 11112 1232 11118 1284
rect 11164 1272 11192 1303
rect 11333 1275 11391 1281
rect 11333 1272 11345 1275
rect 11164 1244 11345 1272
rect 11333 1241 11345 1244
rect 11379 1241 11391 1275
rect 12728 1272 12756 1303
rect 12986 1300 12992 1312
rect 13044 1300 13050 1352
rect 13814 1300 13820 1352
rect 13872 1340 13878 1352
rect 14001 1343 14059 1349
rect 14001 1340 14013 1343
rect 13872 1312 14013 1340
rect 13872 1300 13878 1312
rect 14001 1309 14013 1312
rect 14047 1309 14059 1343
rect 18230 1340 18236 1352
rect 18191 1312 18236 1340
rect 14001 1303 14059 1309
rect 18230 1300 18236 1312
rect 18288 1300 18294 1352
rect 18322 1300 18328 1352
rect 18380 1340 18386 1352
rect 18380 1312 18425 1340
rect 18380 1300 18386 1312
rect 14458 1272 14464 1284
rect 11333 1235 11391 1241
rect 12406 1244 12756 1272
rect 14419 1244 14464 1272
rect 5629 1207 5687 1213
rect 5629 1173 5641 1207
rect 5675 1173 5687 1207
rect 6914 1204 6920 1216
rect 6875 1176 6920 1204
rect 5629 1167 5687 1173
rect 6914 1164 6920 1176
rect 6972 1164 6978 1216
rect 11149 1207 11207 1213
rect 11149 1173 11161 1207
rect 11195 1204 11207 1207
rect 12406 1204 12434 1244
rect 14458 1232 14464 1244
rect 14516 1232 14522 1284
rect 14918 1232 14924 1284
rect 14976 1272 14982 1284
rect 16206 1272 16212 1284
rect 14976 1258 15042 1272
rect 14976 1244 15056 1258
rect 16167 1244 16212 1272
rect 14976 1232 14982 1244
rect 11195 1176 12434 1204
rect 13541 1207 13599 1213
rect 11195 1173 11207 1176
rect 11149 1167 11207 1173
rect 13541 1173 13553 1207
rect 13587 1204 13599 1207
rect 13630 1204 13636 1216
rect 13587 1176 13636 1204
rect 13587 1173 13599 1176
rect 13541 1167 13599 1173
rect 13630 1164 13636 1176
rect 13688 1164 13694 1216
rect 13909 1207 13967 1213
rect 13909 1173 13921 1207
rect 13955 1204 13967 1207
rect 14366 1204 14372 1216
rect 13955 1176 14372 1204
rect 13955 1173 13967 1176
rect 13909 1167 13967 1173
rect 14366 1164 14372 1176
rect 14424 1164 14430 1216
rect 15028 1204 15056 1244
rect 16206 1232 16212 1244
rect 16264 1232 16270 1284
rect 16298 1232 16304 1284
rect 16356 1272 16362 1284
rect 16822 1275 16880 1281
rect 16822 1272 16834 1275
rect 16356 1244 16834 1272
rect 16356 1232 16362 1244
rect 16822 1241 16834 1244
rect 16868 1241 16880 1275
rect 16822 1235 16880 1241
rect 16390 1204 16396 1216
rect 15028 1176 16396 1204
rect 16390 1164 16396 1176
rect 16448 1164 16454 1216
rect 17954 1204 17960 1216
rect 17915 1176 17960 1204
rect 17954 1164 17960 1176
rect 18012 1164 18018 1216
rect 0 1114 18860 1136
rect 0 1062 4660 1114
rect 4712 1062 4724 1114
rect 4776 1062 4788 1114
rect 4840 1062 4852 1114
rect 4904 1062 4916 1114
rect 4968 1062 7760 1114
rect 7812 1062 7824 1114
rect 7876 1062 7888 1114
rect 7940 1062 7952 1114
rect 8004 1062 8016 1114
rect 8068 1062 10860 1114
rect 10912 1062 10924 1114
rect 10976 1062 10988 1114
rect 11040 1062 11052 1114
rect 11104 1062 11116 1114
rect 11168 1062 13960 1114
rect 14012 1062 14024 1114
rect 14076 1062 14088 1114
rect 14140 1062 14152 1114
rect 14204 1062 14216 1114
rect 14268 1062 17060 1114
rect 17112 1062 17124 1114
rect 17176 1062 17188 1114
rect 17240 1062 17252 1114
rect 17304 1062 17316 1114
rect 17368 1062 18860 1114
rect 0 1040 18860 1062
rect 4062 960 4068 1012
rect 4120 1000 4126 1012
rect 5534 1000 5540 1012
rect 4120 972 5540 1000
rect 4120 960 4126 972
rect 5534 960 5540 972
rect 5592 960 5598 1012
rect 5813 1003 5871 1009
rect 5813 969 5825 1003
rect 5859 1000 5871 1003
rect 6365 1003 6423 1009
rect 6365 1000 6377 1003
rect 5859 972 6377 1000
rect 5859 969 5871 972
rect 5813 963 5871 969
rect 6365 969 6377 972
rect 6411 969 6423 1003
rect 6365 963 6423 969
rect 6457 1003 6515 1009
rect 6457 969 6469 1003
rect 6503 1000 6515 1003
rect 6546 1000 6552 1012
rect 6503 972 6552 1000
rect 6503 969 6515 972
rect 6457 963 6515 969
rect 6546 960 6552 972
rect 6604 960 6610 1012
rect 8938 960 8944 1012
rect 8996 1000 9002 1012
rect 9585 1003 9643 1009
rect 9585 1000 9597 1003
rect 8996 972 9597 1000
rect 8996 960 9002 972
rect 9585 969 9597 972
rect 9631 1000 9643 1003
rect 9953 1003 10011 1009
rect 9953 1000 9965 1003
rect 9631 972 9965 1000
rect 9631 969 9643 972
rect 9585 963 9643 969
rect 9953 969 9965 972
rect 9999 969 10011 1003
rect 10134 1000 10140 1012
rect 10095 972 10140 1000
rect 9953 963 10011 969
rect 10134 960 10140 972
rect 10192 960 10198 1012
rect 10505 1003 10563 1009
rect 10505 969 10517 1003
rect 10551 969 10563 1003
rect 10505 963 10563 969
rect 3896 904 5488 932
rect 3237 867 3295 873
rect 3237 833 3249 867
rect 3283 864 3295 867
rect 3418 864 3424 876
rect 3283 836 3424 864
rect 3283 833 3295 836
rect 3237 827 3295 833
rect 3418 824 3424 836
rect 3476 864 3482 876
rect 3896 873 3924 904
rect 5460 876 5488 904
rect 3789 867 3847 873
rect 3789 864 3801 867
rect 3476 836 3801 864
rect 3476 824 3482 836
rect 3789 833 3801 836
rect 3835 833 3847 867
rect 3789 827 3847 833
rect 3881 867 3939 873
rect 3881 833 3893 867
rect 3927 833 3939 867
rect 3881 827 3939 833
rect 3970 824 3976 876
rect 4028 864 4034 876
rect 4154 864 4160 876
rect 4028 836 4073 864
rect 4115 836 4160 864
rect 4028 824 4034 836
rect 4154 824 4160 836
rect 4212 824 4218 876
rect 5442 864 5448 876
rect 5403 836 5448 864
rect 5442 824 5448 836
rect 5500 824 5506 876
rect 5552 805 5580 960
rect 9030 932 9036 944
rect 8602 904 9036 932
rect 9030 892 9036 904
rect 9088 892 9094 944
rect 9493 935 9551 941
rect 9493 901 9505 935
rect 9539 932 9551 935
rect 10520 932 10548 963
rect 11238 960 11244 1012
rect 11296 1000 11302 1012
rect 11425 1003 11483 1009
rect 11425 1000 11437 1003
rect 11296 972 11437 1000
rect 11296 960 11302 972
rect 11425 969 11437 972
rect 11471 969 11483 1003
rect 11425 963 11483 969
rect 12437 1003 12495 1009
rect 12437 969 12449 1003
rect 12483 1000 12495 1003
rect 12529 1003 12587 1009
rect 12529 1000 12541 1003
rect 12483 972 12541 1000
rect 12483 969 12495 972
rect 12437 963 12495 969
rect 12529 969 12541 972
rect 12575 969 12587 1003
rect 13630 1000 13636 1012
rect 12529 963 12587 969
rect 12820 972 13492 1000
rect 13591 972 13636 1000
rect 10778 932 10784 944
rect 9539 904 10548 932
rect 10612 904 10784 932
rect 9539 901 9551 904
rect 9493 895 9551 901
rect 10045 867 10103 873
rect 10045 864 10057 867
rect 9692 836 10057 864
rect 2961 799 3019 805
rect 2961 765 2973 799
rect 3007 796 3019 799
rect 4065 799 4123 805
rect 4065 796 4077 799
rect 3007 768 4077 796
rect 3007 765 3019 768
rect 2961 759 3019 765
rect 4065 765 4077 768
rect 4111 765 4123 799
rect 4065 759 4123 765
rect 5537 799 5595 805
rect 5537 765 5549 799
rect 5583 765 5595 799
rect 5537 759 5595 765
rect 6549 799 6607 805
rect 6549 765 6561 799
rect 6595 765 6607 799
rect 6549 759 6607 765
rect 7193 799 7251 805
rect 7193 765 7205 799
rect 7239 796 7251 799
rect 7374 796 7380 808
rect 7239 768 7380 796
rect 7239 765 7251 768
rect 7193 759 7251 765
rect 3145 731 3203 737
rect 3145 697 3157 731
rect 3191 728 3203 731
rect 3878 728 3884 740
rect 3191 700 3884 728
rect 3191 697 3203 700
rect 3145 691 3203 697
rect 3878 688 3884 700
rect 3936 688 3942 740
rect 5258 688 5264 740
rect 5316 728 5322 740
rect 6564 728 6592 759
rect 7374 756 7380 768
rect 7432 756 7438 808
rect 7561 799 7619 805
rect 7561 765 7573 799
rect 7607 796 7619 799
rect 8110 796 8116 808
rect 7607 768 8116 796
rect 7607 765 7619 768
rect 7561 759 7619 765
rect 8110 756 8116 768
rect 8168 756 8174 808
rect 5316 700 6592 728
rect 8987 731 9045 737
rect 5316 688 5322 700
rect 8987 697 8999 731
rect 9033 728 9045 731
rect 9692 728 9720 836
rect 10045 833 10057 836
rect 10091 833 10103 867
rect 10045 827 10103 833
rect 10229 867 10287 873
rect 10229 833 10241 867
rect 10275 864 10287 867
rect 10612 864 10640 904
rect 10778 892 10784 904
rect 10836 932 10842 944
rect 12345 935 12403 941
rect 12345 932 12357 935
rect 10836 904 12357 932
rect 10836 892 10842 904
rect 12345 901 12357 904
rect 12391 932 12403 935
rect 12820 932 12848 972
rect 12391 904 12848 932
rect 13464 932 13492 972
rect 13630 960 13636 972
rect 13688 960 13694 1012
rect 13725 1003 13783 1009
rect 13725 969 13737 1003
rect 13771 1000 13783 1003
rect 13814 1000 13820 1012
rect 13771 972 13820 1000
rect 13771 969 13783 972
rect 13725 963 13783 969
rect 13814 960 13820 972
rect 13872 960 13878 1012
rect 14185 1003 14243 1009
rect 14185 969 14197 1003
rect 14231 1000 14243 1003
rect 14366 1000 14372 1012
rect 14231 972 14372 1000
rect 14231 969 14243 972
rect 14185 963 14243 969
rect 14366 960 14372 972
rect 14424 960 14430 1012
rect 16025 1003 16083 1009
rect 16025 969 16037 1003
rect 16071 1000 16083 1003
rect 16206 1000 16212 1012
rect 16071 972 16212 1000
rect 16071 969 16083 972
rect 16025 963 16083 969
rect 16206 960 16212 972
rect 16264 960 16270 1012
rect 17313 1003 17371 1009
rect 17313 1000 17325 1003
rect 17052 972 17325 1000
rect 14642 932 14648 944
rect 13464 904 14648 932
rect 12391 901 12403 904
rect 12345 895 12403 901
rect 10870 864 10876 876
rect 10275 836 10640 864
rect 10831 836 10876 864
rect 10275 833 10287 836
rect 10229 827 10287 833
rect 10870 824 10876 836
rect 10928 824 10934 876
rect 11054 824 11060 876
rect 11112 864 11118 876
rect 11333 867 11391 873
rect 11333 864 11345 867
rect 11112 836 11345 864
rect 11112 824 11118 836
rect 11333 833 11345 836
rect 11379 833 11391 867
rect 12158 864 12164 876
rect 12119 836 12164 864
rect 11333 827 11391 833
rect 12158 824 12164 836
rect 12216 824 12222 876
rect 12437 867 12495 873
rect 12437 833 12449 867
rect 12483 864 12495 867
rect 12710 864 12716 876
rect 12483 836 12716 864
rect 12483 833 12495 836
rect 12437 827 12495 833
rect 12710 824 12716 836
rect 12768 824 12774 876
rect 14200 873 14228 904
rect 14642 892 14648 904
rect 14700 892 14706 944
rect 17052 932 17080 972
rect 17313 969 17325 972
rect 17359 969 17371 1003
rect 17313 963 17371 969
rect 16960 904 17080 932
rect 17221 935 17279 941
rect 16960 873 16988 904
rect 17221 901 17233 935
rect 17267 932 17279 935
rect 17954 932 17960 944
rect 17267 904 17960 932
rect 17267 901 17279 904
rect 17221 895 17279 901
rect 17954 892 17960 904
rect 18012 892 18018 944
rect 14185 867 14243 873
rect 12820 836 13676 864
rect 9769 799 9827 805
rect 9769 765 9781 799
rect 9815 796 9827 799
rect 10318 796 10324 808
rect 9815 768 10324 796
rect 9815 765 9827 768
rect 9769 759 9827 765
rect 10318 756 10324 768
rect 10376 756 10382 808
rect 10413 799 10471 805
rect 10413 765 10425 799
rect 10459 796 10471 799
rect 10962 796 10968 808
rect 10459 768 10968 796
rect 10459 765 10471 768
rect 10413 759 10471 765
rect 10962 756 10968 768
rect 11020 756 11026 808
rect 11149 799 11207 805
rect 11149 765 11161 799
rect 11195 796 11207 799
rect 12820 796 12848 836
rect 11195 768 11376 796
rect 11195 765 11207 768
rect 11149 759 11207 765
rect 11348 740 11376 768
rect 12406 768 12848 796
rect 12897 799 12955 805
rect 11054 728 11060 740
rect 9033 700 11060 728
rect 9033 697 9045 700
rect 8987 691 9045 697
rect 11054 688 11060 700
rect 11112 688 11118 740
rect 11330 688 11336 740
rect 11388 688 11394 740
rect 2958 620 2964 672
rect 3016 660 3022 672
rect 3053 663 3111 669
rect 3053 660 3065 663
rect 3016 632 3065 660
rect 3016 620 3022 632
rect 3053 629 3065 632
rect 3099 629 3111 663
rect 5994 660 6000 672
rect 5955 632 6000 660
rect 3053 623 3111 629
rect 5994 620 6000 632
rect 6052 620 6058 672
rect 9122 620 9128 672
rect 9180 660 9186 672
rect 9953 663 10011 669
rect 9180 632 9225 660
rect 9180 620 9186 632
rect 9953 629 9965 663
rect 9999 660 10011 663
rect 10413 663 10471 669
rect 10413 660 10425 663
rect 9999 632 10425 660
rect 9999 629 10011 632
rect 9953 623 10011 629
rect 10413 629 10425 632
rect 10459 629 10471 663
rect 10413 623 10471 629
rect 10502 620 10508 672
rect 10560 660 10566 672
rect 12406 660 12434 768
rect 12897 765 12909 799
rect 12943 765 12955 799
rect 12897 759 12955 765
rect 12912 728 12940 759
rect 12986 756 12992 808
rect 13044 796 13050 808
rect 13648 796 13676 836
rect 14185 833 14197 867
rect 14231 833 14243 867
rect 15841 867 15899 873
rect 15841 864 15853 867
rect 14185 827 14243 833
rect 14568 836 15853 864
rect 13863 799 13921 805
rect 13863 796 13875 799
rect 13044 768 13492 796
rect 13648 768 13875 796
rect 13044 756 13050 768
rect 13265 731 13323 737
rect 13265 728 13277 731
rect 12912 700 13277 728
rect 13265 697 13277 700
rect 13311 697 13323 731
rect 13464 728 13492 768
rect 13863 765 13875 768
rect 13909 796 13921 799
rect 14458 796 14464 808
rect 13909 768 14464 796
rect 13909 765 13921 768
rect 13863 759 13921 765
rect 14458 756 14464 768
rect 14516 756 14522 808
rect 14568 728 14596 836
rect 15841 833 15853 836
rect 15887 833 15899 867
rect 15841 827 15899 833
rect 16945 867 17003 873
rect 16945 833 16957 867
rect 16991 833 17003 867
rect 16945 827 17003 833
rect 17037 867 17095 873
rect 17037 833 17049 867
rect 17083 833 17095 867
rect 17770 864 17776 876
rect 17731 836 17776 864
rect 17037 827 17095 833
rect 15565 799 15623 805
rect 15565 765 15577 799
rect 15611 796 15623 799
rect 17052 796 17080 827
rect 17770 824 17776 836
rect 17828 824 17834 876
rect 18046 824 18052 876
rect 18104 864 18110 876
rect 18325 867 18383 873
rect 18325 864 18337 867
rect 18104 836 18337 864
rect 18104 824 18110 836
rect 18325 833 18337 836
rect 18371 833 18383 867
rect 18325 827 18383 833
rect 17865 799 17923 805
rect 17865 796 17877 799
rect 15611 768 16988 796
rect 17052 768 17877 796
rect 15611 765 15623 768
rect 15565 759 15623 765
rect 13464 700 14596 728
rect 15657 731 15715 737
rect 13265 691 13323 697
rect 15657 697 15669 731
rect 15703 728 15715 731
rect 15838 728 15844 740
rect 15703 700 15844 728
rect 15703 697 15715 700
rect 15657 691 15715 697
rect 15838 688 15844 700
rect 15896 688 15902 740
rect 16960 737 16988 768
rect 17865 765 17877 768
rect 17911 765 17923 799
rect 17865 759 17923 765
rect 16945 731 17003 737
rect 16945 697 16957 731
rect 16991 697 17003 731
rect 16945 691 17003 697
rect 17770 688 17776 740
rect 17828 728 17834 740
rect 17828 700 18092 728
rect 17828 688 17834 700
rect 13170 660 13176 672
rect 10560 632 12434 660
rect 13131 632 13176 660
rect 10560 620 10566 632
rect 13170 620 13176 632
rect 13228 620 13234 672
rect 17681 663 17739 669
rect 17681 629 17693 663
rect 17727 660 17739 663
rect 17954 660 17960 672
rect 17727 632 17960 660
rect 17727 629 17739 632
rect 17681 623 17739 629
rect 17954 620 17960 632
rect 18012 620 18018 672
rect 18064 669 18092 700
rect 18049 663 18107 669
rect 18049 629 18061 663
rect 18095 629 18107 663
rect 18049 623 18107 629
rect 0 570 18860 592
rect 0 518 3110 570
rect 3162 518 3174 570
rect 3226 518 3238 570
rect 3290 518 3302 570
rect 3354 518 3366 570
rect 3418 518 6210 570
rect 6262 518 6274 570
rect 6326 518 6338 570
rect 6390 518 6402 570
rect 6454 518 6466 570
rect 6518 518 9310 570
rect 9362 518 9374 570
rect 9426 518 9438 570
rect 9490 518 9502 570
rect 9554 518 9566 570
rect 9618 518 12410 570
rect 12462 518 12474 570
rect 12526 518 12538 570
rect 12590 518 12602 570
rect 12654 518 12666 570
rect 12718 518 15510 570
rect 15562 518 15574 570
rect 15626 518 15638 570
rect 15690 518 15702 570
rect 15754 518 15766 570
rect 15818 518 18860 570
rect 0 496 18860 518
rect 4154 416 4160 468
rect 4212 456 4218 468
rect 5629 459 5687 465
rect 5629 456 5641 459
rect 4212 428 5641 456
rect 4212 416 4218 428
rect 5629 425 5641 428
rect 5675 425 5687 459
rect 8110 456 8116 468
rect 8071 428 8116 456
rect 5629 419 5687 425
rect 8110 416 8116 428
rect 8168 416 8174 468
rect 10870 456 10876 468
rect 10831 428 10876 456
rect 10870 416 10876 428
rect 10928 416 10934 468
rect 12986 456 12992 468
rect 12406 428 12992 456
rect 4479 391 4537 397
rect 4479 357 4491 391
rect 4525 388 4537 391
rect 5442 388 5448 400
rect 4525 360 5448 388
rect 4525 357 4537 360
rect 4479 351 4537 357
rect 5442 348 5448 360
rect 5500 348 5506 400
rect 6914 388 6920 400
rect 6104 360 6920 388
rect 2958 280 2964 332
rect 3016 320 3022 332
rect 6104 329 6132 360
rect 6914 348 6920 360
rect 6972 348 6978 400
rect 8662 388 8668 400
rect 8312 360 8668 388
rect 3053 323 3111 329
rect 3053 320 3065 323
rect 3016 292 3065 320
rect 3016 280 3022 292
rect 3053 289 3065 292
rect 3099 289 3111 323
rect 3053 283 3111 289
rect 6089 323 6147 329
rect 6089 289 6101 323
rect 6135 289 6147 323
rect 6089 283 6147 289
rect 6273 323 6331 329
rect 6273 289 6285 323
rect 6319 320 6331 323
rect 6638 320 6644 332
rect 6319 292 6644 320
rect 6319 289 6331 292
rect 6273 283 6331 289
rect 6638 280 6644 292
rect 6696 280 6702 332
rect 8312 329 8340 360
rect 8662 348 8668 360
rect 8720 388 8726 400
rect 12406 388 12434 428
rect 12986 416 12992 428
rect 13044 416 13050 468
rect 14642 416 14648 468
rect 14700 456 14706 468
rect 14737 459 14795 465
rect 14737 456 14749 459
rect 14700 428 14749 456
rect 14700 416 14706 428
rect 14737 425 14749 428
rect 14783 425 14795 459
rect 16482 456 16488 468
rect 14737 419 14795 425
rect 16132 428 16488 456
rect 8720 360 12434 388
rect 8720 348 8726 360
rect 8297 323 8355 329
rect 8297 289 8309 323
rect 8343 289 8355 323
rect 8297 283 8355 289
rect 8389 323 8447 329
rect 8389 289 8401 323
rect 8435 320 8447 323
rect 9122 320 9128 332
rect 8435 292 9128 320
rect 8435 289 8447 292
rect 8389 283 8447 289
rect 9122 280 9128 292
rect 9180 280 9186 332
rect 10689 323 10747 329
rect 10689 289 10701 323
rect 10735 320 10747 323
rect 10778 320 10784 332
rect 10735 292 10784 320
rect 10735 289 10747 292
rect 10689 283 10747 289
rect 10778 280 10784 292
rect 10836 280 10842 332
rect 12986 320 12992 332
rect 12947 292 12992 320
rect 12986 280 12992 292
rect 13044 280 13050 332
rect 16132 329 16160 428
rect 16482 416 16488 428
rect 16540 416 16546 468
rect 17497 459 17555 465
rect 17497 425 17509 459
rect 17543 456 17555 459
rect 17770 456 17776 468
rect 17543 428 17776 456
rect 17543 425 17555 428
rect 17497 419 17555 425
rect 17770 416 17776 428
rect 17828 416 17834 468
rect 18322 456 18328 468
rect 18283 428 18328 456
rect 18322 416 18328 428
rect 18380 416 18386 468
rect 16117 323 16175 329
rect 16117 289 16129 323
rect 16163 289 16175 323
rect 16117 283 16175 289
rect 750 212 756 264
rect 808 252 814 264
rect 2317 255 2375 261
rect 2317 252 2329 255
rect 808 224 2329 252
rect 808 212 814 224
rect 2317 221 2329 224
rect 2363 221 2375 255
rect 2317 215 2375 221
rect 2409 255 2467 261
rect 2409 221 2421 255
rect 2455 252 2467 255
rect 2685 255 2743 261
rect 2685 252 2697 255
rect 2455 224 2697 252
rect 2455 221 2467 224
rect 2409 215 2467 221
rect 2685 221 2697 224
rect 2731 221 2743 255
rect 5994 252 6000 264
rect 5955 224 6000 252
rect 2685 215 2743 221
rect 5994 212 6000 224
rect 6052 212 6058 264
rect 8570 212 8576 264
rect 8628 252 8634 264
rect 8849 255 8907 261
rect 8849 252 8861 255
rect 8628 224 8861 252
rect 8628 212 8634 224
rect 8849 221 8861 224
rect 8895 221 8907 255
rect 8849 215 8907 221
rect 8941 255 8999 261
rect 8941 221 8953 255
rect 8987 252 8999 255
rect 10597 255 10655 261
rect 10597 252 10609 255
rect 8987 224 10609 252
rect 8987 221 8999 224
rect 8941 215 8999 221
rect 10597 221 10609 224
rect 10643 252 10655 255
rect 11054 252 11060 264
rect 10643 224 11060 252
rect 10643 221 10655 224
rect 10597 215 10655 221
rect 11054 212 11060 224
rect 11112 212 11118 264
rect 18506 252 18512 264
rect 18467 224 18512 252
rect 18506 212 18512 224
rect 18564 212 18570 264
rect 2682 76 2688 128
rect 2740 116 2746 128
rect 3436 116 3464 170
rect 8202 144 8208 196
rect 8260 184 8266 196
rect 9125 187 9183 193
rect 9125 184 9137 187
rect 8260 156 9137 184
rect 8260 144 8266 156
rect 9125 153 9137 156
rect 9171 153 9183 187
rect 9125 147 9183 153
rect 10962 144 10968 196
rect 11020 144 11026 196
rect 13170 144 13176 196
rect 13228 184 13234 196
rect 13265 187 13323 193
rect 13265 184 13277 187
rect 13228 156 13277 184
rect 13228 144 13234 156
rect 13265 153 13277 156
rect 13311 153 13323 187
rect 14918 184 14924 196
rect 14490 156 14924 184
rect 13265 147 13323 153
rect 14918 144 14924 156
rect 14976 144 14982 196
rect 16362 187 16420 193
rect 16362 184 16374 187
rect 16132 156 16374 184
rect 2740 88 3464 116
rect 8757 119 8815 125
rect 2740 76 2746 88
rect 8757 85 8769 119
rect 8803 116 8815 119
rect 8849 119 8907 125
rect 8849 116 8861 119
rect 8803 88 8861 116
rect 8803 85 8815 88
rect 8757 79 8815 85
rect 8849 85 8861 88
rect 8895 85 8907 119
rect 10980 116 11008 144
rect 16132 116 16160 156
rect 16362 153 16374 156
rect 16408 184 16420 187
rect 17954 184 17960 196
rect 16408 156 17960 184
rect 16408 153 16420 156
rect 16362 147 16420 153
rect 17954 144 17960 156
rect 18012 144 18018 196
rect 10980 88 16160 116
rect 8849 79 8907 85
rect 0 26 18860 48
rect 0 -26 4660 26
rect 4712 -26 4724 26
rect 4776 -26 4788 26
rect 4840 -26 4852 26
rect 4904 -26 4916 26
rect 4968 -26 7760 26
rect 7812 -26 7824 26
rect 7876 -26 7888 26
rect 7940 -26 7952 26
rect 8004 -26 8016 26
rect 8068 -26 10860 26
rect 10912 -26 10924 26
rect 10976 -26 10988 26
rect 11040 -26 11052 26
rect 11104 -26 11116 26
rect 11168 -26 13960 26
rect 14012 -26 14024 26
rect 14076 -26 14088 26
rect 14140 -26 14152 26
rect 14204 -26 14216 26
rect 14268 -26 17060 26
rect 17112 -26 17124 26
rect 17176 -26 17188 26
rect 17240 -26 17252 26
rect 17304 -26 17316 26
rect 17368 -26 18860 26
rect 0 -48 18860 -26
<< via1 >>
rect 4660 10854 4712 10906
rect 4724 10854 4776 10906
rect 4788 10854 4840 10906
rect 4852 10854 4904 10906
rect 4916 10854 4968 10906
rect 7760 10854 7812 10906
rect 7824 10854 7876 10906
rect 7888 10854 7940 10906
rect 7952 10854 8004 10906
rect 8016 10854 8068 10906
rect 10860 10854 10912 10906
rect 10924 10854 10976 10906
rect 10988 10854 11040 10906
rect 11052 10854 11104 10906
rect 11116 10854 11168 10906
rect 13960 10854 14012 10906
rect 14024 10854 14076 10906
rect 14088 10854 14140 10906
rect 14152 10854 14204 10906
rect 14216 10854 14268 10906
rect 17060 10854 17112 10906
rect 17124 10854 17176 10906
rect 17188 10854 17240 10906
rect 17252 10854 17304 10906
rect 17316 10854 17368 10906
rect 2136 10684 2188 10736
rect 3792 10752 3844 10804
rect 7104 10752 7156 10804
rect 9956 10752 10008 10804
rect 1308 10659 1360 10668
rect 1308 10625 1317 10659
rect 1317 10625 1351 10659
rect 1351 10625 1360 10659
rect 1308 10616 1360 10625
rect 2688 10591 2740 10600
rect 2688 10557 2697 10591
rect 2697 10557 2731 10591
rect 2731 10557 2740 10591
rect 2688 10548 2740 10557
rect 2964 10548 3016 10600
rect 6736 10659 6788 10668
rect 6736 10625 6745 10659
rect 6745 10625 6779 10659
rect 6779 10625 6788 10659
rect 6736 10616 6788 10625
rect 7012 10659 7064 10668
rect 7012 10625 7021 10659
rect 7021 10625 7055 10659
rect 7055 10625 7064 10659
rect 7012 10616 7064 10625
rect 9220 10616 9272 10668
rect 10416 10659 10468 10668
rect 6000 10548 6052 10600
rect 7656 10548 7708 10600
rect 10416 10625 10425 10659
rect 10425 10625 10459 10659
rect 10459 10625 10468 10659
rect 10416 10616 10468 10625
rect 2320 10412 2372 10464
rect 4344 10412 4396 10464
rect 4436 10412 4488 10464
rect 5816 10455 5868 10464
rect 5816 10421 5825 10455
rect 5825 10421 5859 10455
rect 5859 10421 5868 10455
rect 5816 10412 5868 10421
rect 7472 10455 7524 10464
rect 7472 10421 7481 10455
rect 7481 10421 7515 10455
rect 7515 10421 7524 10455
rect 7472 10412 7524 10421
rect 9036 10412 9088 10464
rect 9680 10480 9732 10532
rect 13360 10684 13412 10736
rect 15936 10684 15988 10736
rect 12164 10616 12216 10668
rect 13268 10659 13320 10668
rect 13268 10625 13277 10659
rect 13277 10625 13311 10659
rect 13311 10625 13320 10659
rect 13268 10616 13320 10625
rect 13636 10591 13688 10600
rect 9956 10455 10008 10464
rect 9956 10421 9965 10455
rect 9965 10421 9999 10455
rect 9999 10421 10008 10455
rect 9956 10412 10008 10421
rect 12256 10480 12308 10532
rect 10784 10412 10836 10464
rect 12072 10412 12124 10464
rect 13636 10557 13645 10591
rect 13645 10557 13679 10591
rect 13679 10557 13688 10591
rect 13636 10548 13688 10557
rect 18328 10659 18380 10668
rect 18328 10625 18337 10659
rect 18337 10625 18371 10659
rect 18371 10625 18380 10659
rect 18328 10616 18380 10625
rect 14832 10548 14884 10600
rect 16488 10591 16540 10600
rect 16488 10557 16497 10591
rect 16497 10557 16531 10591
rect 16531 10557 16540 10591
rect 16488 10548 16540 10557
rect 15200 10412 15252 10464
rect 15292 10412 15344 10464
rect 3110 10310 3162 10362
rect 3174 10310 3226 10362
rect 3238 10310 3290 10362
rect 3302 10310 3354 10362
rect 3366 10310 3418 10362
rect 6210 10310 6262 10362
rect 6274 10310 6326 10362
rect 6338 10310 6390 10362
rect 6402 10310 6454 10362
rect 6466 10310 6518 10362
rect 9310 10310 9362 10362
rect 9374 10310 9426 10362
rect 9438 10310 9490 10362
rect 9502 10310 9554 10362
rect 9566 10310 9618 10362
rect 12410 10310 12462 10362
rect 12474 10310 12526 10362
rect 12538 10310 12590 10362
rect 12602 10310 12654 10362
rect 12666 10310 12718 10362
rect 15510 10310 15562 10362
rect 15574 10310 15626 10362
rect 15638 10310 15690 10362
rect 15702 10310 15754 10362
rect 15766 10310 15818 10362
rect 2688 10208 2740 10260
rect 296 10115 348 10124
rect 296 10081 305 10115
rect 305 10081 339 10115
rect 339 10081 348 10115
rect 296 10072 348 10081
rect 2964 10072 3016 10124
rect 3424 10072 3476 10124
rect 2320 10047 2372 10056
rect 2320 10013 2329 10047
rect 2329 10013 2363 10047
rect 2363 10013 2372 10047
rect 2320 10004 2372 10013
rect 3240 10047 3292 10056
rect 572 9979 624 9988
rect 572 9945 581 9979
rect 581 9945 615 9979
rect 615 9945 624 9979
rect 572 9936 624 9945
rect 2136 9936 2188 9988
rect 2228 9911 2280 9920
rect 2228 9877 2237 9911
rect 2237 9877 2271 9911
rect 2271 9877 2280 9911
rect 2228 9868 2280 9877
rect 2688 9911 2740 9920
rect 2688 9877 2697 9911
rect 2697 9877 2731 9911
rect 2731 9877 2740 9911
rect 2688 9868 2740 9877
rect 2872 9936 2924 9988
rect 3240 10013 3249 10047
rect 3249 10013 3283 10047
rect 3283 10013 3292 10047
rect 3240 10004 3292 10013
rect 4068 10004 4120 10056
rect 6000 10251 6052 10260
rect 6000 10217 6009 10251
rect 6009 10217 6043 10251
rect 6043 10217 6052 10251
rect 6000 10208 6052 10217
rect 7012 10208 7064 10260
rect 9220 10208 9272 10260
rect 4252 10140 4304 10192
rect 4344 10072 4396 10124
rect 9036 10072 9088 10124
rect 4436 9936 4488 9988
rect 7472 10004 7524 10056
rect 8944 10047 8996 10056
rect 8944 10013 8953 10047
rect 8953 10013 8987 10047
rect 8987 10013 8996 10047
rect 8944 10004 8996 10013
rect 9128 10047 9180 10056
rect 9128 10013 9137 10047
rect 9137 10013 9171 10047
rect 9171 10013 9180 10047
rect 9128 10004 9180 10013
rect 12808 10208 12860 10260
rect 13636 10251 13688 10260
rect 13636 10217 13645 10251
rect 13645 10217 13679 10251
rect 13679 10217 13688 10251
rect 13636 10208 13688 10217
rect 16488 10208 16540 10260
rect 18328 10251 18380 10260
rect 18328 10217 18337 10251
rect 18337 10217 18371 10251
rect 18371 10217 18380 10251
rect 18328 10208 18380 10217
rect 14832 10115 14884 10124
rect 14832 10081 14841 10115
rect 14841 10081 14875 10115
rect 14875 10081 14884 10115
rect 14832 10072 14884 10081
rect 15200 10115 15252 10124
rect 15200 10081 15209 10115
rect 15209 10081 15243 10115
rect 15243 10081 15252 10115
rect 15200 10072 15252 10081
rect 15292 10004 15344 10056
rect 17960 10047 18012 10056
rect 17960 10013 17969 10047
rect 17969 10013 18003 10047
rect 18003 10013 18012 10047
rect 17960 10004 18012 10013
rect 18788 10004 18840 10056
rect 4988 9911 5040 9920
rect 4988 9877 4997 9911
rect 4997 9877 5031 9911
rect 5031 9877 5040 9911
rect 4988 9868 5040 9877
rect 5908 9911 5960 9920
rect 5908 9877 5917 9911
rect 5917 9877 5951 9911
rect 5951 9877 5960 9911
rect 5908 9868 5960 9877
rect 8300 9868 8352 9920
rect 11244 9936 11296 9988
rect 15936 9936 15988 9988
rect 11520 9868 11572 9920
rect 17776 9911 17828 9920
rect 17776 9877 17785 9911
rect 17785 9877 17819 9911
rect 17819 9877 17828 9911
rect 17776 9868 17828 9877
rect 4660 9766 4712 9818
rect 4724 9766 4776 9818
rect 4788 9766 4840 9818
rect 4852 9766 4904 9818
rect 4916 9766 4968 9818
rect 7760 9766 7812 9818
rect 7824 9766 7876 9818
rect 7888 9766 7940 9818
rect 7952 9766 8004 9818
rect 8016 9766 8068 9818
rect 10860 9766 10912 9818
rect 10924 9766 10976 9818
rect 10988 9766 11040 9818
rect 11052 9766 11104 9818
rect 11116 9766 11168 9818
rect 13960 9766 14012 9818
rect 14024 9766 14076 9818
rect 14088 9766 14140 9818
rect 14152 9766 14204 9818
rect 14216 9766 14268 9818
rect 17060 9766 17112 9818
rect 17124 9766 17176 9818
rect 17188 9766 17240 9818
rect 17252 9766 17304 9818
rect 17316 9766 17368 9818
rect 572 9664 624 9716
rect 2780 9664 2832 9716
rect 4344 9664 4396 9716
rect 5816 9664 5868 9716
rect 6736 9664 6788 9716
rect 13268 9664 13320 9716
rect 2228 9596 2280 9648
rect 3240 9596 3292 9648
rect 5632 9596 5684 9648
rect 8300 9596 8352 9648
rect 9956 9639 10008 9648
rect 4620 9528 4672 9580
rect 2964 9392 3016 9444
rect 3240 9392 3292 9444
rect 3424 9392 3476 9444
rect 5448 9460 5500 9512
rect 5908 9528 5960 9580
rect 6828 9503 6880 9512
rect 6828 9469 6837 9503
rect 6837 9469 6871 9503
rect 6871 9469 6880 9503
rect 6828 9460 6880 9469
rect 9956 9605 9965 9639
rect 9965 9605 9999 9639
rect 9999 9605 10008 9639
rect 9956 9596 10008 9605
rect 11336 9596 11388 9648
rect 12532 9596 12584 9648
rect 12164 9528 12216 9580
rect 10876 9503 10928 9512
rect 4988 9324 5040 9376
rect 5908 9324 5960 9376
rect 10232 9324 10284 9376
rect 10600 9324 10652 9376
rect 10876 9469 10885 9503
rect 10885 9469 10919 9503
rect 10919 9469 10928 9503
rect 10876 9460 10928 9469
rect 12532 9460 12584 9512
rect 12900 9503 12952 9512
rect 12900 9469 12909 9503
rect 12909 9469 12943 9503
rect 12943 9469 12952 9503
rect 12900 9460 12952 9469
rect 11980 9392 12032 9444
rect 12072 9392 12124 9444
rect 13544 9460 13596 9512
rect 17776 9596 17828 9648
rect 15936 9528 15988 9580
rect 14372 9460 14424 9512
rect 15844 9460 15896 9512
rect 16488 9460 16540 9512
rect 17960 9503 18012 9512
rect 17960 9469 17969 9503
rect 17969 9469 18003 9503
rect 18003 9469 18012 9503
rect 17960 9460 18012 9469
rect 14464 9324 14516 9376
rect 3110 9222 3162 9274
rect 3174 9222 3226 9274
rect 3238 9222 3290 9274
rect 3302 9222 3354 9274
rect 3366 9222 3418 9274
rect 6210 9222 6262 9274
rect 6274 9222 6326 9274
rect 6338 9222 6390 9274
rect 6402 9222 6454 9274
rect 6466 9222 6518 9274
rect 9310 9222 9362 9274
rect 9374 9222 9426 9274
rect 9438 9222 9490 9274
rect 9502 9222 9554 9274
rect 9566 9222 9618 9274
rect 12410 9222 12462 9274
rect 12474 9222 12526 9274
rect 12538 9222 12590 9274
rect 12602 9222 12654 9274
rect 12666 9222 12718 9274
rect 15510 9222 15562 9274
rect 15574 9222 15626 9274
rect 15638 9222 15690 9274
rect 15702 9222 15754 9274
rect 15766 9222 15818 9274
rect 2872 9120 2924 9172
rect 4068 9120 4120 9172
rect 4620 9120 4672 9172
rect 10416 9120 10468 9172
rect 12164 9120 12216 9172
rect 13360 9120 13412 9172
rect 17960 9120 18012 9172
rect 296 9027 348 9036
rect 296 8993 305 9027
rect 305 8993 339 9027
rect 339 8993 348 9027
rect 296 8984 348 8993
rect 2504 8984 2556 9036
rect 2964 8984 3016 9036
rect 4988 8984 5040 9036
rect 5540 8984 5592 9036
rect 6092 9027 6144 9036
rect 6092 8993 6101 9027
rect 6101 8993 6135 9027
rect 6135 8993 6144 9027
rect 6092 8984 6144 8993
rect 6184 8984 6236 9036
rect 6828 8984 6880 9036
rect 1860 8848 1912 8900
rect 2780 8916 2832 8968
rect 3608 8916 3660 8968
rect 5908 8959 5960 8968
rect 5908 8925 5917 8959
rect 5917 8925 5951 8959
rect 5951 8925 5960 8959
rect 5908 8916 5960 8925
rect 6000 8916 6052 8968
rect 8116 8959 8168 8968
rect 8116 8925 8150 8959
rect 8150 8925 8168 8959
rect 9680 8984 9732 9036
rect 10876 9052 10928 9104
rect 10232 9027 10284 9036
rect 10232 8993 10241 9027
rect 10241 8993 10275 9027
rect 10275 8993 10284 9027
rect 10232 8984 10284 8993
rect 10416 8984 10468 9036
rect 11336 8984 11388 9036
rect 11980 8984 12032 9036
rect 12164 8984 12216 9036
rect 13728 8984 13780 9036
rect 16672 8984 16724 9036
rect 8116 8916 8168 8925
rect 2320 8780 2372 8832
rect 5448 8848 5500 8900
rect 6920 8848 6972 8900
rect 3240 8780 3292 8832
rect 4252 8823 4304 8832
rect 4252 8789 4261 8823
rect 4261 8789 4295 8823
rect 4295 8789 4304 8823
rect 4252 8780 4304 8789
rect 6184 8780 6236 8832
rect 6368 8780 6420 8832
rect 6828 8780 6880 8832
rect 11244 8916 11296 8968
rect 13360 8959 13412 8968
rect 13360 8925 13369 8959
rect 13369 8925 13403 8959
rect 13403 8925 13412 8959
rect 13360 8916 13412 8925
rect 13544 8959 13596 8968
rect 13544 8925 13553 8959
rect 13553 8925 13587 8959
rect 13587 8925 13596 8959
rect 13544 8916 13596 8925
rect 15292 8916 15344 8968
rect 15844 8959 15896 8968
rect 15844 8925 15853 8959
rect 15853 8925 15887 8959
rect 15887 8925 15896 8959
rect 15844 8916 15896 8925
rect 16120 8916 16172 8968
rect 10232 8848 10284 8900
rect 9864 8823 9916 8832
rect 9864 8789 9873 8823
rect 9873 8789 9907 8823
rect 9907 8789 9916 8823
rect 9864 8780 9916 8789
rect 12440 8848 12492 8900
rect 13452 8823 13504 8832
rect 13452 8789 13461 8823
rect 13461 8789 13495 8823
rect 13495 8789 13504 8823
rect 13452 8780 13504 8789
rect 13820 8780 13872 8832
rect 14372 8848 14424 8900
rect 16488 8848 16540 8900
rect 4660 8678 4712 8730
rect 4724 8678 4776 8730
rect 4788 8678 4840 8730
rect 4852 8678 4904 8730
rect 4916 8678 4968 8730
rect 7760 8678 7812 8730
rect 7824 8678 7876 8730
rect 7888 8678 7940 8730
rect 7952 8678 8004 8730
rect 8016 8678 8068 8730
rect 10860 8678 10912 8730
rect 10924 8678 10976 8730
rect 10988 8678 11040 8730
rect 11052 8678 11104 8730
rect 11116 8678 11168 8730
rect 13960 8678 14012 8730
rect 14024 8678 14076 8730
rect 14088 8678 14140 8730
rect 14152 8678 14204 8730
rect 14216 8678 14268 8730
rect 17060 8678 17112 8730
rect 17124 8678 17176 8730
rect 17188 8678 17240 8730
rect 17252 8678 17304 8730
rect 17316 8678 17368 8730
rect 2320 8619 2372 8628
rect 2320 8585 2329 8619
rect 2329 8585 2363 8619
rect 2363 8585 2372 8619
rect 2320 8576 2372 8585
rect 2504 8619 2556 8628
rect 2504 8585 2513 8619
rect 2513 8585 2547 8619
rect 2547 8585 2556 8619
rect 2504 8576 2556 8585
rect 3240 8619 3292 8628
rect 3240 8585 3249 8619
rect 3249 8585 3283 8619
rect 3283 8585 3292 8619
rect 3240 8576 3292 8585
rect 4252 8576 4304 8628
rect 2780 8551 2832 8560
rect 2780 8517 2789 8551
rect 2789 8517 2823 8551
rect 2823 8517 2832 8551
rect 5448 8551 5500 8560
rect 2780 8508 2832 8517
rect 2964 8440 3016 8492
rect 3700 8483 3752 8492
rect 3700 8449 3709 8483
rect 3709 8449 3743 8483
rect 3743 8449 3752 8483
rect 3700 8440 3752 8449
rect 4344 8483 4396 8492
rect 2872 8372 2924 8424
rect 3608 8372 3660 8424
rect 4344 8449 4353 8483
rect 4353 8449 4387 8483
rect 4387 8449 4396 8483
rect 4344 8440 4396 8449
rect 4528 8483 4580 8492
rect 4528 8449 4537 8483
rect 4537 8449 4571 8483
rect 4571 8449 4580 8483
rect 4528 8440 4580 8449
rect 5448 8517 5457 8551
rect 5457 8517 5491 8551
rect 5491 8517 5500 8551
rect 5448 8508 5500 8517
rect 4988 8440 5040 8492
rect 5540 8505 5592 8526
rect 5540 8474 5547 8505
rect 5547 8474 5581 8505
rect 5581 8474 5592 8505
rect 8300 8508 8352 8560
rect 5908 8483 5960 8492
rect 5908 8449 5917 8483
rect 5917 8449 5951 8483
rect 5951 8449 5960 8483
rect 5908 8440 5960 8449
rect 6368 8483 6420 8492
rect 6368 8449 6377 8483
rect 6377 8449 6411 8483
rect 6411 8449 6420 8483
rect 6368 8440 6420 8449
rect 18512 8576 18564 8628
rect 12164 8551 12216 8560
rect 12164 8517 12173 8551
rect 12173 8517 12207 8551
rect 12207 8517 12216 8551
rect 12164 8508 12216 8517
rect 13728 8508 13780 8560
rect 15292 8508 15344 8560
rect 16028 8508 16080 8560
rect 16304 8508 16356 8560
rect 10692 8483 10744 8492
rect 10692 8449 10726 8483
rect 10726 8449 10744 8483
rect 6000 8347 6052 8356
rect 6000 8313 6009 8347
rect 6009 8313 6043 8347
rect 6043 8313 6052 8347
rect 6000 8304 6052 8313
rect 2964 8236 3016 8288
rect 4620 8236 4672 8288
rect 5632 8236 5684 8288
rect 8024 8236 8076 8288
rect 9864 8236 9916 8288
rect 10692 8440 10744 8449
rect 14372 8483 14424 8492
rect 13452 8415 13504 8424
rect 13452 8381 13461 8415
rect 13461 8381 13495 8415
rect 13495 8381 13504 8415
rect 13452 8372 13504 8381
rect 14372 8449 14381 8483
rect 14381 8449 14415 8483
rect 14415 8449 14424 8483
rect 14372 8440 14424 8449
rect 14556 8483 14608 8492
rect 14556 8449 14565 8483
rect 14565 8449 14599 8483
rect 14599 8449 14608 8483
rect 14556 8440 14608 8449
rect 13820 8372 13872 8424
rect 15844 8372 15896 8424
rect 17500 8440 17552 8492
rect 17868 8440 17920 8492
rect 18512 8483 18564 8492
rect 18512 8449 18521 8483
rect 18521 8449 18555 8483
rect 18555 8449 18564 8483
rect 18512 8440 18564 8449
rect 12164 8304 12216 8356
rect 11336 8236 11388 8288
rect 11428 8236 11480 8288
rect 13820 8236 13872 8288
rect 14924 8279 14976 8288
rect 14924 8245 14933 8279
rect 14933 8245 14967 8279
rect 14967 8245 14976 8279
rect 14924 8236 14976 8245
rect 3110 8134 3162 8186
rect 3174 8134 3226 8186
rect 3238 8134 3290 8186
rect 3302 8134 3354 8186
rect 3366 8134 3418 8186
rect 6210 8134 6262 8186
rect 6274 8134 6326 8186
rect 6338 8134 6390 8186
rect 6402 8134 6454 8186
rect 6466 8134 6518 8186
rect 9310 8134 9362 8186
rect 9374 8134 9426 8186
rect 9438 8134 9490 8186
rect 9502 8134 9554 8186
rect 9566 8134 9618 8186
rect 12410 8134 12462 8186
rect 12474 8134 12526 8186
rect 12538 8134 12590 8186
rect 12602 8134 12654 8186
rect 12666 8134 12718 8186
rect 15510 8134 15562 8186
rect 15574 8134 15626 8186
rect 15638 8134 15690 8186
rect 15702 8134 15754 8186
rect 15766 8134 15818 8186
rect 4528 8075 4580 8084
rect 4528 8041 4537 8075
rect 4537 8041 4571 8075
rect 4571 8041 4580 8075
rect 4528 8032 4580 8041
rect 4620 8075 4672 8084
rect 4620 8041 4629 8075
rect 4629 8041 4663 8075
rect 4663 8041 4672 8075
rect 5540 8075 5592 8084
rect 4620 8032 4672 8041
rect 5540 8041 5549 8075
rect 5549 8041 5583 8075
rect 5583 8041 5592 8075
rect 5540 8032 5592 8041
rect 6920 8032 6972 8084
rect 8944 8032 8996 8084
rect 10140 8075 10192 8084
rect 10140 8041 10149 8075
rect 10149 8041 10183 8075
rect 10183 8041 10192 8075
rect 10140 8032 10192 8041
rect 10508 8032 10560 8084
rect 10692 8032 10744 8084
rect 10784 8032 10836 8084
rect 12256 8032 12308 8084
rect 14372 8075 14424 8084
rect 296 7939 348 7948
rect 296 7905 305 7939
rect 305 7905 339 7939
rect 339 7905 348 7939
rect 296 7896 348 7905
rect 6828 7964 6880 8016
rect 9772 8007 9824 8016
rect 9772 7973 9781 8007
rect 9781 7973 9815 8007
rect 9815 7973 9824 8007
rect 9772 7964 9824 7973
rect 572 7803 624 7812
rect 572 7769 581 7803
rect 581 7769 615 7803
rect 615 7769 624 7803
rect 572 7760 624 7769
rect 1860 7760 1912 7812
rect 3516 7828 3568 7880
rect 3608 7871 3660 7880
rect 3608 7837 3617 7871
rect 3617 7837 3651 7871
rect 3651 7837 3660 7871
rect 4068 7871 4120 7880
rect 3608 7828 3660 7837
rect 4068 7837 4077 7871
rect 4077 7837 4111 7871
rect 4111 7837 4120 7871
rect 4068 7828 4120 7837
rect 4252 7828 4304 7880
rect 5724 7896 5776 7948
rect 9864 7896 9916 7948
rect 8024 7871 8076 7880
rect 2412 7760 2464 7812
rect 2044 7735 2096 7744
rect 2044 7701 2053 7735
rect 2053 7701 2087 7735
rect 2087 7701 2096 7735
rect 2044 7692 2096 7701
rect 2504 7692 2556 7744
rect 3700 7735 3752 7744
rect 3700 7701 3709 7735
rect 3709 7701 3743 7735
rect 3743 7701 3752 7735
rect 3700 7692 3752 7701
rect 3884 7735 3936 7744
rect 3884 7701 3893 7735
rect 3893 7701 3927 7735
rect 3927 7701 3936 7735
rect 3884 7692 3936 7701
rect 8024 7837 8033 7871
rect 8033 7837 8067 7871
rect 8067 7837 8076 7871
rect 8024 7828 8076 7837
rect 9588 7828 9640 7880
rect 10232 7939 10284 7948
rect 10232 7905 10241 7939
rect 10241 7905 10275 7939
rect 10275 7905 10284 7939
rect 10232 7896 10284 7905
rect 11428 8007 11480 8016
rect 11428 7973 11437 8007
rect 11437 7973 11471 8007
rect 11471 7973 11480 8007
rect 14372 8041 14381 8075
rect 14381 8041 14415 8075
rect 14415 8041 14424 8075
rect 14372 8032 14424 8041
rect 14556 8032 14608 8084
rect 11428 7964 11480 7973
rect 10508 7871 10560 7880
rect 10508 7837 10517 7871
rect 10517 7837 10551 7871
rect 10551 7837 10560 7871
rect 10508 7828 10560 7837
rect 5816 7803 5868 7812
rect 5816 7769 5825 7803
rect 5825 7769 5859 7803
rect 5859 7769 5868 7803
rect 5816 7760 5868 7769
rect 6184 7803 6236 7812
rect 6184 7769 6193 7803
rect 6193 7769 6227 7803
rect 6227 7769 6236 7803
rect 6184 7760 6236 7769
rect 6552 7760 6604 7812
rect 5908 7735 5960 7744
rect 5908 7701 5917 7735
rect 5917 7701 5951 7735
rect 5951 7701 5960 7735
rect 5908 7692 5960 7701
rect 6736 7692 6788 7744
rect 9036 7760 9088 7812
rect 10140 7760 10192 7812
rect 11244 7939 11296 7948
rect 11244 7905 11253 7939
rect 11253 7905 11287 7939
rect 11287 7905 11296 7939
rect 11244 7896 11296 7905
rect 10876 7871 10928 7880
rect 10876 7837 10885 7871
rect 10885 7837 10919 7871
rect 10919 7837 10928 7871
rect 10876 7828 10928 7837
rect 10968 7871 11020 7880
rect 10968 7837 10977 7871
rect 10977 7837 11011 7871
rect 11011 7837 11020 7871
rect 10968 7828 11020 7837
rect 11152 7871 11204 7880
rect 11152 7837 11161 7871
rect 11161 7837 11195 7871
rect 11195 7837 11204 7871
rect 11152 7828 11204 7837
rect 11796 7828 11848 7880
rect 12348 7871 12400 7880
rect 12348 7837 12357 7871
rect 12357 7837 12391 7871
rect 12391 7837 12400 7871
rect 12348 7828 12400 7837
rect 12992 7871 13044 7880
rect 12992 7837 13001 7871
rect 13001 7837 13035 7871
rect 13035 7837 13044 7871
rect 12992 7828 13044 7837
rect 15844 7896 15896 7948
rect 13820 7871 13872 7880
rect 13820 7837 13829 7871
rect 13829 7837 13863 7871
rect 13863 7837 13872 7871
rect 13820 7828 13872 7837
rect 11520 7760 11572 7812
rect 11704 7803 11756 7812
rect 11704 7769 11713 7803
rect 11713 7769 11747 7803
rect 11747 7769 11756 7803
rect 11704 7760 11756 7769
rect 11888 7803 11940 7812
rect 11888 7769 11897 7803
rect 11897 7769 11931 7803
rect 11931 7769 11940 7803
rect 11888 7760 11940 7769
rect 14740 7828 14792 7880
rect 14924 7871 14976 7880
rect 14924 7837 14933 7871
rect 14933 7837 14967 7871
rect 14967 7837 14976 7871
rect 15200 7871 15252 7880
rect 14924 7828 14976 7837
rect 15200 7837 15209 7871
rect 15209 7837 15243 7871
rect 15243 7837 15252 7871
rect 15200 7828 15252 7837
rect 14740 7735 14792 7744
rect 14740 7701 14749 7735
rect 14749 7701 14783 7735
rect 14783 7701 14792 7735
rect 14740 7692 14792 7701
rect 14924 7692 14976 7744
rect 15568 7760 15620 7812
rect 16304 7760 16356 7812
rect 17592 7760 17644 7812
rect 4660 7590 4712 7642
rect 4724 7590 4776 7642
rect 4788 7590 4840 7642
rect 4852 7590 4904 7642
rect 4916 7590 4968 7642
rect 7760 7590 7812 7642
rect 7824 7590 7876 7642
rect 7888 7590 7940 7642
rect 7952 7590 8004 7642
rect 8016 7590 8068 7642
rect 10860 7590 10912 7642
rect 10924 7590 10976 7642
rect 10988 7590 11040 7642
rect 11052 7590 11104 7642
rect 11116 7590 11168 7642
rect 13960 7590 14012 7642
rect 14024 7590 14076 7642
rect 14088 7590 14140 7642
rect 14152 7590 14204 7642
rect 14216 7590 14268 7642
rect 17060 7590 17112 7642
rect 17124 7590 17176 7642
rect 17188 7590 17240 7642
rect 17252 7590 17304 7642
rect 17316 7590 17368 7642
rect 572 7488 624 7540
rect 1952 7488 2004 7540
rect 3148 7488 3200 7540
rect 3700 7488 3752 7540
rect 2596 7420 2648 7472
rect 3884 7420 3936 7472
rect 2044 7352 2096 7404
rect 2504 7395 2556 7404
rect 2504 7361 2513 7395
rect 2513 7361 2547 7395
rect 2547 7361 2556 7395
rect 2504 7352 2556 7361
rect 2780 7395 2832 7404
rect 2780 7361 2789 7395
rect 2789 7361 2823 7395
rect 2823 7361 2832 7395
rect 3148 7395 3200 7404
rect 2780 7352 2832 7361
rect 3148 7361 3157 7395
rect 3157 7361 3191 7395
rect 3191 7361 3200 7395
rect 3148 7352 3200 7361
rect 2412 7327 2464 7336
rect 2412 7293 2421 7327
rect 2421 7293 2455 7327
rect 2455 7293 2464 7327
rect 3332 7395 3384 7404
rect 3332 7361 3341 7395
rect 3341 7361 3375 7395
rect 3375 7361 3384 7395
rect 3332 7352 3384 7361
rect 3516 7352 3568 7404
rect 5816 7488 5868 7540
rect 5908 7488 5960 7540
rect 6092 7488 6144 7540
rect 6184 7420 6236 7472
rect 5264 7395 5316 7404
rect 5264 7361 5273 7395
rect 5273 7361 5307 7395
rect 5307 7361 5316 7395
rect 5264 7352 5316 7361
rect 5724 7395 5776 7404
rect 5724 7361 5733 7395
rect 5733 7361 5767 7395
rect 5767 7361 5776 7395
rect 5724 7352 5776 7361
rect 5908 7395 5960 7404
rect 5908 7361 5917 7395
rect 5917 7361 5951 7395
rect 5951 7361 5960 7395
rect 5908 7352 5960 7361
rect 5080 7327 5132 7336
rect 2412 7284 2464 7293
rect 5080 7293 5089 7327
rect 5089 7293 5123 7327
rect 5123 7293 5132 7327
rect 5080 7284 5132 7293
rect 6092 7284 6144 7336
rect 2320 7216 2372 7268
rect 2412 7148 2464 7200
rect 2688 7191 2740 7200
rect 2688 7157 2697 7191
rect 2697 7157 2731 7191
rect 2731 7157 2740 7191
rect 2688 7148 2740 7157
rect 4068 7216 4120 7268
rect 5264 7216 5316 7268
rect 4252 7148 4304 7200
rect 9588 7488 9640 7540
rect 10416 7488 10468 7540
rect 6644 7284 6696 7336
rect 6920 7352 6972 7404
rect 8944 7395 8996 7404
rect 8944 7361 8953 7395
rect 8953 7361 8987 7395
rect 8987 7361 8996 7395
rect 8944 7352 8996 7361
rect 9036 7395 9088 7404
rect 9036 7361 9045 7395
rect 9045 7361 9079 7395
rect 9079 7361 9088 7395
rect 9036 7352 9088 7361
rect 9220 7352 9272 7404
rect 6828 7327 6880 7336
rect 6828 7293 6837 7327
rect 6837 7293 6871 7327
rect 6871 7293 6880 7327
rect 6828 7284 6880 7293
rect 8116 7284 8168 7336
rect 10416 7352 10468 7404
rect 11428 7488 11480 7540
rect 15568 7531 15620 7540
rect 15568 7497 15577 7531
rect 15577 7497 15611 7531
rect 15611 7497 15620 7531
rect 15568 7488 15620 7497
rect 17960 7488 18012 7540
rect 11980 7420 12032 7472
rect 16304 7420 16356 7472
rect 18328 7420 18380 7472
rect 8392 7216 8444 7268
rect 9772 7216 9824 7268
rect 10784 7284 10836 7336
rect 12348 7352 12400 7404
rect 14740 7352 14792 7404
rect 15200 7352 15252 7404
rect 17500 7352 17552 7404
rect 11336 7284 11388 7336
rect 17868 7327 17920 7336
rect 17868 7293 17877 7327
rect 17877 7293 17911 7327
rect 17911 7293 17920 7327
rect 17868 7284 17920 7293
rect 10416 7148 10468 7200
rect 15016 7191 15068 7200
rect 15016 7157 15025 7191
rect 15025 7157 15059 7191
rect 15059 7157 15068 7191
rect 17408 7191 17460 7200
rect 15016 7148 15068 7157
rect 17408 7157 17417 7191
rect 17417 7157 17451 7191
rect 17451 7157 17460 7191
rect 17408 7148 17460 7157
rect 3110 7046 3162 7098
rect 3174 7046 3226 7098
rect 3238 7046 3290 7098
rect 3302 7046 3354 7098
rect 3366 7046 3418 7098
rect 6210 7046 6262 7098
rect 6274 7046 6326 7098
rect 6338 7046 6390 7098
rect 6402 7046 6454 7098
rect 6466 7046 6518 7098
rect 9310 7046 9362 7098
rect 9374 7046 9426 7098
rect 9438 7046 9490 7098
rect 9502 7046 9554 7098
rect 9566 7046 9618 7098
rect 12410 7046 12462 7098
rect 12474 7046 12526 7098
rect 12538 7046 12590 7098
rect 12602 7046 12654 7098
rect 12666 7046 12718 7098
rect 15510 7046 15562 7098
rect 15574 7046 15626 7098
rect 15638 7046 15690 7098
rect 15702 7046 15754 7098
rect 15766 7046 15818 7098
rect 5632 6944 5684 6996
rect 6644 6944 6696 6996
rect 10140 6987 10192 6996
rect 10140 6953 10149 6987
rect 10149 6953 10183 6987
rect 10183 6953 10192 6987
rect 10140 6944 10192 6953
rect 10416 6987 10468 6996
rect 10416 6953 10425 6987
rect 10425 6953 10459 6987
rect 10459 6953 10468 6987
rect 10416 6944 10468 6953
rect 2780 6876 2832 6928
rect 3240 6876 3292 6928
rect 3608 6876 3660 6928
rect 5908 6876 5960 6928
rect 1952 6851 2004 6860
rect 1952 6817 1961 6851
rect 1961 6817 1995 6851
rect 1995 6817 2004 6851
rect 1952 6808 2004 6817
rect 2964 6808 3016 6860
rect 2688 6740 2740 6792
rect 2044 6715 2096 6724
rect 2044 6681 2053 6715
rect 2053 6681 2087 6715
rect 2087 6681 2096 6715
rect 3240 6783 3292 6792
rect 3240 6749 3249 6783
rect 3249 6749 3283 6783
rect 3283 6749 3292 6783
rect 3240 6740 3292 6749
rect 6092 6808 6144 6860
rect 3516 6783 3568 6792
rect 3516 6749 3525 6783
rect 3525 6749 3559 6783
rect 3559 6749 3568 6783
rect 3516 6740 3568 6749
rect 4068 6783 4120 6792
rect 4068 6749 4077 6783
rect 4077 6749 4111 6783
rect 4111 6749 4120 6783
rect 4068 6740 4120 6749
rect 8024 6808 8076 6860
rect 8668 6851 8720 6860
rect 8668 6817 8677 6851
rect 8677 6817 8711 6851
rect 8711 6817 8720 6851
rect 8668 6808 8720 6817
rect 10508 6876 10560 6928
rect 8392 6783 8444 6792
rect 2044 6672 2096 6681
rect 4344 6715 4396 6724
rect 4344 6681 4353 6715
rect 4353 6681 4387 6715
rect 4387 6681 4396 6715
rect 4344 6672 4396 6681
rect 4436 6672 4488 6724
rect 572 6604 624 6656
rect 2412 6604 2464 6656
rect 2596 6604 2648 6656
rect 5908 6604 5960 6656
rect 6092 6604 6144 6656
rect 6828 6647 6880 6656
rect 6828 6613 6837 6647
rect 6837 6613 6871 6647
rect 6871 6613 6880 6647
rect 6828 6604 6880 6613
rect 8392 6749 8401 6783
rect 8401 6749 8435 6783
rect 8435 6749 8444 6783
rect 8392 6740 8444 6749
rect 8576 6740 8628 6792
rect 9220 6740 9272 6792
rect 9772 6808 9824 6860
rect 12992 6944 13044 6996
rect 15200 6987 15252 6996
rect 15200 6953 15209 6987
rect 15209 6953 15243 6987
rect 15243 6953 15252 6987
rect 15200 6944 15252 6953
rect 17868 6944 17920 6996
rect 18328 6987 18380 6996
rect 18328 6953 18337 6987
rect 18337 6953 18371 6987
rect 18371 6953 18380 6987
rect 18328 6944 18380 6953
rect 9864 6740 9916 6792
rect 10232 6740 10284 6792
rect 10324 6740 10376 6792
rect 11244 6740 11296 6792
rect 11888 6808 11940 6860
rect 14832 6808 14884 6860
rect 15016 6851 15068 6860
rect 15016 6817 15025 6851
rect 15025 6817 15059 6851
rect 15059 6817 15068 6851
rect 15016 6808 15068 6817
rect 15568 6851 15620 6860
rect 15568 6817 15577 6851
rect 15577 6817 15611 6851
rect 15611 6817 15620 6851
rect 15568 6808 15620 6817
rect 10692 6672 10744 6724
rect 11520 6740 11572 6792
rect 13544 6740 13596 6792
rect 15200 6740 15252 6792
rect 15476 6783 15528 6792
rect 15476 6749 15485 6783
rect 15485 6749 15519 6783
rect 15519 6749 15528 6783
rect 15476 6740 15528 6749
rect 9588 6647 9640 6656
rect 9588 6613 9597 6647
rect 9597 6613 9631 6647
rect 9631 6613 9640 6647
rect 9588 6604 9640 6613
rect 10784 6647 10836 6656
rect 10784 6613 10793 6647
rect 10793 6613 10827 6647
rect 10827 6613 10836 6647
rect 10784 6604 10836 6613
rect 17592 6808 17644 6860
rect 17408 6740 17460 6792
rect 17776 6783 17828 6792
rect 17776 6749 17785 6783
rect 17785 6749 17819 6783
rect 17819 6749 17828 6783
rect 17776 6740 17828 6749
rect 18512 6783 18564 6792
rect 18512 6749 18521 6783
rect 18521 6749 18555 6783
rect 18555 6749 18564 6783
rect 18512 6740 18564 6749
rect 11520 6604 11572 6656
rect 13176 6604 13228 6656
rect 13820 6604 13872 6656
rect 14832 6647 14884 6656
rect 14832 6613 14841 6647
rect 14841 6613 14875 6647
rect 14875 6613 14884 6647
rect 14832 6604 14884 6613
rect 16396 6604 16448 6656
rect 4660 6502 4712 6554
rect 4724 6502 4776 6554
rect 4788 6502 4840 6554
rect 4852 6502 4904 6554
rect 4916 6502 4968 6554
rect 7760 6502 7812 6554
rect 7824 6502 7876 6554
rect 7888 6502 7940 6554
rect 7952 6502 8004 6554
rect 8016 6502 8068 6554
rect 10860 6502 10912 6554
rect 10924 6502 10976 6554
rect 10988 6502 11040 6554
rect 11052 6502 11104 6554
rect 11116 6502 11168 6554
rect 13960 6502 14012 6554
rect 14024 6502 14076 6554
rect 14088 6502 14140 6554
rect 14152 6502 14204 6554
rect 14216 6502 14268 6554
rect 17060 6502 17112 6554
rect 17124 6502 17176 6554
rect 17188 6502 17240 6554
rect 17252 6502 17304 6554
rect 17316 6502 17368 6554
rect 2044 6443 2096 6452
rect 2044 6409 2053 6443
rect 2053 6409 2087 6443
rect 2087 6409 2096 6443
rect 2044 6400 2096 6409
rect 4344 6400 4396 6452
rect 6828 6443 6880 6452
rect 6828 6409 6837 6443
rect 6837 6409 6871 6443
rect 6871 6409 6880 6443
rect 6828 6400 6880 6409
rect 572 6375 624 6384
rect 572 6341 581 6375
rect 581 6341 615 6375
rect 615 6341 624 6375
rect 572 6332 624 6341
rect 9036 6400 9088 6452
rect 8668 6332 8720 6384
rect 9588 6332 9640 6384
rect 2320 6307 2372 6316
rect 296 6239 348 6248
rect 296 6205 305 6239
rect 305 6205 339 6239
rect 339 6205 348 6239
rect 296 6196 348 6205
rect 2320 6273 2329 6307
rect 2329 6273 2363 6307
rect 2363 6273 2372 6307
rect 2320 6264 2372 6273
rect 2412 6307 2464 6316
rect 2412 6273 2421 6307
rect 2421 6273 2455 6307
rect 2455 6273 2464 6307
rect 2412 6264 2464 6273
rect 5080 6264 5132 6316
rect 5724 6307 5776 6316
rect 5724 6273 5733 6307
rect 5733 6273 5767 6307
rect 5767 6273 5776 6307
rect 5724 6264 5776 6273
rect 5908 6264 5960 6316
rect 6276 6307 6328 6316
rect 2596 6239 2648 6248
rect 2596 6205 2605 6239
rect 2605 6205 2639 6239
rect 2639 6205 2648 6239
rect 2596 6196 2648 6205
rect 5816 6239 5868 6248
rect 1860 6128 1912 6180
rect 2412 6128 2464 6180
rect 4436 6128 4488 6180
rect 5816 6205 5825 6239
rect 5825 6205 5859 6239
rect 5859 6205 5868 6239
rect 5816 6196 5868 6205
rect 6276 6273 6285 6307
rect 6285 6273 6319 6307
rect 6319 6273 6328 6307
rect 6276 6264 6328 6273
rect 6552 6307 6604 6316
rect 6552 6273 6561 6307
rect 6561 6273 6595 6307
rect 6595 6273 6604 6307
rect 6552 6264 6604 6273
rect 6736 6307 6788 6316
rect 6736 6273 6745 6307
rect 6745 6273 6779 6307
rect 6779 6273 6788 6307
rect 6920 6307 6972 6316
rect 6736 6264 6788 6273
rect 6920 6273 6929 6307
rect 6929 6273 6963 6307
rect 6963 6273 6972 6307
rect 6920 6264 6972 6273
rect 8392 6307 8444 6316
rect 8392 6273 8401 6307
rect 8401 6273 8435 6307
rect 8435 6273 8444 6307
rect 8392 6264 8444 6273
rect 7472 6196 7524 6248
rect 9956 6307 10008 6316
rect 9956 6273 9965 6307
rect 9965 6273 9999 6307
rect 9999 6273 10008 6307
rect 9956 6264 10008 6273
rect 6276 6128 6328 6180
rect 2964 6060 3016 6112
rect 9772 6196 9824 6248
rect 6736 6060 6788 6112
rect 10232 6307 10284 6316
rect 10232 6273 10241 6307
rect 10241 6273 10275 6307
rect 10275 6273 10284 6307
rect 10784 6307 10836 6316
rect 10232 6264 10284 6273
rect 10784 6273 10793 6307
rect 10793 6273 10827 6307
rect 10827 6273 10836 6307
rect 10784 6264 10836 6273
rect 11244 6400 11296 6452
rect 11520 6443 11572 6452
rect 11520 6409 11529 6443
rect 11529 6409 11563 6443
rect 11563 6409 11572 6443
rect 11520 6400 11572 6409
rect 11888 6400 11940 6452
rect 13820 6400 13872 6452
rect 11336 6332 11388 6384
rect 11796 6332 11848 6384
rect 14832 6400 14884 6452
rect 10508 6196 10560 6248
rect 13820 6264 13872 6316
rect 15476 6332 15528 6384
rect 12992 6196 13044 6248
rect 15568 6264 15620 6316
rect 16396 6307 16448 6316
rect 16396 6273 16405 6307
rect 16405 6273 16439 6307
rect 16439 6273 16448 6307
rect 16396 6264 16448 6273
rect 17776 6400 17828 6452
rect 17408 6332 17460 6384
rect 14924 6196 14976 6248
rect 16672 6239 16724 6248
rect 16672 6205 16681 6239
rect 16681 6205 16715 6239
rect 16715 6205 16724 6239
rect 16672 6196 16724 6205
rect 11612 6128 11664 6180
rect 11520 6060 11572 6112
rect 14924 6103 14976 6112
rect 14924 6069 14933 6103
rect 14933 6069 14967 6103
rect 14967 6069 14976 6103
rect 14924 6060 14976 6069
rect 3110 5958 3162 6010
rect 3174 5958 3226 6010
rect 3238 5958 3290 6010
rect 3302 5958 3354 6010
rect 3366 5958 3418 6010
rect 6210 5958 6262 6010
rect 6274 5958 6326 6010
rect 6338 5958 6390 6010
rect 6402 5958 6454 6010
rect 6466 5958 6518 6010
rect 9310 5958 9362 6010
rect 9374 5958 9426 6010
rect 9438 5958 9490 6010
rect 9502 5958 9554 6010
rect 9566 5958 9618 6010
rect 12410 5958 12462 6010
rect 12474 5958 12526 6010
rect 12538 5958 12590 6010
rect 12602 5958 12654 6010
rect 12666 5958 12718 6010
rect 15510 5958 15562 6010
rect 15574 5958 15626 6010
rect 15638 5958 15690 6010
rect 15702 5958 15754 6010
rect 15766 5958 15818 6010
rect 3516 5856 3568 5908
rect 6920 5856 6972 5908
rect 8208 5856 8260 5908
rect 9956 5856 10008 5908
rect 12992 5899 13044 5908
rect 12992 5865 13001 5899
rect 13001 5865 13035 5899
rect 13035 5865 13044 5899
rect 12992 5856 13044 5865
rect 296 5720 348 5772
rect 4068 5720 4120 5772
rect 6000 5720 6052 5772
rect 6092 5720 6144 5772
rect 15384 5788 15436 5840
rect 2964 5652 3016 5704
rect 14924 5720 14976 5772
rect 15200 5763 15252 5772
rect 15200 5729 15209 5763
rect 15209 5729 15243 5763
rect 15243 5729 15252 5763
rect 15200 5720 15252 5729
rect 16672 5720 16724 5772
rect 11796 5695 11848 5704
rect 11796 5661 11805 5695
rect 11805 5661 11839 5695
rect 11839 5661 11848 5695
rect 13176 5695 13228 5704
rect 11796 5652 11848 5661
rect 13176 5661 13185 5695
rect 13185 5661 13219 5695
rect 13219 5661 13228 5695
rect 13176 5652 13228 5661
rect 18512 5695 18564 5704
rect 18512 5661 18521 5695
rect 18521 5661 18555 5695
rect 18555 5661 18564 5695
rect 18512 5652 18564 5661
rect 3792 5584 3844 5636
rect 11520 5627 11572 5636
rect 2412 5516 2464 5568
rect 8300 5516 8352 5568
rect 8852 5516 8904 5568
rect 11520 5593 11529 5627
rect 11529 5593 11563 5627
rect 11563 5593 11572 5627
rect 11520 5584 11572 5593
rect 15108 5584 15160 5636
rect 13820 5516 13872 5568
rect 18236 5516 18288 5568
rect 4660 5414 4712 5466
rect 4724 5414 4776 5466
rect 4788 5414 4840 5466
rect 4852 5414 4904 5466
rect 4916 5414 4968 5466
rect 7760 5414 7812 5466
rect 7824 5414 7876 5466
rect 7888 5414 7940 5466
rect 7952 5414 8004 5466
rect 8016 5414 8068 5466
rect 10860 5414 10912 5466
rect 10924 5414 10976 5466
rect 10988 5414 11040 5466
rect 11052 5414 11104 5466
rect 11116 5414 11168 5466
rect 13960 5414 14012 5466
rect 14024 5414 14076 5466
rect 14088 5414 14140 5466
rect 14152 5414 14204 5466
rect 14216 5414 14268 5466
rect 17060 5414 17112 5466
rect 17124 5414 17176 5466
rect 17188 5414 17240 5466
rect 17252 5414 17304 5466
rect 17316 5414 17368 5466
rect 7472 5244 7524 5296
rect 5080 5176 5132 5228
rect 6920 5176 6972 5228
rect 6920 4972 6972 5024
rect 7840 5176 7892 5228
rect 8208 5244 8260 5296
rect 10600 5312 10652 5364
rect 9128 5244 9180 5296
rect 13820 5244 13872 5296
rect 15108 5244 15160 5296
rect 16304 5244 16356 5296
rect 17408 5312 17460 5364
rect 17960 5244 18012 5296
rect 8944 5209 8996 5218
rect 8944 5175 8953 5209
rect 8953 5175 8987 5209
rect 8987 5175 8996 5209
rect 9772 5219 9824 5228
rect 8944 5166 8996 5175
rect 8392 5151 8444 5160
rect 8392 5117 8401 5151
rect 8401 5117 8435 5151
rect 8435 5117 8444 5151
rect 8392 5108 8444 5117
rect 9772 5185 9781 5219
rect 9781 5185 9815 5219
rect 9815 5185 9824 5219
rect 9772 5176 9824 5185
rect 12256 5151 12308 5160
rect 8484 5040 8536 5092
rect 12256 5117 12265 5151
rect 12265 5117 12299 5151
rect 12299 5117 12308 5151
rect 12256 5108 12308 5117
rect 14556 5151 14608 5160
rect 14556 5117 14565 5151
rect 14565 5117 14599 5151
rect 14599 5117 14608 5151
rect 14556 5108 14608 5117
rect 18236 5151 18288 5160
rect 18236 5117 18245 5151
rect 18245 5117 18279 5151
rect 18279 5117 18288 5151
rect 18236 5108 18288 5117
rect 12808 5083 12860 5092
rect 12808 5049 12817 5083
rect 12817 5049 12851 5083
rect 12851 5049 12860 5083
rect 12808 5040 12860 5049
rect 10048 4972 10100 5024
rect 17684 4972 17736 5024
rect 3110 4870 3162 4922
rect 3174 4870 3226 4922
rect 3238 4870 3290 4922
rect 3302 4870 3354 4922
rect 3366 4870 3418 4922
rect 6210 4870 6262 4922
rect 6274 4870 6326 4922
rect 6338 4870 6390 4922
rect 6402 4870 6454 4922
rect 6466 4870 6518 4922
rect 9310 4870 9362 4922
rect 9374 4870 9426 4922
rect 9438 4870 9490 4922
rect 9502 4870 9554 4922
rect 9566 4870 9618 4922
rect 12410 4870 12462 4922
rect 12474 4870 12526 4922
rect 12538 4870 12590 4922
rect 12602 4870 12654 4922
rect 12666 4870 12718 4922
rect 15510 4870 15562 4922
rect 15574 4870 15626 4922
rect 15638 4870 15690 4922
rect 15702 4870 15754 4922
rect 15766 4870 15818 4922
rect 5080 4811 5132 4820
rect 5080 4777 5089 4811
rect 5089 4777 5123 4811
rect 5123 4777 5132 4811
rect 5080 4768 5132 4777
rect 9864 4768 9916 4820
rect 12256 4811 12308 4820
rect 12256 4777 12265 4811
rect 12265 4777 12299 4811
rect 12299 4777 12308 4811
rect 12256 4768 12308 4777
rect 14464 4768 14516 4820
rect 2320 4607 2372 4616
rect 2320 4573 2329 4607
rect 2329 4573 2363 4607
rect 2363 4573 2372 4607
rect 2320 4564 2372 4573
rect 3056 4607 3108 4616
rect 3056 4573 3065 4607
rect 3065 4573 3099 4607
rect 3099 4573 3108 4607
rect 3056 4564 3108 4573
rect 4988 4564 5040 4616
rect 8760 4632 8812 4684
rect 10600 4632 10652 4684
rect 12072 4632 12124 4684
rect 7656 4564 7708 4616
rect 8208 4607 8260 4616
rect 8208 4573 8217 4607
rect 8217 4573 8251 4607
rect 8251 4573 8260 4607
rect 8208 4564 8260 4573
rect 2412 4428 2464 4480
rect 5172 4428 5224 4480
rect 5632 4428 5684 4480
rect 7380 4496 7432 4548
rect 8484 4496 8536 4548
rect 9036 4564 9088 4616
rect 14556 4632 14608 4684
rect 17684 4675 17736 4684
rect 17684 4641 17693 4675
rect 17693 4641 17727 4675
rect 17727 4641 17736 4675
rect 17684 4632 17736 4641
rect 9634 4540 9686 4592
rect 10048 4539 10100 4548
rect 10048 4505 10057 4539
rect 10057 4505 10091 4539
rect 10091 4505 10100 4539
rect 10048 4496 10100 4505
rect 11336 4496 11388 4548
rect 11428 4496 11480 4548
rect 12256 4496 12308 4548
rect 12808 4564 12860 4616
rect 17960 4607 18012 4616
rect 17960 4573 17969 4607
rect 17969 4573 18003 4607
rect 18003 4573 18012 4607
rect 18512 4607 18564 4616
rect 17960 4564 18012 4573
rect 18512 4573 18521 4607
rect 18521 4573 18555 4607
rect 18555 4573 18564 4607
rect 18512 4564 18564 4573
rect 9128 4428 9180 4480
rect 11520 4471 11572 4480
rect 11520 4437 11529 4471
rect 11529 4437 11563 4471
rect 11563 4437 11572 4471
rect 15108 4496 15160 4548
rect 15936 4539 15988 4548
rect 12624 4471 12676 4480
rect 11520 4428 11572 4437
rect 12624 4437 12633 4471
rect 12633 4437 12667 4471
rect 12667 4437 12676 4471
rect 12624 4428 12676 4437
rect 15936 4505 15945 4539
rect 15945 4505 15979 4539
rect 15979 4505 15988 4539
rect 15936 4496 15988 4505
rect 16304 4496 16356 4548
rect 18236 4496 18288 4548
rect 17408 4428 17460 4480
rect 4660 4326 4712 4378
rect 4724 4326 4776 4378
rect 4788 4326 4840 4378
rect 4852 4326 4904 4378
rect 4916 4326 4968 4378
rect 7760 4326 7812 4378
rect 7824 4326 7876 4378
rect 7888 4326 7940 4378
rect 7952 4326 8004 4378
rect 8016 4326 8068 4378
rect 10860 4326 10912 4378
rect 10924 4326 10976 4378
rect 10988 4326 11040 4378
rect 11052 4326 11104 4378
rect 11116 4326 11168 4378
rect 13960 4326 14012 4378
rect 14024 4326 14076 4378
rect 14088 4326 14140 4378
rect 14152 4326 14204 4378
rect 14216 4326 14268 4378
rect 17060 4326 17112 4378
rect 17124 4326 17176 4378
rect 17188 4326 17240 4378
rect 17252 4326 17304 4378
rect 17316 4326 17368 4378
rect 3056 4224 3108 4276
rect 8208 4224 8260 4276
rect 9772 4224 9824 4276
rect 15936 4224 15988 4276
rect 4988 4156 5040 4208
rect 5448 4156 5500 4208
rect 8944 4156 8996 4208
rect 11612 4199 11664 4208
rect 11612 4165 11621 4199
rect 11621 4165 11655 4199
rect 11655 4165 11664 4199
rect 11612 4156 11664 4165
rect 5080 4131 5132 4140
rect 5080 4097 5089 4131
rect 5089 4097 5123 4131
rect 5123 4097 5132 4131
rect 5080 4088 5132 4097
rect 5172 4088 5224 4140
rect 6920 4131 6972 4140
rect 6920 4097 6929 4131
rect 6929 4097 6963 4131
rect 6963 4097 6972 4131
rect 6920 4088 6972 4097
rect 7472 4131 7524 4140
rect 6552 4020 6604 4072
rect 6644 4063 6696 4072
rect 6644 4029 6653 4063
rect 6653 4029 6687 4063
rect 6687 4029 6696 4063
rect 7104 4063 7156 4072
rect 6644 4020 6696 4029
rect 7104 4029 7113 4063
rect 7113 4029 7147 4063
rect 7147 4029 7156 4063
rect 7104 4020 7156 4029
rect 3976 3952 4028 4004
rect 4528 3952 4580 4004
rect 5908 3952 5960 4004
rect 7472 4097 7481 4131
rect 7481 4097 7515 4131
rect 7515 4097 7524 4131
rect 7472 4088 7524 4097
rect 9772 4088 9824 4140
rect 8760 4020 8812 4072
rect 9680 4063 9732 4072
rect 3516 3884 3568 3936
rect 5540 3884 5592 3936
rect 6828 3927 6880 3936
rect 6828 3893 6837 3927
rect 6837 3893 6871 3927
rect 6871 3893 6880 3927
rect 6828 3884 6880 3893
rect 9680 4029 9689 4063
rect 9689 4029 9723 4063
rect 9723 4029 9732 4063
rect 9680 4020 9732 4029
rect 10784 4088 10836 4140
rect 10876 4131 10928 4140
rect 10876 4097 10885 4131
rect 10885 4097 10919 4131
rect 10919 4097 10928 4131
rect 10876 4088 10928 4097
rect 11520 4088 11572 4140
rect 12072 4131 12124 4140
rect 12072 4097 12081 4131
rect 12081 4097 12115 4131
rect 12115 4097 12124 4131
rect 12072 4088 12124 4097
rect 11428 4020 11480 4072
rect 11704 4063 11756 4072
rect 11704 4029 11713 4063
rect 11713 4029 11747 4063
rect 11747 4029 11756 4063
rect 11704 4020 11756 4029
rect 10784 3952 10836 4004
rect 12348 4088 12400 4140
rect 12624 4131 12676 4140
rect 12624 4097 12629 4131
rect 12629 4097 12663 4131
rect 12663 4097 12676 4131
rect 13360 4131 13412 4140
rect 12624 4088 12676 4097
rect 13360 4097 13369 4131
rect 13369 4097 13403 4131
rect 13403 4097 13412 4131
rect 13360 4088 13412 4097
rect 15200 4088 15252 4140
rect 18144 4088 18196 4140
rect 12624 3952 12676 4004
rect 17592 3952 17644 4004
rect 18328 4020 18380 4072
rect 12808 3884 12860 3936
rect 14188 3884 14240 3936
rect 14648 3884 14700 3936
rect 16948 3884 17000 3936
rect 18052 3927 18104 3936
rect 18052 3893 18061 3927
rect 18061 3893 18095 3927
rect 18095 3893 18104 3927
rect 18052 3884 18104 3893
rect 3110 3782 3162 3834
rect 3174 3782 3226 3834
rect 3238 3782 3290 3834
rect 3302 3782 3354 3834
rect 3366 3782 3418 3834
rect 6210 3782 6262 3834
rect 6274 3782 6326 3834
rect 6338 3782 6390 3834
rect 6402 3782 6454 3834
rect 6466 3782 6518 3834
rect 9310 3782 9362 3834
rect 9374 3782 9426 3834
rect 9438 3782 9490 3834
rect 9502 3782 9554 3834
rect 9566 3782 9618 3834
rect 12410 3782 12462 3834
rect 12474 3782 12526 3834
rect 12538 3782 12590 3834
rect 12602 3782 12654 3834
rect 12666 3782 12718 3834
rect 15510 3782 15562 3834
rect 15574 3782 15626 3834
rect 15638 3782 15690 3834
rect 15702 3782 15754 3834
rect 15766 3782 15818 3834
rect 756 3587 808 3596
rect 756 3553 765 3587
rect 765 3553 799 3587
rect 799 3553 808 3587
rect 756 3544 808 3553
rect 2320 3544 2372 3596
rect 2412 3476 2464 3528
rect 5356 3680 5408 3732
rect 5632 3723 5684 3732
rect 5632 3689 5641 3723
rect 5641 3689 5675 3723
rect 5675 3689 5684 3723
rect 5632 3680 5684 3689
rect 6828 3680 6880 3732
rect 7472 3680 7524 3732
rect 9680 3680 9732 3732
rect 11704 3680 11756 3732
rect 3884 3655 3936 3664
rect 3884 3621 3893 3655
rect 3893 3621 3927 3655
rect 3927 3621 3936 3655
rect 3884 3612 3936 3621
rect 4068 3612 4120 3664
rect 6368 3612 6420 3664
rect 6644 3612 6696 3664
rect 12808 3680 12860 3732
rect 12900 3680 12952 3732
rect 2872 3519 2924 3528
rect 2872 3485 2881 3519
rect 2881 3485 2915 3519
rect 2915 3485 2924 3519
rect 2872 3476 2924 3485
rect 3608 3519 3660 3528
rect 3608 3485 3617 3519
rect 3617 3485 3651 3519
rect 3651 3485 3660 3519
rect 3608 3476 3660 3485
rect 3884 3519 3936 3528
rect 3884 3485 3893 3519
rect 3893 3485 3927 3519
rect 3927 3485 3936 3519
rect 3884 3476 3936 3485
rect 4160 3476 4212 3528
rect 4344 3519 4396 3528
rect 4344 3485 4353 3519
rect 4353 3485 4387 3519
rect 4387 3485 4396 3519
rect 4344 3476 4396 3485
rect 4528 3519 4580 3528
rect 4528 3485 4537 3519
rect 4537 3485 4571 3519
rect 4571 3485 4580 3519
rect 7104 3587 7156 3596
rect 7104 3553 7113 3587
rect 7113 3553 7147 3587
rect 7147 3553 7156 3587
rect 7104 3544 7156 3553
rect 18144 3655 18196 3664
rect 18144 3621 18153 3655
rect 18153 3621 18187 3655
rect 18187 3621 18196 3655
rect 18144 3612 18196 3621
rect 4528 3476 4580 3485
rect 5080 3476 5132 3528
rect 5356 3476 5408 3528
rect 5908 3519 5960 3528
rect 5908 3485 5917 3519
rect 5917 3485 5951 3519
rect 5951 3485 5960 3519
rect 5908 3476 5960 3485
rect 3976 3408 4028 3460
rect 3884 3340 3936 3392
rect 5448 3408 5500 3460
rect 7288 3476 7340 3528
rect 9128 3519 9180 3528
rect 9128 3485 9137 3519
rect 9137 3485 9171 3519
rect 9171 3485 9180 3519
rect 9772 3519 9824 3528
rect 9128 3476 9180 3485
rect 9772 3485 9781 3519
rect 9781 3485 9815 3519
rect 9815 3485 9824 3519
rect 10876 3544 10928 3596
rect 9772 3476 9824 3485
rect 5632 3340 5684 3392
rect 8760 3408 8812 3460
rect 10692 3476 10744 3528
rect 13084 3476 13136 3528
rect 14556 3544 14608 3596
rect 15844 3587 15896 3596
rect 15844 3553 15853 3587
rect 15853 3553 15887 3587
rect 15887 3553 15896 3587
rect 15844 3544 15896 3553
rect 17592 3587 17644 3596
rect 17592 3553 17601 3587
rect 17601 3553 17635 3587
rect 17635 3553 17644 3587
rect 17592 3544 17644 3553
rect 14188 3519 14240 3528
rect 14188 3485 14197 3519
rect 14197 3485 14231 3519
rect 14231 3485 14240 3519
rect 14188 3476 14240 3485
rect 15108 3476 15160 3528
rect 16212 3519 16264 3528
rect 12072 3408 12124 3460
rect 12256 3408 12308 3460
rect 13820 3408 13872 3460
rect 16212 3485 16221 3519
rect 16221 3485 16255 3519
rect 16255 3485 16264 3519
rect 16212 3476 16264 3485
rect 18328 3519 18380 3528
rect 18328 3485 18337 3519
rect 18337 3485 18371 3519
rect 18371 3485 18380 3519
rect 18328 3476 18380 3485
rect 6644 3383 6696 3392
rect 6644 3349 6653 3383
rect 6653 3349 6687 3383
rect 6687 3349 6696 3383
rect 6644 3340 6696 3349
rect 6736 3383 6788 3392
rect 6736 3349 6745 3383
rect 6745 3349 6779 3383
rect 6779 3349 6788 3383
rect 6736 3340 6788 3349
rect 7104 3340 7156 3392
rect 8668 3340 8720 3392
rect 13360 3340 13412 3392
rect 16304 3340 16356 3392
rect 4660 3238 4712 3290
rect 4724 3238 4776 3290
rect 4788 3238 4840 3290
rect 4852 3238 4904 3290
rect 4916 3238 4968 3290
rect 7760 3238 7812 3290
rect 7824 3238 7876 3290
rect 7888 3238 7940 3290
rect 7952 3238 8004 3290
rect 8016 3238 8068 3290
rect 10860 3238 10912 3290
rect 10924 3238 10976 3290
rect 10988 3238 11040 3290
rect 11052 3238 11104 3290
rect 11116 3238 11168 3290
rect 13960 3238 14012 3290
rect 14024 3238 14076 3290
rect 14088 3238 14140 3290
rect 14152 3238 14204 3290
rect 14216 3238 14268 3290
rect 17060 3238 17112 3290
rect 17124 3238 17176 3290
rect 17188 3238 17240 3290
rect 17252 3238 17304 3290
rect 17316 3238 17368 3290
rect 3516 3136 3568 3188
rect 3608 3179 3660 3188
rect 3608 3145 3617 3179
rect 3617 3145 3651 3179
rect 3651 3145 3660 3179
rect 3608 3136 3660 3145
rect 2872 3068 2924 3120
rect 4436 3136 4488 3188
rect 14556 3179 14608 3188
rect 5816 3068 5868 3120
rect 3884 3000 3936 3052
rect 4160 3000 4212 3052
rect 4528 3000 4580 3052
rect 4804 3043 4856 3052
rect 4804 3009 4813 3043
rect 4813 3009 4847 3043
rect 4847 3009 4856 3043
rect 4804 3000 4856 3009
rect 5540 3043 5592 3052
rect 5540 3009 5549 3043
rect 5549 3009 5583 3043
rect 5583 3009 5592 3043
rect 5540 3000 5592 3009
rect 5908 3043 5960 3052
rect 5908 3009 5917 3043
rect 5917 3009 5951 3043
rect 5951 3009 5960 3043
rect 5908 3000 5960 3009
rect 4344 2932 4396 2984
rect 5632 2975 5684 2984
rect 5632 2941 5641 2975
rect 5641 2941 5675 2975
rect 5675 2941 5684 2975
rect 5632 2932 5684 2941
rect 6368 3068 6420 3120
rect 4436 2864 4488 2916
rect 7196 3000 7248 3052
rect 7472 3068 7524 3120
rect 8300 3111 8352 3120
rect 8300 3077 8309 3111
rect 8309 3077 8343 3111
rect 8343 3077 8352 3111
rect 8300 3068 8352 3077
rect 9128 3068 9180 3120
rect 11336 3068 11388 3120
rect 7564 3043 7616 3052
rect 7564 3009 7573 3043
rect 7573 3009 7607 3043
rect 7607 3009 7616 3043
rect 7564 3000 7616 3009
rect 7656 3043 7708 3052
rect 7656 3009 7665 3043
rect 7665 3009 7699 3043
rect 7699 3009 7708 3043
rect 7840 3043 7892 3052
rect 7656 3000 7708 3009
rect 7840 3009 7849 3043
rect 7849 3009 7883 3043
rect 7883 3009 7892 3043
rect 7840 3000 7892 3009
rect 8668 3000 8720 3052
rect 14556 3145 14565 3179
rect 14565 3145 14599 3179
rect 14599 3145 14608 3179
rect 14556 3136 14608 3145
rect 15384 3136 15436 3188
rect 16212 3136 16264 3188
rect 18328 3179 18380 3188
rect 18328 3145 18337 3179
rect 18337 3145 18371 3179
rect 18371 3145 18380 3179
rect 18328 3136 18380 3145
rect 12900 3111 12952 3120
rect 12900 3077 12909 3111
rect 12909 3077 12943 3111
rect 12943 3077 12952 3111
rect 12900 3068 12952 3077
rect 13360 3068 13412 3120
rect 16396 3068 16448 3120
rect 12808 3043 12860 3052
rect 10600 2932 10652 2984
rect 12256 2932 12308 2984
rect 12808 3009 12817 3043
rect 12817 3009 12851 3043
rect 12851 3009 12860 3043
rect 12808 3000 12860 3009
rect 12900 2932 12952 2984
rect 13820 3000 13872 3052
rect 14648 2975 14700 2984
rect 14648 2941 14657 2975
rect 14657 2941 14691 2975
rect 14691 2941 14700 2975
rect 14648 2932 14700 2941
rect 15844 2932 15896 2984
rect 17960 3000 18012 3052
rect 17408 2975 17460 2984
rect 17408 2941 17417 2975
rect 17417 2941 17451 2975
rect 17451 2941 17460 2975
rect 17408 2932 17460 2941
rect 17592 2932 17644 2984
rect 6644 2796 6696 2848
rect 8760 2796 8812 2848
rect 10232 2796 10284 2848
rect 11796 2796 11848 2848
rect 3110 2694 3162 2746
rect 3174 2694 3226 2746
rect 3238 2694 3290 2746
rect 3302 2694 3354 2746
rect 3366 2694 3418 2746
rect 6210 2694 6262 2746
rect 6274 2694 6326 2746
rect 6338 2694 6390 2746
rect 6402 2694 6454 2746
rect 6466 2694 6518 2746
rect 9310 2694 9362 2746
rect 9374 2694 9426 2746
rect 9438 2694 9490 2746
rect 9502 2694 9554 2746
rect 9566 2694 9618 2746
rect 12410 2694 12462 2746
rect 12474 2694 12526 2746
rect 12538 2694 12590 2746
rect 12602 2694 12654 2746
rect 12666 2694 12718 2746
rect 15510 2694 15562 2746
rect 15574 2694 15626 2746
rect 15638 2694 15690 2746
rect 15702 2694 15754 2746
rect 15766 2694 15818 2746
rect 7564 2592 7616 2644
rect 12256 2635 12308 2644
rect 12256 2601 12265 2635
rect 12265 2601 12299 2635
rect 12299 2601 12308 2635
rect 12256 2592 12308 2601
rect 756 2499 808 2508
rect 756 2465 765 2499
rect 765 2465 799 2499
rect 799 2465 808 2499
rect 756 2456 808 2465
rect 3884 2524 3936 2576
rect 3700 2456 3752 2508
rect 5632 2524 5684 2576
rect 7656 2524 7708 2576
rect 12808 2524 12860 2576
rect 16488 2524 16540 2576
rect 5264 2456 5316 2508
rect 4436 2431 4488 2440
rect 2412 2320 2464 2372
rect 2688 2320 2740 2372
rect 4436 2397 4445 2431
rect 4445 2397 4479 2431
rect 4479 2397 4488 2431
rect 4436 2388 4488 2397
rect 5724 2456 5776 2508
rect 5816 2431 5868 2440
rect 5816 2397 5825 2431
rect 5825 2397 5859 2431
rect 5859 2397 5868 2431
rect 5816 2388 5868 2397
rect 15384 2499 15436 2508
rect 7104 2388 7156 2440
rect 7196 2388 7248 2440
rect 8300 2388 8352 2440
rect 8576 2431 8628 2440
rect 8576 2397 8585 2431
rect 8585 2397 8619 2431
rect 8619 2397 8628 2431
rect 8576 2388 8628 2397
rect 8668 2431 8720 2440
rect 8668 2397 8677 2431
rect 8677 2397 8711 2431
rect 8711 2397 8720 2431
rect 10232 2431 10284 2440
rect 8668 2388 8720 2397
rect 10232 2397 10241 2431
rect 10241 2397 10275 2431
rect 10275 2397 10284 2431
rect 10232 2388 10284 2397
rect 11796 2431 11848 2440
rect 11796 2397 11805 2431
rect 11805 2397 11839 2431
rect 11839 2397 11848 2431
rect 12256 2431 12308 2440
rect 11796 2388 11848 2397
rect 12256 2397 12265 2431
rect 12265 2397 12299 2431
rect 12299 2397 12308 2431
rect 12256 2388 12308 2397
rect 15384 2465 15393 2499
rect 15393 2465 15427 2499
rect 15427 2465 15436 2499
rect 15384 2456 15436 2465
rect 15752 2499 15804 2508
rect 15752 2465 15761 2499
rect 15761 2465 15795 2499
rect 15795 2465 15804 2499
rect 17960 2499 18012 2508
rect 15752 2456 15804 2465
rect 17960 2465 17969 2499
rect 17969 2465 18003 2499
rect 18003 2465 18012 2499
rect 17960 2456 18012 2465
rect 14556 2388 14608 2440
rect 15568 2431 15620 2440
rect 15568 2397 15577 2431
rect 15577 2397 15611 2431
rect 15611 2397 15620 2431
rect 18512 2431 18564 2440
rect 15568 2388 15620 2397
rect 18512 2397 18521 2431
rect 18521 2397 18555 2431
rect 18555 2397 18564 2431
rect 18512 2388 18564 2397
rect 3516 2320 3568 2372
rect 5264 2320 5316 2372
rect 7840 2320 7892 2372
rect 2964 2252 3016 2304
rect 3608 2252 3660 2304
rect 4068 2252 4120 2304
rect 4344 2252 4396 2304
rect 8208 2252 8260 2304
rect 12164 2320 12216 2372
rect 13176 2320 13228 2372
rect 15200 2320 15252 2372
rect 15384 2320 15436 2372
rect 16304 2320 16356 2372
rect 16396 2320 16448 2372
rect 17408 2320 17460 2372
rect 9128 2252 9180 2304
rect 12716 2295 12768 2304
rect 12716 2261 12725 2295
rect 12725 2261 12759 2295
rect 12759 2261 12768 2295
rect 12716 2252 12768 2261
rect 14372 2252 14424 2304
rect 15752 2295 15804 2304
rect 15752 2261 15761 2295
rect 15761 2261 15795 2295
rect 15795 2261 15804 2295
rect 15752 2252 15804 2261
rect 16028 2252 16080 2304
rect 4660 2150 4712 2202
rect 4724 2150 4776 2202
rect 4788 2150 4840 2202
rect 4852 2150 4904 2202
rect 4916 2150 4968 2202
rect 7760 2150 7812 2202
rect 7824 2150 7876 2202
rect 7888 2150 7940 2202
rect 7952 2150 8004 2202
rect 8016 2150 8068 2202
rect 10860 2150 10912 2202
rect 10924 2150 10976 2202
rect 10988 2150 11040 2202
rect 11052 2150 11104 2202
rect 11116 2150 11168 2202
rect 13960 2150 14012 2202
rect 14024 2150 14076 2202
rect 14088 2150 14140 2202
rect 14152 2150 14204 2202
rect 14216 2150 14268 2202
rect 17060 2150 17112 2202
rect 17124 2150 17176 2202
rect 17188 2150 17240 2202
rect 17252 2150 17304 2202
rect 17316 2150 17368 2202
rect 3516 2091 3568 2100
rect 3516 2057 3525 2091
rect 3525 2057 3559 2091
rect 3559 2057 3568 2091
rect 3516 2048 3568 2057
rect 3700 2091 3752 2100
rect 3700 2057 3709 2091
rect 3709 2057 3743 2091
rect 3743 2057 3752 2091
rect 3700 2048 3752 2057
rect 4344 2091 4396 2100
rect 4344 2057 4353 2091
rect 4353 2057 4387 2091
rect 4387 2057 4396 2091
rect 4344 2048 4396 2057
rect 5908 2048 5960 2100
rect 7288 2048 7340 2100
rect 8668 2048 8720 2100
rect 3608 1955 3660 1964
rect 3608 1921 3617 1955
rect 3617 1921 3651 1955
rect 3651 1921 3660 1955
rect 3608 1912 3660 1921
rect 4436 1980 4488 2032
rect 5264 1980 5316 2032
rect 5172 1912 5224 1964
rect 4528 1887 4580 1896
rect 4528 1853 4537 1887
rect 4537 1853 4571 1887
rect 4571 1853 4580 1887
rect 5540 1887 5592 1896
rect 4528 1844 4580 1853
rect 5540 1853 5549 1887
rect 5549 1853 5583 1887
rect 5583 1853 5592 1887
rect 5540 1844 5592 1853
rect 9036 1980 9088 2032
rect 11612 2048 11664 2100
rect 12256 2091 12308 2100
rect 12256 2057 12265 2091
rect 12265 2057 12299 2091
rect 12299 2057 12308 2091
rect 12256 2048 12308 2057
rect 7380 1955 7432 1964
rect 7380 1921 7389 1955
rect 7389 1921 7423 1955
rect 7423 1921 7432 1955
rect 7380 1912 7432 1921
rect 7656 1887 7708 1896
rect 7656 1853 7665 1887
rect 7665 1853 7699 1887
rect 7699 1853 7708 1887
rect 7656 1844 7708 1853
rect 5632 1776 5684 1828
rect 6000 1751 6052 1760
rect 6000 1717 6009 1751
rect 6009 1717 6043 1751
rect 6043 1717 6052 1751
rect 6000 1708 6052 1717
rect 7288 1708 7340 1760
rect 10876 1955 10928 1964
rect 10876 1921 10885 1955
rect 10885 1921 10919 1955
rect 10919 1921 10928 1955
rect 10876 1912 10928 1921
rect 12716 2048 12768 2100
rect 13176 2048 13228 2100
rect 14556 2048 14608 2100
rect 15568 2048 15620 2100
rect 17408 2091 17460 2100
rect 17408 2057 17417 2091
rect 17417 2057 17451 2091
rect 17451 2057 17460 2091
rect 17408 2048 17460 2057
rect 9220 1708 9272 1760
rect 10324 1844 10376 1896
rect 11336 1844 11388 1896
rect 12900 1912 12952 1964
rect 12992 1955 13044 1964
rect 12992 1921 13001 1955
rect 13001 1921 13035 1955
rect 13035 1921 13044 1955
rect 13820 1980 13872 2032
rect 12992 1912 13044 1921
rect 14372 1955 14424 1964
rect 14372 1921 14381 1955
rect 14381 1921 14415 1955
rect 14415 1921 14424 1955
rect 15384 1980 15436 2032
rect 15844 1980 15896 2032
rect 16028 1980 16080 2032
rect 16396 1980 16448 2032
rect 14372 1912 14424 1921
rect 15200 1844 15252 1896
rect 15660 1776 15712 1828
rect 16948 1708 17000 1760
rect 3110 1606 3162 1658
rect 3174 1606 3226 1658
rect 3238 1606 3290 1658
rect 3302 1606 3354 1658
rect 3366 1606 3418 1658
rect 6210 1606 6262 1658
rect 6274 1606 6326 1658
rect 6338 1606 6390 1658
rect 6402 1606 6454 1658
rect 6466 1606 6518 1658
rect 9310 1606 9362 1658
rect 9374 1606 9426 1658
rect 9438 1606 9490 1658
rect 9502 1606 9554 1658
rect 9566 1606 9618 1658
rect 12410 1606 12462 1658
rect 12474 1606 12526 1658
rect 12538 1606 12590 1658
rect 12602 1606 12654 1658
rect 12666 1606 12718 1658
rect 15510 1606 15562 1658
rect 15574 1606 15626 1658
rect 15638 1606 15690 1658
rect 15702 1606 15754 1658
rect 15766 1606 15818 1658
rect 3884 1504 3936 1556
rect 5540 1547 5592 1556
rect 5540 1513 5549 1547
rect 5549 1513 5583 1547
rect 5583 1513 5592 1547
rect 5540 1504 5592 1513
rect 10876 1504 10928 1556
rect 756 1411 808 1420
rect 756 1377 765 1411
rect 765 1377 799 1411
rect 799 1377 808 1411
rect 756 1368 808 1377
rect 5724 1436 5776 1488
rect 8668 1436 8720 1488
rect 2688 1232 2740 1284
rect 2964 1232 3016 1284
rect 3424 1275 3476 1284
rect 3424 1241 3433 1275
rect 3433 1241 3467 1275
rect 3467 1241 3476 1275
rect 3424 1232 3476 1241
rect 3884 1343 3936 1352
rect 3884 1309 3893 1343
rect 3893 1309 3927 1343
rect 3927 1309 3936 1343
rect 3884 1300 3936 1309
rect 4160 1300 4212 1352
rect 5080 1300 5132 1352
rect 5908 1368 5960 1420
rect 5356 1343 5408 1352
rect 5356 1309 5365 1343
rect 5365 1309 5399 1343
rect 5399 1309 5408 1343
rect 5356 1300 5408 1309
rect 5540 1343 5592 1352
rect 5540 1309 5549 1343
rect 5549 1309 5583 1343
rect 5583 1309 5592 1343
rect 5540 1300 5592 1309
rect 6000 1343 6052 1352
rect 6000 1309 6009 1343
rect 6009 1309 6043 1343
rect 6043 1309 6052 1343
rect 6000 1300 6052 1309
rect 9220 1368 9272 1420
rect 6552 1300 6604 1352
rect 7656 1300 7708 1352
rect 8668 1343 8720 1352
rect 8668 1309 8677 1343
rect 8677 1309 8711 1343
rect 8711 1309 8720 1343
rect 8668 1300 8720 1309
rect 9128 1343 9180 1352
rect 9128 1309 9137 1343
rect 9137 1309 9171 1343
rect 9171 1309 9180 1343
rect 9128 1300 9180 1309
rect 10140 1411 10192 1420
rect 10140 1377 10149 1411
rect 10149 1377 10183 1411
rect 10183 1377 10192 1411
rect 10140 1368 10192 1377
rect 11336 1368 11388 1420
rect 16488 1411 16540 1420
rect 16488 1377 16497 1411
rect 16497 1377 16531 1411
rect 16531 1377 16540 1411
rect 16488 1368 16540 1377
rect 5080 1164 5132 1216
rect 5264 1164 5316 1216
rect 6644 1232 6696 1284
rect 10324 1232 10376 1284
rect 10784 1232 10836 1284
rect 11060 1275 11112 1284
rect 11060 1241 11069 1275
rect 11069 1241 11103 1275
rect 11103 1241 11112 1275
rect 11060 1232 11112 1241
rect 12992 1300 13044 1352
rect 13820 1300 13872 1352
rect 18236 1343 18288 1352
rect 18236 1309 18245 1343
rect 18245 1309 18279 1343
rect 18279 1309 18288 1343
rect 18236 1300 18288 1309
rect 18328 1343 18380 1352
rect 18328 1309 18337 1343
rect 18337 1309 18371 1343
rect 18371 1309 18380 1343
rect 18328 1300 18380 1309
rect 14464 1275 14516 1284
rect 6920 1207 6972 1216
rect 6920 1173 6929 1207
rect 6929 1173 6963 1207
rect 6963 1173 6972 1207
rect 6920 1164 6972 1173
rect 14464 1241 14473 1275
rect 14473 1241 14507 1275
rect 14507 1241 14516 1275
rect 14464 1232 14516 1241
rect 14924 1232 14976 1284
rect 16212 1275 16264 1284
rect 13636 1164 13688 1216
rect 14372 1164 14424 1216
rect 16212 1241 16221 1275
rect 16221 1241 16255 1275
rect 16255 1241 16264 1275
rect 16212 1232 16264 1241
rect 16304 1232 16356 1284
rect 16396 1164 16448 1216
rect 17960 1207 18012 1216
rect 17960 1173 17969 1207
rect 17969 1173 18003 1207
rect 18003 1173 18012 1207
rect 17960 1164 18012 1173
rect 4660 1062 4712 1114
rect 4724 1062 4776 1114
rect 4788 1062 4840 1114
rect 4852 1062 4904 1114
rect 4916 1062 4968 1114
rect 7760 1062 7812 1114
rect 7824 1062 7876 1114
rect 7888 1062 7940 1114
rect 7952 1062 8004 1114
rect 8016 1062 8068 1114
rect 10860 1062 10912 1114
rect 10924 1062 10976 1114
rect 10988 1062 11040 1114
rect 11052 1062 11104 1114
rect 11116 1062 11168 1114
rect 13960 1062 14012 1114
rect 14024 1062 14076 1114
rect 14088 1062 14140 1114
rect 14152 1062 14204 1114
rect 14216 1062 14268 1114
rect 17060 1062 17112 1114
rect 17124 1062 17176 1114
rect 17188 1062 17240 1114
rect 17252 1062 17304 1114
rect 17316 1062 17368 1114
rect 4068 960 4120 1012
rect 5540 960 5592 1012
rect 6552 960 6604 1012
rect 8944 960 8996 1012
rect 10140 1003 10192 1012
rect 10140 969 10149 1003
rect 10149 969 10183 1003
rect 10183 969 10192 1003
rect 10140 960 10192 969
rect 3424 824 3476 876
rect 3976 867 4028 876
rect 3976 833 3985 867
rect 3985 833 4019 867
rect 4019 833 4028 867
rect 4160 867 4212 876
rect 3976 824 4028 833
rect 4160 833 4169 867
rect 4169 833 4203 867
rect 4203 833 4212 867
rect 4160 824 4212 833
rect 5448 867 5500 876
rect 5448 833 5457 867
rect 5457 833 5491 867
rect 5491 833 5500 867
rect 5448 824 5500 833
rect 9036 892 9088 944
rect 11244 960 11296 1012
rect 13636 1003 13688 1012
rect 3884 688 3936 740
rect 5264 688 5316 740
rect 7380 756 7432 808
rect 8116 756 8168 808
rect 10784 892 10836 944
rect 13636 969 13645 1003
rect 13645 969 13679 1003
rect 13679 969 13688 1003
rect 13636 960 13688 969
rect 13820 960 13872 1012
rect 14372 960 14424 1012
rect 16212 960 16264 1012
rect 10876 867 10928 876
rect 10876 833 10885 867
rect 10885 833 10919 867
rect 10919 833 10928 867
rect 10876 824 10928 833
rect 11060 824 11112 876
rect 12164 867 12216 876
rect 12164 833 12173 867
rect 12173 833 12207 867
rect 12207 833 12216 867
rect 12164 824 12216 833
rect 12716 824 12768 876
rect 14648 892 14700 944
rect 17960 892 18012 944
rect 10324 756 10376 808
rect 10968 799 11020 808
rect 10968 765 10977 799
rect 10977 765 11011 799
rect 11011 765 11020 799
rect 10968 756 11020 765
rect 11060 688 11112 740
rect 11336 688 11388 740
rect 2964 620 3016 672
rect 6000 663 6052 672
rect 6000 629 6009 663
rect 6009 629 6043 663
rect 6043 629 6052 663
rect 6000 620 6052 629
rect 9128 663 9180 672
rect 9128 629 9137 663
rect 9137 629 9171 663
rect 9171 629 9180 663
rect 9128 620 9180 629
rect 10508 620 10560 672
rect 12992 799 13044 808
rect 12992 765 13001 799
rect 13001 765 13035 799
rect 13035 765 13044 799
rect 12992 756 13044 765
rect 14464 756 14516 808
rect 17776 867 17828 876
rect 17776 833 17785 867
rect 17785 833 17819 867
rect 17819 833 17828 867
rect 17776 824 17828 833
rect 18052 824 18104 876
rect 15844 688 15896 740
rect 17776 688 17828 740
rect 13176 663 13228 672
rect 13176 629 13185 663
rect 13185 629 13219 663
rect 13219 629 13228 663
rect 13176 620 13228 629
rect 17960 620 18012 672
rect 3110 518 3162 570
rect 3174 518 3226 570
rect 3238 518 3290 570
rect 3302 518 3354 570
rect 3366 518 3418 570
rect 6210 518 6262 570
rect 6274 518 6326 570
rect 6338 518 6390 570
rect 6402 518 6454 570
rect 6466 518 6518 570
rect 9310 518 9362 570
rect 9374 518 9426 570
rect 9438 518 9490 570
rect 9502 518 9554 570
rect 9566 518 9618 570
rect 12410 518 12462 570
rect 12474 518 12526 570
rect 12538 518 12590 570
rect 12602 518 12654 570
rect 12666 518 12718 570
rect 15510 518 15562 570
rect 15574 518 15626 570
rect 15638 518 15690 570
rect 15702 518 15754 570
rect 15766 518 15818 570
rect 4160 416 4212 468
rect 8116 459 8168 468
rect 8116 425 8125 459
rect 8125 425 8159 459
rect 8159 425 8168 459
rect 8116 416 8168 425
rect 10876 459 10928 468
rect 10876 425 10885 459
rect 10885 425 10919 459
rect 10919 425 10928 459
rect 10876 416 10928 425
rect 5448 348 5500 400
rect 2964 280 3016 332
rect 6920 348 6972 400
rect 6644 280 6696 332
rect 8668 348 8720 400
rect 12992 416 13044 468
rect 14648 416 14700 468
rect 9128 280 9180 332
rect 10784 280 10836 332
rect 12992 323 13044 332
rect 12992 289 13001 323
rect 13001 289 13035 323
rect 13035 289 13044 323
rect 12992 280 13044 289
rect 16488 416 16540 468
rect 17776 416 17828 468
rect 18328 459 18380 468
rect 18328 425 18337 459
rect 18337 425 18371 459
rect 18371 425 18380 459
rect 18328 416 18380 425
rect 756 212 808 264
rect 6000 255 6052 264
rect 6000 221 6009 255
rect 6009 221 6043 255
rect 6043 221 6052 255
rect 6000 212 6052 221
rect 8576 212 8628 264
rect 11060 212 11112 264
rect 18512 255 18564 264
rect 18512 221 18521 255
rect 18521 221 18555 255
rect 18555 221 18564 255
rect 18512 212 18564 221
rect 2688 76 2740 128
rect 8208 144 8260 196
rect 10968 144 11020 196
rect 13176 144 13228 196
rect 14924 144 14976 196
rect 17960 144 18012 196
rect 4660 -26 4712 26
rect 4724 -26 4776 26
rect 4788 -26 4840 26
rect 4852 -26 4904 26
rect 4916 -26 4968 26
rect 7760 -26 7812 26
rect 7824 -26 7876 26
rect 7888 -26 7940 26
rect 7952 -26 8004 26
rect 8016 -26 8068 26
rect 10860 -26 10912 26
rect 10924 -26 10976 26
rect 10988 -26 11040 26
rect 11052 -26 11104 26
rect 11116 -26 11168 26
rect 13960 -26 14012 26
rect 14024 -26 14076 26
rect 14088 -26 14140 26
rect 14152 -26 14204 26
rect 14216 -26 14268 26
rect 17060 -26 17112 26
rect 17124 -26 17176 26
rect 17188 -26 17240 26
rect 17252 -26 17304 26
rect 17316 -26 17368 26
<< metal2 >>
rect 1398 11200 1454 12000
rect 4250 11200 4306 12000
rect 7102 11200 7158 12000
rect 9954 11200 10010 12000
rect 12806 11200 12862 12000
rect 15396 11206 15608 11234
rect 1308 10668 1360 10674
rect 1412 10656 1440 11200
rect 3792 10804 3844 10810
rect 3792 10746 3844 10752
rect 2136 10736 2188 10742
rect 2136 10678 2188 10684
rect 1360 10628 1440 10656
rect 1308 10610 1360 10616
rect 296 10124 348 10130
rect 296 10066 348 10072
rect 308 9042 336 10066
rect 2148 9994 2176 10678
rect 2688 10600 2740 10606
rect 2688 10542 2740 10548
rect 2964 10600 3016 10606
rect 2964 10542 3016 10548
rect 2320 10464 2372 10470
rect 2320 10406 2372 10412
rect 2332 10062 2360 10406
rect 2700 10266 2728 10542
rect 2688 10260 2740 10266
rect 2688 10202 2740 10208
rect 2976 10130 3004 10542
rect 3110 10364 3418 10384
rect 3110 10362 3116 10364
rect 3172 10362 3196 10364
rect 3252 10362 3276 10364
rect 3332 10362 3356 10364
rect 3412 10362 3418 10364
rect 3172 10310 3174 10362
rect 3354 10310 3356 10362
rect 3110 10308 3116 10310
rect 3172 10308 3196 10310
rect 3252 10308 3276 10310
rect 3332 10308 3356 10310
rect 3412 10308 3418 10310
rect 3110 10288 3418 10308
rect 2964 10124 3016 10130
rect 2964 10066 3016 10072
rect 3424 10124 3476 10130
rect 3424 10066 3476 10072
rect 2320 10056 2372 10062
rect 2320 9998 2372 10004
rect 3240 10056 3292 10062
rect 3240 9998 3292 10004
rect 572 9988 624 9994
rect 572 9930 624 9936
rect 2136 9988 2188 9994
rect 2136 9930 2188 9936
rect 2872 9988 2924 9994
rect 2872 9930 2924 9936
rect 584 9722 612 9930
rect 2228 9920 2280 9926
rect 2228 9862 2280 9868
rect 2688 9920 2740 9926
rect 2688 9862 2740 9868
rect 572 9716 624 9722
rect 572 9658 624 9664
rect 2240 9654 2268 9862
rect 2700 9704 2728 9862
rect 2780 9716 2832 9722
rect 2700 9676 2780 9704
rect 2780 9658 2832 9664
rect 2228 9648 2280 9654
rect 2228 9590 2280 9596
rect 2884 9178 2912 9930
rect 3252 9654 3280 9998
rect 3240 9648 3292 9654
rect 3240 9590 3292 9596
rect 3252 9450 3280 9590
rect 3436 9450 3464 10066
rect 2964 9444 3016 9450
rect 2964 9386 3016 9392
rect 3240 9444 3292 9450
rect 3240 9386 3292 9392
rect 3424 9444 3476 9450
rect 3424 9386 3476 9392
rect 2872 9172 2924 9178
rect 2872 9114 2924 9120
rect 296 9036 348 9042
rect 296 8978 348 8984
rect 2504 9036 2556 9042
rect 2504 8978 2556 8984
rect 308 7954 336 8978
rect 1860 8900 1912 8906
rect 1860 8842 1912 8848
rect 296 7948 348 7954
rect 296 7890 348 7896
rect 308 6254 336 7890
rect 1872 7818 1900 8842
rect 2320 8832 2372 8838
rect 2320 8774 2372 8780
rect 2332 8634 2360 8774
rect 2516 8634 2544 8978
rect 2780 8968 2832 8974
rect 2780 8910 2832 8916
rect 2320 8628 2372 8634
rect 2320 8570 2372 8576
rect 2504 8628 2556 8634
rect 2504 8570 2556 8576
rect 2792 8566 2820 8910
rect 2780 8560 2832 8566
rect 2780 8502 2832 8508
rect 2884 8430 2912 9114
rect 2976 9042 3004 9386
rect 3110 9276 3418 9296
rect 3110 9274 3116 9276
rect 3172 9274 3196 9276
rect 3252 9274 3276 9276
rect 3332 9274 3356 9276
rect 3412 9274 3418 9276
rect 3172 9222 3174 9274
rect 3354 9222 3356 9274
rect 3110 9220 3116 9222
rect 3172 9220 3196 9222
rect 3252 9220 3276 9222
rect 3332 9220 3356 9222
rect 3412 9220 3418 9222
rect 3110 9200 3418 9220
rect 2964 9036 3016 9042
rect 2964 8978 3016 8984
rect 3608 8968 3660 8974
rect 3608 8910 3660 8916
rect 3240 8832 3292 8838
rect 3240 8774 3292 8780
rect 3252 8634 3280 8774
rect 3240 8628 3292 8634
rect 3240 8570 3292 8576
rect 2964 8492 3016 8498
rect 2964 8434 3016 8440
rect 2872 8424 2924 8430
rect 2872 8366 2924 8372
rect 2976 8294 3004 8434
rect 3620 8430 3648 8910
rect 3700 8492 3752 8498
rect 3700 8434 3752 8440
rect 3608 8424 3660 8430
rect 3608 8366 3660 8372
rect 2964 8288 3016 8294
rect 2964 8230 3016 8236
rect 3110 8188 3418 8208
rect 3110 8186 3116 8188
rect 3172 8186 3196 8188
rect 3252 8186 3276 8188
rect 3332 8186 3356 8188
rect 3412 8186 3418 8188
rect 3172 8134 3174 8186
rect 3354 8134 3356 8186
rect 3110 8132 3116 8134
rect 3172 8132 3196 8134
rect 3252 8132 3276 8134
rect 3332 8132 3356 8134
rect 3412 8132 3418 8134
rect 3110 8112 3418 8132
rect 3620 7886 3648 8366
rect 3516 7880 3568 7886
rect 3516 7822 3568 7828
rect 3608 7880 3660 7886
rect 3608 7822 3660 7828
rect 572 7812 624 7818
rect 572 7754 624 7760
rect 1860 7812 1912 7818
rect 1860 7754 1912 7760
rect 2412 7812 2464 7818
rect 2412 7754 2464 7760
rect 584 7546 612 7754
rect 572 7540 624 7546
rect 572 7482 624 7488
rect 572 6656 624 6662
rect 572 6598 624 6604
rect 584 6390 612 6598
rect 572 6384 624 6390
rect 572 6326 624 6332
rect 296 6248 348 6254
rect 296 6190 348 6196
rect 308 5778 336 6190
rect 1872 6186 1900 7754
rect 2044 7744 2096 7750
rect 2044 7686 2096 7692
rect 1952 7540 2004 7546
rect 1952 7482 2004 7488
rect 1964 6866 1992 7482
rect 2056 7410 2084 7686
rect 2044 7404 2096 7410
rect 2044 7346 2096 7352
rect 2424 7342 2452 7754
rect 2504 7744 2556 7750
rect 2504 7686 2556 7692
rect 2516 7410 2544 7686
rect 3148 7540 3200 7546
rect 3148 7482 3200 7488
rect 2596 7472 2648 7478
rect 2596 7414 2648 7420
rect 2504 7404 2556 7410
rect 2504 7346 2556 7352
rect 2412 7336 2464 7342
rect 2412 7278 2464 7284
rect 2320 7268 2372 7274
rect 2320 7210 2372 7216
rect 1952 6860 2004 6866
rect 1952 6802 2004 6808
rect 2044 6724 2096 6730
rect 2044 6666 2096 6672
rect 2056 6458 2084 6666
rect 2044 6452 2096 6458
rect 2044 6394 2096 6400
rect 2332 6322 2360 7210
rect 2424 7206 2452 7278
rect 2412 7200 2464 7206
rect 2412 7142 2464 7148
rect 2608 6662 2636 7414
rect 3160 7410 3188 7482
rect 3528 7410 3556 7822
rect 2780 7404 2832 7410
rect 2780 7346 2832 7352
rect 3148 7404 3200 7410
rect 3148 7346 3200 7352
rect 3332 7404 3384 7410
rect 3332 7346 3384 7352
rect 3516 7404 3568 7410
rect 3516 7346 3568 7352
rect 2688 7200 2740 7206
rect 2688 7142 2740 7148
rect 2700 6798 2728 7142
rect 2792 6934 2820 7346
rect 3344 7188 3372 7346
rect 2976 7160 3372 7188
rect 2780 6928 2832 6934
rect 2780 6870 2832 6876
rect 2976 6866 3004 7160
rect 3110 7100 3418 7120
rect 3110 7098 3116 7100
rect 3172 7098 3196 7100
rect 3252 7098 3276 7100
rect 3332 7098 3356 7100
rect 3412 7098 3418 7100
rect 3172 7046 3174 7098
rect 3354 7046 3356 7098
rect 3110 7044 3116 7046
rect 3172 7044 3196 7046
rect 3252 7044 3276 7046
rect 3332 7044 3356 7046
rect 3412 7044 3418 7046
rect 3110 7024 3418 7044
rect 3240 6928 3292 6934
rect 3240 6870 3292 6876
rect 2964 6860 3016 6866
rect 2964 6802 3016 6808
rect 3252 6798 3280 6870
rect 3528 6798 3556 7346
rect 3620 6934 3648 7822
rect 3712 7750 3740 8434
rect 3700 7744 3752 7750
rect 3700 7686 3752 7692
rect 3712 7546 3740 7686
rect 3700 7540 3752 7546
rect 3700 7482 3752 7488
rect 3608 6928 3660 6934
rect 3608 6870 3660 6876
rect 2688 6792 2740 6798
rect 2688 6734 2740 6740
rect 3240 6792 3292 6798
rect 3240 6734 3292 6740
rect 3516 6792 3568 6798
rect 3516 6734 3568 6740
rect 2412 6656 2464 6662
rect 2412 6598 2464 6604
rect 2596 6656 2648 6662
rect 2596 6598 2648 6604
rect 2424 6322 2452 6598
rect 2320 6316 2372 6322
rect 2320 6258 2372 6264
rect 2412 6316 2464 6322
rect 2412 6258 2464 6264
rect 2608 6254 2636 6598
rect 2596 6248 2648 6254
rect 2596 6190 2648 6196
rect 1860 6180 1912 6186
rect 1860 6122 1912 6128
rect 2412 6180 2464 6186
rect 2412 6122 2464 6128
rect 296 5772 348 5778
rect 296 5714 348 5720
rect 2424 5574 2452 6122
rect 2964 6112 3016 6118
rect 2964 6054 3016 6060
rect 2976 5710 3004 6054
rect 3110 6012 3418 6032
rect 3110 6010 3116 6012
rect 3172 6010 3196 6012
rect 3252 6010 3276 6012
rect 3332 6010 3356 6012
rect 3412 6010 3418 6012
rect 3172 5958 3174 6010
rect 3354 5958 3356 6010
rect 3110 5956 3116 5958
rect 3172 5956 3196 5958
rect 3252 5956 3276 5958
rect 3332 5956 3356 5958
rect 3412 5956 3418 5958
rect 3110 5936 3418 5956
rect 3528 5914 3556 6734
rect 3516 5908 3568 5914
rect 3516 5850 3568 5856
rect 2964 5704 3016 5710
rect 2964 5646 3016 5652
rect 3804 5642 3832 10746
rect 4264 10198 4292 11200
rect 4660 10908 4968 10928
rect 4660 10906 4666 10908
rect 4722 10906 4746 10908
rect 4802 10906 4826 10908
rect 4882 10906 4906 10908
rect 4962 10906 4968 10908
rect 4722 10854 4724 10906
rect 4904 10854 4906 10906
rect 4660 10852 4666 10854
rect 4722 10852 4746 10854
rect 4802 10852 4826 10854
rect 4882 10852 4906 10854
rect 4962 10852 4968 10854
rect 4660 10832 4968 10852
rect 7116 10810 7144 11200
rect 7760 10908 8068 10928
rect 7760 10906 7766 10908
rect 7822 10906 7846 10908
rect 7902 10906 7926 10908
rect 7982 10906 8006 10908
rect 8062 10906 8068 10908
rect 7822 10854 7824 10906
rect 8004 10854 8006 10906
rect 7760 10852 7766 10854
rect 7822 10852 7846 10854
rect 7902 10852 7926 10854
rect 7982 10852 8006 10854
rect 8062 10852 8068 10854
rect 7760 10832 8068 10852
rect 9968 10810 9996 11200
rect 10860 10908 11168 10928
rect 10860 10906 10866 10908
rect 10922 10906 10946 10908
rect 11002 10906 11026 10908
rect 11082 10906 11106 10908
rect 11162 10906 11168 10908
rect 10922 10854 10924 10906
rect 11104 10854 11106 10906
rect 10860 10852 10866 10854
rect 10922 10852 10946 10854
rect 11002 10852 11026 10854
rect 11082 10852 11106 10854
rect 11162 10852 11168 10854
rect 10860 10832 11168 10852
rect 7104 10804 7156 10810
rect 7104 10746 7156 10752
rect 9956 10804 10008 10810
rect 9956 10746 10008 10752
rect 6736 10668 6788 10674
rect 6736 10610 6788 10616
rect 7012 10668 7064 10674
rect 7012 10610 7064 10616
rect 9220 10668 9272 10674
rect 9220 10610 9272 10616
rect 10416 10668 10468 10674
rect 10416 10610 10468 10616
rect 12164 10668 12216 10674
rect 12164 10610 12216 10616
rect 6000 10600 6052 10606
rect 6000 10542 6052 10548
rect 4344 10464 4396 10470
rect 4344 10406 4396 10412
rect 4436 10464 4488 10470
rect 4436 10406 4488 10412
rect 5816 10464 5868 10470
rect 5816 10406 5868 10412
rect 4252 10192 4304 10198
rect 4252 10134 4304 10140
rect 4356 10130 4384 10406
rect 4344 10124 4396 10130
rect 4344 10066 4396 10072
rect 4068 10056 4120 10062
rect 4068 9998 4120 10004
rect 4080 9178 4108 9998
rect 4448 9994 4476 10406
rect 4436 9988 4488 9994
rect 4436 9930 4488 9936
rect 4988 9920 5040 9926
rect 4988 9862 5040 9868
rect 4660 9820 4968 9840
rect 4660 9818 4666 9820
rect 4722 9818 4746 9820
rect 4802 9818 4826 9820
rect 4882 9818 4906 9820
rect 4962 9818 4968 9820
rect 4722 9766 4724 9818
rect 4904 9766 4906 9818
rect 4660 9764 4666 9766
rect 4722 9764 4746 9766
rect 4802 9764 4826 9766
rect 4882 9764 4906 9766
rect 4962 9764 4968 9766
rect 4660 9744 4968 9764
rect 4344 9716 4396 9722
rect 4344 9658 4396 9664
rect 4068 9172 4120 9178
rect 4068 9114 4120 9120
rect 4252 8832 4304 8838
rect 4252 8774 4304 8780
rect 4264 8634 4292 8774
rect 4252 8628 4304 8634
rect 4252 8570 4304 8576
rect 4264 7886 4292 8570
rect 4356 8498 4384 9658
rect 4620 9580 4672 9586
rect 4620 9522 4672 9528
rect 4632 9178 4660 9522
rect 5000 9382 5028 9862
rect 5828 9722 5856 10406
rect 6012 10266 6040 10542
rect 6210 10364 6518 10384
rect 6210 10362 6216 10364
rect 6272 10362 6296 10364
rect 6352 10362 6376 10364
rect 6432 10362 6456 10364
rect 6512 10362 6518 10364
rect 6272 10310 6274 10362
rect 6454 10310 6456 10362
rect 6210 10308 6216 10310
rect 6272 10308 6296 10310
rect 6352 10308 6376 10310
rect 6432 10308 6456 10310
rect 6512 10308 6518 10310
rect 6210 10288 6518 10308
rect 6000 10260 6052 10266
rect 6000 10202 6052 10208
rect 5908 9920 5960 9926
rect 5908 9862 5960 9868
rect 5816 9716 5868 9722
rect 5816 9658 5868 9664
rect 5632 9648 5684 9654
rect 5632 9590 5684 9596
rect 5448 9512 5500 9518
rect 5500 9460 5580 9466
rect 5448 9454 5580 9460
rect 5460 9438 5580 9454
rect 4988 9376 5040 9382
rect 4988 9318 5040 9324
rect 4620 9172 4672 9178
rect 4620 9114 4672 9120
rect 5000 9042 5028 9318
rect 5552 9042 5580 9438
rect 4988 9036 5040 9042
rect 4988 8978 5040 8984
rect 5540 9036 5592 9042
rect 5540 8978 5592 8984
rect 4660 8732 4968 8752
rect 4660 8730 4666 8732
rect 4722 8730 4746 8732
rect 4802 8730 4826 8732
rect 4882 8730 4906 8732
rect 4962 8730 4968 8732
rect 4722 8678 4724 8730
rect 4904 8678 4906 8730
rect 4660 8676 4666 8678
rect 4722 8676 4746 8678
rect 4802 8676 4826 8678
rect 4882 8676 4906 8678
rect 4962 8676 4968 8678
rect 4660 8656 4968 8676
rect 5000 8498 5028 8978
rect 5448 8900 5500 8906
rect 5448 8842 5500 8848
rect 5460 8566 5488 8842
rect 5448 8560 5500 8566
rect 5448 8502 5500 8508
rect 5540 8526 5592 8532
rect 4344 8492 4396 8498
rect 4344 8434 4396 8440
rect 4528 8492 4580 8498
rect 4528 8434 4580 8440
rect 4988 8492 5040 8498
rect 5540 8468 5592 8474
rect 4988 8434 5040 8440
rect 4540 8090 4568 8434
rect 4620 8288 4672 8294
rect 4620 8230 4672 8236
rect 4632 8090 4660 8230
rect 5552 8090 5580 8468
rect 5644 8294 5672 9590
rect 5920 9586 5948 9862
rect 6748 9722 6776 10610
rect 7024 10266 7052 10610
rect 7656 10600 7708 10606
rect 7656 10542 7708 10548
rect 7472 10464 7524 10470
rect 7472 10406 7524 10412
rect 7012 10260 7064 10266
rect 7012 10202 7064 10208
rect 7484 10062 7512 10406
rect 7472 10056 7524 10062
rect 7472 9998 7524 10004
rect 6736 9716 6788 9722
rect 6736 9658 6788 9664
rect 5908 9580 5960 9586
rect 5908 9522 5960 9528
rect 6828 9512 6880 9518
rect 6828 9454 6880 9460
rect 5908 9376 5960 9382
rect 5908 9318 5960 9324
rect 5920 8974 5948 9318
rect 6210 9276 6518 9296
rect 6210 9274 6216 9276
rect 6272 9274 6296 9276
rect 6352 9274 6376 9276
rect 6432 9274 6456 9276
rect 6512 9274 6518 9276
rect 6272 9222 6274 9274
rect 6454 9222 6456 9274
rect 6210 9220 6216 9222
rect 6272 9220 6296 9222
rect 6352 9220 6376 9222
rect 6432 9220 6456 9222
rect 6512 9220 6518 9222
rect 6210 9200 6518 9220
rect 6840 9042 6868 9454
rect 6092 9036 6144 9042
rect 6092 8978 6144 8984
rect 6184 9036 6236 9042
rect 6184 8978 6236 8984
rect 6828 9036 6880 9042
rect 6828 8978 6880 8984
rect 5908 8968 5960 8974
rect 5908 8910 5960 8916
rect 6000 8968 6052 8974
rect 6000 8910 6052 8916
rect 5908 8492 5960 8498
rect 5908 8434 5960 8440
rect 5632 8288 5684 8294
rect 5632 8230 5684 8236
rect 4528 8084 4580 8090
rect 4528 8026 4580 8032
rect 4620 8084 4672 8090
rect 4620 8026 4672 8032
rect 5540 8084 5592 8090
rect 5540 8026 5592 8032
rect 4068 7880 4120 7886
rect 4068 7822 4120 7828
rect 4252 7880 4304 7886
rect 4252 7822 4304 7828
rect 3884 7744 3936 7750
rect 3884 7686 3936 7692
rect 3896 7478 3924 7686
rect 3884 7472 3936 7478
rect 3884 7414 3936 7420
rect 4080 7274 4108 7822
rect 4068 7268 4120 7274
rect 4068 7210 4120 7216
rect 4264 7206 4292 7822
rect 4660 7644 4968 7664
rect 4660 7642 4666 7644
rect 4722 7642 4746 7644
rect 4802 7642 4826 7644
rect 4882 7642 4906 7644
rect 4962 7642 4968 7644
rect 4722 7590 4724 7642
rect 4904 7590 4906 7642
rect 4660 7588 4666 7590
rect 4722 7588 4746 7590
rect 4802 7588 4826 7590
rect 4882 7588 4906 7590
rect 4962 7588 4968 7590
rect 4660 7568 4968 7588
rect 5264 7404 5316 7410
rect 5264 7346 5316 7352
rect 5080 7336 5132 7342
rect 5080 7278 5132 7284
rect 4252 7200 4304 7206
rect 4252 7142 4304 7148
rect 4068 6792 4120 6798
rect 4068 6734 4120 6740
rect 4080 5778 4108 6734
rect 4344 6724 4396 6730
rect 4344 6666 4396 6672
rect 4436 6724 4488 6730
rect 4436 6666 4488 6672
rect 4356 6458 4384 6666
rect 4344 6452 4396 6458
rect 4344 6394 4396 6400
rect 4448 6186 4476 6666
rect 4660 6556 4968 6576
rect 4660 6554 4666 6556
rect 4722 6554 4746 6556
rect 4802 6554 4826 6556
rect 4882 6554 4906 6556
rect 4962 6554 4968 6556
rect 4722 6502 4724 6554
rect 4904 6502 4906 6554
rect 4660 6500 4666 6502
rect 4722 6500 4746 6502
rect 4802 6500 4826 6502
rect 4882 6500 4906 6502
rect 4962 6500 4968 6502
rect 4660 6480 4968 6500
rect 5092 6322 5120 7278
rect 5276 7274 5304 7346
rect 5264 7268 5316 7274
rect 5264 7210 5316 7216
rect 5644 7002 5672 8230
rect 5724 7948 5776 7954
rect 5724 7890 5776 7896
rect 5736 7410 5764 7890
rect 5816 7812 5868 7818
rect 5816 7754 5868 7760
rect 5828 7546 5856 7754
rect 5920 7750 5948 8434
rect 6012 8362 6040 8910
rect 6000 8356 6052 8362
rect 6000 8298 6052 8304
rect 5908 7744 5960 7750
rect 5908 7686 5960 7692
rect 5816 7540 5868 7546
rect 5816 7482 5868 7488
rect 5908 7540 5960 7546
rect 5908 7482 5960 7488
rect 5920 7410 5948 7482
rect 5724 7404 5776 7410
rect 5724 7346 5776 7352
rect 5908 7404 5960 7410
rect 5908 7346 5960 7352
rect 5632 6996 5684 7002
rect 5632 6938 5684 6944
rect 5080 6316 5132 6322
rect 5644 6304 5672 6938
rect 5920 6934 5948 7346
rect 5908 6928 5960 6934
rect 5828 6876 5908 6882
rect 5828 6870 5960 6876
rect 5828 6854 5948 6870
rect 5724 6316 5776 6322
rect 5644 6276 5724 6304
rect 5080 6258 5132 6264
rect 5724 6258 5776 6264
rect 5828 6254 5856 6854
rect 5908 6656 5960 6662
rect 5908 6598 5960 6604
rect 5920 6322 5948 6598
rect 5908 6316 5960 6322
rect 5908 6258 5960 6264
rect 5816 6248 5868 6254
rect 5816 6190 5868 6196
rect 4436 6180 4488 6186
rect 4436 6122 4488 6128
rect 6012 5778 6040 8298
rect 6104 7546 6132 8978
rect 6196 8838 6224 8978
rect 6840 8838 6868 8978
rect 6920 8900 6972 8906
rect 6920 8842 6972 8848
rect 6184 8832 6236 8838
rect 6184 8774 6236 8780
rect 6368 8832 6420 8838
rect 6368 8774 6420 8780
rect 6828 8832 6880 8838
rect 6828 8774 6880 8780
rect 6380 8498 6408 8774
rect 6368 8492 6420 8498
rect 6368 8434 6420 8440
rect 6210 8188 6518 8208
rect 6210 8186 6216 8188
rect 6272 8186 6296 8188
rect 6352 8186 6376 8188
rect 6432 8186 6456 8188
rect 6512 8186 6518 8188
rect 6272 8134 6274 8186
rect 6454 8134 6456 8186
rect 6210 8132 6216 8134
rect 6272 8132 6296 8134
rect 6352 8132 6376 8134
rect 6432 8132 6456 8134
rect 6512 8132 6518 8134
rect 6210 8112 6518 8132
rect 6840 8022 6868 8774
rect 6932 8090 6960 8842
rect 6920 8084 6972 8090
rect 6920 8026 6972 8032
rect 6828 8016 6880 8022
rect 6828 7958 6880 7964
rect 6184 7812 6236 7818
rect 6184 7754 6236 7760
rect 6552 7812 6604 7818
rect 6552 7754 6604 7760
rect 6092 7540 6144 7546
rect 6092 7482 6144 7488
rect 6196 7478 6224 7754
rect 6184 7472 6236 7478
rect 6184 7414 6236 7420
rect 6092 7336 6144 7342
rect 6092 7278 6144 7284
rect 6104 6866 6132 7278
rect 6210 7100 6518 7120
rect 6210 7098 6216 7100
rect 6272 7098 6296 7100
rect 6352 7098 6376 7100
rect 6432 7098 6456 7100
rect 6512 7098 6518 7100
rect 6272 7046 6274 7098
rect 6454 7046 6456 7098
rect 6210 7044 6216 7046
rect 6272 7044 6296 7046
rect 6352 7044 6376 7046
rect 6432 7044 6456 7046
rect 6512 7044 6518 7046
rect 6210 7024 6518 7044
rect 6092 6860 6144 6866
rect 6092 6802 6144 6808
rect 6092 6656 6144 6662
rect 6092 6598 6144 6604
rect 6104 5778 6132 6598
rect 6564 6322 6592 7754
rect 6736 7744 6788 7750
rect 6736 7686 6788 7692
rect 6644 7336 6696 7342
rect 6644 7278 6696 7284
rect 6656 7002 6684 7278
rect 6644 6996 6696 7002
rect 6644 6938 6696 6944
rect 6748 6322 6776 7686
rect 6840 7342 6868 7958
rect 6920 7404 6972 7410
rect 6920 7346 6972 7352
rect 6828 7336 6880 7342
rect 6828 7278 6880 7284
rect 6828 6656 6880 6662
rect 6828 6598 6880 6604
rect 6840 6458 6868 6598
rect 6828 6452 6880 6458
rect 6828 6394 6880 6400
rect 6932 6322 6960 7346
rect 6276 6316 6328 6322
rect 6276 6258 6328 6264
rect 6552 6316 6604 6322
rect 6552 6258 6604 6264
rect 6736 6316 6788 6322
rect 6736 6258 6788 6264
rect 6920 6316 6972 6322
rect 6920 6258 6972 6264
rect 6288 6186 6316 6258
rect 6276 6180 6328 6186
rect 6276 6122 6328 6128
rect 6748 6118 6776 6258
rect 6736 6112 6788 6118
rect 6736 6054 6788 6060
rect 6210 6012 6518 6032
rect 6210 6010 6216 6012
rect 6272 6010 6296 6012
rect 6352 6010 6376 6012
rect 6432 6010 6456 6012
rect 6512 6010 6518 6012
rect 6272 5958 6274 6010
rect 6454 5958 6456 6010
rect 6210 5956 6216 5958
rect 6272 5956 6296 5958
rect 6352 5956 6376 5958
rect 6432 5956 6456 5958
rect 6512 5956 6518 5958
rect 6210 5936 6518 5956
rect 6932 5914 6960 6258
rect 7472 6248 7524 6254
rect 7472 6190 7524 6196
rect 6920 5908 6972 5914
rect 6920 5850 6972 5856
rect 4068 5772 4120 5778
rect 4068 5714 4120 5720
rect 6000 5772 6052 5778
rect 6000 5714 6052 5720
rect 6092 5772 6144 5778
rect 6092 5714 6144 5720
rect 3792 5636 3844 5642
rect 3792 5578 3844 5584
rect 2412 5568 2464 5574
rect 2412 5510 2464 5516
rect 2320 4616 2372 4622
rect 2320 4558 2372 4564
rect 2332 3602 2360 4558
rect 2424 4486 2452 5510
rect 4660 5468 4968 5488
rect 4660 5466 4666 5468
rect 4722 5466 4746 5468
rect 4802 5466 4826 5468
rect 4882 5466 4906 5468
rect 4962 5466 4968 5468
rect 4722 5414 4724 5466
rect 4904 5414 4906 5466
rect 4660 5412 4666 5414
rect 4722 5412 4746 5414
rect 4802 5412 4826 5414
rect 4882 5412 4906 5414
rect 4962 5412 4968 5414
rect 4660 5392 4968 5412
rect 6932 5234 6960 5850
rect 7484 5302 7512 6190
rect 7472 5296 7524 5302
rect 7470 5264 7472 5273
rect 7524 5264 7526 5273
rect 5080 5228 5132 5234
rect 5080 5170 5132 5176
rect 6920 5228 6972 5234
rect 7470 5199 7526 5208
rect 6920 5170 6972 5176
rect 3110 4924 3418 4944
rect 3110 4922 3116 4924
rect 3172 4922 3196 4924
rect 3252 4922 3276 4924
rect 3332 4922 3356 4924
rect 3412 4922 3418 4924
rect 3172 4870 3174 4922
rect 3354 4870 3356 4922
rect 3110 4868 3116 4870
rect 3172 4868 3196 4870
rect 3252 4868 3276 4870
rect 3332 4868 3356 4870
rect 3412 4868 3418 4870
rect 3110 4848 3418 4868
rect 5092 4826 5120 5170
rect 6920 5024 6972 5030
rect 6920 4966 6972 4972
rect 6210 4924 6518 4944
rect 6210 4922 6216 4924
rect 6272 4922 6296 4924
rect 6352 4922 6376 4924
rect 6432 4922 6456 4924
rect 6512 4922 6518 4924
rect 6272 4870 6274 4922
rect 6454 4870 6456 4922
rect 6210 4868 6216 4870
rect 6272 4868 6296 4870
rect 6352 4868 6376 4870
rect 6432 4868 6456 4870
rect 6512 4868 6518 4870
rect 6210 4848 6518 4868
rect 5080 4820 5132 4826
rect 5080 4762 5132 4768
rect 3056 4616 3108 4622
rect 3056 4558 3108 4564
rect 4988 4616 5040 4622
rect 4988 4558 5040 4564
rect 2412 4480 2464 4486
rect 2412 4422 2464 4428
rect 756 3596 808 3602
rect 756 3538 808 3544
rect 2320 3596 2372 3602
rect 2320 3538 2372 3544
rect 768 2514 796 3538
rect 2424 3534 2452 4422
rect 3068 4282 3096 4558
rect 4660 4380 4968 4400
rect 4660 4378 4666 4380
rect 4722 4378 4746 4380
rect 4802 4378 4826 4380
rect 4882 4378 4906 4380
rect 4962 4378 4968 4380
rect 4722 4326 4724 4378
rect 4904 4326 4906 4378
rect 4660 4324 4666 4326
rect 4722 4324 4746 4326
rect 4802 4324 4826 4326
rect 4882 4324 4906 4326
rect 4962 4324 4968 4326
rect 4660 4304 4968 4324
rect 3056 4276 3108 4282
rect 3056 4218 3108 4224
rect 5000 4214 5028 4558
rect 4988 4208 5040 4214
rect 4988 4150 5040 4156
rect 5092 4146 5120 4762
rect 5172 4480 5224 4486
rect 5172 4422 5224 4428
rect 5632 4480 5684 4486
rect 5632 4422 5684 4428
rect 5184 4146 5212 4422
rect 5448 4208 5500 4214
rect 5448 4150 5500 4156
rect 5080 4140 5132 4146
rect 5080 4082 5132 4088
rect 5172 4140 5224 4146
rect 5172 4082 5224 4088
rect 3976 4004 4028 4010
rect 3976 3946 4028 3952
rect 4528 4004 4580 4010
rect 4528 3946 4580 3952
rect 3516 3936 3568 3942
rect 3516 3878 3568 3884
rect 3110 3836 3418 3856
rect 3110 3834 3116 3836
rect 3172 3834 3196 3836
rect 3252 3834 3276 3836
rect 3332 3834 3356 3836
rect 3412 3834 3418 3836
rect 3172 3782 3174 3834
rect 3354 3782 3356 3834
rect 3110 3780 3116 3782
rect 3172 3780 3196 3782
rect 3252 3780 3276 3782
rect 3332 3780 3356 3782
rect 3412 3780 3418 3782
rect 3110 3760 3418 3780
rect 2412 3528 2464 3534
rect 2412 3470 2464 3476
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 756 2508 808 2514
rect 756 2450 808 2456
rect 768 1426 796 2450
rect 2424 2378 2452 3470
rect 2884 3126 2912 3470
rect 3528 3194 3556 3878
rect 3884 3664 3936 3670
rect 3988 3652 4016 3946
rect 3936 3624 4016 3652
rect 3884 3606 3936 3612
rect 3608 3528 3660 3534
rect 3884 3528 3936 3534
rect 3608 3470 3660 3476
rect 3882 3496 3884 3505
rect 3936 3496 3938 3505
rect 3620 3194 3648 3470
rect 3988 3466 4016 3624
rect 4068 3664 4120 3670
rect 4068 3606 4120 3612
rect 4080 3505 4108 3606
rect 4540 3534 4568 3946
rect 5092 3534 5120 4082
rect 5356 3732 5408 3738
rect 5356 3674 5408 3680
rect 5368 3534 5396 3674
rect 4160 3528 4212 3534
rect 4066 3496 4122 3505
rect 3882 3431 3938 3440
rect 3976 3460 4028 3466
rect 4160 3470 4212 3476
rect 4344 3528 4396 3534
rect 4528 3528 4580 3534
rect 4344 3470 4396 3476
rect 4448 3488 4528 3516
rect 4066 3431 4122 3440
rect 3976 3402 4028 3408
rect 3884 3392 3936 3398
rect 3884 3334 3936 3340
rect 3516 3188 3568 3194
rect 3516 3130 3568 3136
rect 3608 3188 3660 3194
rect 3608 3130 3660 3136
rect 2872 3120 2924 3126
rect 2872 3062 2924 3068
rect 3896 3058 3924 3334
rect 4172 3058 4200 3470
rect 3884 3052 3936 3058
rect 3884 2994 3936 3000
rect 4160 3052 4212 3058
rect 4160 2994 4212 3000
rect 4356 2990 4384 3470
rect 4448 3194 4476 3488
rect 4528 3470 4580 3476
rect 5080 3528 5132 3534
rect 5080 3470 5132 3476
rect 5356 3528 5408 3534
rect 5356 3470 5408 3476
rect 5460 3466 5488 4150
rect 5540 3936 5592 3942
rect 5540 3878 5592 3884
rect 5448 3460 5500 3466
rect 5448 3402 5500 3408
rect 4660 3292 4968 3312
rect 4660 3290 4666 3292
rect 4722 3290 4746 3292
rect 4802 3290 4826 3292
rect 4882 3290 4906 3292
rect 4962 3290 4968 3292
rect 4722 3238 4724 3290
rect 4904 3238 4906 3290
rect 4660 3236 4666 3238
rect 4722 3236 4746 3238
rect 4802 3236 4826 3238
rect 4882 3236 4906 3238
rect 4962 3236 4968 3238
rect 4660 3216 4968 3236
rect 4436 3188 4488 3194
rect 4436 3130 4488 3136
rect 4802 3088 4858 3097
rect 4528 3052 4580 3058
rect 5552 3058 5580 3878
rect 5644 3738 5672 4422
rect 6932 4146 6960 4966
rect 7668 4622 7696 10542
rect 9036 10464 9088 10470
rect 9036 10406 9088 10412
rect 9048 10130 9076 10406
rect 9232 10266 9260 10610
rect 9680 10532 9732 10538
rect 9680 10474 9732 10480
rect 9310 10364 9618 10384
rect 9310 10362 9316 10364
rect 9372 10362 9396 10364
rect 9452 10362 9476 10364
rect 9532 10362 9556 10364
rect 9612 10362 9618 10364
rect 9372 10310 9374 10362
rect 9554 10310 9556 10362
rect 9310 10308 9316 10310
rect 9372 10308 9396 10310
rect 9452 10308 9476 10310
rect 9532 10308 9556 10310
rect 9612 10308 9618 10310
rect 9310 10288 9618 10308
rect 9220 10260 9272 10266
rect 9220 10202 9272 10208
rect 9036 10124 9088 10130
rect 9036 10066 9088 10072
rect 8944 10056 8996 10062
rect 8944 9998 8996 10004
rect 9128 10056 9180 10062
rect 9128 9998 9180 10004
rect 8300 9920 8352 9926
rect 8300 9862 8352 9868
rect 7760 9820 8068 9840
rect 7760 9818 7766 9820
rect 7822 9818 7846 9820
rect 7902 9818 7926 9820
rect 7982 9818 8006 9820
rect 8062 9818 8068 9820
rect 7822 9766 7824 9818
rect 8004 9766 8006 9818
rect 7760 9764 7766 9766
rect 7822 9764 7846 9766
rect 7902 9764 7926 9766
rect 7982 9764 8006 9766
rect 8062 9764 8068 9766
rect 7760 9744 8068 9764
rect 8312 9654 8340 9862
rect 8300 9648 8352 9654
rect 8300 9590 8352 9596
rect 8116 8968 8168 8974
rect 8116 8910 8168 8916
rect 7760 8732 8068 8752
rect 7760 8730 7766 8732
rect 7822 8730 7846 8732
rect 7902 8730 7926 8732
rect 7982 8730 8006 8732
rect 8062 8730 8068 8732
rect 7822 8678 7824 8730
rect 8004 8678 8006 8730
rect 7760 8676 7766 8678
rect 7822 8676 7846 8678
rect 7902 8676 7926 8678
rect 7982 8676 8006 8678
rect 8062 8676 8068 8678
rect 7760 8656 8068 8676
rect 8024 8288 8076 8294
rect 8024 8230 8076 8236
rect 8036 7886 8064 8230
rect 8024 7880 8076 7886
rect 8024 7822 8076 7828
rect 7760 7644 8068 7664
rect 7760 7642 7766 7644
rect 7822 7642 7846 7644
rect 7902 7642 7926 7644
rect 7982 7642 8006 7644
rect 8062 7642 8068 7644
rect 7822 7590 7824 7642
rect 8004 7590 8006 7642
rect 7760 7588 7766 7590
rect 7822 7588 7846 7590
rect 7902 7588 7926 7590
rect 7982 7588 8006 7590
rect 8062 7588 8068 7590
rect 7760 7568 8068 7588
rect 8128 7426 8156 8910
rect 8312 8566 8340 9590
rect 8300 8560 8352 8566
rect 8300 8502 8352 8508
rect 8036 7398 8156 7426
rect 8036 6866 8064 7398
rect 8116 7336 8168 7342
rect 8168 7296 8248 7324
rect 8116 7278 8168 7284
rect 8024 6860 8076 6866
rect 8024 6802 8076 6808
rect 7760 6556 8068 6576
rect 7760 6554 7766 6556
rect 7822 6554 7846 6556
rect 7902 6554 7926 6556
rect 7982 6554 8006 6556
rect 8062 6554 8068 6556
rect 7822 6502 7824 6554
rect 8004 6502 8006 6554
rect 7760 6500 7766 6502
rect 7822 6500 7846 6502
rect 7902 6500 7926 6502
rect 7982 6500 8006 6502
rect 8062 6500 8068 6502
rect 7760 6480 8068 6500
rect 8220 5914 8248 7296
rect 8208 5908 8260 5914
rect 8208 5850 8260 5856
rect 7760 5468 8068 5488
rect 7760 5466 7766 5468
rect 7822 5466 7846 5468
rect 7902 5466 7926 5468
rect 7982 5466 8006 5468
rect 8062 5466 8068 5468
rect 7822 5414 7824 5466
rect 8004 5414 8006 5466
rect 7760 5412 7766 5414
rect 7822 5412 7846 5414
rect 7902 5412 7926 5414
rect 7982 5412 8006 5414
rect 8062 5412 8068 5414
rect 7760 5392 8068 5412
rect 8220 5302 8248 5850
rect 8312 5574 8340 8502
rect 8956 8090 8984 9998
rect 8944 8084 8996 8090
rect 8944 8026 8996 8032
rect 8956 7410 8984 8026
rect 9140 7970 9168 9998
rect 9310 9276 9618 9296
rect 9310 9274 9316 9276
rect 9372 9274 9396 9276
rect 9452 9274 9476 9276
rect 9532 9274 9556 9276
rect 9612 9274 9618 9276
rect 9372 9222 9374 9274
rect 9554 9222 9556 9274
rect 9310 9220 9316 9222
rect 9372 9220 9396 9222
rect 9452 9220 9476 9222
rect 9532 9220 9556 9222
rect 9612 9220 9618 9222
rect 9310 9200 9618 9220
rect 9692 9042 9720 10474
rect 9956 10464 10008 10470
rect 9956 10406 10008 10412
rect 9968 9654 9996 10406
rect 9956 9648 10008 9654
rect 9956 9590 10008 9596
rect 10232 9376 10284 9382
rect 10232 9318 10284 9324
rect 10244 9042 10272 9318
rect 10428 9178 10456 10610
rect 10784 10464 10836 10470
rect 10784 10406 10836 10412
rect 12072 10464 12124 10470
rect 12072 10406 12124 10412
rect 10600 9376 10652 9382
rect 10600 9318 10652 9324
rect 10416 9172 10468 9178
rect 10416 9114 10468 9120
rect 9680 9036 9732 9042
rect 9680 8978 9732 8984
rect 10232 9036 10284 9042
rect 10416 9036 10468 9042
rect 10232 8978 10284 8984
rect 10336 8996 10416 9024
rect 10232 8900 10284 8906
rect 10232 8842 10284 8848
rect 9864 8832 9916 8838
rect 9864 8774 9916 8780
rect 9876 8537 9904 8774
rect 9862 8528 9918 8537
rect 9862 8463 9918 8472
rect 9864 8288 9916 8294
rect 9864 8230 9916 8236
rect 9310 8188 9618 8208
rect 9310 8186 9316 8188
rect 9372 8186 9396 8188
rect 9452 8186 9476 8188
rect 9532 8186 9556 8188
rect 9612 8186 9618 8188
rect 9372 8134 9374 8186
rect 9554 8134 9556 8186
rect 9310 8132 9316 8134
rect 9372 8132 9396 8134
rect 9452 8132 9476 8134
rect 9532 8132 9556 8134
rect 9612 8132 9618 8134
rect 9310 8112 9618 8132
rect 9772 8016 9824 8022
rect 9048 7942 9168 7970
rect 9770 7984 9772 7993
rect 9824 7984 9826 7993
rect 9048 7818 9076 7942
rect 9876 7954 9904 8230
rect 10140 8084 10192 8090
rect 10140 8026 10192 8032
rect 9770 7919 9826 7928
rect 9864 7948 9916 7954
rect 9588 7880 9640 7886
rect 9588 7822 9640 7828
rect 9036 7812 9088 7818
rect 9036 7754 9088 7760
rect 9048 7410 9076 7754
rect 9600 7546 9628 7822
rect 9588 7540 9640 7546
rect 9588 7482 9640 7488
rect 8944 7404 8996 7410
rect 8944 7346 8996 7352
rect 9036 7404 9088 7410
rect 9036 7346 9088 7352
rect 9220 7404 9272 7410
rect 9220 7346 9272 7352
rect 8392 7268 8444 7274
rect 8392 7210 8444 7216
rect 8404 6798 8432 7210
rect 8668 6860 8720 6866
rect 8668 6802 8720 6808
rect 8392 6792 8444 6798
rect 8392 6734 8444 6740
rect 8576 6792 8628 6798
rect 8576 6734 8628 6740
rect 8588 6338 8616 6734
rect 8680 6390 8708 6802
rect 9048 6458 9076 7346
rect 9232 6798 9260 7346
rect 9784 7274 9812 7919
rect 9864 7890 9916 7896
rect 10152 7818 10180 8026
rect 10244 7954 10272 8842
rect 10232 7948 10284 7954
rect 10232 7890 10284 7896
rect 10140 7812 10192 7818
rect 10140 7754 10192 7760
rect 10152 7313 10180 7754
rect 10138 7304 10194 7313
rect 9772 7268 9824 7274
rect 10138 7239 10194 7248
rect 9772 7210 9824 7216
rect 9310 7100 9618 7120
rect 9310 7098 9316 7100
rect 9372 7098 9396 7100
rect 9452 7098 9476 7100
rect 9532 7098 9556 7100
rect 9612 7098 9618 7100
rect 9372 7046 9374 7098
rect 9554 7046 9556 7098
rect 9310 7044 9316 7046
rect 9372 7044 9396 7046
rect 9452 7044 9476 7046
rect 9532 7044 9556 7046
rect 9612 7044 9618 7046
rect 9310 7024 9618 7044
rect 10138 7032 10194 7041
rect 10138 6967 10140 6976
rect 10192 6967 10194 6976
rect 10140 6938 10192 6944
rect 10336 6882 10364 8996
rect 10416 8978 10468 8984
rect 10506 8392 10562 8401
rect 10506 8327 10562 8336
rect 10520 8090 10548 8327
rect 10508 8084 10560 8090
rect 10508 8026 10560 8032
rect 10508 7880 10560 7886
rect 10414 7848 10470 7857
rect 10508 7822 10560 7828
rect 10414 7783 10470 7792
rect 10428 7546 10456 7783
rect 10416 7540 10468 7546
rect 10416 7482 10468 7488
rect 10416 7404 10468 7410
rect 10416 7346 10468 7352
rect 10428 7206 10456 7346
rect 10416 7200 10468 7206
rect 10416 7142 10468 7148
rect 10428 7002 10456 7142
rect 10416 6996 10468 7002
rect 10416 6938 10468 6944
rect 10520 6934 10548 7822
rect 9772 6860 9824 6866
rect 9772 6802 9824 6808
rect 9876 6854 10364 6882
rect 10508 6928 10560 6934
rect 10508 6870 10560 6876
rect 9220 6792 9272 6798
rect 9220 6734 9272 6740
rect 9588 6656 9640 6662
rect 9588 6598 9640 6604
rect 9036 6452 9088 6458
rect 9036 6394 9088 6400
rect 9600 6390 9628 6598
rect 8392 6316 8444 6322
rect 8392 6258 8444 6264
rect 8496 6310 8616 6338
rect 8668 6384 8720 6390
rect 8668 6326 8720 6332
rect 9588 6384 9640 6390
rect 9588 6326 9640 6332
rect 8300 5568 8352 5574
rect 8300 5510 8352 5516
rect 8208 5296 8260 5302
rect 7852 5244 8208 5250
rect 7852 5238 8260 5244
rect 7852 5234 8248 5238
rect 7840 5228 8248 5234
rect 7892 5222 8248 5228
rect 7840 5170 7892 5176
rect 8312 4842 8340 5510
rect 8404 5166 8432 6258
rect 8392 5160 8444 5166
rect 8392 5102 8444 5108
rect 8496 5098 8524 6310
rect 9784 6254 9812 6802
rect 9876 6798 9904 6854
rect 10336 6798 10364 6854
rect 9864 6792 9916 6798
rect 10232 6792 10284 6798
rect 9864 6734 9916 6740
rect 9954 6760 10010 6769
rect 10232 6734 10284 6740
rect 10324 6792 10376 6798
rect 10324 6734 10376 6740
rect 9954 6695 10010 6704
rect 9968 6322 9996 6695
rect 10244 6322 10272 6734
rect 9956 6316 10008 6322
rect 9956 6258 10008 6264
rect 10232 6316 10284 6322
rect 10232 6258 10284 6264
rect 9772 6248 9824 6254
rect 9772 6190 9824 6196
rect 9310 6012 9618 6032
rect 9310 6010 9316 6012
rect 9372 6010 9396 6012
rect 9452 6010 9476 6012
rect 9532 6010 9556 6012
rect 9612 6010 9618 6012
rect 9372 5958 9374 6010
rect 9554 5958 9556 6010
rect 9310 5956 9316 5958
rect 9372 5956 9396 5958
rect 9452 5956 9476 5958
rect 9532 5956 9556 5958
rect 9612 5956 9618 5958
rect 9310 5936 9618 5956
rect 9968 5914 9996 6258
rect 10520 6254 10548 6870
rect 10508 6248 10560 6254
rect 10508 6190 10560 6196
rect 9956 5908 10008 5914
rect 9956 5850 10008 5856
rect 8852 5568 8904 5574
rect 8772 5516 8852 5534
rect 8904 5516 9168 5534
rect 8772 5506 9168 5516
rect 8484 5092 8536 5098
rect 8484 5034 8536 5040
rect 8312 4814 8524 4842
rect 7656 4616 7708 4622
rect 7656 4558 7708 4564
rect 8208 4616 8260 4622
rect 8208 4558 8260 4564
rect 7380 4548 7432 4554
rect 7380 4490 7432 4496
rect 6920 4140 6972 4146
rect 6920 4082 6972 4088
rect 6552 4072 6604 4078
rect 6552 4014 6604 4020
rect 6644 4072 6696 4078
rect 6644 4014 6696 4020
rect 7104 4072 7156 4078
rect 7104 4014 7156 4020
rect 5908 4004 5960 4010
rect 5908 3946 5960 3952
rect 5632 3732 5684 3738
rect 5632 3674 5684 3680
rect 5920 3534 5948 3946
rect 6210 3836 6518 3856
rect 6210 3834 6216 3836
rect 6272 3834 6296 3836
rect 6352 3834 6376 3836
rect 6432 3834 6456 3836
rect 6512 3834 6518 3836
rect 6272 3782 6274 3834
rect 6454 3782 6456 3834
rect 6210 3780 6216 3782
rect 6272 3780 6296 3782
rect 6352 3780 6376 3782
rect 6432 3780 6456 3782
rect 6512 3780 6518 3782
rect 6210 3760 6518 3780
rect 6368 3664 6420 3670
rect 6368 3606 6420 3612
rect 5908 3528 5960 3534
rect 5908 3470 5960 3476
rect 5632 3392 5684 3398
rect 5632 3334 5684 3340
rect 4802 3023 4804 3032
rect 4528 2994 4580 3000
rect 4856 3023 4858 3032
rect 5540 3052 5592 3058
rect 4804 2994 4856 3000
rect 5540 2994 5592 3000
rect 4344 2984 4396 2990
rect 4344 2926 4396 2932
rect 4436 2916 4488 2922
rect 4436 2858 4488 2864
rect 3110 2748 3418 2768
rect 3110 2746 3116 2748
rect 3172 2746 3196 2748
rect 3252 2746 3276 2748
rect 3332 2746 3356 2748
rect 3412 2746 3418 2748
rect 3172 2694 3174 2746
rect 3354 2694 3356 2746
rect 3110 2692 3116 2694
rect 3172 2692 3196 2694
rect 3252 2692 3276 2694
rect 3332 2692 3356 2694
rect 3412 2692 3418 2694
rect 3110 2672 3418 2692
rect 3884 2576 3936 2582
rect 3884 2518 3936 2524
rect 3700 2508 3752 2514
rect 3700 2450 3752 2456
rect 2412 2372 2464 2378
rect 2412 2314 2464 2320
rect 2688 2372 2740 2378
rect 2688 2314 2740 2320
rect 3516 2372 3568 2378
rect 3516 2314 3568 2320
rect 756 1420 808 1426
rect 756 1362 808 1368
rect 768 270 796 1362
rect 2700 1290 2728 2314
rect 2964 2304 3016 2310
rect 2964 2246 3016 2252
rect 2976 1290 3004 2246
rect 3528 2106 3556 2314
rect 3608 2304 3660 2310
rect 3608 2246 3660 2252
rect 3516 2100 3568 2106
rect 3516 2042 3568 2048
rect 3620 1970 3648 2246
rect 3712 2106 3740 2450
rect 3700 2100 3752 2106
rect 3700 2042 3752 2048
rect 3608 1964 3660 1970
rect 3608 1906 3660 1912
rect 3110 1660 3418 1680
rect 3110 1658 3116 1660
rect 3172 1658 3196 1660
rect 3252 1658 3276 1660
rect 3332 1658 3356 1660
rect 3412 1658 3418 1660
rect 3172 1606 3174 1658
rect 3354 1606 3356 1658
rect 3110 1604 3116 1606
rect 3172 1604 3196 1606
rect 3252 1604 3276 1606
rect 3332 1604 3356 1606
rect 3412 1604 3418 1606
rect 3110 1584 3418 1604
rect 3896 1562 3924 2518
rect 4448 2446 4476 2858
rect 4436 2440 4488 2446
rect 4436 2382 4488 2388
rect 4068 2304 4120 2310
rect 4068 2246 4120 2252
rect 4344 2304 4396 2310
rect 4344 2246 4396 2252
rect 3884 1556 3936 1562
rect 3884 1498 3936 1504
rect 3896 1358 3924 1498
rect 3884 1352 3936 1358
rect 3884 1294 3936 1300
rect 4080 1306 4108 2246
rect 4356 2106 4384 2246
rect 4344 2100 4396 2106
rect 4344 2042 4396 2048
rect 4448 2038 4476 2382
rect 4436 2032 4488 2038
rect 4436 1974 4488 1980
rect 4540 1902 4568 2994
rect 5644 2990 5672 3334
rect 6380 3126 6408 3606
rect 5816 3120 5868 3126
rect 5816 3062 5868 3068
rect 6368 3120 6420 3126
rect 6368 3062 6420 3068
rect 5632 2984 5684 2990
rect 5632 2926 5684 2932
rect 5644 2582 5672 2926
rect 5632 2576 5684 2582
rect 5632 2518 5684 2524
rect 5264 2508 5316 2514
rect 5264 2450 5316 2456
rect 5276 2378 5304 2450
rect 5264 2372 5316 2378
rect 5264 2314 5316 2320
rect 4660 2204 4968 2224
rect 4660 2202 4666 2204
rect 4722 2202 4746 2204
rect 4802 2202 4826 2204
rect 4882 2202 4906 2204
rect 4962 2202 4968 2204
rect 4722 2150 4724 2202
rect 4904 2150 4906 2202
rect 4660 2148 4666 2150
rect 4722 2148 4746 2150
rect 4802 2148 4826 2150
rect 4882 2148 4906 2150
rect 4962 2148 4968 2150
rect 4660 2128 4968 2148
rect 5276 2038 5304 2314
rect 5264 2032 5316 2038
rect 5264 1974 5316 1980
rect 5172 1964 5224 1970
rect 5172 1906 5224 1912
rect 4528 1896 4580 1902
rect 5184 1850 5212 1906
rect 4528 1838 4580 1844
rect 5092 1822 5212 1850
rect 5092 1358 5120 1822
rect 4160 1352 4212 1358
rect 4080 1300 4160 1306
rect 4080 1294 4212 1300
rect 5080 1352 5132 1358
rect 5080 1294 5132 1300
rect 2688 1284 2740 1290
rect 2688 1226 2740 1232
rect 2964 1284 3016 1290
rect 2964 1226 3016 1232
rect 3424 1284 3476 1290
rect 3424 1226 3476 1232
rect 756 264 808 270
rect 756 206 808 212
rect 2700 134 2728 1226
rect 3436 882 3464 1226
rect 3424 876 3476 882
rect 3424 818 3476 824
rect 3896 864 3924 1294
rect 4080 1278 4200 1294
rect 4080 1018 4108 1278
rect 5092 1222 5120 1294
rect 5276 1222 5304 1974
rect 5540 1896 5592 1902
rect 5540 1838 5592 1844
rect 5552 1562 5580 1838
rect 5644 1834 5672 2518
rect 5724 2508 5776 2514
rect 5724 2450 5776 2456
rect 5632 1828 5684 1834
rect 5632 1770 5684 1776
rect 5540 1556 5592 1562
rect 5540 1498 5592 1504
rect 5736 1494 5764 2450
rect 5828 2446 5856 3062
rect 5908 3052 5960 3058
rect 5908 2994 5960 3000
rect 5816 2440 5868 2446
rect 5816 2382 5868 2388
rect 5920 2106 5948 2994
rect 6210 2748 6518 2768
rect 6210 2746 6216 2748
rect 6272 2746 6296 2748
rect 6352 2746 6376 2748
rect 6432 2746 6456 2748
rect 6512 2746 6518 2748
rect 6272 2694 6274 2746
rect 6454 2694 6456 2746
rect 6210 2692 6216 2694
rect 6272 2692 6296 2694
rect 6352 2692 6376 2694
rect 6432 2692 6456 2694
rect 6512 2692 6518 2694
rect 6210 2672 6518 2692
rect 5908 2100 5960 2106
rect 5908 2042 5960 2048
rect 5724 1488 5776 1494
rect 5724 1430 5776 1436
rect 5920 1426 5948 2042
rect 6000 1760 6052 1766
rect 6000 1702 6052 1708
rect 5908 1420 5960 1426
rect 5908 1362 5960 1368
rect 6012 1358 6040 1702
rect 6210 1660 6518 1680
rect 6210 1658 6216 1660
rect 6272 1658 6296 1660
rect 6352 1658 6376 1660
rect 6432 1658 6456 1660
rect 6512 1658 6518 1660
rect 6272 1606 6274 1658
rect 6454 1606 6456 1658
rect 6210 1604 6216 1606
rect 6272 1604 6296 1606
rect 6352 1604 6376 1606
rect 6432 1604 6456 1606
rect 6512 1604 6518 1606
rect 6210 1584 6518 1604
rect 6564 1358 6592 4014
rect 6656 3670 6684 4014
rect 6828 3936 6880 3942
rect 6828 3878 6880 3884
rect 6840 3738 6868 3878
rect 6828 3732 6880 3738
rect 6828 3674 6880 3680
rect 6644 3664 6696 3670
rect 6644 3606 6696 3612
rect 7116 3602 7144 4014
rect 7104 3596 7156 3602
rect 7104 3538 7156 3544
rect 7288 3528 7340 3534
rect 7288 3470 7340 3476
rect 6644 3392 6696 3398
rect 6644 3334 6696 3340
rect 6736 3392 6788 3398
rect 6736 3334 6788 3340
rect 7104 3392 7156 3398
rect 7104 3334 7156 3340
rect 6656 2854 6684 3334
rect 6748 3097 6776 3334
rect 6734 3088 6790 3097
rect 6734 3023 6790 3032
rect 6644 2848 6696 2854
rect 6644 2790 6696 2796
rect 5356 1352 5408 1358
rect 5356 1294 5408 1300
rect 5540 1352 5592 1358
rect 5540 1294 5592 1300
rect 6000 1352 6052 1358
rect 6000 1294 6052 1300
rect 6552 1352 6604 1358
rect 6552 1294 6604 1300
rect 5080 1216 5132 1222
rect 5080 1158 5132 1164
rect 5264 1216 5316 1222
rect 5264 1158 5316 1164
rect 4660 1116 4968 1136
rect 4660 1114 4666 1116
rect 4722 1114 4746 1116
rect 4802 1114 4826 1116
rect 4882 1114 4906 1116
rect 4962 1114 4968 1116
rect 4722 1062 4724 1114
rect 4904 1062 4906 1114
rect 4660 1060 4666 1062
rect 4722 1060 4746 1062
rect 4802 1060 4826 1062
rect 4882 1060 4906 1062
rect 4962 1060 4968 1062
rect 4660 1040 4968 1060
rect 4068 1012 4120 1018
rect 4068 954 4120 960
rect 3976 876 4028 882
rect 3896 836 3976 864
rect 3896 746 3924 836
rect 3976 818 4028 824
rect 4160 876 4212 882
rect 4160 818 4212 824
rect 3884 740 3936 746
rect 3884 682 3936 688
rect 2964 672 3016 678
rect 2964 614 3016 620
rect 2976 338 3004 614
rect 3110 572 3418 592
rect 3110 570 3116 572
rect 3172 570 3196 572
rect 3252 570 3276 572
rect 3332 570 3356 572
rect 3412 570 3418 572
rect 3172 518 3174 570
rect 3354 518 3356 570
rect 3110 516 3116 518
rect 3172 516 3196 518
rect 3252 516 3276 518
rect 3332 516 3356 518
rect 3412 516 3418 518
rect 3110 496 3418 516
rect 4172 474 4200 818
rect 5276 746 5304 1158
rect 5368 864 5396 1294
rect 5552 1018 5580 1294
rect 6564 1018 6592 1294
rect 6644 1284 6696 1290
rect 6748 1272 6776 3023
rect 7116 2446 7144 3334
rect 7196 3052 7248 3058
rect 7196 2994 7248 3000
rect 7208 2446 7236 2994
rect 7104 2440 7156 2446
rect 7104 2382 7156 2388
rect 7196 2440 7248 2446
rect 7196 2382 7248 2388
rect 7300 2106 7328 3470
rect 7288 2100 7340 2106
rect 7288 2042 7340 2048
rect 7300 1766 7328 2042
rect 7392 1970 7420 4490
rect 7760 4380 8068 4400
rect 7760 4378 7766 4380
rect 7822 4378 7846 4380
rect 7902 4378 7926 4380
rect 7982 4378 8006 4380
rect 8062 4378 8068 4380
rect 7822 4326 7824 4378
rect 8004 4326 8006 4378
rect 7760 4324 7766 4326
rect 7822 4324 7846 4326
rect 7902 4324 7926 4326
rect 7982 4324 8006 4326
rect 8062 4324 8068 4326
rect 7760 4304 8068 4324
rect 8220 4282 8248 4558
rect 8496 4554 8524 4814
rect 8772 4690 8800 5506
rect 9140 5302 9168 5506
rect 10612 5370 10640 9318
rect 10796 8616 10824 10406
rect 11244 9988 11296 9994
rect 11244 9930 11296 9936
rect 10860 9820 11168 9840
rect 10860 9818 10866 9820
rect 10922 9818 10946 9820
rect 11002 9818 11026 9820
rect 11082 9818 11106 9820
rect 11162 9818 11168 9820
rect 10922 9766 10924 9818
rect 11104 9766 11106 9818
rect 10860 9764 10866 9766
rect 10922 9764 10946 9766
rect 11002 9764 11026 9766
rect 11082 9764 11106 9766
rect 11162 9764 11168 9766
rect 10860 9744 11168 9764
rect 10876 9512 10928 9518
rect 10876 9454 10928 9460
rect 10888 9110 10916 9454
rect 10876 9104 10928 9110
rect 10876 9046 10928 9052
rect 11256 8974 11284 9930
rect 11520 9920 11572 9926
rect 11520 9862 11572 9868
rect 11336 9648 11388 9654
rect 11336 9590 11388 9596
rect 11348 9042 11376 9590
rect 11336 9036 11388 9042
rect 11336 8978 11388 8984
rect 11244 8968 11296 8974
rect 11244 8910 11296 8916
rect 10860 8732 11168 8752
rect 10860 8730 10866 8732
rect 10922 8730 10946 8732
rect 11002 8730 11026 8732
rect 11082 8730 11106 8732
rect 11162 8730 11168 8732
rect 10922 8678 10924 8730
rect 11104 8678 11106 8730
rect 10860 8676 10866 8678
rect 10922 8676 10946 8678
rect 11002 8676 11026 8678
rect 11082 8676 11106 8678
rect 11162 8676 11168 8678
rect 10860 8656 11168 8676
rect 10796 8588 11008 8616
rect 10874 8528 10930 8537
rect 10692 8492 10744 8498
rect 10874 8463 10930 8472
rect 10692 8434 10744 8440
rect 10704 8090 10732 8434
rect 10692 8084 10744 8090
rect 10692 8026 10744 8032
rect 10784 8084 10836 8090
rect 10784 8026 10836 8032
rect 10704 6730 10732 8026
rect 10796 7342 10824 8026
rect 10888 7886 10916 8463
rect 10980 7886 11008 8588
rect 11164 8350 11468 8378
rect 11164 7886 11192 8350
rect 11440 8294 11468 8350
rect 11336 8288 11388 8294
rect 11336 8230 11388 8236
rect 11428 8288 11480 8294
rect 11428 8230 11480 8236
rect 11242 7984 11298 7993
rect 11242 7919 11244 7928
rect 11296 7919 11298 7928
rect 11244 7890 11296 7896
rect 10876 7880 10928 7886
rect 10876 7822 10928 7828
rect 10968 7880 11020 7886
rect 10968 7822 11020 7828
rect 11152 7880 11204 7886
rect 11152 7822 11204 7828
rect 10860 7644 11168 7664
rect 10860 7642 10866 7644
rect 10922 7642 10946 7644
rect 11002 7642 11026 7644
rect 11082 7642 11106 7644
rect 11162 7642 11168 7644
rect 10922 7590 10924 7642
rect 11104 7590 11106 7642
rect 10860 7588 10866 7590
rect 10922 7588 10946 7590
rect 11002 7588 11026 7590
rect 11082 7588 11106 7590
rect 11162 7588 11168 7590
rect 10860 7568 11168 7588
rect 11348 7342 11376 8230
rect 11428 8016 11480 8022
rect 11428 7958 11480 7964
rect 11440 7546 11468 7958
rect 11532 7818 11560 9862
rect 12084 9450 12112 10406
rect 12176 9586 12204 10610
rect 12256 10532 12308 10538
rect 12256 10474 12308 10480
rect 12164 9580 12216 9586
rect 12164 9522 12216 9528
rect 11980 9444 12032 9450
rect 11980 9386 12032 9392
rect 12072 9444 12124 9450
rect 12072 9386 12124 9392
rect 11992 9042 12020 9386
rect 12176 9178 12204 9522
rect 12164 9172 12216 9178
rect 12164 9114 12216 9120
rect 11980 9036 12032 9042
rect 11980 8978 12032 8984
rect 12164 9036 12216 9042
rect 12164 8978 12216 8984
rect 11796 7880 11848 7886
rect 11794 7848 11796 7857
rect 11848 7848 11850 7857
rect 11520 7812 11572 7818
rect 11520 7754 11572 7760
rect 11704 7812 11756 7818
rect 11794 7783 11850 7792
rect 11888 7812 11940 7818
rect 11704 7754 11756 7760
rect 11888 7754 11940 7760
rect 11428 7540 11480 7546
rect 11428 7482 11480 7488
rect 10784 7336 10836 7342
rect 10784 7278 10836 7284
rect 11336 7336 11388 7342
rect 11336 7278 11388 7284
rect 11244 6792 11296 6798
rect 11244 6734 11296 6740
rect 10692 6724 10744 6730
rect 10692 6666 10744 6672
rect 10784 6656 10836 6662
rect 10784 6598 10836 6604
rect 10796 6322 10824 6598
rect 10860 6556 11168 6576
rect 10860 6554 10866 6556
rect 10922 6554 10946 6556
rect 11002 6554 11026 6556
rect 11082 6554 11106 6556
rect 11162 6554 11168 6556
rect 10922 6502 10924 6554
rect 11104 6502 11106 6554
rect 10860 6500 10866 6502
rect 10922 6500 10946 6502
rect 11002 6500 11026 6502
rect 11082 6500 11106 6502
rect 11162 6500 11168 6502
rect 10860 6480 11168 6500
rect 11256 6458 11284 6734
rect 11244 6452 11296 6458
rect 11244 6394 11296 6400
rect 11348 6390 11376 7278
rect 11520 6792 11572 6798
rect 11518 6760 11520 6769
rect 11572 6760 11574 6769
rect 11518 6695 11574 6704
rect 11520 6656 11572 6662
rect 11520 6598 11572 6604
rect 11532 6458 11560 6598
rect 11520 6452 11572 6458
rect 11520 6394 11572 6400
rect 11336 6384 11388 6390
rect 11336 6326 11388 6332
rect 10784 6316 10836 6322
rect 10784 6258 10836 6264
rect 11612 6180 11664 6186
rect 11716 6168 11744 7754
rect 11900 7041 11928 7754
rect 11992 7478 12020 8978
rect 12176 8566 12204 8978
rect 12164 8560 12216 8566
rect 12164 8502 12216 8508
rect 12176 8362 12204 8502
rect 12164 8356 12216 8362
rect 12164 8298 12216 8304
rect 12268 8090 12296 10474
rect 12410 10364 12718 10384
rect 12410 10362 12416 10364
rect 12472 10362 12496 10364
rect 12552 10362 12576 10364
rect 12632 10362 12656 10364
rect 12712 10362 12718 10364
rect 12472 10310 12474 10362
rect 12654 10310 12656 10362
rect 12410 10308 12416 10310
rect 12472 10308 12496 10310
rect 12552 10308 12576 10310
rect 12632 10308 12656 10310
rect 12712 10308 12718 10310
rect 12410 10288 12718 10308
rect 12820 10266 12848 11200
rect 13960 10908 14268 10928
rect 13960 10906 13966 10908
rect 14022 10906 14046 10908
rect 14102 10906 14126 10908
rect 14182 10906 14206 10908
rect 14262 10906 14268 10908
rect 14022 10854 14024 10906
rect 14204 10854 14206 10906
rect 13960 10852 13966 10854
rect 14022 10852 14046 10854
rect 14102 10852 14126 10854
rect 14182 10852 14206 10854
rect 14262 10852 14268 10854
rect 13960 10832 14268 10852
rect 13360 10736 13412 10742
rect 13360 10678 13412 10684
rect 13268 10668 13320 10674
rect 13268 10610 13320 10616
rect 12808 10260 12860 10266
rect 12808 10202 12860 10208
rect 13280 9722 13308 10610
rect 13268 9716 13320 9722
rect 13268 9658 13320 9664
rect 12532 9648 12584 9654
rect 12532 9590 12584 9596
rect 12544 9518 12572 9590
rect 12532 9512 12584 9518
rect 12532 9454 12584 9460
rect 12900 9512 12952 9518
rect 12900 9454 12952 9460
rect 12410 9276 12718 9296
rect 12410 9274 12416 9276
rect 12472 9274 12496 9276
rect 12552 9274 12576 9276
rect 12632 9274 12656 9276
rect 12712 9274 12718 9276
rect 12472 9222 12474 9274
rect 12654 9222 12656 9274
rect 12410 9220 12416 9222
rect 12472 9220 12496 9222
rect 12552 9220 12576 9222
rect 12632 9220 12656 9222
rect 12712 9220 12718 9222
rect 12410 9200 12718 9220
rect 12440 8900 12492 8906
rect 12440 8842 12492 8848
rect 12452 8401 12480 8842
rect 12438 8392 12494 8401
rect 12438 8327 12494 8336
rect 12410 8188 12718 8208
rect 12410 8186 12416 8188
rect 12472 8186 12496 8188
rect 12552 8186 12576 8188
rect 12632 8186 12656 8188
rect 12712 8186 12718 8188
rect 12472 8134 12474 8186
rect 12654 8134 12656 8186
rect 12410 8132 12416 8134
rect 12472 8132 12496 8134
rect 12552 8132 12576 8134
rect 12632 8132 12656 8134
rect 12712 8132 12718 8134
rect 12410 8112 12718 8132
rect 12256 8084 12308 8090
rect 12256 8026 12308 8032
rect 12348 7880 12400 7886
rect 12348 7822 12400 7828
rect 11980 7472 12032 7478
rect 11980 7414 12032 7420
rect 12360 7410 12388 7822
rect 12348 7404 12400 7410
rect 12348 7346 12400 7352
rect 12410 7100 12718 7120
rect 12410 7098 12416 7100
rect 12472 7098 12496 7100
rect 12552 7098 12576 7100
rect 12632 7098 12656 7100
rect 12712 7098 12718 7100
rect 12472 7046 12474 7098
rect 12654 7046 12656 7098
rect 12410 7044 12416 7046
rect 12472 7044 12496 7046
rect 12552 7044 12576 7046
rect 12632 7044 12656 7046
rect 12712 7044 12718 7046
rect 11886 7032 11942 7041
rect 12410 7024 12718 7044
rect 11886 6967 11942 6976
rect 11888 6860 11940 6866
rect 11888 6802 11940 6808
rect 11900 6458 11928 6802
rect 11888 6452 11940 6458
rect 11888 6394 11940 6400
rect 11796 6384 11848 6390
rect 11796 6326 11848 6332
rect 11664 6140 11744 6168
rect 11612 6122 11664 6128
rect 11520 6112 11572 6118
rect 11520 6054 11572 6060
rect 11532 5642 11560 6054
rect 11808 5710 11836 6326
rect 12410 6012 12718 6032
rect 12410 6010 12416 6012
rect 12472 6010 12496 6012
rect 12552 6010 12576 6012
rect 12632 6010 12656 6012
rect 12712 6010 12718 6012
rect 12472 5958 12474 6010
rect 12654 5958 12656 6010
rect 12410 5956 12416 5958
rect 12472 5956 12496 5958
rect 12552 5956 12576 5958
rect 12632 5956 12656 5958
rect 12712 5956 12718 5958
rect 12410 5936 12718 5956
rect 11796 5704 11848 5710
rect 11796 5646 11848 5652
rect 11520 5636 11572 5642
rect 11520 5578 11572 5584
rect 10860 5468 11168 5488
rect 10860 5466 10866 5468
rect 10922 5466 10946 5468
rect 11002 5466 11026 5468
rect 11082 5466 11106 5468
rect 11162 5466 11168 5468
rect 10922 5414 10924 5466
rect 11104 5414 11106 5466
rect 10860 5412 10866 5414
rect 10922 5412 10946 5414
rect 11002 5412 11026 5414
rect 11082 5412 11106 5414
rect 11162 5412 11168 5414
rect 10860 5392 11168 5412
rect 10600 5364 10652 5370
rect 10600 5306 10652 5312
rect 9128 5296 9180 5302
rect 8942 5264 8998 5273
rect 9128 5238 9180 5244
rect 8942 5199 8944 5208
rect 8996 5199 8998 5208
rect 9772 5228 9824 5234
rect 9772 5170 9824 5176
rect 8944 5160 8996 5166
rect 9310 4924 9618 4944
rect 9310 4922 9316 4924
rect 9372 4922 9396 4924
rect 9452 4922 9476 4924
rect 9532 4922 9556 4924
rect 9612 4922 9618 4924
rect 9372 4870 9374 4922
rect 9554 4870 9556 4922
rect 9310 4868 9316 4870
rect 9372 4868 9396 4870
rect 9452 4868 9476 4870
rect 9532 4868 9556 4870
rect 9612 4868 9618 4870
rect 9310 4848 9618 4868
rect 8760 4684 8812 4690
rect 8760 4626 8812 4632
rect 9036 4616 9088 4622
rect 9646 4598 9720 4604
rect 9036 4558 9088 4564
rect 9634 4593 9720 4598
rect 9634 4592 9734 4593
rect 9686 4584 9734 4592
rect 8484 4548 8536 4554
rect 8484 4490 8536 4496
rect 8208 4276 8260 4282
rect 8208 4218 8260 4224
rect 8944 4208 8996 4214
rect 8944 4150 8996 4156
rect 7472 4140 7524 4146
rect 7472 4082 7524 4088
rect 7484 3738 7512 4082
rect 8760 4072 8812 4078
rect 8760 4014 8812 4020
rect 7472 3732 7524 3738
rect 7472 3674 7524 3680
rect 7484 3126 7512 3674
rect 8772 3466 8800 4014
rect 8760 3460 8812 3466
rect 8760 3402 8812 3408
rect 8668 3392 8720 3398
rect 8668 3334 8720 3340
rect 7760 3292 8068 3312
rect 7760 3290 7766 3292
rect 7822 3290 7846 3292
rect 7902 3290 7926 3292
rect 7982 3290 8006 3292
rect 8062 3290 8068 3292
rect 7822 3238 7824 3290
rect 8004 3238 8006 3290
rect 7760 3236 7766 3238
rect 7822 3236 7846 3238
rect 7902 3236 7926 3238
rect 7982 3236 8006 3238
rect 8062 3236 8068 3238
rect 7760 3216 8068 3236
rect 7472 3120 7524 3126
rect 7472 3062 7524 3068
rect 8300 3120 8352 3126
rect 8300 3062 8352 3068
rect 7564 3052 7616 3058
rect 7564 2994 7616 3000
rect 7656 3052 7708 3058
rect 7656 2994 7708 3000
rect 7840 3052 7892 3058
rect 7840 2994 7892 3000
rect 7576 2650 7604 2994
rect 7564 2644 7616 2650
rect 7564 2586 7616 2592
rect 7668 2582 7696 2994
rect 7656 2576 7708 2582
rect 7656 2518 7708 2524
rect 7852 2378 7880 2994
rect 8312 2446 8340 3062
rect 8680 3058 8708 3334
rect 8668 3052 8720 3058
rect 8668 2994 8720 3000
rect 8760 2848 8812 2854
rect 8760 2790 8812 2796
rect 8300 2440 8352 2446
rect 8300 2382 8352 2388
rect 8576 2440 8628 2446
rect 8576 2382 8628 2388
rect 8668 2440 8720 2446
rect 8668 2382 8720 2388
rect 7840 2372 7892 2378
rect 7840 2314 7892 2320
rect 8208 2304 8260 2310
rect 8208 2246 8260 2252
rect 7760 2204 8068 2224
rect 7760 2202 7766 2204
rect 7822 2202 7846 2204
rect 7902 2202 7926 2204
rect 7982 2202 8006 2204
rect 8062 2202 8068 2204
rect 7822 2150 7824 2202
rect 8004 2150 8006 2202
rect 7760 2148 7766 2150
rect 7822 2148 7846 2150
rect 7902 2148 7926 2150
rect 7982 2148 8006 2150
rect 8062 2148 8068 2150
rect 7760 2128 8068 2148
rect 7380 1964 7432 1970
rect 7380 1906 7432 1912
rect 7288 1760 7340 1766
rect 7288 1702 7340 1708
rect 6696 1244 6776 1272
rect 6644 1226 6696 1232
rect 5540 1012 5592 1018
rect 5540 954 5592 960
rect 6552 1012 6604 1018
rect 6552 954 6604 960
rect 5448 876 5500 882
rect 5368 836 5448 864
rect 5448 818 5500 824
rect 5264 740 5316 746
rect 5264 682 5316 688
rect 4160 468 4212 474
rect 4160 410 4212 416
rect 5460 406 5488 818
rect 6000 672 6052 678
rect 6000 614 6052 620
rect 5448 400 5500 406
rect 5448 342 5500 348
rect 2964 332 3016 338
rect 2964 274 3016 280
rect 6012 270 6040 614
rect 6210 572 6518 592
rect 6210 570 6216 572
rect 6272 570 6296 572
rect 6352 570 6376 572
rect 6432 570 6456 572
rect 6512 570 6518 572
rect 6272 518 6274 570
rect 6454 518 6456 570
rect 6210 516 6216 518
rect 6272 516 6296 518
rect 6352 516 6376 518
rect 6432 516 6456 518
rect 6512 516 6518 518
rect 6210 496 6518 516
rect 6656 338 6684 1226
rect 6920 1216 6972 1222
rect 6920 1158 6972 1164
rect 6932 406 6960 1158
rect 7392 814 7420 1906
rect 7656 1896 7708 1902
rect 7656 1838 7708 1844
rect 7668 1358 7696 1838
rect 7656 1352 7708 1358
rect 7656 1294 7708 1300
rect 7760 1116 8068 1136
rect 7760 1114 7766 1116
rect 7822 1114 7846 1116
rect 7902 1114 7926 1116
rect 7982 1114 8006 1116
rect 8062 1114 8068 1116
rect 7822 1062 7824 1114
rect 8004 1062 8006 1114
rect 7760 1060 7766 1062
rect 7822 1060 7846 1062
rect 7902 1060 7926 1062
rect 7982 1060 8006 1062
rect 8062 1060 8068 1062
rect 7760 1040 8068 1060
rect 7380 808 7432 814
rect 7380 750 7432 756
rect 8116 808 8168 814
rect 8116 750 8168 756
rect 8128 474 8156 750
rect 8116 468 8168 474
rect 8116 410 8168 416
rect 6920 400 6972 406
rect 6920 342 6972 348
rect 6644 332 6696 338
rect 6644 274 6696 280
rect 6000 264 6052 270
rect 6000 206 6052 212
rect 8220 202 8248 2246
rect 8588 270 8616 2382
rect 8680 2106 8708 2382
rect 8668 2100 8720 2106
rect 8668 2042 8720 2048
rect 8680 1494 8708 2042
rect 8668 1488 8720 1494
rect 8668 1430 8720 1436
rect 8668 1352 8720 1358
rect 8772 1306 8800 2790
rect 8720 1300 8800 1306
rect 8668 1294 8800 1300
rect 8680 1278 8800 1294
rect 8680 406 8708 1278
rect 8956 1018 8984 4150
rect 9048 3346 9076 4558
rect 9634 4534 9678 4540
rect 9678 4519 9734 4528
rect 9128 4480 9180 4486
rect 9128 4422 9180 4428
rect 9140 3534 9168 4422
rect 9784 4282 9812 5170
rect 10048 5024 10100 5030
rect 10048 4966 10100 4972
rect 9864 4820 9916 4826
rect 9864 4762 9916 4768
rect 9772 4276 9824 4282
rect 9772 4218 9824 4224
rect 9772 4140 9824 4146
rect 9876 4128 9904 4762
rect 10060 4554 10088 4966
rect 10612 4690 10640 5306
rect 12256 5160 12308 5166
rect 12256 5102 12308 5108
rect 12268 4826 12296 5102
rect 12808 5092 12860 5098
rect 12808 5034 12860 5040
rect 12410 4924 12718 4944
rect 12410 4922 12416 4924
rect 12472 4922 12496 4924
rect 12552 4922 12576 4924
rect 12632 4922 12656 4924
rect 12712 4922 12718 4924
rect 12472 4870 12474 4922
rect 12654 4870 12656 4922
rect 12410 4868 12416 4870
rect 12472 4868 12496 4870
rect 12552 4868 12576 4870
rect 12632 4868 12656 4870
rect 12712 4868 12718 4870
rect 12410 4848 12718 4868
rect 12256 4820 12308 4826
rect 12256 4762 12308 4768
rect 10600 4684 10652 4690
rect 10600 4626 10652 4632
rect 12072 4684 12124 4690
rect 12072 4626 12124 4632
rect 10048 4548 10100 4554
rect 10048 4490 10100 4496
rect 9824 4100 9904 4128
rect 9772 4082 9824 4088
rect 9680 4072 9732 4078
rect 9680 4014 9732 4020
rect 9310 3836 9618 3856
rect 9310 3834 9316 3836
rect 9372 3834 9396 3836
rect 9452 3834 9476 3836
rect 9532 3834 9556 3836
rect 9612 3834 9618 3836
rect 9372 3782 9374 3834
rect 9554 3782 9556 3834
rect 9310 3780 9316 3782
rect 9372 3780 9396 3782
rect 9452 3780 9476 3782
rect 9532 3780 9556 3782
rect 9612 3780 9618 3782
rect 9310 3760 9618 3780
rect 9692 3738 9720 4014
rect 9680 3732 9732 3738
rect 9680 3674 9732 3680
rect 9784 3534 9812 4082
rect 9128 3528 9180 3534
rect 9128 3470 9180 3476
rect 9772 3528 9824 3534
rect 9772 3470 9824 3476
rect 10612 3516 10640 4626
rect 11334 4584 11390 4593
rect 11334 4519 11336 4528
rect 11388 4519 11390 4528
rect 11428 4548 11480 4554
rect 11336 4490 11388 4496
rect 11428 4490 11480 4496
rect 10860 4380 11168 4400
rect 10860 4378 10866 4380
rect 10922 4378 10946 4380
rect 11002 4378 11026 4380
rect 11082 4378 11106 4380
rect 11162 4378 11168 4380
rect 10922 4326 10924 4378
rect 11104 4326 11106 4378
rect 10860 4324 10866 4326
rect 10922 4324 10946 4326
rect 11002 4324 11026 4326
rect 11082 4324 11106 4326
rect 11162 4324 11168 4326
rect 10860 4304 11168 4324
rect 10784 4140 10836 4146
rect 10784 4082 10836 4088
rect 10876 4140 10928 4146
rect 10876 4082 10928 4088
rect 10796 4010 10824 4082
rect 10784 4004 10836 4010
rect 10784 3946 10836 3952
rect 10888 3602 10916 4082
rect 10876 3596 10928 3602
rect 10876 3538 10928 3544
rect 10692 3528 10744 3534
rect 10612 3488 10692 3516
rect 9048 3318 9168 3346
rect 9140 3126 9168 3318
rect 9128 3120 9180 3126
rect 9128 3062 9180 3068
rect 9140 2394 9168 3062
rect 10612 2990 10640 3488
rect 10692 3470 10744 3476
rect 10860 3292 11168 3312
rect 10860 3290 10866 3292
rect 10922 3290 10946 3292
rect 11002 3290 11026 3292
rect 11082 3290 11106 3292
rect 11162 3290 11168 3292
rect 10922 3238 10924 3290
rect 11104 3238 11106 3290
rect 10860 3236 10866 3238
rect 10922 3236 10946 3238
rect 11002 3236 11026 3238
rect 11082 3236 11106 3238
rect 11162 3236 11168 3238
rect 10860 3216 11168 3236
rect 11348 3126 11376 4490
rect 11440 4078 11468 4490
rect 11520 4480 11572 4486
rect 11520 4422 11572 4428
rect 11532 4146 11560 4422
rect 11612 4208 11664 4214
rect 11612 4150 11664 4156
rect 11520 4140 11572 4146
rect 11520 4082 11572 4088
rect 11428 4072 11480 4078
rect 11428 4014 11480 4020
rect 11336 3120 11388 3126
rect 11336 3062 11388 3068
rect 10600 2984 10652 2990
rect 10600 2926 10652 2932
rect 10232 2848 10284 2854
rect 10232 2790 10284 2796
rect 9310 2748 9618 2768
rect 9310 2746 9316 2748
rect 9372 2746 9396 2748
rect 9452 2746 9476 2748
rect 9532 2746 9556 2748
rect 9612 2746 9618 2748
rect 9372 2694 9374 2746
rect 9554 2694 9556 2746
rect 9310 2692 9316 2694
rect 9372 2692 9396 2694
rect 9452 2692 9476 2694
rect 9532 2692 9556 2694
rect 9612 2692 9618 2694
rect 9310 2672 9618 2692
rect 10244 2446 10272 2790
rect 9048 2366 9168 2394
rect 10232 2440 10284 2446
rect 10232 2382 10284 2388
rect 9048 2038 9076 2366
rect 9128 2304 9180 2310
rect 9128 2246 9180 2252
rect 9036 2032 9088 2038
rect 9036 1974 9088 1980
rect 8944 1012 8996 1018
rect 8944 954 8996 960
rect 9048 950 9076 1974
rect 9140 1358 9168 2246
rect 10860 2204 11168 2224
rect 10860 2202 10866 2204
rect 10922 2202 10946 2204
rect 11002 2202 11026 2204
rect 11082 2202 11106 2204
rect 11162 2202 11168 2204
rect 10922 2150 10924 2202
rect 11104 2150 11106 2202
rect 10860 2148 10866 2150
rect 10922 2148 10946 2150
rect 11002 2148 11026 2150
rect 11082 2148 11106 2150
rect 11162 2148 11168 2150
rect 10860 2128 11168 2148
rect 11624 2106 11652 4150
rect 12084 4146 12112 4626
rect 12820 4622 12848 5034
rect 12808 4616 12860 4622
rect 12808 4558 12860 4564
rect 12256 4548 12308 4554
rect 12256 4490 12308 4496
rect 12072 4140 12124 4146
rect 12072 4082 12124 4088
rect 12268 4128 12296 4490
rect 12624 4480 12676 4486
rect 12624 4422 12676 4428
rect 12636 4146 12664 4422
rect 12348 4140 12400 4146
rect 12268 4100 12348 4128
rect 11704 4072 11756 4078
rect 11704 4014 11756 4020
rect 11716 3738 11744 4014
rect 11704 3732 11756 3738
rect 11704 3674 11756 3680
rect 12084 3466 12112 4082
rect 12268 3466 12296 4100
rect 12348 4082 12400 4088
rect 12624 4140 12676 4146
rect 12624 4082 12676 4088
rect 12636 4010 12664 4082
rect 12624 4004 12676 4010
rect 12624 3946 12676 3952
rect 12808 3936 12860 3942
rect 12808 3878 12860 3884
rect 12410 3836 12718 3856
rect 12410 3834 12416 3836
rect 12472 3834 12496 3836
rect 12552 3834 12576 3836
rect 12632 3834 12656 3836
rect 12712 3834 12718 3836
rect 12472 3782 12474 3834
rect 12654 3782 12656 3834
rect 12410 3780 12416 3782
rect 12472 3780 12496 3782
rect 12552 3780 12576 3782
rect 12632 3780 12656 3782
rect 12712 3780 12718 3782
rect 12410 3760 12718 3780
rect 12820 3738 12848 3878
rect 12912 3738 12940 9454
rect 13372 9178 13400 10678
rect 13636 10600 13688 10606
rect 13636 10542 13688 10548
rect 14832 10600 14884 10606
rect 14832 10542 14884 10548
rect 13648 10266 13676 10542
rect 13636 10260 13688 10266
rect 13636 10202 13688 10208
rect 14844 10130 14872 10542
rect 15200 10464 15252 10470
rect 15200 10406 15252 10412
rect 15292 10464 15344 10470
rect 15292 10406 15344 10412
rect 15212 10130 15240 10406
rect 14832 10124 14884 10130
rect 14832 10066 14884 10072
rect 15200 10124 15252 10130
rect 15200 10066 15252 10072
rect 15304 10062 15332 10406
rect 15292 10056 15344 10062
rect 15292 9998 15344 10004
rect 13960 9820 14268 9840
rect 13960 9818 13966 9820
rect 14022 9818 14046 9820
rect 14102 9818 14126 9820
rect 14182 9818 14206 9820
rect 14262 9818 14268 9820
rect 14022 9766 14024 9818
rect 14204 9766 14206 9818
rect 13960 9764 13966 9766
rect 14022 9764 14046 9766
rect 14102 9764 14126 9766
rect 14182 9764 14206 9766
rect 14262 9764 14268 9766
rect 13960 9744 14268 9764
rect 13544 9512 13596 9518
rect 13544 9454 13596 9460
rect 14372 9512 14424 9518
rect 14372 9454 14424 9460
rect 13360 9172 13412 9178
rect 13360 9114 13412 9120
rect 13372 8974 13400 9114
rect 13556 8974 13584 9454
rect 13728 9036 13780 9042
rect 13728 8978 13780 8984
rect 13360 8968 13412 8974
rect 13360 8910 13412 8916
rect 13544 8968 13596 8974
rect 13544 8910 13596 8916
rect 13452 8832 13504 8838
rect 13452 8774 13504 8780
rect 13464 8430 13492 8774
rect 13452 8424 13504 8430
rect 13452 8366 13504 8372
rect 12992 7880 13044 7886
rect 12992 7822 13044 7828
rect 13004 7002 13032 7822
rect 13556 7313 13584 8910
rect 13740 8566 13768 8978
rect 14384 8906 14412 9454
rect 14464 9376 14516 9382
rect 14464 9318 14516 9324
rect 14372 8900 14424 8906
rect 14372 8842 14424 8848
rect 13820 8832 13872 8838
rect 13820 8774 13872 8780
rect 13728 8560 13780 8566
rect 13728 8502 13780 8508
rect 13832 8430 13860 8774
rect 13960 8732 14268 8752
rect 13960 8730 13966 8732
rect 14022 8730 14046 8732
rect 14102 8730 14126 8732
rect 14182 8730 14206 8732
rect 14262 8730 14268 8732
rect 14022 8678 14024 8730
rect 14204 8678 14206 8730
rect 13960 8676 13966 8678
rect 14022 8676 14046 8678
rect 14102 8676 14126 8678
rect 14182 8676 14206 8678
rect 14262 8676 14268 8678
rect 13960 8656 14268 8676
rect 14372 8492 14424 8498
rect 14372 8434 14424 8440
rect 13820 8424 13872 8430
rect 13820 8366 13872 8372
rect 13820 8288 13872 8294
rect 13820 8230 13872 8236
rect 13832 7886 13860 8230
rect 14384 8090 14412 8434
rect 14372 8084 14424 8090
rect 14372 8026 14424 8032
rect 13820 7880 13872 7886
rect 13820 7822 13872 7828
rect 13960 7644 14268 7664
rect 13960 7642 13966 7644
rect 14022 7642 14046 7644
rect 14102 7642 14126 7644
rect 14182 7642 14206 7644
rect 14262 7642 14268 7644
rect 14022 7590 14024 7642
rect 14204 7590 14206 7642
rect 13960 7588 13966 7590
rect 14022 7588 14046 7590
rect 14102 7588 14126 7590
rect 14182 7588 14206 7590
rect 14262 7588 14268 7590
rect 13960 7568 14268 7588
rect 13542 7304 13598 7313
rect 13542 7239 13598 7248
rect 12992 6996 13044 7002
rect 12992 6938 13044 6944
rect 13556 6798 13584 7239
rect 13544 6792 13596 6798
rect 13544 6734 13596 6740
rect 13176 6656 13228 6662
rect 13176 6598 13228 6604
rect 13820 6656 13872 6662
rect 13820 6598 13872 6604
rect 12992 6248 13044 6254
rect 12992 6190 13044 6196
rect 13004 5914 13032 6190
rect 12992 5908 13044 5914
rect 12992 5850 13044 5856
rect 13188 5710 13216 6598
rect 13832 6458 13860 6598
rect 13960 6556 14268 6576
rect 13960 6554 13966 6556
rect 14022 6554 14046 6556
rect 14102 6554 14126 6556
rect 14182 6554 14206 6556
rect 14262 6554 14268 6556
rect 14022 6502 14024 6554
rect 14204 6502 14206 6554
rect 13960 6500 13966 6502
rect 14022 6500 14046 6502
rect 14102 6500 14126 6502
rect 14182 6500 14206 6502
rect 14262 6500 14268 6502
rect 13960 6480 14268 6500
rect 13820 6452 13872 6458
rect 13820 6394 13872 6400
rect 13820 6316 13872 6322
rect 13820 6258 13872 6264
rect 13176 5704 13228 5710
rect 13176 5646 13228 5652
rect 13832 5574 13860 6258
rect 13820 5568 13872 5574
rect 13820 5510 13872 5516
rect 13832 5302 13860 5510
rect 13960 5468 14268 5488
rect 13960 5466 13966 5468
rect 14022 5466 14046 5468
rect 14102 5466 14126 5468
rect 14182 5466 14206 5468
rect 14262 5466 14268 5468
rect 14022 5414 14024 5466
rect 14204 5414 14206 5466
rect 13960 5412 13966 5414
rect 14022 5412 14046 5414
rect 14102 5412 14126 5414
rect 14182 5412 14206 5414
rect 14262 5412 14268 5414
rect 13960 5392 14268 5412
rect 13820 5296 13872 5302
rect 13820 5238 13872 5244
rect 14476 4826 14504 9318
rect 15292 8968 15344 8974
rect 15292 8910 15344 8916
rect 15304 8566 15332 8910
rect 15292 8560 15344 8566
rect 15292 8502 15344 8508
rect 14556 8492 14608 8498
rect 14556 8434 14608 8440
rect 14568 8090 14596 8434
rect 14924 8288 14976 8294
rect 14924 8230 14976 8236
rect 14556 8084 14608 8090
rect 14556 8026 14608 8032
rect 14936 7886 14964 8230
rect 14740 7880 14792 7886
rect 14924 7880 14976 7886
rect 14792 7840 14924 7868
rect 14740 7822 14792 7828
rect 14924 7822 14976 7828
rect 15200 7880 15252 7886
rect 15200 7822 15252 7828
rect 14740 7744 14792 7750
rect 14740 7686 14792 7692
rect 14924 7744 14976 7750
rect 14924 7686 14976 7692
rect 14752 7410 14780 7686
rect 14740 7404 14792 7410
rect 14740 7346 14792 7352
rect 14832 6860 14884 6866
rect 14936 6848 14964 7686
rect 15212 7410 15240 7822
rect 15200 7404 15252 7410
rect 15200 7346 15252 7352
rect 15016 7200 15068 7206
rect 15016 7142 15068 7148
rect 15028 6866 15056 7142
rect 15212 7002 15240 7346
rect 15200 6996 15252 7002
rect 15200 6938 15252 6944
rect 14884 6820 14964 6848
rect 14832 6802 14884 6808
rect 14832 6656 14884 6662
rect 14832 6598 14884 6604
rect 14844 6458 14872 6598
rect 14832 6452 14884 6458
rect 14832 6394 14884 6400
rect 14936 6254 14964 6820
rect 15016 6860 15068 6866
rect 15016 6802 15068 6808
rect 15200 6792 15252 6798
rect 15200 6734 15252 6740
rect 14924 6248 14976 6254
rect 14924 6190 14976 6196
rect 14924 6112 14976 6118
rect 14924 6054 14976 6060
rect 14936 5778 14964 6054
rect 15212 5778 15240 6734
rect 15396 5846 15424 11206
rect 15580 11098 15608 11206
rect 15658 11200 15714 12000
rect 18510 11200 18566 12000
rect 18786 11248 18842 11257
rect 15672 11098 15700 11200
rect 15580 11070 15700 11098
rect 17060 10908 17368 10928
rect 17060 10906 17066 10908
rect 17122 10906 17146 10908
rect 17202 10906 17226 10908
rect 17282 10906 17306 10908
rect 17362 10906 17368 10908
rect 17122 10854 17124 10906
rect 17304 10854 17306 10906
rect 17060 10852 17066 10854
rect 17122 10852 17146 10854
rect 17202 10852 17226 10854
rect 17282 10852 17306 10854
rect 17362 10852 17368 10854
rect 17060 10832 17368 10852
rect 15936 10736 15988 10742
rect 15936 10678 15988 10684
rect 15510 10364 15818 10384
rect 15510 10362 15516 10364
rect 15572 10362 15596 10364
rect 15652 10362 15676 10364
rect 15732 10362 15756 10364
rect 15812 10362 15818 10364
rect 15572 10310 15574 10362
rect 15754 10310 15756 10362
rect 15510 10308 15516 10310
rect 15572 10308 15596 10310
rect 15652 10308 15676 10310
rect 15732 10308 15756 10310
rect 15812 10308 15818 10310
rect 15510 10288 15818 10308
rect 15948 9994 15976 10678
rect 18328 10668 18380 10674
rect 18328 10610 18380 10616
rect 16488 10600 16540 10606
rect 16488 10542 16540 10548
rect 16500 10266 16528 10542
rect 18340 10266 18368 10610
rect 16488 10260 16540 10266
rect 16488 10202 16540 10208
rect 18328 10260 18380 10266
rect 18328 10202 18380 10208
rect 17960 10056 18012 10062
rect 17960 9998 18012 10004
rect 15936 9988 15988 9994
rect 15936 9930 15988 9936
rect 15948 9586 15976 9930
rect 17776 9920 17828 9926
rect 17776 9862 17828 9868
rect 17060 9820 17368 9840
rect 17060 9818 17066 9820
rect 17122 9818 17146 9820
rect 17202 9818 17226 9820
rect 17282 9818 17306 9820
rect 17362 9818 17368 9820
rect 17122 9766 17124 9818
rect 17304 9766 17306 9818
rect 17060 9764 17066 9766
rect 17122 9764 17146 9766
rect 17202 9764 17226 9766
rect 17282 9764 17306 9766
rect 17362 9764 17368 9766
rect 17060 9744 17368 9764
rect 17788 9654 17816 9862
rect 17972 9761 18000 9998
rect 17958 9752 18014 9761
rect 17958 9687 18014 9696
rect 17776 9648 17828 9654
rect 17776 9590 17828 9596
rect 15936 9580 15988 9586
rect 15936 9522 15988 9528
rect 15844 9512 15896 9518
rect 15844 9454 15896 9460
rect 16488 9512 16540 9518
rect 17960 9512 18012 9518
rect 16488 9454 16540 9460
rect 17880 9472 17960 9500
rect 15510 9276 15818 9296
rect 15510 9274 15516 9276
rect 15572 9274 15596 9276
rect 15652 9274 15676 9276
rect 15732 9274 15756 9276
rect 15812 9274 15818 9276
rect 15572 9222 15574 9274
rect 15754 9222 15756 9274
rect 15510 9220 15516 9222
rect 15572 9220 15596 9222
rect 15652 9220 15676 9222
rect 15732 9220 15756 9222
rect 15812 9220 15818 9222
rect 15510 9200 15818 9220
rect 15856 8974 15884 9454
rect 15844 8968 15896 8974
rect 15844 8910 15896 8916
rect 16120 8968 16172 8974
rect 16120 8910 16172 8916
rect 15856 8430 15884 8910
rect 16132 8650 16160 8910
rect 16500 8906 16528 9454
rect 16672 9036 16724 9042
rect 16672 8978 16724 8984
rect 16488 8900 16540 8906
rect 16488 8842 16540 8848
rect 16040 8622 16160 8650
rect 16040 8566 16068 8622
rect 16028 8560 16080 8566
rect 16028 8502 16080 8508
rect 16304 8560 16356 8566
rect 16500 8548 16528 8842
rect 16356 8520 16528 8548
rect 16304 8502 16356 8508
rect 15844 8424 15896 8430
rect 15844 8366 15896 8372
rect 15510 8188 15818 8208
rect 15510 8186 15516 8188
rect 15572 8186 15596 8188
rect 15652 8186 15676 8188
rect 15732 8186 15756 8188
rect 15812 8186 15818 8188
rect 15572 8134 15574 8186
rect 15754 8134 15756 8186
rect 15510 8132 15516 8134
rect 15572 8132 15596 8134
rect 15652 8132 15676 8134
rect 15732 8132 15756 8134
rect 15812 8132 15818 8134
rect 15510 8112 15818 8132
rect 15856 7954 15884 8366
rect 15844 7948 15896 7954
rect 15844 7890 15896 7896
rect 16316 7818 16344 8502
rect 15568 7812 15620 7818
rect 15568 7754 15620 7760
rect 16304 7812 16356 7818
rect 16304 7754 16356 7760
rect 15580 7546 15608 7754
rect 15568 7540 15620 7546
rect 15568 7482 15620 7488
rect 16316 7478 16344 7754
rect 16304 7472 16356 7478
rect 16304 7414 16356 7420
rect 15510 7100 15818 7120
rect 15510 7098 15516 7100
rect 15572 7098 15596 7100
rect 15652 7098 15676 7100
rect 15732 7098 15756 7100
rect 15812 7098 15818 7100
rect 15572 7046 15574 7098
rect 15754 7046 15756 7098
rect 15510 7044 15516 7046
rect 15572 7044 15596 7046
rect 15652 7044 15676 7046
rect 15732 7044 15756 7046
rect 15812 7044 15818 7046
rect 15510 7024 15818 7044
rect 15568 6860 15620 6866
rect 15568 6802 15620 6808
rect 15476 6792 15528 6798
rect 15476 6734 15528 6740
rect 15488 6390 15516 6734
rect 15476 6384 15528 6390
rect 15476 6326 15528 6332
rect 15580 6322 15608 6802
rect 15568 6316 15620 6322
rect 15568 6258 15620 6264
rect 15510 6012 15818 6032
rect 15510 6010 15516 6012
rect 15572 6010 15596 6012
rect 15652 6010 15676 6012
rect 15732 6010 15756 6012
rect 15812 6010 15818 6012
rect 15572 5958 15574 6010
rect 15754 5958 15756 6010
rect 15510 5956 15516 5958
rect 15572 5956 15596 5958
rect 15652 5956 15676 5958
rect 15732 5956 15756 5958
rect 15812 5956 15818 5958
rect 15510 5936 15818 5956
rect 15384 5840 15436 5846
rect 15384 5782 15436 5788
rect 14924 5772 14976 5778
rect 14924 5714 14976 5720
rect 15200 5772 15252 5778
rect 15200 5714 15252 5720
rect 15108 5636 15160 5642
rect 15108 5578 15160 5584
rect 15120 5302 15148 5578
rect 16316 5302 16344 7414
rect 16396 6656 16448 6662
rect 16396 6598 16448 6604
rect 16408 6322 16436 6598
rect 16396 6316 16448 6322
rect 16396 6258 16448 6264
rect 16684 6254 16712 8978
rect 17060 8732 17368 8752
rect 17060 8730 17066 8732
rect 17122 8730 17146 8732
rect 17202 8730 17226 8732
rect 17282 8730 17306 8732
rect 17362 8730 17368 8732
rect 17122 8678 17124 8730
rect 17304 8678 17306 8730
rect 17060 8676 17066 8678
rect 17122 8676 17146 8678
rect 17202 8676 17226 8678
rect 17282 8676 17306 8678
rect 17362 8676 17368 8678
rect 17060 8656 17368 8676
rect 17880 8498 17908 9472
rect 17960 9454 18012 9460
rect 17960 9172 18012 9178
rect 17960 9114 18012 9120
rect 17500 8492 17552 8498
rect 17500 8434 17552 8440
rect 17868 8492 17920 8498
rect 17868 8434 17920 8440
rect 17060 7644 17368 7664
rect 17060 7642 17066 7644
rect 17122 7642 17146 7644
rect 17202 7642 17226 7644
rect 17282 7642 17306 7644
rect 17362 7642 17368 7644
rect 17122 7590 17124 7642
rect 17304 7590 17306 7642
rect 17060 7588 17066 7590
rect 17122 7588 17146 7590
rect 17202 7588 17226 7590
rect 17282 7588 17306 7590
rect 17362 7588 17368 7590
rect 17060 7568 17368 7588
rect 17512 7410 17540 8434
rect 17592 7812 17644 7818
rect 17592 7754 17644 7760
rect 17500 7404 17552 7410
rect 17500 7346 17552 7352
rect 17408 7200 17460 7206
rect 17408 7142 17460 7148
rect 17420 6798 17448 7142
rect 17604 6866 17632 7754
rect 17972 7546 18000 9114
rect 18524 8634 18552 11200
rect 18786 11183 18842 11192
rect 18800 10062 18828 11183
rect 18788 10056 18840 10062
rect 18788 9998 18840 10004
rect 18512 8628 18564 8634
rect 18512 8570 18564 8576
rect 18512 8492 18564 8498
rect 18512 8434 18564 8440
rect 18524 8265 18552 8434
rect 18510 8256 18566 8265
rect 18510 8191 18566 8200
rect 17960 7540 18012 7546
rect 17960 7482 18012 7488
rect 18328 7472 18380 7478
rect 18328 7414 18380 7420
rect 17868 7336 17920 7342
rect 17868 7278 17920 7284
rect 17880 7002 17908 7278
rect 18340 7002 18368 7414
rect 17868 6996 17920 7002
rect 17868 6938 17920 6944
rect 18328 6996 18380 7002
rect 18328 6938 18380 6944
rect 17592 6860 17644 6866
rect 17592 6802 17644 6808
rect 17408 6792 17460 6798
rect 17408 6734 17460 6740
rect 17776 6792 17828 6798
rect 18512 6792 18564 6798
rect 17776 6734 17828 6740
rect 18510 6760 18512 6769
rect 18564 6760 18566 6769
rect 17060 6556 17368 6576
rect 17060 6554 17066 6556
rect 17122 6554 17146 6556
rect 17202 6554 17226 6556
rect 17282 6554 17306 6556
rect 17362 6554 17368 6556
rect 17122 6502 17124 6554
rect 17304 6502 17306 6554
rect 17060 6500 17066 6502
rect 17122 6500 17146 6502
rect 17202 6500 17226 6502
rect 17282 6500 17306 6502
rect 17362 6500 17368 6502
rect 17060 6480 17368 6500
rect 17788 6458 17816 6734
rect 18510 6695 18566 6704
rect 17776 6452 17828 6458
rect 17776 6394 17828 6400
rect 17408 6384 17460 6390
rect 17408 6326 17460 6332
rect 16672 6248 16724 6254
rect 16672 6190 16724 6196
rect 16684 5778 16712 6190
rect 16672 5772 16724 5778
rect 16672 5714 16724 5720
rect 17060 5468 17368 5488
rect 17060 5466 17066 5468
rect 17122 5466 17146 5468
rect 17202 5466 17226 5468
rect 17282 5466 17306 5468
rect 17362 5466 17368 5468
rect 17122 5414 17124 5466
rect 17304 5414 17306 5466
rect 17060 5412 17066 5414
rect 17122 5412 17146 5414
rect 17202 5412 17226 5414
rect 17282 5412 17306 5414
rect 17362 5412 17368 5414
rect 17060 5392 17368 5412
rect 17420 5370 17448 6326
rect 18512 5704 18564 5710
rect 18512 5646 18564 5652
rect 18236 5568 18288 5574
rect 18236 5510 18288 5516
rect 17408 5364 17460 5370
rect 17408 5306 17460 5312
rect 15108 5296 15160 5302
rect 15108 5238 15160 5244
rect 16304 5296 16356 5302
rect 16304 5238 16356 5244
rect 17960 5296 18012 5302
rect 17960 5238 18012 5244
rect 14556 5160 14608 5166
rect 14556 5102 14608 5108
rect 14464 4820 14516 4826
rect 14464 4762 14516 4768
rect 14568 4690 14596 5102
rect 14556 4684 14608 4690
rect 14556 4626 14608 4632
rect 13960 4380 14268 4400
rect 13960 4378 13966 4380
rect 14022 4378 14046 4380
rect 14102 4378 14126 4380
rect 14182 4378 14206 4380
rect 14262 4378 14268 4380
rect 14022 4326 14024 4378
rect 14204 4326 14206 4378
rect 13960 4324 13966 4326
rect 14022 4324 14046 4326
rect 14102 4324 14126 4326
rect 14182 4324 14206 4326
rect 14262 4324 14268 4326
rect 13960 4304 14268 4324
rect 13360 4140 13412 4146
rect 13360 4082 13412 4088
rect 12808 3732 12860 3738
rect 12808 3674 12860 3680
rect 12900 3732 12952 3738
rect 12900 3674 12952 3680
rect 12072 3460 12124 3466
rect 12072 3402 12124 3408
rect 12256 3460 12308 3466
rect 12256 3402 12308 3408
rect 12912 3126 12940 3674
rect 13084 3528 13136 3534
rect 13084 3470 13136 3476
rect 12900 3120 12952 3126
rect 12900 3062 12952 3068
rect 12808 3052 12860 3058
rect 12808 2994 12860 3000
rect 12256 2984 12308 2990
rect 12256 2926 12308 2932
rect 11796 2848 11848 2854
rect 11796 2790 11848 2796
rect 11808 2446 11836 2790
rect 12268 2650 12296 2926
rect 12410 2748 12718 2768
rect 12410 2746 12416 2748
rect 12472 2746 12496 2748
rect 12552 2746 12576 2748
rect 12632 2746 12656 2748
rect 12712 2746 12718 2748
rect 12472 2694 12474 2746
rect 12654 2694 12656 2746
rect 12410 2692 12416 2694
rect 12472 2692 12496 2694
rect 12552 2692 12576 2694
rect 12632 2692 12656 2694
rect 12712 2692 12718 2694
rect 12410 2672 12718 2692
rect 12256 2644 12308 2650
rect 12256 2586 12308 2592
rect 12820 2582 12848 2994
rect 12900 2984 12952 2990
rect 12900 2926 12952 2932
rect 12808 2576 12860 2582
rect 12808 2518 12860 2524
rect 11796 2440 11848 2446
rect 11796 2382 11848 2388
rect 12256 2440 12308 2446
rect 12256 2382 12308 2388
rect 12164 2372 12216 2378
rect 12164 2314 12216 2320
rect 11612 2100 11664 2106
rect 11612 2042 11664 2048
rect 10876 1964 10928 1970
rect 10876 1906 10928 1912
rect 10324 1896 10376 1902
rect 10324 1838 10376 1844
rect 9220 1760 9272 1766
rect 9220 1702 9272 1708
rect 9232 1426 9260 1702
rect 9310 1660 9618 1680
rect 9310 1658 9316 1660
rect 9372 1658 9396 1660
rect 9452 1658 9476 1660
rect 9532 1658 9556 1660
rect 9612 1658 9618 1660
rect 9372 1606 9374 1658
rect 9554 1606 9556 1658
rect 9310 1604 9316 1606
rect 9372 1604 9396 1606
rect 9452 1604 9476 1606
rect 9532 1604 9556 1606
rect 9612 1604 9618 1606
rect 9310 1584 9618 1604
rect 9220 1420 9272 1426
rect 9220 1362 9272 1368
rect 10140 1420 10192 1426
rect 10140 1362 10192 1368
rect 9128 1352 9180 1358
rect 9128 1294 9180 1300
rect 10152 1018 10180 1362
rect 10336 1290 10364 1838
rect 10888 1562 10916 1906
rect 11336 1896 11388 1902
rect 11336 1838 11388 1844
rect 10876 1556 10928 1562
rect 10876 1498 10928 1504
rect 11348 1426 11376 1838
rect 11336 1420 11388 1426
rect 11336 1362 11388 1368
rect 10324 1284 10376 1290
rect 10324 1226 10376 1232
rect 10784 1284 10836 1290
rect 10784 1226 10836 1232
rect 11060 1284 11112 1290
rect 11112 1244 11284 1272
rect 11060 1226 11112 1232
rect 10140 1012 10192 1018
rect 10140 954 10192 960
rect 9036 944 9088 950
rect 9036 886 9088 892
rect 10336 814 10364 1226
rect 10796 950 10824 1226
rect 10860 1116 11168 1136
rect 10860 1114 10866 1116
rect 10922 1114 10946 1116
rect 11002 1114 11026 1116
rect 11082 1114 11106 1116
rect 11162 1114 11168 1116
rect 10922 1062 10924 1114
rect 11104 1062 11106 1114
rect 10860 1060 10866 1062
rect 10922 1060 10946 1062
rect 11002 1060 11026 1062
rect 11082 1060 11106 1062
rect 11162 1060 11168 1062
rect 10860 1040 11168 1060
rect 11256 1018 11284 1244
rect 11244 1012 11296 1018
rect 11244 954 11296 960
rect 10784 944 10836 950
rect 10784 886 10836 892
rect 10324 808 10376 814
rect 10376 756 10548 762
rect 10324 750 10548 756
rect 10336 734 10548 750
rect 10520 678 10548 734
rect 9128 672 9180 678
rect 9128 614 9180 620
rect 10508 672 10560 678
rect 10508 614 10560 620
rect 8668 400 8720 406
rect 8668 342 8720 348
rect 9140 338 9168 614
rect 9310 572 9618 592
rect 9310 570 9316 572
rect 9372 570 9396 572
rect 9452 570 9476 572
rect 9532 570 9556 572
rect 9612 570 9618 572
rect 9372 518 9374 570
rect 9554 518 9556 570
rect 9310 516 9316 518
rect 9372 516 9396 518
rect 9452 516 9476 518
rect 9532 516 9556 518
rect 9612 516 9618 518
rect 9310 496 9618 516
rect 10796 338 10824 886
rect 10876 876 10928 882
rect 10876 818 10928 824
rect 11060 876 11112 882
rect 11060 818 11112 824
rect 10888 474 10916 818
rect 10968 808 11020 814
rect 10968 750 11020 756
rect 10876 468 10928 474
rect 10876 410 10928 416
rect 9128 332 9180 338
rect 9128 274 9180 280
rect 10784 332 10836 338
rect 10784 274 10836 280
rect 8576 264 8628 270
rect 8576 206 8628 212
rect 10980 202 11008 750
rect 11072 746 11100 818
rect 11348 746 11376 1362
rect 12176 882 12204 2314
rect 12268 2106 12296 2382
rect 12716 2304 12768 2310
rect 12716 2246 12768 2252
rect 12728 2106 12756 2246
rect 12256 2100 12308 2106
rect 12256 2042 12308 2048
rect 12716 2100 12768 2106
rect 12716 2042 12768 2048
rect 12912 1970 12940 2926
rect 12900 1964 12952 1970
rect 12900 1906 12952 1912
rect 12992 1964 13044 1970
rect 12992 1906 13044 1912
rect 12410 1660 12718 1680
rect 12410 1658 12416 1660
rect 12472 1658 12496 1660
rect 12552 1658 12576 1660
rect 12632 1658 12656 1660
rect 12712 1658 12718 1660
rect 12472 1606 12474 1658
rect 12654 1606 12656 1658
rect 12410 1604 12416 1606
rect 12472 1604 12496 1606
rect 12552 1604 12576 1606
rect 12632 1604 12656 1606
rect 12712 1604 12718 1606
rect 12410 1584 12718 1604
rect 12164 876 12216 882
rect 12164 818 12216 824
rect 12716 876 12768 882
rect 12912 864 12940 1906
rect 13004 1358 13032 1906
rect 12992 1352 13044 1358
rect 12992 1294 13044 1300
rect 12768 836 12940 864
rect 12716 818 12768 824
rect 12992 808 13044 814
rect 12992 750 13044 756
rect 11060 740 11112 746
rect 11060 682 11112 688
rect 11336 740 11388 746
rect 11336 682 11388 688
rect 11072 270 11100 682
rect 12410 572 12718 592
rect 12410 570 12416 572
rect 12472 570 12496 572
rect 12552 570 12576 572
rect 12632 570 12656 572
rect 12712 570 12718 572
rect 12472 518 12474 570
rect 12654 518 12656 570
rect 12410 516 12416 518
rect 12472 516 12496 518
rect 12552 516 12576 518
rect 12632 516 12656 518
rect 12712 516 12718 518
rect 12410 496 12718 516
rect 13004 474 13032 750
rect 12992 468 13044 474
rect 12992 410 13044 416
rect 12992 332 13044 338
rect 13096 320 13124 3470
rect 13372 3398 13400 4082
rect 14188 3936 14240 3942
rect 14188 3878 14240 3884
rect 14200 3534 14228 3878
rect 14568 3602 14596 4626
rect 15120 4554 15148 5238
rect 15510 4924 15818 4944
rect 15510 4922 15516 4924
rect 15572 4922 15596 4924
rect 15652 4922 15676 4924
rect 15732 4922 15756 4924
rect 15812 4922 15818 4924
rect 15572 4870 15574 4922
rect 15754 4870 15756 4922
rect 15510 4868 15516 4870
rect 15572 4868 15596 4870
rect 15652 4868 15676 4870
rect 15732 4868 15756 4870
rect 15812 4868 15818 4870
rect 15510 4848 15818 4868
rect 16316 4554 16344 5238
rect 17684 5024 17736 5030
rect 17684 4966 17736 4972
rect 17696 4690 17724 4966
rect 17684 4684 17736 4690
rect 17684 4626 17736 4632
rect 17972 4622 18000 5238
rect 18248 5166 18276 5510
rect 18524 5273 18552 5646
rect 18510 5264 18566 5273
rect 18510 5199 18566 5208
rect 18236 5160 18288 5166
rect 18236 5102 18288 5108
rect 17960 4616 18012 4622
rect 17960 4558 18012 4564
rect 18512 4616 18564 4622
rect 18512 4558 18564 4564
rect 15108 4548 15160 4554
rect 15108 4490 15160 4496
rect 15936 4548 15988 4554
rect 15936 4490 15988 4496
rect 16304 4548 16356 4554
rect 16304 4490 16356 4496
rect 14648 3936 14700 3942
rect 14648 3878 14700 3884
rect 14556 3596 14608 3602
rect 14556 3538 14608 3544
rect 14188 3528 14240 3534
rect 14188 3470 14240 3476
rect 13820 3460 13872 3466
rect 13820 3402 13872 3408
rect 13360 3392 13412 3398
rect 13360 3334 13412 3340
rect 13372 3126 13400 3334
rect 13360 3120 13412 3126
rect 13360 3062 13412 3068
rect 13832 3058 13860 3402
rect 13960 3292 14268 3312
rect 13960 3290 13966 3292
rect 14022 3290 14046 3292
rect 14102 3290 14126 3292
rect 14182 3290 14206 3292
rect 14262 3290 14268 3292
rect 14022 3238 14024 3290
rect 14204 3238 14206 3290
rect 13960 3236 13966 3238
rect 14022 3236 14046 3238
rect 14102 3236 14126 3238
rect 14182 3236 14206 3238
rect 14262 3236 14268 3238
rect 13960 3216 14268 3236
rect 14568 3194 14596 3538
rect 14556 3188 14608 3194
rect 14556 3130 14608 3136
rect 13820 3052 13872 3058
rect 13820 2994 13872 3000
rect 13176 2372 13228 2378
rect 13176 2314 13228 2320
rect 13188 2106 13216 2314
rect 13176 2100 13228 2106
rect 13176 2042 13228 2048
rect 13832 2038 13860 2994
rect 14660 2990 14688 3878
rect 15120 3534 15148 4490
rect 15948 4282 15976 4490
rect 15936 4276 15988 4282
rect 15936 4218 15988 4224
rect 15200 4140 15252 4146
rect 15200 4082 15252 4088
rect 15108 3528 15160 3534
rect 15108 3470 15160 3476
rect 14648 2984 14700 2990
rect 14648 2926 14700 2932
rect 14556 2440 14608 2446
rect 14556 2382 14608 2388
rect 14372 2304 14424 2310
rect 14372 2246 14424 2252
rect 13960 2204 14268 2224
rect 13960 2202 13966 2204
rect 14022 2202 14046 2204
rect 14102 2202 14126 2204
rect 14182 2202 14206 2204
rect 14262 2202 14268 2204
rect 14022 2150 14024 2202
rect 14204 2150 14206 2202
rect 13960 2148 13966 2150
rect 14022 2148 14046 2150
rect 14102 2148 14126 2150
rect 14182 2148 14206 2150
rect 14262 2148 14268 2150
rect 13960 2128 14268 2148
rect 13820 2032 13872 2038
rect 13820 1974 13872 1980
rect 13832 1358 13860 1974
rect 14384 1970 14412 2246
rect 14568 2106 14596 2382
rect 15212 2378 15240 4082
rect 15510 3836 15818 3856
rect 15510 3834 15516 3836
rect 15572 3834 15596 3836
rect 15652 3834 15676 3836
rect 15732 3834 15756 3836
rect 15812 3834 15818 3836
rect 15572 3782 15574 3834
rect 15754 3782 15756 3834
rect 15510 3780 15516 3782
rect 15572 3780 15596 3782
rect 15652 3780 15676 3782
rect 15732 3780 15756 3782
rect 15812 3780 15818 3782
rect 15510 3760 15818 3780
rect 15844 3596 15896 3602
rect 15844 3538 15896 3544
rect 15384 3188 15436 3194
rect 15384 3130 15436 3136
rect 15396 2514 15424 3130
rect 15856 2990 15884 3538
rect 16212 3528 16264 3534
rect 16212 3470 16264 3476
rect 16224 3194 16252 3470
rect 16316 3398 16344 4490
rect 17408 4480 17460 4486
rect 17408 4422 17460 4428
rect 17060 4380 17368 4400
rect 17060 4378 17066 4380
rect 17122 4378 17146 4380
rect 17202 4378 17226 4380
rect 17282 4378 17306 4380
rect 17362 4378 17368 4380
rect 17122 4326 17124 4378
rect 17304 4326 17306 4378
rect 17060 4324 17066 4326
rect 17122 4324 17146 4326
rect 17202 4324 17226 4326
rect 17282 4324 17306 4326
rect 17362 4324 17368 4326
rect 17060 4304 17368 4324
rect 16948 3936 17000 3942
rect 16948 3878 17000 3884
rect 16304 3392 16356 3398
rect 16304 3334 16356 3340
rect 16212 3188 16264 3194
rect 16212 3130 16264 3136
rect 16316 3108 16344 3334
rect 16396 3120 16448 3126
rect 16316 3080 16396 3108
rect 16396 3062 16448 3068
rect 15844 2984 15896 2990
rect 15844 2926 15896 2932
rect 15510 2748 15818 2768
rect 15510 2746 15516 2748
rect 15572 2746 15596 2748
rect 15652 2746 15676 2748
rect 15732 2746 15756 2748
rect 15812 2746 15818 2748
rect 15572 2694 15574 2746
rect 15754 2694 15756 2746
rect 15510 2692 15516 2694
rect 15572 2692 15596 2694
rect 15652 2692 15676 2694
rect 15732 2692 15756 2694
rect 15812 2692 15818 2694
rect 15510 2672 15818 2692
rect 15384 2508 15436 2514
rect 15384 2450 15436 2456
rect 15752 2508 15804 2514
rect 15752 2450 15804 2456
rect 15568 2440 15620 2446
rect 15764 2394 15792 2450
rect 15568 2382 15620 2388
rect 15200 2372 15252 2378
rect 15200 2314 15252 2320
rect 15384 2372 15436 2378
rect 15384 2314 15436 2320
rect 14556 2100 14608 2106
rect 14556 2042 14608 2048
rect 14372 1964 14424 1970
rect 14372 1906 14424 1912
rect 15212 1902 15240 2314
rect 15396 2038 15424 2314
rect 15580 2106 15608 2382
rect 15672 2366 15792 2394
rect 15568 2100 15620 2106
rect 15568 2042 15620 2048
rect 15384 2032 15436 2038
rect 15384 1974 15436 1980
rect 15200 1896 15252 1902
rect 15200 1838 15252 1844
rect 15672 1834 15700 2366
rect 15752 2304 15804 2310
rect 15752 2246 15804 2252
rect 15764 1850 15792 2246
rect 15856 2038 15884 2926
rect 16408 2378 16436 3062
rect 16488 2576 16540 2582
rect 16488 2518 16540 2524
rect 16304 2372 16356 2378
rect 16304 2314 16356 2320
rect 16396 2372 16448 2378
rect 16396 2314 16448 2320
rect 16028 2304 16080 2310
rect 16028 2246 16080 2252
rect 16040 2038 16068 2246
rect 15844 2032 15896 2038
rect 15844 1974 15896 1980
rect 16028 2032 16080 2038
rect 16028 1974 16080 1980
rect 15660 1828 15712 1834
rect 15764 1822 15884 1850
rect 15660 1770 15712 1776
rect 15510 1660 15818 1680
rect 15510 1658 15516 1660
rect 15572 1658 15596 1660
rect 15652 1658 15676 1660
rect 15732 1658 15756 1660
rect 15812 1658 15818 1660
rect 15572 1606 15574 1658
rect 15754 1606 15756 1658
rect 15510 1604 15516 1606
rect 15572 1604 15596 1606
rect 15652 1604 15676 1606
rect 15732 1604 15756 1606
rect 15812 1604 15818 1606
rect 15510 1584 15818 1604
rect 13820 1352 13872 1358
rect 13820 1294 13872 1300
rect 13636 1216 13688 1222
rect 13636 1158 13688 1164
rect 13648 1018 13676 1158
rect 13832 1018 13860 1294
rect 14464 1284 14516 1290
rect 14464 1226 14516 1232
rect 14924 1284 14976 1290
rect 14924 1226 14976 1232
rect 14372 1216 14424 1222
rect 14372 1158 14424 1164
rect 13960 1116 14268 1136
rect 13960 1114 13966 1116
rect 14022 1114 14046 1116
rect 14102 1114 14126 1116
rect 14182 1114 14206 1116
rect 14262 1114 14268 1116
rect 14022 1062 14024 1114
rect 14204 1062 14206 1114
rect 13960 1060 13966 1062
rect 14022 1060 14046 1062
rect 14102 1060 14126 1062
rect 14182 1060 14206 1062
rect 14262 1060 14268 1062
rect 13960 1040 14268 1060
rect 14384 1018 14412 1158
rect 13636 1012 13688 1018
rect 13636 954 13688 960
rect 13820 1012 13872 1018
rect 13820 954 13872 960
rect 14372 1012 14424 1018
rect 14372 954 14424 960
rect 14476 814 14504 1226
rect 14648 944 14700 950
rect 14648 886 14700 892
rect 14464 808 14516 814
rect 14464 750 14516 756
rect 13176 672 13228 678
rect 13176 614 13228 620
rect 13044 292 13124 320
rect 12992 274 13044 280
rect 11060 264 11112 270
rect 11060 206 11112 212
rect 13188 202 13216 614
rect 14660 474 14688 886
rect 14648 468 14700 474
rect 14648 410 14700 416
rect 14936 202 14964 1226
rect 15856 746 15884 1822
rect 16316 1290 16344 2314
rect 16408 2038 16436 2314
rect 16396 2032 16448 2038
rect 16396 1974 16448 1980
rect 16212 1284 16264 1290
rect 16212 1226 16264 1232
rect 16304 1284 16356 1290
rect 16304 1226 16356 1232
rect 16224 1018 16252 1226
rect 16408 1222 16436 1974
rect 16500 1426 16528 2518
rect 16960 1766 16988 3878
rect 17060 3292 17368 3312
rect 17060 3290 17066 3292
rect 17122 3290 17146 3292
rect 17202 3290 17226 3292
rect 17282 3290 17306 3292
rect 17362 3290 17368 3292
rect 17122 3238 17124 3290
rect 17304 3238 17306 3290
rect 17060 3236 17066 3238
rect 17122 3236 17146 3238
rect 17202 3236 17226 3238
rect 17282 3236 17306 3238
rect 17362 3236 17368 3238
rect 17060 3216 17368 3236
rect 17420 2990 17448 4422
rect 17592 4004 17644 4010
rect 17592 3946 17644 3952
rect 17604 3602 17632 3946
rect 17592 3596 17644 3602
rect 17592 3538 17644 3544
rect 17604 2990 17632 3538
rect 17972 3058 18000 4558
rect 18236 4548 18288 4554
rect 18236 4490 18288 4496
rect 18144 4140 18196 4146
rect 18144 4082 18196 4088
rect 18052 3936 18104 3942
rect 18052 3878 18104 3884
rect 17960 3052 18012 3058
rect 17960 2994 18012 3000
rect 17408 2984 17460 2990
rect 17408 2926 17460 2932
rect 17592 2984 17644 2990
rect 17592 2926 17644 2932
rect 17972 2514 18000 2994
rect 17960 2508 18012 2514
rect 17960 2450 18012 2456
rect 17408 2372 17460 2378
rect 17408 2314 17460 2320
rect 17060 2204 17368 2224
rect 17060 2202 17066 2204
rect 17122 2202 17146 2204
rect 17202 2202 17226 2204
rect 17282 2202 17306 2204
rect 17362 2202 17368 2204
rect 17122 2150 17124 2202
rect 17304 2150 17306 2202
rect 17060 2148 17066 2150
rect 17122 2148 17146 2150
rect 17202 2148 17226 2150
rect 17282 2148 17306 2150
rect 17362 2148 17368 2150
rect 17060 2128 17368 2148
rect 17420 2106 17448 2314
rect 17408 2100 17460 2106
rect 17408 2042 17460 2048
rect 16948 1760 17000 1766
rect 16948 1702 17000 1708
rect 16488 1420 16540 1426
rect 16488 1362 16540 1368
rect 16396 1216 16448 1222
rect 16396 1158 16448 1164
rect 16212 1012 16264 1018
rect 16212 954 16264 960
rect 15844 740 15896 746
rect 15844 682 15896 688
rect 15510 572 15818 592
rect 15510 570 15516 572
rect 15572 570 15596 572
rect 15652 570 15676 572
rect 15732 570 15756 572
rect 15812 570 15818 572
rect 15572 518 15574 570
rect 15754 518 15756 570
rect 15510 516 15516 518
rect 15572 516 15596 518
rect 15652 516 15676 518
rect 15732 516 15756 518
rect 15812 516 15818 518
rect 15510 496 15818 516
rect 16500 474 16528 1362
rect 17960 1216 18012 1222
rect 17960 1158 18012 1164
rect 17060 1116 17368 1136
rect 17060 1114 17066 1116
rect 17122 1114 17146 1116
rect 17202 1114 17226 1116
rect 17282 1114 17306 1116
rect 17362 1114 17368 1116
rect 17122 1062 17124 1114
rect 17304 1062 17306 1114
rect 17060 1060 17066 1062
rect 17122 1060 17146 1062
rect 17202 1060 17226 1062
rect 17282 1060 17306 1062
rect 17362 1060 17368 1062
rect 17060 1040 17368 1060
rect 17972 950 18000 1158
rect 17960 944 18012 950
rect 17960 886 18012 892
rect 18064 882 18092 3878
rect 18156 3670 18184 4082
rect 18144 3664 18196 3670
rect 18144 3606 18196 3612
rect 17776 876 17828 882
rect 17776 818 17828 824
rect 18052 876 18104 882
rect 18052 818 18104 824
rect 17788 746 17816 818
rect 18156 762 18184 3606
rect 18248 1358 18276 4490
rect 18328 4072 18380 4078
rect 18328 4014 18380 4020
rect 18340 3534 18368 4014
rect 18524 3777 18552 4558
rect 18510 3768 18566 3777
rect 18510 3703 18566 3712
rect 18328 3528 18380 3534
rect 18328 3470 18380 3476
rect 18340 3194 18368 3470
rect 18328 3188 18380 3194
rect 18328 3130 18380 3136
rect 18512 2440 18564 2446
rect 18512 2382 18564 2388
rect 18524 2281 18552 2382
rect 18510 2272 18566 2281
rect 18510 2207 18566 2216
rect 18236 1352 18288 1358
rect 18236 1294 18288 1300
rect 18328 1352 18380 1358
rect 18328 1294 18380 1300
rect 17776 740 17828 746
rect 17776 682 17828 688
rect 17972 734 18184 762
rect 17788 474 17816 682
rect 17972 678 18000 734
rect 17960 672 18012 678
rect 17960 614 18012 620
rect 16488 468 16540 474
rect 16488 410 16540 416
rect 17776 468 17828 474
rect 17776 410 17828 416
rect 17972 202 18000 614
rect 18340 474 18368 1294
rect 18510 776 18566 785
rect 18510 711 18566 720
rect 18328 468 18380 474
rect 18328 410 18380 416
rect 18524 270 18552 711
rect 18512 264 18564 270
rect 18512 206 18564 212
rect 8208 196 8260 202
rect 8208 138 8260 144
rect 10968 196 11020 202
rect 10968 138 11020 144
rect 13176 196 13228 202
rect 13176 138 13228 144
rect 14924 196 14976 202
rect 14924 138 14976 144
rect 17960 196 18012 202
rect 17960 138 18012 144
rect 2688 128 2740 134
rect 2688 70 2740 76
rect 4660 28 4968 48
rect 4660 26 4666 28
rect 4722 26 4746 28
rect 4802 26 4826 28
rect 4882 26 4906 28
rect 4962 26 4968 28
rect 4722 -26 4724 26
rect 4904 -26 4906 26
rect 4660 -28 4666 -26
rect 4722 -28 4746 -26
rect 4802 -28 4826 -26
rect 4882 -28 4906 -26
rect 4962 -28 4968 -26
rect 4660 -48 4968 -28
rect 7760 28 8068 48
rect 7760 26 7766 28
rect 7822 26 7846 28
rect 7902 26 7926 28
rect 7982 26 8006 28
rect 8062 26 8068 28
rect 7822 -26 7824 26
rect 8004 -26 8006 26
rect 7760 -28 7766 -26
rect 7822 -28 7846 -26
rect 7902 -28 7926 -26
rect 7982 -28 8006 -26
rect 8062 -28 8068 -26
rect 7760 -48 8068 -28
rect 10860 28 11168 48
rect 10860 26 10866 28
rect 10922 26 10946 28
rect 11002 26 11026 28
rect 11082 26 11106 28
rect 11162 26 11168 28
rect 10922 -26 10924 26
rect 11104 -26 11106 26
rect 10860 -28 10866 -26
rect 10922 -28 10946 -26
rect 11002 -28 11026 -26
rect 11082 -28 11106 -26
rect 11162 -28 11168 -26
rect 10860 -48 11168 -28
rect 13960 28 14268 48
rect 13960 26 13966 28
rect 14022 26 14046 28
rect 14102 26 14126 28
rect 14182 26 14206 28
rect 14262 26 14268 28
rect 14022 -26 14024 26
rect 14204 -26 14206 26
rect 13960 -28 13966 -26
rect 14022 -28 14046 -26
rect 14102 -28 14126 -26
rect 14182 -28 14206 -26
rect 14262 -28 14268 -26
rect 13960 -48 14268 -28
rect 17060 28 17368 48
rect 17060 26 17066 28
rect 17122 26 17146 28
rect 17202 26 17226 28
rect 17282 26 17306 28
rect 17362 26 17368 28
rect 17122 -26 17124 26
rect 17304 -26 17306 26
rect 17060 -28 17066 -26
rect 17122 -28 17146 -26
rect 17202 -28 17226 -26
rect 17282 -28 17306 -26
rect 17362 -28 17368 -26
rect 17060 -48 17368 -28
<< via2 >>
rect 3116 10362 3172 10364
rect 3196 10362 3252 10364
rect 3276 10362 3332 10364
rect 3356 10362 3412 10364
rect 3116 10310 3162 10362
rect 3162 10310 3172 10362
rect 3196 10310 3226 10362
rect 3226 10310 3238 10362
rect 3238 10310 3252 10362
rect 3276 10310 3290 10362
rect 3290 10310 3302 10362
rect 3302 10310 3332 10362
rect 3356 10310 3366 10362
rect 3366 10310 3412 10362
rect 3116 10308 3172 10310
rect 3196 10308 3252 10310
rect 3276 10308 3332 10310
rect 3356 10308 3412 10310
rect 3116 9274 3172 9276
rect 3196 9274 3252 9276
rect 3276 9274 3332 9276
rect 3356 9274 3412 9276
rect 3116 9222 3162 9274
rect 3162 9222 3172 9274
rect 3196 9222 3226 9274
rect 3226 9222 3238 9274
rect 3238 9222 3252 9274
rect 3276 9222 3290 9274
rect 3290 9222 3302 9274
rect 3302 9222 3332 9274
rect 3356 9222 3366 9274
rect 3366 9222 3412 9274
rect 3116 9220 3172 9222
rect 3196 9220 3252 9222
rect 3276 9220 3332 9222
rect 3356 9220 3412 9222
rect 3116 8186 3172 8188
rect 3196 8186 3252 8188
rect 3276 8186 3332 8188
rect 3356 8186 3412 8188
rect 3116 8134 3162 8186
rect 3162 8134 3172 8186
rect 3196 8134 3226 8186
rect 3226 8134 3238 8186
rect 3238 8134 3252 8186
rect 3276 8134 3290 8186
rect 3290 8134 3302 8186
rect 3302 8134 3332 8186
rect 3356 8134 3366 8186
rect 3366 8134 3412 8186
rect 3116 8132 3172 8134
rect 3196 8132 3252 8134
rect 3276 8132 3332 8134
rect 3356 8132 3412 8134
rect 3116 7098 3172 7100
rect 3196 7098 3252 7100
rect 3276 7098 3332 7100
rect 3356 7098 3412 7100
rect 3116 7046 3162 7098
rect 3162 7046 3172 7098
rect 3196 7046 3226 7098
rect 3226 7046 3238 7098
rect 3238 7046 3252 7098
rect 3276 7046 3290 7098
rect 3290 7046 3302 7098
rect 3302 7046 3332 7098
rect 3356 7046 3366 7098
rect 3366 7046 3412 7098
rect 3116 7044 3172 7046
rect 3196 7044 3252 7046
rect 3276 7044 3332 7046
rect 3356 7044 3412 7046
rect 3116 6010 3172 6012
rect 3196 6010 3252 6012
rect 3276 6010 3332 6012
rect 3356 6010 3412 6012
rect 3116 5958 3162 6010
rect 3162 5958 3172 6010
rect 3196 5958 3226 6010
rect 3226 5958 3238 6010
rect 3238 5958 3252 6010
rect 3276 5958 3290 6010
rect 3290 5958 3302 6010
rect 3302 5958 3332 6010
rect 3356 5958 3366 6010
rect 3366 5958 3412 6010
rect 3116 5956 3172 5958
rect 3196 5956 3252 5958
rect 3276 5956 3332 5958
rect 3356 5956 3412 5958
rect 4666 10906 4722 10908
rect 4746 10906 4802 10908
rect 4826 10906 4882 10908
rect 4906 10906 4962 10908
rect 4666 10854 4712 10906
rect 4712 10854 4722 10906
rect 4746 10854 4776 10906
rect 4776 10854 4788 10906
rect 4788 10854 4802 10906
rect 4826 10854 4840 10906
rect 4840 10854 4852 10906
rect 4852 10854 4882 10906
rect 4906 10854 4916 10906
rect 4916 10854 4962 10906
rect 4666 10852 4722 10854
rect 4746 10852 4802 10854
rect 4826 10852 4882 10854
rect 4906 10852 4962 10854
rect 7766 10906 7822 10908
rect 7846 10906 7902 10908
rect 7926 10906 7982 10908
rect 8006 10906 8062 10908
rect 7766 10854 7812 10906
rect 7812 10854 7822 10906
rect 7846 10854 7876 10906
rect 7876 10854 7888 10906
rect 7888 10854 7902 10906
rect 7926 10854 7940 10906
rect 7940 10854 7952 10906
rect 7952 10854 7982 10906
rect 8006 10854 8016 10906
rect 8016 10854 8062 10906
rect 7766 10852 7822 10854
rect 7846 10852 7902 10854
rect 7926 10852 7982 10854
rect 8006 10852 8062 10854
rect 10866 10906 10922 10908
rect 10946 10906 11002 10908
rect 11026 10906 11082 10908
rect 11106 10906 11162 10908
rect 10866 10854 10912 10906
rect 10912 10854 10922 10906
rect 10946 10854 10976 10906
rect 10976 10854 10988 10906
rect 10988 10854 11002 10906
rect 11026 10854 11040 10906
rect 11040 10854 11052 10906
rect 11052 10854 11082 10906
rect 11106 10854 11116 10906
rect 11116 10854 11162 10906
rect 10866 10852 10922 10854
rect 10946 10852 11002 10854
rect 11026 10852 11082 10854
rect 11106 10852 11162 10854
rect 4666 9818 4722 9820
rect 4746 9818 4802 9820
rect 4826 9818 4882 9820
rect 4906 9818 4962 9820
rect 4666 9766 4712 9818
rect 4712 9766 4722 9818
rect 4746 9766 4776 9818
rect 4776 9766 4788 9818
rect 4788 9766 4802 9818
rect 4826 9766 4840 9818
rect 4840 9766 4852 9818
rect 4852 9766 4882 9818
rect 4906 9766 4916 9818
rect 4916 9766 4962 9818
rect 4666 9764 4722 9766
rect 4746 9764 4802 9766
rect 4826 9764 4882 9766
rect 4906 9764 4962 9766
rect 6216 10362 6272 10364
rect 6296 10362 6352 10364
rect 6376 10362 6432 10364
rect 6456 10362 6512 10364
rect 6216 10310 6262 10362
rect 6262 10310 6272 10362
rect 6296 10310 6326 10362
rect 6326 10310 6338 10362
rect 6338 10310 6352 10362
rect 6376 10310 6390 10362
rect 6390 10310 6402 10362
rect 6402 10310 6432 10362
rect 6456 10310 6466 10362
rect 6466 10310 6512 10362
rect 6216 10308 6272 10310
rect 6296 10308 6352 10310
rect 6376 10308 6432 10310
rect 6456 10308 6512 10310
rect 4666 8730 4722 8732
rect 4746 8730 4802 8732
rect 4826 8730 4882 8732
rect 4906 8730 4962 8732
rect 4666 8678 4712 8730
rect 4712 8678 4722 8730
rect 4746 8678 4776 8730
rect 4776 8678 4788 8730
rect 4788 8678 4802 8730
rect 4826 8678 4840 8730
rect 4840 8678 4852 8730
rect 4852 8678 4882 8730
rect 4906 8678 4916 8730
rect 4916 8678 4962 8730
rect 4666 8676 4722 8678
rect 4746 8676 4802 8678
rect 4826 8676 4882 8678
rect 4906 8676 4962 8678
rect 6216 9274 6272 9276
rect 6296 9274 6352 9276
rect 6376 9274 6432 9276
rect 6456 9274 6512 9276
rect 6216 9222 6262 9274
rect 6262 9222 6272 9274
rect 6296 9222 6326 9274
rect 6326 9222 6338 9274
rect 6338 9222 6352 9274
rect 6376 9222 6390 9274
rect 6390 9222 6402 9274
rect 6402 9222 6432 9274
rect 6456 9222 6466 9274
rect 6466 9222 6512 9274
rect 6216 9220 6272 9222
rect 6296 9220 6352 9222
rect 6376 9220 6432 9222
rect 6456 9220 6512 9222
rect 4666 7642 4722 7644
rect 4746 7642 4802 7644
rect 4826 7642 4882 7644
rect 4906 7642 4962 7644
rect 4666 7590 4712 7642
rect 4712 7590 4722 7642
rect 4746 7590 4776 7642
rect 4776 7590 4788 7642
rect 4788 7590 4802 7642
rect 4826 7590 4840 7642
rect 4840 7590 4852 7642
rect 4852 7590 4882 7642
rect 4906 7590 4916 7642
rect 4916 7590 4962 7642
rect 4666 7588 4722 7590
rect 4746 7588 4802 7590
rect 4826 7588 4882 7590
rect 4906 7588 4962 7590
rect 4666 6554 4722 6556
rect 4746 6554 4802 6556
rect 4826 6554 4882 6556
rect 4906 6554 4962 6556
rect 4666 6502 4712 6554
rect 4712 6502 4722 6554
rect 4746 6502 4776 6554
rect 4776 6502 4788 6554
rect 4788 6502 4802 6554
rect 4826 6502 4840 6554
rect 4840 6502 4852 6554
rect 4852 6502 4882 6554
rect 4906 6502 4916 6554
rect 4916 6502 4962 6554
rect 4666 6500 4722 6502
rect 4746 6500 4802 6502
rect 4826 6500 4882 6502
rect 4906 6500 4962 6502
rect 6216 8186 6272 8188
rect 6296 8186 6352 8188
rect 6376 8186 6432 8188
rect 6456 8186 6512 8188
rect 6216 8134 6262 8186
rect 6262 8134 6272 8186
rect 6296 8134 6326 8186
rect 6326 8134 6338 8186
rect 6338 8134 6352 8186
rect 6376 8134 6390 8186
rect 6390 8134 6402 8186
rect 6402 8134 6432 8186
rect 6456 8134 6466 8186
rect 6466 8134 6512 8186
rect 6216 8132 6272 8134
rect 6296 8132 6352 8134
rect 6376 8132 6432 8134
rect 6456 8132 6512 8134
rect 6216 7098 6272 7100
rect 6296 7098 6352 7100
rect 6376 7098 6432 7100
rect 6456 7098 6512 7100
rect 6216 7046 6262 7098
rect 6262 7046 6272 7098
rect 6296 7046 6326 7098
rect 6326 7046 6338 7098
rect 6338 7046 6352 7098
rect 6376 7046 6390 7098
rect 6390 7046 6402 7098
rect 6402 7046 6432 7098
rect 6456 7046 6466 7098
rect 6466 7046 6512 7098
rect 6216 7044 6272 7046
rect 6296 7044 6352 7046
rect 6376 7044 6432 7046
rect 6456 7044 6512 7046
rect 6216 6010 6272 6012
rect 6296 6010 6352 6012
rect 6376 6010 6432 6012
rect 6456 6010 6512 6012
rect 6216 5958 6262 6010
rect 6262 5958 6272 6010
rect 6296 5958 6326 6010
rect 6326 5958 6338 6010
rect 6338 5958 6352 6010
rect 6376 5958 6390 6010
rect 6390 5958 6402 6010
rect 6402 5958 6432 6010
rect 6456 5958 6466 6010
rect 6466 5958 6512 6010
rect 6216 5956 6272 5958
rect 6296 5956 6352 5958
rect 6376 5956 6432 5958
rect 6456 5956 6512 5958
rect 4666 5466 4722 5468
rect 4746 5466 4802 5468
rect 4826 5466 4882 5468
rect 4906 5466 4962 5468
rect 4666 5414 4712 5466
rect 4712 5414 4722 5466
rect 4746 5414 4776 5466
rect 4776 5414 4788 5466
rect 4788 5414 4802 5466
rect 4826 5414 4840 5466
rect 4840 5414 4852 5466
rect 4852 5414 4882 5466
rect 4906 5414 4916 5466
rect 4916 5414 4962 5466
rect 4666 5412 4722 5414
rect 4746 5412 4802 5414
rect 4826 5412 4882 5414
rect 4906 5412 4962 5414
rect 7470 5244 7472 5264
rect 7472 5244 7524 5264
rect 7524 5244 7526 5264
rect 7470 5208 7526 5244
rect 3116 4922 3172 4924
rect 3196 4922 3252 4924
rect 3276 4922 3332 4924
rect 3356 4922 3412 4924
rect 3116 4870 3162 4922
rect 3162 4870 3172 4922
rect 3196 4870 3226 4922
rect 3226 4870 3238 4922
rect 3238 4870 3252 4922
rect 3276 4870 3290 4922
rect 3290 4870 3302 4922
rect 3302 4870 3332 4922
rect 3356 4870 3366 4922
rect 3366 4870 3412 4922
rect 3116 4868 3172 4870
rect 3196 4868 3252 4870
rect 3276 4868 3332 4870
rect 3356 4868 3412 4870
rect 6216 4922 6272 4924
rect 6296 4922 6352 4924
rect 6376 4922 6432 4924
rect 6456 4922 6512 4924
rect 6216 4870 6262 4922
rect 6262 4870 6272 4922
rect 6296 4870 6326 4922
rect 6326 4870 6338 4922
rect 6338 4870 6352 4922
rect 6376 4870 6390 4922
rect 6390 4870 6402 4922
rect 6402 4870 6432 4922
rect 6456 4870 6466 4922
rect 6466 4870 6512 4922
rect 6216 4868 6272 4870
rect 6296 4868 6352 4870
rect 6376 4868 6432 4870
rect 6456 4868 6512 4870
rect 4666 4378 4722 4380
rect 4746 4378 4802 4380
rect 4826 4378 4882 4380
rect 4906 4378 4962 4380
rect 4666 4326 4712 4378
rect 4712 4326 4722 4378
rect 4746 4326 4776 4378
rect 4776 4326 4788 4378
rect 4788 4326 4802 4378
rect 4826 4326 4840 4378
rect 4840 4326 4852 4378
rect 4852 4326 4882 4378
rect 4906 4326 4916 4378
rect 4916 4326 4962 4378
rect 4666 4324 4722 4326
rect 4746 4324 4802 4326
rect 4826 4324 4882 4326
rect 4906 4324 4962 4326
rect 3116 3834 3172 3836
rect 3196 3834 3252 3836
rect 3276 3834 3332 3836
rect 3356 3834 3412 3836
rect 3116 3782 3162 3834
rect 3162 3782 3172 3834
rect 3196 3782 3226 3834
rect 3226 3782 3238 3834
rect 3238 3782 3252 3834
rect 3276 3782 3290 3834
rect 3290 3782 3302 3834
rect 3302 3782 3332 3834
rect 3356 3782 3366 3834
rect 3366 3782 3412 3834
rect 3116 3780 3172 3782
rect 3196 3780 3252 3782
rect 3276 3780 3332 3782
rect 3356 3780 3412 3782
rect 3882 3476 3884 3496
rect 3884 3476 3936 3496
rect 3936 3476 3938 3496
rect 3882 3440 3938 3476
rect 4066 3440 4122 3496
rect 4666 3290 4722 3292
rect 4746 3290 4802 3292
rect 4826 3290 4882 3292
rect 4906 3290 4962 3292
rect 4666 3238 4712 3290
rect 4712 3238 4722 3290
rect 4746 3238 4776 3290
rect 4776 3238 4788 3290
rect 4788 3238 4802 3290
rect 4826 3238 4840 3290
rect 4840 3238 4852 3290
rect 4852 3238 4882 3290
rect 4906 3238 4916 3290
rect 4916 3238 4962 3290
rect 4666 3236 4722 3238
rect 4746 3236 4802 3238
rect 4826 3236 4882 3238
rect 4906 3236 4962 3238
rect 4802 3052 4858 3088
rect 9316 10362 9372 10364
rect 9396 10362 9452 10364
rect 9476 10362 9532 10364
rect 9556 10362 9612 10364
rect 9316 10310 9362 10362
rect 9362 10310 9372 10362
rect 9396 10310 9426 10362
rect 9426 10310 9438 10362
rect 9438 10310 9452 10362
rect 9476 10310 9490 10362
rect 9490 10310 9502 10362
rect 9502 10310 9532 10362
rect 9556 10310 9566 10362
rect 9566 10310 9612 10362
rect 9316 10308 9372 10310
rect 9396 10308 9452 10310
rect 9476 10308 9532 10310
rect 9556 10308 9612 10310
rect 7766 9818 7822 9820
rect 7846 9818 7902 9820
rect 7926 9818 7982 9820
rect 8006 9818 8062 9820
rect 7766 9766 7812 9818
rect 7812 9766 7822 9818
rect 7846 9766 7876 9818
rect 7876 9766 7888 9818
rect 7888 9766 7902 9818
rect 7926 9766 7940 9818
rect 7940 9766 7952 9818
rect 7952 9766 7982 9818
rect 8006 9766 8016 9818
rect 8016 9766 8062 9818
rect 7766 9764 7822 9766
rect 7846 9764 7902 9766
rect 7926 9764 7982 9766
rect 8006 9764 8062 9766
rect 7766 8730 7822 8732
rect 7846 8730 7902 8732
rect 7926 8730 7982 8732
rect 8006 8730 8062 8732
rect 7766 8678 7812 8730
rect 7812 8678 7822 8730
rect 7846 8678 7876 8730
rect 7876 8678 7888 8730
rect 7888 8678 7902 8730
rect 7926 8678 7940 8730
rect 7940 8678 7952 8730
rect 7952 8678 7982 8730
rect 8006 8678 8016 8730
rect 8016 8678 8062 8730
rect 7766 8676 7822 8678
rect 7846 8676 7902 8678
rect 7926 8676 7982 8678
rect 8006 8676 8062 8678
rect 7766 7642 7822 7644
rect 7846 7642 7902 7644
rect 7926 7642 7982 7644
rect 8006 7642 8062 7644
rect 7766 7590 7812 7642
rect 7812 7590 7822 7642
rect 7846 7590 7876 7642
rect 7876 7590 7888 7642
rect 7888 7590 7902 7642
rect 7926 7590 7940 7642
rect 7940 7590 7952 7642
rect 7952 7590 7982 7642
rect 8006 7590 8016 7642
rect 8016 7590 8062 7642
rect 7766 7588 7822 7590
rect 7846 7588 7902 7590
rect 7926 7588 7982 7590
rect 8006 7588 8062 7590
rect 7766 6554 7822 6556
rect 7846 6554 7902 6556
rect 7926 6554 7982 6556
rect 8006 6554 8062 6556
rect 7766 6502 7812 6554
rect 7812 6502 7822 6554
rect 7846 6502 7876 6554
rect 7876 6502 7888 6554
rect 7888 6502 7902 6554
rect 7926 6502 7940 6554
rect 7940 6502 7952 6554
rect 7952 6502 7982 6554
rect 8006 6502 8016 6554
rect 8016 6502 8062 6554
rect 7766 6500 7822 6502
rect 7846 6500 7902 6502
rect 7926 6500 7982 6502
rect 8006 6500 8062 6502
rect 7766 5466 7822 5468
rect 7846 5466 7902 5468
rect 7926 5466 7982 5468
rect 8006 5466 8062 5468
rect 7766 5414 7812 5466
rect 7812 5414 7822 5466
rect 7846 5414 7876 5466
rect 7876 5414 7888 5466
rect 7888 5414 7902 5466
rect 7926 5414 7940 5466
rect 7940 5414 7952 5466
rect 7952 5414 7982 5466
rect 8006 5414 8016 5466
rect 8016 5414 8062 5466
rect 7766 5412 7822 5414
rect 7846 5412 7902 5414
rect 7926 5412 7982 5414
rect 8006 5412 8062 5414
rect 9316 9274 9372 9276
rect 9396 9274 9452 9276
rect 9476 9274 9532 9276
rect 9556 9274 9612 9276
rect 9316 9222 9362 9274
rect 9362 9222 9372 9274
rect 9396 9222 9426 9274
rect 9426 9222 9438 9274
rect 9438 9222 9452 9274
rect 9476 9222 9490 9274
rect 9490 9222 9502 9274
rect 9502 9222 9532 9274
rect 9556 9222 9566 9274
rect 9566 9222 9612 9274
rect 9316 9220 9372 9222
rect 9396 9220 9452 9222
rect 9476 9220 9532 9222
rect 9556 9220 9612 9222
rect 9862 8472 9918 8528
rect 9316 8186 9372 8188
rect 9396 8186 9452 8188
rect 9476 8186 9532 8188
rect 9556 8186 9612 8188
rect 9316 8134 9362 8186
rect 9362 8134 9372 8186
rect 9396 8134 9426 8186
rect 9426 8134 9438 8186
rect 9438 8134 9452 8186
rect 9476 8134 9490 8186
rect 9490 8134 9502 8186
rect 9502 8134 9532 8186
rect 9556 8134 9566 8186
rect 9566 8134 9612 8186
rect 9316 8132 9372 8134
rect 9396 8132 9452 8134
rect 9476 8132 9532 8134
rect 9556 8132 9612 8134
rect 9770 7964 9772 7984
rect 9772 7964 9824 7984
rect 9824 7964 9826 7984
rect 9770 7928 9826 7964
rect 10138 7248 10194 7304
rect 9316 7098 9372 7100
rect 9396 7098 9452 7100
rect 9476 7098 9532 7100
rect 9556 7098 9612 7100
rect 9316 7046 9362 7098
rect 9362 7046 9372 7098
rect 9396 7046 9426 7098
rect 9426 7046 9438 7098
rect 9438 7046 9452 7098
rect 9476 7046 9490 7098
rect 9490 7046 9502 7098
rect 9502 7046 9532 7098
rect 9556 7046 9566 7098
rect 9566 7046 9612 7098
rect 9316 7044 9372 7046
rect 9396 7044 9452 7046
rect 9476 7044 9532 7046
rect 9556 7044 9612 7046
rect 10138 6996 10194 7032
rect 10138 6976 10140 6996
rect 10140 6976 10192 6996
rect 10192 6976 10194 6996
rect 10506 8336 10562 8392
rect 10414 7792 10470 7848
rect 9954 6704 10010 6760
rect 9316 6010 9372 6012
rect 9396 6010 9452 6012
rect 9476 6010 9532 6012
rect 9556 6010 9612 6012
rect 9316 5958 9362 6010
rect 9362 5958 9372 6010
rect 9396 5958 9426 6010
rect 9426 5958 9438 6010
rect 9438 5958 9452 6010
rect 9476 5958 9490 6010
rect 9490 5958 9502 6010
rect 9502 5958 9532 6010
rect 9556 5958 9566 6010
rect 9566 5958 9612 6010
rect 9316 5956 9372 5958
rect 9396 5956 9452 5958
rect 9476 5956 9532 5958
rect 9556 5956 9612 5958
rect 6216 3834 6272 3836
rect 6296 3834 6352 3836
rect 6376 3834 6432 3836
rect 6456 3834 6512 3836
rect 6216 3782 6262 3834
rect 6262 3782 6272 3834
rect 6296 3782 6326 3834
rect 6326 3782 6338 3834
rect 6338 3782 6352 3834
rect 6376 3782 6390 3834
rect 6390 3782 6402 3834
rect 6402 3782 6432 3834
rect 6456 3782 6466 3834
rect 6466 3782 6512 3834
rect 6216 3780 6272 3782
rect 6296 3780 6352 3782
rect 6376 3780 6432 3782
rect 6456 3780 6512 3782
rect 4802 3032 4804 3052
rect 4804 3032 4856 3052
rect 4856 3032 4858 3052
rect 3116 2746 3172 2748
rect 3196 2746 3252 2748
rect 3276 2746 3332 2748
rect 3356 2746 3412 2748
rect 3116 2694 3162 2746
rect 3162 2694 3172 2746
rect 3196 2694 3226 2746
rect 3226 2694 3238 2746
rect 3238 2694 3252 2746
rect 3276 2694 3290 2746
rect 3290 2694 3302 2746
rect 3302 2694 3332 2746
rect 3356 2694 3366 2746
rect 3366 2694 3412 2746
rect 3116 2692 3172 2694
rect 3196 2692 3252 2694
rect 3276 2692 3332 2694
rect 3356 2692 3412 2694
rect 3116 1658 3172 1660
rect 3196 1658 3252 1660
rect 3276 1658 3332 1660
rect 3356 1658 3412 1660
rect 3116 1606 3162 1658
rect 3162 1606 3172 1658
rect 3196 1606 3226 1658
rect 3226 1606 3238 1658
rect 3238 1606 3252 1658
rect 3276 1606 3290 1658
rect 3290 1606 3302 1658
rect 3302 1606 3332 1658
rect 3356 1606 3366 1658
rect 3366 1606 3412 1658
rect 3116 1604 3172 1606
rect 3196 1604 3252 1606
rect 3276 1604 3332 1606
rect 3356 1604 3412 1606
rect 4666 2202 4722 2204
rect 4746 2202 4802 2204
rect 4826 2202 4882 2204
rect 4906 2202 4962 2204
rect 4666 2150 4712 2202
rect 4712 2150 4722 2202
rect 4746 2150 4776 2202
rect 4776 2150 4788 2202
rect 4788 2150 4802 2202
rect 4826 2150 4840 2202
rect 4840 2150 4852 2202
rect 4852 2150 4882 2202
rect 4906 2150 4916 2202
rect 4916 2150 4962 2202
rect 4666 2148 4722 2150
rect 4746 2148 4802 2150
rect 4826 2148 4882 2150
rect 4906 2148 4962 2150
rect 6216 2746 6272 2748
rect 6296 2746 6352 2748
rect 6376 2746 6432 2748
rect 6456 2746 6512 2748
rect 6216 2694 6262 2746
rect 6262 2694 6272 2746
rect 6296 2694 6326 2746
rect 6326 2694 6338 2746
rect 6338 2694 6352 2746
rect 6376 2694 6390 2746
rect 6390 2694 6402 2746
rect 6402 2694 6432 2746
rect 6456 2694 6466 2746
rect 6466 2694 6512 2746
rect 6216 2692 6272 2694
rect 6296 2692 6352 2694
rect 6376 2692 6432 2694
rect 6456 2692 6512 2694
rect 6216 1658 6272 1660
rect 6296 1658 6352 1660
rect 6376 1658 6432 1660
rect 6456 1658 6512 1660
rect 6216 1606 6262 1658
rect 6262 1606 6272 1658
rect 6296 1606 6326 1658
rect 6326 1606 6338 1658
rect 6338 1606 6352 1658
rect 6376 1606 6390 1658
rect 6390 1606 6402 1658
rect 6402 1606 6432 1658
rect 6456 1606 6466 1658
rect 6466 1606 6512 1658
rect 6216 1604 6272 1606
rect 6296 1604 6352 1606
rect 6376 1604 6432 1606
rect 6456 1604 6512 1606
rect 6734 3032 6790 3088
rect 4666 1114 4722 1116
rect 4746 1114 4802 1116
rect 4826 1114 4882 1116
rect 4906 1114 4962 1116
rect 4666 1062 4712 1114
rect 4712 1062 4722 1114
rect 4746 1062 4776 1114
rect 4776 1062 4788 1114
rect 4788 1062 4802 1114
rect 4826 1062 4840 1114
rect 4840 1062 4852 1114
rect 4852 1062 4882 1114
rect 4906 1062 4916 1114
rect 4916 1062 4962 1114
rect 4666 1060 4722 1062
rect 4746 1060 4802 1062
rect 4826 1060 4882 1062
rect 4906 1060 4962 1062
rect 3116 570 3172 572
rect 3196 570 3252 572
rect 3276 570 3332 572
rect 3356 570 3412 572
rect 3116 518 3162 570
rect 3162 518 3172 570
rect 3196 518 3226 570
rect 3226 518 3238 570
rect 3238 518 3252 570
rect 3276 518 3290 570
rect 3290 518 3302 570
rect 3302 518 3332 570
rect 3356 518 3366 570
rect 3366 518 3412 570
rect 3116 516 3172 518
rect 3196 516 3252 518
rect 3276 516 3332 518
rect 3356 516 3412 518
rect 7766 4378 7822 4380
rect 7846 4378 7902 4380
rect 7926 4378 7982 4380
rect 8006 4378 8062 4380
rect 7766 4326 7812 4378
rect 7812 4326 7822 4378
rect 7846 4326 7876 4378
rect 7876 4326 7888 4378
rect 7888 4326 7902 4378
rect 7926 4326 7940 4378
rect 7940 4326 7952 4378
rect 7952 4326 7982 4378
rect 8006 4326 8016 4378
rect 8016 4326 8062 4378
rect 7766 4324 7822 4326
rect 7846 4324 7902 4326
rect 7926 4324 7982 4326
rect 8006 4324 8062 4326
rect 10866 9818 10922 9820
rect 10946 9818 11002 9820
rect 11026 9818 11082 9820
rect 11106 9818 11162 9820
rect 10866 9766 10912 9818
rect 10912 9766 10922 9818
rect 10946 9766 10976 9818
rect 10976 9766 10988 9818
rect 10988 9766 11002 9818
rect 11026 9766 11040 9818
rect 11040 9766 11052 9818
rect 11052 9766 11082 9818
rect 11106 9766 11116 9818
rect 11116 9766 11162 9818
rect 10866 9764 10922 9766
rect 10946 9764 11002 9766
rect 11026 9764 11082 9766
rect 11106 9764 11162 9766
rect 10866 8730 10922 8732
rect 10946 8730 11002 8732
rect 11026 8730 11082 8732
rect 11106 8730 11162 8732
rect 10866 8678 10912 8730
rect 10912 8678 10922 8730
rect 10946 8678 10976 8730
rect 10976 8678 10988 8730
rect 10988 8678 11002 8730
rect 11026 8678 11040 8730
rect 11040 8678 11052 8730
rect 11052 8678 11082 8730
rect 11106 8678 11116 8730
rect 11116 8678 11162 8730
rect 10866 8676 10922 8678
rect 10946 8676 11002 8678
rect 11026 8676 11082 8678
rect 11106 8676 11162 8678
rect 10874 8472 10930 8528
rect 11242 7948 11298 7984
rect 11242 7928 11244 7948
rect 11244 7928 11296 7948
rect 11296 7928 11298 7948
rect 10866 7642 10922 7644
rect 10946 7642 11002 7644
rect 11026 7642 11082 7644
rect 11106 7642 11162 7644
rect 10866 7590 10912 7642
rect 10912 7590 10922 7642
rect 10946 7590 10976 7642
rect 10976 7590 10988 7642
rect 10988 7590 11002 7642
rect 11026 7590 11040 7642
rect 11040 7590 11052 7642
rect 11052 7590 11082 7642
rect 11106 7590 11116 7642
rect 11116 7590 11162 7642
rect 10866 7588 10922 7590
rect 10946 7588 11002 7590
rect 11026 7588 11082 7590
rect 11106 7588 11162 7590
rect 11794 7828 11796 7848
rect 11796 7828 11848 7848
rect 11848 7828 11850 7848
rect 11794 7792 11850 7828
rect 10866 6554 10922 6556
rect 10946 6554 11002 6556
rect 11026 6554 11082 6556
rect 11106 6554 11162 6556
rect 10866 6502 10912 6554
rect 10912 6502 10922 6554
rect 10946 6502 10976 6554
rect 10976 6502 10988 6554
rect 10988 6502 11002 6554
rect 11026 6502 11040 6554
rect 11040 6502 11052 6554
rect 11052 6502 11082 6554
rect 11106 6502 11116 6554
rect 11116 6502 11162 6554
rect 10866 6500 10922 6502
rect 10946 6500 11002 6502
rect 11026 6500 11082 6502
rect 11106 6500 11162 6502
rect 11518 6740 11520 6760
rect 11520 6740 11572 6760
rect 11572 6740 11574 6760
rect 11518 6704 11574 6740
rect 12416 10362 12472 10364
rect 12496 10362 12552 10364
rect 12576 10362 12632 10364
rect 12656 10362 12712 10364
rect 12416 10310 12462 10362
rect 12462 10310 12472 10362
rect 12496 10310 12526 10362
rect 12526 10310 12538 10362
rect 12538 10310 12552 10362
rect 12576 10310 12590 10362
rect 12590 10310 12602 10362
rect 12602 10310 12632 10362
rect 12656 10310 12666 10362
rect 12666 10310 12712 10362
rect 12416 10308 12472 10310
rect 12496 10308 12552 10310
rect 12576 10308 12632 10310
rect 12656 10308 12712 10310
rect 13966 10906 14022 10908
rect 14046 10906 14102 10908
rect 14126 10906 14182 10908
rect 14206 10906 14262 10908
rect 13966 10854 14012 10906
rect 14012 10854 14022 10906
rect 14046 10854 14076 10906
rect 14076 10854 14088 10906
rect 14088 10854 14102 10906
rect 14126 10854 14140 10906
rect 14140 10854 14152 10906
rect 14152 10854 14182 10906
rect 14206 10854 14216 10906
rect 14216 10854 14262 10906
rect 13966 10852 14022 10854
rect 14046 10852 14102 10854
rect 14126 10852 14182 10854
rect 14206 10852 14262 10854
rect 12416 9274 12472 9276
rect 12496 9274 12552 9276
rect 12576 9274 12632 9276
rect 12656 9274 12712 9276
rect 12416 9222 12462 9274
rect 12462 9222 12472 9274
rect 12496 9222 12526 9274
rect 12526 9222 12538 9274
rect 12538 9222 12552 9274
rect 12576 9222 12590 9274
rect 12590 9222 12602 9274
rect 12602 9222 12632 9274
rect 12656 9222 12666 9274
rect 12666 9222 12712 9274
rect 12416 9220 12472 9222
rect 12496 9220 12552 9222
rect 12576 9220 12632 9222
rect 12656 9220 12712 9222
rect 12438 8336 12494 8392
rect 12416 8186 12472 8188
rect 12496 8186 12552 8188
rect 12576 8186 12632 8188
rect 12656 8186 12712 8188
rect 12416 8134 12462 8186
rect 12462 8134 12472 8186
rect 12496 8134 12526 8186
rect 12526 8134 12538 8186
rect 12538 8134 12552 8186
rect 12576 8134 12590 8186
rect 12590 8134 12602 8186
rect 12602 8134 12632 8186
rect 12656 8134 12666 8186
rect 12666 8134 12712 8186
rect 12416 8132 12472 8134
rect 12496 8132 12552 8134
rect 12576 8132 12632 8134
rect 12656 8132 12712 8134
rect 12416 7098 12472 7100
rect 12496 7098 12552 7100
rect 12576 7098 12632 7100
rect 12656 7098 12712 7100
rect 12416 7046 12462 7098
rect 12462 7046 12472 7098
rect 12496 7046 12526 7098
rect 12526 7046 12538 7098
rect 12538 7046 12552 7098
rect 12576 7046 12590 7098
rect 12590 7046 12602 7098
rect 12602 7046 12632 7098
rect 12656 7046 12666 7098
rect 12666 7046 12712 7098
rect 12416 7044 12472 7046
rect 12496 7044 12552 7046
rect 12576 7044 12632 7046
rect 12656 7044 12712 7046
rect 11886 6976 11942 7032
rect 12416 6010 12472 6012
rect 12496 6010 12552 6012
rect 12576 6010 12632 6012
rect 12656 6010 12712 6012
rect 12416 5958 12462 6010
rect 12462 5958 12472 6010
rect 12496 5958 12526 6010
rect 12526 5958 12538 6010
rect 12538 5958 12552 6010
rect 12576 5958 12590 6010
rect 12590 5958 12602 6010
rect 12602 5958 12632 6010
rect 12656 5958 12666 6010
rect 12666 5958 12712 6010
rect 12416 5956 12472 5958
rect 12496 5956 12552 5958
rect 12576 5956 12632 5958
rect 12656 5956 12712 5958
rect 10866 5466 10922 5468
rect 10946 5466 11002 5468
rect 11026 5466 11082 5468
rect 11106 5466 11162 5468
rect 10866 5414 10912 5466
rect 10912 5414 10922 5466
rect 10946 5414 10976 5466
rect 10976 5414 10988 5466
rect 10988 5414 11002 5466
rect 11026 5414 11040 5466
rect 11040 5414 11052 5466
rect 11052 5414 11082 5466
rect 11106 5414 11116 5466
rect 11116 5414 11162 5466
rect 10866 5412 10922 5414
rect 10946 5412 11002 5414
rect 11026 5412 11082 5414
rect 11106 5412 11162 5414
rect 8942 5218 8998 5264
rect 8942 5208 8944 5218
rect 8944 5208 8996 5218
rect 8996 5208 8998 5218
rect 9316 4922 9372 4924
rect 9396 4922 9452 4924
rect 9476 4922 9532 4924
rect 9556 4922 9612 4924
rect 9316 4870 9362 4922
rect 9362 4870 9372 4922
rect 9396 4870 9426 4922
rect 9426 4870 9438 4922
rect 9438 4870 9452 4922
rect 9476 4870 9490 4922
rect 9490 4870 9502 4922
rect 9502 4870 9532 4922
rect 9556 4870 9566 4922
rect 9566 4870 9612 4922
rect 9316 4868 9372 4870
rect 9396 4868 9452 4870
rect 9476 4868 9532 4870
rect 9556 4868 9612 4870
rect 7766 3290 7822 3292
rect 7846 3290 7902 3292
rect 7926 3290 7982 3292
rect 8006 3290 8062 3292
rect 7766 3238 7812 3290
rect 7812 3238 7822 3290
rect 7846 3238 7876 3290
rect 7876 3238 7888 3290
rect 7888 3238 7902 3290
rect 7926 3238 7940 3290
rect 7940 3238 7952 3290
rect 7952 3238 7982 3290
rect 8006 3238 8016 3290
rect 8016 3238 8062 3290
rect 7766 3236 7822 3238
rect 7846 3236 7902 3238
rect 7926 3236 7982 3238
rect 8006 3236 8062 3238
rect 7766 2202 7822 2204
rect 7846 2202 7902 2204
rect 7926 2202 7982 2204
rect 8006 2202 8062 2204
rect 7766 2150 7812 2202
rect 7812 2150 7822 2202
rect 7846 2150 7876 2202
rect 7876 2150 7888 2202
rect 7888 2150 7902 2202
rect 7926 2150 7940 2202
rect 7940 2150 7952 2202
rect 7952 2150 7982 2202
rect 8006 2150 8016 2202
rect 8016 2150 8062 2202
rect 7766 2148 7822 2150
rect 7846 2148 7902 2150
rect 7926 2148 7982 2150
rect 8006 2148 8062 2150
rect 6216 570 6272 572
rect 6296 570 6352 572
rect 6376 570 6432 572
rect 6456 570 6512 572
rect 6216 518 6262 570
rect 6262 518 6272 570
rect 6296 518 6326 570
rect 6326 518 6338 570
rect 6338 518 6352 570
rect 6376 518 6390 570
rect 6390 518 6402 570
rect 6402 518 6432 570
rect 6456 518 6466 570
rect 6466 518 6512 570
rect 6216 516 6272 518
rect 6296 516 6352 518
rect 6376 516 6432 518
rect 6456 516 6512 518
rect 7766 1114 7822 1116
rect 7846 1114 7902 1116
rect 7926 1114 7982 1116
rect 8006 1114 8062 1116
rect 7766 1062 7812 1114
rect 7812 1062 7822 1114
rect 7846 1062 7876 1114
rect 7876 1062 7888 1114
rect 7888 1062 7902 1114
rect 7926 1062 7940 1114
rect 7940 1062 7952 1114
rect 7952 1062 7982 1114
rect 8006 1062 8016 1114
rect 8016 1062 8062 1114
rect 7766 1060 7822 1062
rect 7846 1060 7902 1062
rect 7926 1060 7982 1062
rect 8006 1060 8062 1062
rect 9678 4540 9686 4584
rect 9686 4540 9734 4584
rect 9678 4528 9734 4540
rect 12416 4922 12472 4924
rect 12496 4922 12552 4924
rect 12576 4922 12632 4924
rect 12656 4922 12712 4924
rect 12416 4870 12462 4922
rect 12462 4870 12472 4922
rect 12496 4870 12526 4922
rect 12526 4870 12538 4922
rect 12538 4870 12552 4922
rect 12576 4870 12590 4922
rect 12590 4870 12602 4922
rect 12602 4870 12632 4922
rect 12656 4870 12666 4922
rect 12666 4870 12712 4922
rect 12416 4868 12472 4870
rect 12496 4868 12552 4870
rect 12576 4868 12632 4870
rect 12656 4868 12712 4870
rect 9316 3834 9372 3836
rect 9396 3834 9452 3836
rect 9476 3834 9532 3836
rect 9556 3834 9612 3836
rect 9316 3782 9362 3834
rect 9362 3782 9372 3834
rect 9396 3782 9426 3834
rect 9426 3782 9438 3834
rect 9438 3782 9452 3834
rect 9476 3782 9490 3834
rect 9490 3782 9502 3834
rect 9502 3782 9532 3834
rect 9556 3782 9566 3834
rect 9566 3782 9612 3834
rect 9316 3780 9372 3782
rect 9396 3780 9452 3782
rect 9476 3780 9532 3782
rect 9556 3780 9612 3782
rect 11334 4548 11390 4584
rect 11334 4528 11336 4548
rect 11336 4528 11388 4548
rect 11388 4528 11390 4548
rect 10866 4378 10922 4380
rect 10946 4378 11002 4380
rect 11026 4378 11082 4380
rect 11106 4378 11162 4380
rect 10866 4326 10912 4378
rect 10912 4326 10922 4378
rect 10946 4326 10976 4378
rect 10976 4326 10988 4378
rect 10988 4326 11002 4378
rect 11026 4326 11040 4378
rect 11040 4326 11052 4378
rect 11052 4326 11082 4378
rect 11106 4326 11116 4378
rect 11116 4326 11162 4378
rect 10866 4324 10922 4326
rect 10946 4324 11002 4326
rect 11026 4324 11082 4326
rect 11106 4324 11162 4326
rect 10866 3290 10922 3292
rect 10946 3290 11002 3292
rect 11026 3290 11082 3292
rect 11106 3290 11162 3292
rect 10866 3238 10912 3290
rect 10912 3238 10922 3290
rect 10946 3238 10976 3290
rect 10976 3238 10988 3290
rect 10988 3238 11002 3290
rect 11026 3238 11040 3290
rect 11040 3238 11052 3290
rect 11052 3238 11082 3290
rect 11106 3238 11116 3290
rect 11116 3238 11162 3290
rect 10866 3236 10922 3238
rect 10946 3236 11002 3238
rect 11026 3236 11082 3238
rect 11106 3236 11162 3238
rect 9316 2746 9372 2748
rect 9396 2746 9452 2748
rect 9476 2746 9532 2748
rect 9556 2746 9612 2748
rect 9316 2694 9362 2746
rect 9362 2694 9372 2746
rect 9396 2694 9426 2746
rect 9426 2694 9438 2746
rect 9438 2694 9452 2746
rect 9476 2694 9490 2746
rect 9490 2694 9502 2746
rect 9502 2694 9532 2746
rect 9556 2694 9566 2746
rect 9566 2694 9612 2746
rect 9316 2692 9372 2694
rect 9396 2692 9452 2694
rect 9476 2692 9532 2694
rect 9556 2692 9612 2694
rect 10866 2202 10922 2204
rect 10946 2202 11002 2204
rect 11026 2202 11082 2204
rect 11106 2202 11162 2204
rect 10866 2150 10912 2202
rect 10912 2150 10922 2202
rect 10946 2150 10976 2202
rect 10976 2150 10988 2202
rect 10988 2150 11002 2202
rect 11026 2150 11040 2202
rect 11040 2150 11052 2202
rect 11052 2150 11082 2202
rect 11106 2150 11116 2202
rect 11116 2150 11162 2202
rect 10866 2148 10922 2150
rect 10946 2148 11002 2150
rect 11026 2148 11082 2150
rect 11106 2148 11162 2150
rect 12416 3834 12472 3836
rect 12496 3834 12552 3836
rect 12576 3834 12632 3836
rect 12656 3834 12712 3836
rect 12416 3782 12462 3834
rect 12462 3782 12472 3834
rect 12496 3782 12526 3834
rect 12526 3782 12538 3834
rect 12538 3782 12552 3834
rect 12576 3782 12590 3834
rect 12590 3782 12602 3834
rect 12602 3782 12632 3834
rect 12656 3782 12666 3834
rect 12666 3782 12712 3834
rect 12416 3780 12472 3782
rect 12496 3780 12552 3782
rect 12576 3780 12632 3782
rect 12656 3780 12712 3782
rect 13966 9818 14022 9820
rect 14046 9818 14102 9820
rect 14126 9818 14182 9820
rect 14206 9818 14262 9820
rect 13966 9766 14012 9818
rect 14012 9766 14022 9818
rect 14046 9766 14076 9818
rect 14076 9766 14088 9818
rect 14088 9766 14102 9818
rect 14126 9766 14140 9818
rect 14140 9766 14152 9818
rect 14152 9766 14182 9818
rect 14206 9766 14216 9818
rect 14216 9766 14262 9818
rect 13966 9764 14022 9766
rect 14046 9764 14102 9766
rect 14126 9764 14182 9766
rect 14206 9764 14262 9766
rect 13966 8730 14022 8732
rect 14046 8730 14102 8732
rect 14126 8730 14182 8732
rect 14206 8730 14262 8732
rect 13966 8678 14012 8730
rect 14012 8678 14022 8730
rect 14046 8678 14076 8730
rect 14076 8678 14088 8730
rect 14088 8678 14102 8730
rect 14126 8678 14140 8730
rect 14140 8678 14152 8730
rect 14152 8678 14182 8730
rect 14206 8678 14216 8730
rect 14216 8678 14262 8730
rect 13966 8676 14022 8678
rect 14046 8676 14102 8678
rect 14126 8676 14182 8678
rect 14206 8676 14262 8678
rect 13966 7642 14022 7644
rect 14046 7642 14102 7644
rect 14126 7642 14182 7644
rect 14206 7642 14262 7644
rect 13966 7590 14012 7642
rect 14012 7590 14022 7642
rect 14046 7590 14076 7642
rect 14076 7590 14088 7642
rect 14088 7590 14102 7642
rect 14126 7590 14140 7642
rect 14140 7590 14152 7642
rect 14152 7590 14182 7642
rect 14206 7590 14216 7642
rect 14216 7590 14262 7642
rect 13966 7588 14022 7590
rect 14046 7588 14102 7590
rect 14126 7588 14182 7590
rect 14206 7588 14262 7590
rect 13542 7248 13598 7304
rect 13966 6554 14022 6556
rect 14046 6554 14102 6556
rect 14126 6554 14182 6556
rect 14206 6554 14262 6556
rect 13966 6502 14012 6554
rect 14012 6502 14022 6554
rect 14046 6502 14076 6554
rect 14076 6502 14088 6554
rect 14088 6502 14102 6554
rect 14126 6502 14140 6554
rect 14140 6502 14152 6554
rect 14152 6502 14182 6554
rect 14206 6502 14216 6554
rect 14216 6502 14262 6554
rect 13966 6500 14022 6502
rect 14046 6500 14102 6502
rect 14126 6500 14182 6502
rect 14206 6500 14262 6502
rect 13966 5466 14022 5468
rect 14046 5466 14102 5468
rect 14126 5466 14182 5468
rect 14206 5466 14262 5468
rect 13966 5414 14012 5466
rect 14012 5414 14022 5466
rect 14046 5414 14076 5466
rect 14076 5414 14088 5466
rect 14088 5414 14102 5466
rect 14126 5414 14140 5466
rect 14140 5414 14152 5466
rect 14152 5414 14182 5466
rect 14206 5414 14216 5466
rect 14216 5414 14262 5466
rect 13966 5412 14022 5414
rect 14046 5412 14102 5414
rect 14126 5412 14182 5414
rect 14206 5412 14262 5414
rect 17066 10906 17122 10908
rect 17146 10906 17202 10908
rect 17226 10906 17282 10908
rect 17306 10906 17362 10908
rect 17066 10854 17112 10906
rect 17112 10854 17122 10906
rect 17146 10854 17176 10906
rect 17176 10854 17188 10906
rect 17188 10854 17202 10906
rect 17226 10854 17240 10906
rect 17240 10854 17252 10906
rect 17252 10854 17282 10906
rect 17306 10854 17316 10906
rect 17316 10854 17362 10906
rect 17066 10852 17122 10854
rect 17146 10852 17202 10854
rect 17226 10852 17282 10854
rect 17306 10852 17362 10854
rect 15516 10362 15572 10364
rect 15596 10362 15652 10364
rect 15676 10362 15732 10364
rect 15756 10362 15812 10364
rect 15516 10310 15562 10362
rect 15562 10310 15572 10362
rect 15596 10310 15626 10362
rect 15626 10310 15638 10362
rect 15638 10310 15652 10362
rect 15676 10310 15690 10362
rect 15690 10310 15702 10362
rect 15702 10310 15732 10362
rect 15756 10310 15766 10362
rect 15766 10310 15812 10362
rect 15516 10308 15572 10310
rect 15596 10308 15652 10310
rect 15676 10308 15732 10310
rect 15756 10308 15812 10310
rect 17066 9818 17122 9820
rect 17146 9818 17202 9820
rect 17226 9818 17282 9820
rect 17306 9818 17362 9820
rect 17066 9766 17112 9818
rect 17112 9766 17122 9818
rect 17146 9766 17176 9818
rect 17176 9766 17188 9818
rect 17188 9766 17202 9818
rect 17226 9766 17240 9818
rect 17240 9766 17252 9818
rect 17252 9766 17282 9818
rect 17306 9766 17316 9818
rect 17316 9766 17362 9818
rect 17066 9764 17122 9766
rect 17146 9764 17202 9766
rect 17226 9764 17282 9766
rect 17306 9764 17362 9766
rect 17958 9696 18014 9752
rect 15516 9274 15572 9276
rect 15596 9274 15652 9276
rect 15676 9274 15732 9276
rect 15756 9274 15812 9276
rect 15516 9222 15562 9274
rect 15562 9222 15572 9274
rect 15596 9222 15626 9274
rect 15626 9222 15638 9274
rect 15638 9222 15652 9274
rect 15676 9222 15690 9274
rect 15690 9222 15702 9274
rect 15702 9222 15732 9274
rect 15756 9222 15766 9274
rect 15766 9222 15812 9274
rect 15516 9220 15572 9222
rect 15596 9220 15652 9222
rect 15676 9220 15732 9222
rect 15756 9220 15812 9222
rect 15516 8186 15572 8188
rect 15596 8186 15652 8188
rect 15676 8186 15732 8188
rect 15756 8186 15812 8188
rect 15516 8134 15562 8186
rect 15562 8134 15572 8186
rect 15596 8134 15626 8186
rect 15626 8134 15638 8186
rect 15638 8134 15652 8186
rect 15676 8134 15690 8186
rect 15690 8134 15702 8186
rect 15702 8134 15732 8186
rect 15756 8134 15766 8186
rect 15766 8134 15812 8186
rect 15516 8132 15572 8134
rect 15596 8132 15652 8134
rect 15676 8132 15732 8134
rect 15756 8132 15812 8134
rect 15516 7098 15572 7100
rect 15596 7098 15652 7100
rect 15676 7098 15732 7100
rect 15756 7098 15812 7100
rect 15516 7046 15562 7098
rect 15562 7046 15572 7098
rect 15596 7046 15626 7098
rect 15626 7046 15638 7098
rect 15638 7046 15652 7098
rect 15676 7046 15690 7098
rect 15690 7046 15702 7098
rect 15702 7046 15732 7098
rect 15756 7046 15766 7098
rect 15766 7046 15812 7098
rect 15516 7044 15572 7046
rect 15596 7044 15652 7046
rect 15676 7044 15732 7046
rect 15756 7044 15812 7046
rect 15516 6010 15572 6012
rect 15596 6010 15652 6012
rect 15676 6010 15732 6012
rect 15756 6010 15812 6012
rect 15516 5958 15562 6010
rect 15562 5958 15572 6010
rect 15596 5958 15626 6010
rect 15626 5958 15638 6010
rect 15638 5958 15652 6010
rect 15676 5958 15690 6010
rect 15690 5958 15702 6010
rect 15702 5958 15732 6010
rect 15756 5958 15766 6010
rect 15766 5958 15812 6010
rect 15516 5956 15572 5958
rect 15596 5956 15652 5958
rect 15676 5956 15732 5958
rect 15756 5956 15812 5958
rect 17066 8730 17122 8732
rect 17146 8730 17202 8732
rect 17226 8730 17282 8732
rect 17306 8730 17362 8732
rect 17066 8678 17112 8730
rect 17112 8678 17122 8730
rect 17146 8678 17176 8730
rect 17176 8678 17188 8730
rect 17188 8678 17202 8730
rect 17226 8678 17240 8730
rect 17240 8678 17252 8730
rect 17252 8678 17282 8730
rect 17306 8678 17316 8730
rect 17316 8678 17362 8730
rect 17066 8676 17122 8678
rect 17146 8676 17202 8678
rect 17226 8676 17282 8678
rect 17306 8676 17362 8678
rect 17066 7642 17122 7644
rect 17146 7642 17202 7644
rect 17226 7642 17282 7644
rect 17306 7642 17362 7644
rect 17066 7590 17112 7642
rect 17112 7590 17122 7642
rect 17146 7590 17176 7642
rect 17176 7590 17188 7642
rect 17188 7590 17202 7642
rect 17226 7590 17240 7642
rect 17240 7590 17252 7642
rect 17252 7590 17282 7642
rect 17306 7590 17316 7642
rect 17316 7590 17362 7642
rect 17066 7588 17122 7590
rect 17146 7588 17202 7590
rect 17226 7588 17282 7590
rect 17306 7588 17362 7590
rect 18786 11192 18842 11248
rect 18510 8200 18566 8256
rect 18510 6740 18512 6760
rect 18512 6740 18564 6760
rect 18564 6740 18566 6760
rect 17066 6554 17122 6556
rect 17146 6554 17202 6556
rect 17226 6554 17282 6556
rect 17306 6554 17362 6556
rect 17066 6502 17112 6554
rect 17112 6502 17122 6554
rect 17146 6502 17176 6554
rect 17176 6502 17188 6554
rect 17188 6502 17202 6554
rect 17226 6502 17240 6554
rect 17240 6502 17252 6554
rect 17252 6502 17282 6554
rect 17306 6502 17316 6554
rect 17316 6502 17362 6554
rect 17066 6500 17122 6502
rect 17146 6500 17202 6502
rect 17226 6500 17282 6502
rect 17306 6500 17362 6502
rect 18510 6704 18566 6740
rect 17066 5466 17122 5468
rect 17146 5466 17202 5468
rect 17226 5466 17282 5468
rect 17306 5466 17362 5468
rect 17066 5414 17112 5466
rect 17112 5414 17122 5466
rect 17146 5414 17176 5466
rect 17176 5414 17188 5466
rect 17188 5414 17202 5466
rect 17226 5414 17240 5466
rect 17240 5414 17252 5466
rect 17252 5414 17282 5466
rect 17306 5414 17316 5466
rect 17316 5414 17362 5466
rect 17066 5412 17122 5414
rect 17146 5412 17202 5414
rect 17226 5412 17282 5414
rect 17306 5412 17362 5414
rect 13966 4378 14022 4380
rect 14046 4378 14102 4380
rect 14126 4378 14182 4380
rect 14206 4378 14262 4380
rect 13966 4326 14012 4378
rect 14012 4326 14022 4378
rect 14046 4326 14076 4378
rect 14076 4326 14088 4378
rect 14088 4326 14102 4378
rect 14126 4326 14140 4378
rect 14140 4326 14152 4378
rect 14152 4326 14182 4378
rect 14206 4326 14216 4378
rect 14216 4326 14262 4378
rect 13966 4324 14022 4326
rect 14046 4324 14102 4326
rect 14126 4324 14182 4326
rect 14206 4324 14262 4326
rect 12416 2746 12472 2748
rect 12496 2746 12552 2748
rect 12576 2746 12632 2748
rect 12656 2746 12712 2748
rect 12416 2694 12462 2746
rect 12462 2694 12472 2746
rect 12496 2694 12526 2746
rect 12526 2694 12538 2746
rect 12538 2694 12552 2746
rect 12576 2694 12590 2746
rect 12590 2694 12602 2746
rect 12602 2694 12632 2746
rect 12656 2694 12666 2746
rect 12666 2694 12712 2746
rect 12416 2692 12472 2694
rect 12496 2692 12552 2694
rect 12576 2692 12632 2694
rect 12656 2692 12712 2694
rect 9316 1658 9372 1660
rect 9396 1658 9452 1660
rect 9476 1658 9532 1660
rect 9556 1658 9612 1660
rect 9316 1606 9362 1658
rect 9362 1606 9372 1658
rect 9396 1606 9426 1658
rect 9426 1606 9438 1658
rect 9438 1606 9452 1658
rect 9476 1606 9490 1658
rect 9490 1606 9502 1658
rect 9502 1606 9532 1658
rect 9556 1606 9566 1658
rect 9566 1606 9612 1658
rect 9316 1604 9372 1606
rect 9396 1604 9452 1606
rect 9476 1604 9532 1606
rect 9556 1604 9612 1606
rect 10866 1114 10922 1116
rect 10946 1114 11002 1116
rect 11026 1114 11082 1116
rect 11106 1114 11162 1116
rect 10866 1062 10912 1114
rect 10912 1062 10922 1114
rect 10946 1062 10976 1114
rect 10976 1062 10988 1114
rect 10988 1062 11002 1114
rect 11026 1062 11040 1114
rect 11040 1062 11052 1114
rect 11052 1062 11082 1114
rect 11106 1062 11116 1114
rect 11116 1062 11162 1114
rect 10866 1060 10922 1062
rect 10946 1060 11002 1062
rect 11026 1060 11082 1062
rect 11106 1060 11162 1062
rect 9316 570 9372 572
rect 9396 570 9452 572
rect 9476 570 9532 572
rect 9556 570 9612 572
rect 9316 518 9362 570
rect 9362 518 9372 570
rect 9396 518 9426 570
rect 9426 518 9438 570
rect 9438 518 9452 570
rect 9476 518 9490 570
rect 9490 518 9502 570
rect 9502 518 9532 570
rect 9556 518 9566 570
rect 9566 518 9612 570
rect 9316 516 9372 518
rect 9396 516 9452 518
rect 9476 516 9532 518
rect 9556 516 9612 518
rect 12416 1658 12472 1660
rect 12496 1658 12552 1660
rect 12576 1658 12632 1660
rect 12656 1658 12712 1660
rect 12416 1606 12462 1658
rect 12462 1606 12472 1658
rect 12496 1606 12526 1658
rect 12526 1606 12538 1658
rect 12538 1606 12552 1658
rect 12576 1606 12590 1658
rect 12590 1606 12602 1658
rect 12602 1606 12632 1658
rect 12656 1606 12666 1658
rect 12666 1606 12712 1658
rect 12416 1604 12472 1606
rect 12496 1604 12552 1606
rect 12576 1604 12632 1606
rect 12656 1604 12712 1606
rect 12416 570 12472 572
rect 12496 570 12552 572
rect 12576 570 12632 572
rect 12656 570 12712 572
rect 12416 518 12462 570
rect 12462 518 12472 570
rect 12496 518 12526 570
rect 12526 518 12538 570
rect 12538 518 12552 570
rect 12576 518 12590 570
rect 12590 518 12602 570
rect 12602 518 12632 570
rect 12656 518 12666 570
rect 12666 518 12712 570
rect 12416 516 12472 518
rect 12496 516 12552 518
rect 12576 516 12632 518
rect 12656 516 12712 518
rect 15516 4922 15572 4924
rect 15596 4922 15652 4924
rect 15676 4922 15732 4924
rect 15756 4922 15812 4924
rect 15516 4870 15562 4922
rect 15562 4870 15572 4922
rect 15596 4870 15626 4922
rect 15626 4870 15638 4922
rect 15638 4870 15652 4922
rect 15676 4870 15690 4922
rect 15690 4870 15702 4922
rect 15702 4870 15732 4922
rect 15756 4870 15766 4922
rect 15766 4870 15812 4922
rect 15516 4868 15572 4870
rect 15596 4868 15652 4870
rect 15676 4868 15732 4870
rect 15756 4868 15812 4870
rect 18510 5208 18566 5264
rect 13966 3290 14022 3292
rect 14046 3290 14102 3292
rect 14126 3290 14182 3292
rect 14206 3290 14262 3292
rect 13966 3238 14012 3290
rect 14012 3238 14022 3290
rect 14046 3238 14076 3290
rect 14076 3238 14088 3290
rect 14088 3238 14102 3290
rect 14126 3238 14140 3290
rect 14140 3238 14152 3290
rect 14152 3238 14182 3290
rect 14206 3238 14216 3290
rect 14216 3238 14262 3290
rect 13966 3236 14022 3238
rect 14046 3236 14102 3238
rect 14126 3236 14182 3238
rect 14206 3236 14262 3238
rect 13966 2202 14022 2204
rect 14046 2202 14102 2204
rect 14126 2202 14182 2204
rect 14206 2202 14262 2204
rect 13966 2150 14012 2202
rect 14012 2150 14022 2202
rect 14046 2150 14076 2202
rect 14076 2150 14088 2202
rect 14088 2150 14102 2202
rect 14126 2150 14140 2202
rect 14140 2150 14152 2202
rect 14152 2150 14182 2202
rect 14206 2150 14216 2202
rect 14216 2150 14262 2202
rect 13966 2148 14022 2150
rect 14046 2148 14102 2150
rect 14126 2148 14182 2150
rect 14206 2148 14262 2150
rect 15516 3834 15572 3836
rect 15596 3834 15652 3836
rect 15676 3834 15732 3836
rect 15756 3834 15812 3836
rect 15516 3782 15562 3834
rect 15562 3782 15572 3834
rect 15596 3782 15626 3834
rect 15626 3782 15638 3834
rect 15638 3782 15652 3834
rect 15676 3782 15690 3834
rect 15690 3782 15702 3834
rect 15702 3782 15732 3834
rect 15756 3782 15766 3834
rect 15766 3782 15812 3834
rect 15516 3780 15572 3782
rect 15596 3780 15652 3782
rect 15676 3780 15732 3782
rect 15756 3780 15812 3782
rect 17066 4378 17122 4380
rect 17146 4378 17202 4380
rect 17226 4378 17282 4380
rect 17306 4378 17362 4380
rect 17066 4326 17112 4378
rect 17112 4326 17122 4378
rect 17146 4326 17176 4378
rect 17176 4326 17188 4378
rect 17188 4326 17202 4378
rect 17226 4326 17240 4378
rect 17240 4326 17252 4378
rect 17252 4326 17282 4378
rect 17306 4326 17316 4378
rect 17316 4326 17362 4378
rect 17066 4324 17122 4326
rect 17146 4324 17202 4326
rect 17226 4324 17282 4326
rect 17306 4324 17362 4326
rect 15516 2746 15572 2748
rect 15596 2746 15652 2748
rect 15676 2746 15732 2748
rect 15756 2746 15812 2748
rect 15516 2694 15562 2746
rect 15562 2694 15572 2746
rect 15596 2694 15626 2746
rect 15626 2694 15638 2746
rect 15638 2694 15652 2746
rect 15676 2694 15690 2746
rect 15690 2694 15702 2746
rect 15702 2694 15732 2746
rect 15756 2694 15766 2746
rect 15766 2694 15812 2746
rect 15516 2692 15572 2694
rect 15596 2692 15652 2694
rect 15676 2692 15732 2694
rect 15756 2692 15812 2694
rect 15516 1658 15572 1660
rect 15596 1658 15652 1660
rect 15676 1658 15732 1660
rect 15756 1658 15812 1660
rect 15516 1606 15562 1658
rect 15562 1606 15572 1658
rect 15596 1606 15626 1658
rect 15626 1606 15638 1658
rect 15638 1606 15652 1658
rect 15676 1606 15690 1658
rect 15690 1606 15702 1658
rect 15702 1606 15732 1658
rect 15756 1606 15766 1658
rect 15766 1606 15812 1658
rect 15516 1604 15572 1606
rect 15596 1604 15652 1606
rect 15676 1604 15732 1606
rect 15756 1604 15812 1606
rect 13966 1114 14022 1116
rect 14046 1114 14102 1116
rect 14126 1114 14182 1116
rect 14206 1114 14262 1116
rect 13966 1062 14012 1114
rect 14012 1062 14022 1114
rect 14046 1062 14076 1114
rect 14076 1062 14088 1114
rect 14088 1062 14102 1114
rect 14126 1062 14140 1114
rect 14140 1062 14152 1114
rect 14152 1062 14182 1114
rect 14206 1062 14216 1114
rect 14216 1062 14262 1114
rect 13966 1060 14022 1062
rect 14046 1060 14102 1062
rect 14126 1060 14182 1062
rect 14206 1060 14262 1062
rect 17066 3290 17122 3292
rect 17146 3290 17202 3292
rect 17226 3290 17282 3292
rect 17306 3290 17362 3292
rect 17066 3238 17112 3290
rect 17112 3238 17122 3290
rect 17146 3238 17176 3290
rect 17176 3238 17188 3290
rect 17188 3238 17202 3290
rect 17226 3238 17240 3290
rect 17240 3238 17252 3290
rect 17252 3238 17282 3290
rect 17306 3238 17316 3290
rect 17316 3238 17362 3290
rect 17066 3236 17122 3238
rect 17146 3236 17202 3238
rect 17226 3236 17282 3238
rect 17306 3236 17362 3238
rect 17066 2202 17122 2204
rect 17146 2202 17202 2204
rect 17226 2202 17282 2204
rect 17306 2202 17362 2204
rect 17066 2150 17112 2202
rect 17112 2150 17122 2202
rect 17146 2150 17176 2202
rect 17176 2150 17188 2202
rect 17188 2150 17202 2202
rect 17226 2150 17240 2202
rect 17240 2150 17252 2202
rect 17252 2150 17282 2202
rect 17306 2150 17316 2202
rect 17316 2150 17362 2202
rect 17066 2148 17122 2150
rect 17146 2148 17202 2150
rect 17226 2148 17282 2150
rect 17306 2148 17362 2150
rect 15516 570 15572 572
rect 15596 570 15652 572
rect 15676 570 15732 572
rect 15756 570 15812 572
rect 15516 518 15562 570
rect 15562 518 15572 570
rect 15596 518 15626 570
rect 15626 518 15638 570
rect 15638 518 15652 570
rect 15676 518 15690 570
rect 15690 518 15702 570
rect 15702 518 15732 570
rect 15756 518 15766 570
rect 15766 518 15812 570
rect 15516 516 15572 518
rect 15596 516 15652 518
rect 15676 516 15732 518
rect 15756 516 15812 518
rect 17066 1114 17122 1116
rect 17146 1114 17202 1116
rect 17226 1114 17282 1116
rect 17306 1114 17362 1116
rect 17066 1062 17112 1114
rect 17112 1062 17122 1114
rect 17146 1062 17176 1114
rect 17176 1062 17188 1114
rect 17188 1062 17202 1114
rect 17226 1062 17240 1114
rect 17240 1062 17252 1114
rect 17252 1062 17282 1114
rect 17306 1062 17316 1114
rect 17316 1062 17362 1114
rect 17066 1060 17122 1062
rect 17146 1060 17202 1062
rect 17226 1060 17282 1062
rect 17306 1060 17362 1062
rect 18510 3712 18566 3768
rect 18510 2216 18566 2272
rect 18510 720 18566 776
rect 4666 26 4722 28
rect 4746 26 4802 28
rect 4826 26 4882 28
rect 4906 26 4962 28
rect 4666 -26 4712 26
rect 4712 -26 4722 26
rect 4746 -26 4776 26
rect 4776 -26 4788 26
rect 4788 -26 4802 26
rect 4826 -26 4840 26
rect 4840 -26 4852 26
rect 4852 -26 4882 26
rect 4906 -26 4916 26
rect 4916 -26 4962 26
rect 4666 -28 4722 -26
rect 4746 -28 4802 -26
rect 4826 -28 4882 -26
rect 4906 -28 4962 -26
rect 7766 26 7822 28
rect 7846 26 7902 28
rect 7926 26 7982 28
rect 8006 26 8062 28
rect 7766 -26 7812 26
rect 7812 -26 7822 26
rect 7846 -26 7876 26
rect 7876 -26 7888 26
rect 7888 -26 7902 26
rect 7926 -26 7940 26
rect 7940 -26 7952 26
rect 7952 -26 7982 26
rect 8006 -26 8016 26
rect 8016 -26 8062 26
rect 7766 -28 7822 -26
rect 7846 -28 7902 -26
rect 7926 -28 7982 -26
rect 8006 -28 8062 -26
rect 10866 26 10922 28
rect 10946 26 11002 28
rect 11026 26 11082 28
rect 11106 26 11162 28
rect 10866 -26 10912 26
rect 10912 -26 10922 26
rect 10946 -26 10976 26
rect 10976 -26 10988 26
rect 10988 -26 11002 26
rect 11026 -26 11040 26
rect 11040 -26 11052 26
rect 11052 -26 11082 26
rect 11106 -26 11116 26
rect 11116 -26 11162 26
rect 10866 -28 10922 -26
rect 10946 -28 11002 -26
rect 11026 -28 11082 -26
rect 11106 -28 11162 -26
rect 13966 26 14022 28
rect 14046 26 14102 28
rect 14126 26 14182 28
rect 14206 26 14262 28
rect 13966 -26 14012 26
rect 14012 -26 14022 26
rect 14046 -26 14076 26
rect 14076 -26 14088 26
rect 14088 -26 14102 26
rect 14126 -26 14140 26
rect 14140 -26 14152 26
rect 14152 -26 14182 26
rect 14206 -26 14216 26
rect 14216 -26 14262 26
rect 13966 -28 14022 -26
rect 14046 -28 14102 -26
rect 14126 -28 14182 -26
rect 14206 -28 14262 -26
rect 17066 26 17122 28
rect 17146 26 17202 28
rect 17226 26 17282 28
rect 17306 26 17362 28
rect 17066 -26 17112 26
rect 17112 -26 17122 26
rect 17146 -26 17176 26
rect 17176 -26 17188 26
rect 17188 -26 17202 26
rect 17226 -26 17240 26
rect 17240 -26 17252 26
rect 17252 -26 17282 26
rect 17306 -26 17316 26
rect 17316 -26 17362 26
rect 17066 -28 17122 -26
rect 17146 -28 17202 -26
rect 17226 -28 17282 -26
rect 17306 -28 17362 -26
<< metal3 >>
rect 18781 11250 18847 11253
rect 19200 11250 20000 11280
rect 18781 11248 20000 11250
rect 18781 11192 18786 11248
rect 18842 11192 20000 11248
rect 18781 11190 20000 11192
rect 18781 11187 18847 11190
rect 19200 11160 20000 11190
rect 4654 10912 4974 10913
rect 4654 10848 4662 10912
rect 4726 10848 4742 10912
rect 4806 10848 4822 10912
rect 4886 10848 4902 10912
rect 4966 10848 4974 10912
rect 4654 10847 4974 10848
rect 7754 10912 8074 10913
rect 7754 10848 7762 10912
rect 7826 10848 7842 10912
rect 7906 10848 7922 10912
rect 7986 10848 8002 10912
rect 8066 10848 8074 10912
rect 7754 10847 8074 10848
rect 10854 10912 11174 10913
rect 10854 10848 10862 10912
rect 10926 10848 10942 10912
rect 11006 10848 11022 10912
rect 11086 10848 11102 10912
rect 11166 10848 11174 10912
rect 10854 10847 11174 10848
rect 13954 10912 14274 10913
rect 13954 10848 13962 10912
rect 14026 10848 14042 10912
rect 14106 10848 14122 10912
rect 14186 10848 14202 10912
rect 14266 10848 14274 10912
rect 13954 10847 14274 10848
rect 17054 10912 17374 10913
rect 17054 10848 17062 10912
rect 17126 10848 17142 10912
rect 17206 10848 17222 10912
rect 17286 10848 17302 10912
rect 17366 10848 17374 10912
rect 17054 10847 17374 10848
rect 3104 10368 3424 10369
rect 3104 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3272 10368
rect 3336 10304 3352 10368
rect 3416 10304 3424 10368
rect 3104 10303 3424 10304
rect 6204 10368 6524 10369
rect 6204 10304 6212 10368
rect 6276 10304 6292 10368
rect 6356 10304 6372 10368
rect 6436 10304 6452 10368
rect 6516 10304 6524 10368
rect 6204 10303 6524 10304
rect 9304 10368 9624 10369
rect 9304 10304 9312 10368
rect 9376 10304 9392 10368
rect 9456 10304 9472 10368
rect 9536 10304 9552 10368
rect 9616 10304 9624 10368
rect 9304 10303 9624 10304
rect 12404 10368 12724 10369
rect 12404 10304 12412 10368
rect 12476 10304 12492 10368
rect 12556 10304 12572 10368
rect 12636 10304 12652 10368
rect 12716 10304 12724 10368
rect 12404 10303 12724 10304
rect 15504 10368 15824 10369
rect 15504 10304 15512 10368
rect 15576 10304 15592 10368
rect 15656 10304 15672 10368
rect 15736 10304 15752 10368
rect 15816 10304 15824 10368
rect 15504 10303 15824 10304
rect 4654 9824 4974 9825
rect 4654 9760 4662 9824
rect 4726 9760 4742 9824
rect 4806 9760 4822 9824
rect 4886 9760 4902 9824
rect 4966 9760 4974 9824
rect 4654 9759 4974 9760
rect 7754 9824 8074 9825
rect 7754 9760 7762 9824
rect 7826 9760 7842 9824
rect 7906 9760 7922 9824
rect 7986 9760 8002 9824
rect 8066 9760 8074 9824
rect 7754 9759 8074 9760
rect 10854 9824 11174 9825
rect 10854 9760 10862 9824
rect 10926 9760 10942 9824
rect 11006 9760 11022 9824
rect 11086 9760 11102 9824
rect 11166 9760 11174 9824
rect 10854 9759 11174 9760
rect 13954 9824 14274 9825
rect 13954 9760 13962 9824
rect 14026 9760 14042 9824
rect 14106 9760 14122 9824
rect 14186 9760 14202 9824
rect 14266 9760 14274 9824
rect 13954 9759 14274 9760
rect 17054 9824 17374 9825
rect 17054 9760 17062 9824
rect 17126 9760 17142 9824
rect 17206 9760 17222 9824
rect 17286 9760 17302 9824
rect 17366 9760 17374 9824
rect 17054 9759 17374 9760
rect 17953 9754 18019 9757
rect 19200 9754 20000 9784
rect 17953 9752 20000 9754
rect 17953 9696 17958 9752
rect 18014 9696 20000 9752
rect 17953 9694 20000 9696
rect 17953 9691 18019 9694
rect 19200 9664 20000 9694
rect 3104 9280 3424 9281
rect 3104 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3272 9280
rect 3336 9216 3352 9280
rect 3416 9216 3424 9280
rect 3104 9215 3424 9216
rect 6204 9280 6524 9281
rect 6204 9216 6212 9280
rect 6276 9216 6292 9280
rect 6356 9216 6372 9280
rect 6436 9216 6452 9280
rect 6516 9216 6524 9280
rect 6204 9215 6524 9216
rect 9304 9280 9624 9281
rect 9304 9216 9312 9280
rect 9376 9216 9392 9280
rect 9456 9216 9472 9280
rect 9536 9216 9552 9280
rect 9616 9216 9624 9280
rect 9304 9215 9624 9216
rect 12404 9280 12724 9281
rect 12404 9216 12412 9280
rect 12476 9216 12492 9280
rect 12556 9216 12572 9280
rect 12636 9216 12652 9280
rect 12716 9216 12724 9280
rect 12404 9215 12724 9216
rect 15504 9280 15824 9281
rect 15504 9216 15512 9280
rect 15576 9216 15592 9280
rect 15656 9216 15672 9280
rect 15736 9216 15752 9280
rect 15816 9216 15824 9280
rect 15504 9215 15824 9216
rect 4654 8736 4974 8737
rect 4654 8672 4662 8736
rect 4726 8672 4742 8736
rect 4806 8672 4822 8736
rect 4886 8672 4902 8736
rect 4966 8672 4974 8736
rect 4654 8671 4974 8672
rect 7754 8736 8074 8737
rect 7754 8672 7762 8736
rect 7826 8672 7842 8736
rect 7906 8672 7922 8736
rect 7986 8672 8002 8736
rect 8066 8672 8074 8736
rect 7754 8671 8074 8672
rect 10854 8736 11174 8737
rect 10854 8672 10862 8736
rect 10926 8672 10942 8736
rect 11006 8672 11022 8736
rect 11086 8672 11102 8736
rect 11166 8672 11174 8736
rect 10854 8671 11174 8672
rect 13954 8736 14274 8737
rect 13954 8672 13962 8736
rect 14026 8672 14042 8736
rect 14106 8672 14122 8736
rect 14186 8672 14202 8736
rect 14266 8672 14274 8736
rect 13954 8671 14274 8672
rect 17054 8736 17374 8737
rect 17054 8672 17062 8736
rect 17126 8672 17142 8736
rect 17206 8672 17222 8736
rect 17286 8672 17302 8736
rect 17366 8672 17374 8736
rect 17054 8671 17374 8672
rect 9857 8530 9923 8533
rect 10869 8530 10935 8533
rect 9857 8528 10935 8530
rect 9857 8472 9862 8528
rect 9918 8472 10874 8528
rect 10930 8472 10935 8528
rect 9857 8470 10935 8472
rect 9857 8467 9923 8470
rect 10869 8467 10935 8470
rect 10501 8394 10567 8397
rect 12433 8394 12499 8397
rect 10501 8392 12499 8394
rect 10501 8336 10506 8392
rect 10562 8336 12438 8392
rect 12494 8336 12499 8392
rect 10501 8334 12499 8336
rect 10501 8331 10567 8334
rect 12433 8331 12499 8334
rect 18505 8258 18571 8261
rect 19200 8258 20000 8288
rect 18505 8256 20000 8258
rect 18505 8200 18510 8256
rect 18566 8200 20000 8256
rect 18505 8198 20000 8200
rect 18505 8195 18571 8198
rect 3104 8192 3424 8193
rect 3104 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3272 8192
rect 3336 8128 3352 8192
rect 3416 8128 3424 8192
rect 3104 8127 3424 8128
rect 6204 8192 6524 8193
rect 6204 8128 6212 8192
rect 6276 8128 6292 8192
rect 6356 8128 6372 8192
rect 6436 8128 6452 8192
rect 6516 8128 6524 8192
rect 6204 8127 6524 8128
rect 9304 8192 9624 8193
rect 9304 8128 9312 8192
rect 9376 8128 9392 8192
rect 9456 8128 9472 8192
rect 9536 8128 9552 8192
rect 9616 8128 9624 8192
rect 9304 8127 9624 8128
rect 12404 8192 12724 8193
rect 12404 8128 12412 8192
rect 12476 8128 12492 8192
rect 12556 8128 12572 8192
rect 12636 8128 12652 8192
rect 12716 8128 12724 8192
rect 12404 8127 12724 8128
rect 15504 8192 15824 8193
rect 15504 8128 15512 8192
rect 15576 8128 15592 8192
rect 15656 8128 15672 8192
rect 15736 8128 15752 8192
rect 15816 8128 15824 8192
rect 19200 8168 20000 8198
rect 15504 8127 15824 8128
rect 9765 7986 9831 7989
rect 11237 7986 11303 7989
rect 9765 7984 11303 7986
rect 9765 7928 9770 7984
rect 9826 7928 11242 7984
rect 11298 7928 11303 7984
rect 9765 7926 11303 7928
rect 9765 7923 9831 7926
rect 11237 7923 11303 7926
rect 10409 7850 10475 7853
rect 11789 7850 11855 7853
rect 10409 7848 11855 7850
rect 10409 7792 10414 7848
rect 10470 7792 11794 7848
rect 11850 7792 11855 7848
rect 10409 7790 11855 7792
rect 10409 7787 10475 7790
rect 11789 7787 11855 7790
rect 4654 7648 4974 7649
rect 4654 7584 4662 7648
rect 4726 7584 4742 7648
rect 4806 7584 4822 7648
rect 4886 7584 4902 7648
rect 4966 7584 4974 7648
rect 4654 7583 4974 7584
rect 7754 7648 8074 7649
rect 7754 7584 7762 7648
rect 7826 7584 7842 7648
rect 7906 7584 7922 7648
rect 7986 7584 8002 7648
rect 8066 7584 8074 7648
rect 7754 7583 8074 7584
rect 10854 7648 11174 7649
rect 10854 7584 10862 7648
rect 10926 7584 10942 7648
rect 11006 7584 11022 7648
rect 11086 7584 11102 7648
rect 11166 7584 11174 7648
rect 10854 7583 11174 7584
rect 13954 7648 14274 7649
rect 13954 7584 13962 7648
rect 14026 7584 14042 7648
rect 14106 7584 14122 7648
rect 14186 7584 14202 7648
rect 14266 7584 14274 7648
rect 13954 7583 14274 7584
rect 17054 7648 17374 7649
rect 17054 7584 17062 7648
rect 17126 7584 17142 7648
rect 17206 7584 17222 7648
rect 17286 7584 17302 7648
rect 17366 7584 17374 7648
rect 17054 7583 17374 7584
rect 10133 7306 10199 7309
rect 13537 7306 13603 7309
rect 10133 7304 13603 7306
rect 10133 7248 10138 7304
rect 10194 7248 13542 7304
rect 13598 7248 13603 7304
rect 10133 7246 13603 7248
rect 10133 7243 10199 7246
rect 13537 7243 13603 7246
rect 3104 7104 3424 7105
rect 3104 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3272 7104
rect 3336 7040 3352 7104
rect 3416 7040 3424 7104
rect 3104 7039 3424 7040
rect 6204 7104 6524 7105
rect 6204 7040 6212 7104
rect 6276 7040 6292 7104
rect 6356 7040 6372 7104
rect 6436 7040 6452 7104
rect 6516 7040 6524 7104
rect 6204 7039 6524 7040
rect 9304 7104 9624 7105
rect 9304 7040 9312 7104
rect 9376 7040 9392 7104
rect 9456 7040 9472 7104
rect 9536 7040 9552 7104
rect 9616 7040 9624 7104
rect 9304 7039 9624 7040
rect 12404 7104 12724 7105
rect 12404 7040 12412 7104
rect 12476 7040 12492 7104
rect 12556 7040 12572 7104
rect 12636 7040 12652 7104
rect 12716 7040 12724 7104
rect 12404 7039 12724 7040
rect 15504 7104 15824 7105
rect 15504 7040 15512 7104
rect 15576 7040 15592 7104
rect 15656 7040 15672 7104
rect 15736 7040 15752 7104
rect 15816 7040 15824 7104
rect 15504 7039 15824 7040
rect 10133 7034 10199 7037
rect 11881 7034 11947 7037
rect 10133 7032 11947 7034
rect 10133 6976 10138 7032
rect 10194 6976 11886 7032
rect 11942 6976 11947 7032
rect 10133 6974 11947 6976
rect 10133 6971 10199 6974
rect 11881 6971 11947 6974
rect 9949 6762 10015 6765
rect 11513 6762 11579 6765
rect 9949 6760 11579 6762
rect 9949 6704 9954 6760
rect 10010 6704 11518 6760
rect 11574 6704 11579 6760
rect 9949 6702 11579 6704
rect 9949 6699 10015 6702
rect 11513 6699 11579 6702
rect 18505 6762 18571 6765
rect 19200 6762 20000 6792
rect 18505 6760 20000 6762
rect 18505 6704 18510 6760
rect 18566 6704 20000 6760
rect 18505 6702 20000 6704
rect 18505 6699 18571 6702
rect 19200 6672 20000 6702
rect 4654 6560 4974 6561
rect 4654 6496 4662 6560
rect 4726 6496 4742 6560
rect 4806 6496 4822 6560
rect 4886 6496 4902 6560
rect 4966 6496 4974 6560
rect 4654 6495 4974 6496
rect 7754 6560 8074 6561
rect 7754 6496 7762 6560
rect 7826 6496 7842 6560
rect 7906 6496 7922 6560
rect 7986 6496 8002 6560
rect 8066 6496 8074 6560
rect 7754 6495 8074 6496
rect 10854 6560 11174 6561
rect 10854 6496 10862 6560
rect 10926 6496 10942 6560
rect 11006 6496 11022 6560
rect 11086 6496 11102 6560
rect 11166 6496 11174 6560
rect 10854 6495 11174 6496
rect 13954 6560 14274 6561
rect 13954 6496 13962 6560
rect 14026 6496 14042 6560
rect 14106 6496 14122 6560
rect 14186 6496 14202 6560
rect 14266 6496 14274 6560
rect 13954 6495 14274 6496
rect 17054 6560 17374 6561
rect 17054 6496 17062 6560
rect 17126 6496 17142 6560
rect 17206 6496 17222 6560
rect 17286 6496 17302 6560
rect 17366 6496 17374 6560
rect 17054 6495 17374 6496
rect 3104 6016 3424 6017
rect 3104 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3272 6016
rect 3336 5952 3352 6016
rect 3416 5952 3424 6016
rect 3104 5951 3424 5952
rect 6204 6016 6524 6017
rect 6204 5952 6212 6016
rect 6276 5952 6292 6016
rect 6356 5952 6372 6016
rect 6436 5952 6452 6016
rect 6516 5952 6524 6016
rect 6204 5951 6524 5952
rect 9304 6016 9624 6017
rect 9304 5952 9312 6016
rect 9376 5952 9392 6016
rect 9456 5952 9472 6016
rect 9536 5952 9552 6016
rect 9616 5952 9624 6016
rect 9304 5951 9624 5952
rect 12404 6016 12724 6017
rect 12404 5952 12412 6016
rect 12476 5952 12492 6016
rect 12556 5952 12572 6016
rect 12636 5952 12652 6016
rect 12716 5952 12724 6016
rect 12404 5951 12724 5952
rect 15504 6016 15824 6017
rect 15504 5952 15512 6016
rect 15576 5952 15592 6016
rect 15656 5952 15672 6016
rect 15736 5952 15752 6016
rect 15816 5952 15824 6016
rect 15504 5951 15824 5952
rect 4654 5472 4974 5473
rect 4654 5408 4662 5472
rect 4726 5408 4742 5472
rect 4806 5408 4822 5472
rect 4886 5408 4902 5472
rect 4966 5408 4974 5472
rect 4654 5407 4974 5408
rect 7754 5472 8074 5473
rect 7754 5408 7762 5472
rect 7826 5408 7842 5472
rect 7906 5408 7922 5472
rect 7986 5408 8002 5472
rect 8066 5408 8074 5472
rect 7754 5407 8074 5408
rect 10854 5472 11174 5473
rect 10854 5408 10862 5472
rect 10926 5408 10942 5472
rect 11006 5408 11022 5472
rect 11086 5408 11102 5472
rect 11166 5408 11174 5472
rect 10854 5407 11174 5408
rect 13954 5472 14274 5473
rect 13954 5408 13962 5472
rect 14026 5408 14042 5472
rect 14106 5408 14122 5472
rect 14186 5408 14202 5472
rect 14266 5408 14274 5472
rect 13954 5407 14274 5408
rect 17054 5472 17374 5473
rect 17054 5408 17062 5472
rect 17126 5408 17142 5472
rect 17206 5408 17222 5472
rect 17286 5408 17302 5472
rect 17366 5408 17374 5472
rect 17054 5407 17374 5408
rect 7465 5266 7531 5269
rect 8937 5266 9003 5269
rect 7465 5264 9003 5266
rect 7465 5208 7470 5264
rect 7526 5208 8942 5264
rect 8998 5208 9003 5264
rect 7465 5206 9003 5208
rect 7465 5203 7531 5206
rect 8937 5203 9003 5206
rect 18505 5266 18571 5269
rect 19200 5266 20000 5296
rect 18505 5264 20000 5266
rect 18505 5208 18510 5264
rect 18566 5208 20000 5264
rect 18505 5206 20000 5208
rect 18505 5203 18571 5206
rect 19200 5176 20000 5206
rect 3104 4928 3424 4929
rect 3104 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3272 4928
rect 3336 4864 3352 4928
rect 3416 4864 3424 4928
rect 3104 4863 3424 4864
rect 6204 4928 6524 4929
rect 6204 4864 6212 4928
rect 6276 4864 6292 4928
rect 6356 4864 6372 4928
rect 6436 4864 6452 4928
rect 6516 4864 6524 4928
rect 6204 4863 6524 4864
rect 9304 4928 9624 4929
rect 9304 4864 9312 4928
rect 9376 4864 9392 4928
rect 9456 4864 9472 4928
rect 9536 4864 9552 4928
rect 9616 4864 9624 4928
rect 9304 4863 9624 4864
rect 12404 4928 12724 4929
rect 12404 4864 12412 4928
rect 12476 4864 12492 4928
rect 12556 4864 12572 4928
rect 12636 4864 12652 4928
rect 12716 4864 12724 4928
rect 12404 4863 12724 4864
rect 15504 4928 15824 4929
rect 15504 4864 15512 4928
rect 15576 4864 15592 4928
rect 15656 4864 15672 4928
rect 15736 4864 15752 4928
rect 15816 4864 15824 4928
rect 15504 4863 15824 4864
rect 9673 4586 9739 4589
rect 11329 4586 11395 4589
rect 9673 4584 11395 4586
rect 9673 4528 9678 4584
rect 9734 4528 11334 4584
rect 11390 4528 11395 4584
rect 9673 4526 11395 4528
rect 9673 4523 9739 4526
rect 11329 4523 11395 4526
rect 4654 4384 4974 4385
rect 4654 4320 4662 4384
rect 4726 4320 4742 4384
rect 4806 4320 4822 4384
rect 4886 4320 4902 4384
rect 4966 4320 4974 4384
rect 4654 4319 4974 4320
rect 7754 4384 8074 4385
rect 7754 4320 7762 4384
rect 7826 4320 7842 4384
rect 7906 4320 7922 4384
rect 7986 4320 8002 4384
rect 8066 4320 8074 4384
rect 7754 4319 8074 4320
rect 10854 4384 11174 4385
rect 10854 4320 10862 4384
rect 10926 4320 10942 4384
rect 11006 4320 11022 4384
rect 11086 4320 11102 4384
rect 11166 4320 11174 4384
rect 10854 4319 11174 4320
rect 13954 4384 14274 4385
rect 13954 4320 13962 4384
rect 14026 4320 14042 4384
rect 14106 4320 14122 4384
rect 14186 4320 14202 4384
rect 14266 4320 14274 4384
rect 13954 4319 14274 4320
rect 17054 4384 17374 4385
rect 17054 4320 17062 4384
rect 17126 4320 17142 4384
rect 17206 4320 17222 4384
rect 17286 4320 17302 4384
rect 17366 4320 17374 4384
rect 17054 4319 17374 4320
rect 3104 3840 3424 3841
rect 3104 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3272 3840
rect 3336 3776 3352 3840
rect 3416 3776 3424 3840
rect 3104 3775 3424 3776
rect 6204 3840 6524 3841
rect 6204 3776 6212 3840
rect 6276 3776 6292 3840
rect 6356 3776 6372 3840
rect 6436 3776 6452 3840
rect 6516 3776 6524 3840
rect 6204 3775 6524 3776
rect 9304 3840 9624 3841
rect 9304 3776 9312 3840
rect 9376 3776 9392 3840
rect 9456 3776 9472 3840
rect 9536 3776 9552 3840
rect 9616 3776 9624 3840
rect 9304 3775 9624 3776
rect 12404 3840 12724 3841
rect 12404 3776 12412 3840
rect 12476 3776 12492 3840
rect 12556 3776 12572 3840
rect 12636 3776 12652 3840
rect 12716 3776 12724 3840
rect 12404 3775 12724 3776
rect 15504 3840 15824 3841
rect 15504 3776 15512 3840
rect 15576 3776 15592 3840
rect 15656 3776 15672 3840
rect 15736 3776 15752 3840
rect 15816 3776 15824 3840
rect 15504 3775 15824 3776
rect 18505 3770 18571 3773
rect 19200 3770 20000 3800
rect 18505 3768 20000 3770
rect 18505 3712 18510 3768
rect 18566 3712 20000 3768
rect 18505 3710 20000 3712
rect 18505 3707 18571 3710
rect 19200 3680 20000 3710
rect 3877 3498 3943 3501
rect 4061 3498 4127 3501
rect 3877 3496 4127 3498
rect 3877 3440 3882 3496
rect 3938 3440 4066 3496
rect 4122 3440 4127 3496
rect 3877 3438 4127 3440
rect 3877 3435 3943 3438
rect 4061 3435 4127 3438
rect 4654 3296 4974 3297
rect 4654 3232 4662 3296
rect 4726 3232 4742 3296
rect 4806 3232 4822 3296
rect 4886 3232 4902 3296
rect 4966 3232 4974 3296
rect 4654 3231 4974 3232
rect 7754 3296 8074 3297
rect 7754 3232 7762 3296
rect 7826 3232 7842 3296
rect 7906 3232 7922 3296
rect 7986 3232 8002 3296
rect 8066 3232 8074 3296
rect 7754 3231 8074 3232
rect 10854 3296 11174 3297
rect 10854 3232 10862 3296
rect 10926 3232 10942 3296
rect 11006 3232 11022 3296
rect 11086 3232 11102 3296
rect 11166 3232 11174 3296
rect 10854 3231 11174 3232
rect 13954 3296 14274 3297
rect 13954 3232 13962 3296
rect 14026 3232 14042 3296
rect 14106 3232 14122 3296
rect 14186 3232 14202 3296
rect 14266 3232 14274 3296
rect 13954 3231 14274 3232
rect 17054 3296 17374 3297
rect 17054 3232 17062 3296
rect 17126 3232 17142 3296
rect 17206 3232 17222 3296
rect 17286 3232 17302 3296
rect 17366 3232 17374 3296
rect 17054 3231 17374 3232
rect 4797 3090 4863 3093
rect 6729 3090 6795 3093
rect 4797 3088 6795 3090
rect 4797 3032 4802 3088
rect 4858 3032 6734 3088
rect 6790 3032 6795 3088
rect 4797 3030 6795 3032
rect 4797 3027 4863 3030
rect 6729 3027 6795 3030
rect 3104 2752 3424 2753
rect 3104 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3272 2752
rect 3336 2688 3352 2752
rect 3416 2688 3424 2752
rect 3104 2687 3424 2688
rect 6204 2752 6524 2753
rect 6204 2688 6212 2752
rect 6276 2688 6292 2752
rect 6356 2688 6372 2752
rect 6436 2688 6452 2752
rect 6516 2688 6524 2752
rect 6204 2687 6524 2688
rect 9304 2752 9624 2753
rect 9304 2688 9312 2752
rect 9376 2688 9392 2752
rect 9456 2688 9472 2752
rect 9536 2688 9552 2752
rect 9616 2688 9624 2752
rect 9304 2687 9624 2688
rect 12404 2752 12724 2753
rect 12404 2688 12412 2752
rect 12476 2688 12492 2752
rect 12556 2688 12572 2752
rect 12636 2688 12652 2752
rect 12716 2688 12724 2752
rect 12404 2687 12724 2688
rect 15504 2752 15824 2753
rect 15504 2688 15512 2752
rect 15576 2688 15592 2752
rect 15656 2688 15672 2752
rect 15736 2688 15752 2752
rect 15816 2688 15824 2752
rect 15504 2687 15824 2688
rect 18505 2274 18571 2277
rect 19200 2274 20000 2304
rect 18505 2272 20000 2274
rect 18505 2216 18510 2272
rect 18566 2216 20000 2272
rect 18505 2214 20000 2216
rect 18505 2211 18571 2214
rect 4654 2208 4974 2209
rect 4654 2144 4662 2208
rect 4726 2144 4742 2208
rect 4806 2144 4822 2208
rect 4886 2144 4902 2208
rect 4966 2144 4974 2208
rect 4654 2143 4974 2144
rect 7754 2208 8074 2209
rect 7754 2144 7762 2208
rect 7826 2144 7842 2208
rect 7906 2144 7922 2208
rect 7986 2144 8002 2208
rect 8066 2144 8074 2208
rect 7754 2143 8074 2144
rect 10854 2208 11174 2209
rect 10854 2144 10862 2208
rect 10926 2144 10942 2208
rect 11006 2144 11022 2208
rect 11086 2144 11102 2208
rect 11166 2144 11174 2208
rect 10854 2143 11174 2144
rect 13954 2208 14274 2209
rect 13954 2144 13962 2208
rect 14026 2144 14042 2208
rect 14106 2144 14122 2208
rect 14186 2144 14202 2208
rect 14266 2144 14274 2208
rect 13954 2143 14274 2144
rect 17054 2208 17374 2209
rect 17054 2144 17062 2208
rect 17126 2144 17142 2208
rect 17206 2144 17222 2208
rect 17286 2144 17302 2208
rect 17366 2144 17374 2208
rect 19200 2184 20000 2214
rect 17054 2143 17374 2144
rect 3104 1664 3424 1665
rect 3104 1600 3112 1664
rect 3176 1600 3192 1664
rect 3256 1600 3272 1664
rect 3336 1600 3352 1664
rect 3416 1600 3424 1664
rect 3104 1599 3424 1600
rect 6204 1664 6524 1665
rect 6204 1600 6212 1664
rect 6276 1600 6292 1664
rect 6356 1600 6372 1664
rect 6436 1600 6452 1664
rect 6516 1600 6524 1664
rect 6204 1599 6524 1600
rect 9304 1664 9624 1665
rect 9304 1600 9312 1664
rect 9376 1600 9392 1664
rect 9456 1600 9472 1664
rect 9536 1600 9552 1664
rect 9616 1600 9624 1664
rect 9304 1599 9624 1600
rect 12404 1664 12724 1665
rect 12404 1600 12412 1664
rect 12476 1600 12492 1664
rect 12556 1600 12572 1664
rect 12636 1600 12652 1664
rect 12716 1600 12724 1664
rect 12404 1599 12724 1600
rect 15504 1664 15824 1665
rect 15504 1600 15512 1664
rect 15576 1600 15592 1664
rect 15656 1600 15672 1664
rect 15736 1600 15752 1664
rect 15816 1600 15824 1664
rect 15504 1599 15824 1600
rect 4654 1120 4974 1121
rect 4654 1056 4662 1120
rect 4726 1056 4742 1120
rect 4806 1056 4822 1120
rect 4886 1056 4902 1120
rect 4966 1056 4974 1120
rect 4654 1055 4974 1056
rect 7754 1120 8074 1121
rect 7754 1056 7762 1120
rect 7826 1056 7842 1120
rect 7906 1056 7922 1120
rect 7986 1056 8002 1120
rect 8066 1056 8074 1120
rect 7754 1055 8074 1056
rect 10854 1120 11174 1121
rect 10854 1056 10862 1120
rect 10926 1056 10942 1120
rect 11006 1056 11022 1120
rect 11086 1056 11102 1120
rect 11166 1056 11174 1120
rect 10854 1055 11174 1056
rect 13954 1120 14274 1121
rect 13954 1056 13962 1120
rect 14026 1056 14042 1120
rect 14106 1056 14122 1120
rect 14186 1056 14202 1120
rect 14266 1056 14274 1120
rect 13954 1055 14274 1056
rect 17054 1120 17374 1121
rect 17054 1056 17062 1120
rect 17126 1056 17142 1120
rect 17206 1056 17222 1120
rect 17286 1056 17302 1120
rect 17366 1056 17374 1120
rect 17054 1055 17374 1056
rect 18505 778 18571 781
rect 19200 778 20000 808
rect 18505 776 20000 778
rect 18505 720 18510 776
rect 18566 720 20000 776
rect 18505 718 20000 720
rect 18505 715 18571 718
rect 19200 688 20000 718
rect 3104 576 3424 577
rect 3104 512 3112 576
rect 3176 512 3192 576
rect 3256 512 3272 576
rect 3336 512 3352 576
rect 3416 512 3424 576
rect 3104 511 3424 512
rect 6204 576 6524 577
rect 6204 512 6212 576
rect 6276 512 6292 576
rect 6356 512 6372 576
rect 6436 512 6452 576
rect 6516 512 6524 576
rect 6204 511 6524 512
rect 9304 576 9624 577
rect 9304 512 9312 576
rect 9376 512 9392 576
rect 9456 512 9472 576
rect 9536 512 9552 576
rect 9616 512 9624 576
rect 9304 511 9624 512
rect 12404 576 12724 577
rect 12404 512 12412 576
rect 12476 512 12492 576
rect 12556 512 12572 576
rect 12636 512 12652 576
rect 12716 512 12724 576
rect 12404 511 12724 512
rect 15504 576 15824 577
rect 15504 512 15512 576
rect 15576 512 15592 576
rect 15656 512 15672 576
rect 15736 512 15752 576
rect 15816 512 15824 576
rect 15504 511 15824 512
rect 4654 32 4974 33
rect 4654 -32 4662 32
rect 4726 -32 4742 32
rect 4806 -32 4822 32
rect 4886 -32 4902 32
rect 4966 -32 4974 32
rect 4654 -33 4974 -32
rect 7754 32 8074 33
rect 7754 -32 7762 32
rect 7826 -32 7842 32
rect 7906 -32 7922 32
rect 7986 -32 8002 32
rect 8066 -32 8074 32
rect 7754 -33 8074 -32
rect 10854 32 11174 33
rect 10854 -32 10862 32
rect 10926 -32 10942 32
rect 11006 -32 11022 32
rect 11086 -32 11102 32
rect 11166 -32 11174 32
rect 10854 -33 11174 -32
rect 13954 32 14274 33
rect 13954 -32 13962 32
rect 14026 -32 14042 32
rect 14106 -32 14122 32
rect 14186 -32 14202 32
rect 14266 -32 14274 32
rect 13954 -33 14274 -32
rect 17054 32 17374 33
rect 17054 -32 17062 32
rect 17126 -32 17142 32
rect 17206 -32 17222 32
rect 17286 -32 17302 32
rect 17366 -32 17374 32
rect 17054 -33 17374 -32
<< via3 >>
rect 4662 10908 4726 10912
rect 4662 10852 4666 10908
rect 4666 10852 4722 10908
rect 4722 10852 4726 10908
rect 4662 10848 4726 10852
rect 4742 10908 4806 10912
rect 4742 10852 4746 10908
rect 4746 10852 4802 10908
rect 4802 10852 4806 10908
rect 4742 10848 4806 10852
rect 4822 10908 4886 10912
rect 4822 10852 4826 10908
rect 4826 10852 4882 10908
rect 4882 10852 4886 10908
rect 4822 10848 4886 10852
rect 4902 10908 4966 10912
rect 4902 10852 4906 10908
rect 4906 10852 4962 10908
rect 4962 10852 4966 10908
rect 4902 10848 4966 10852
rect 7762 10908 7826 10912
rect 7762 10852 7766 10908
rect 7766 10852 7822 10908
rect 7822 10852 7826 10908
rect 7762 10848 7826 10852
rect 7842 10908 7906 10912
rect 7842 10852 7846 10908
rect 7846 10852 7902 10908
rect 7902 10852 7906 10908
rect 7842 10848 7906 10852
rect 7922 10908 7986 10912
rect 7922 10852 7926 10908
rect 7926 10852 7982 10908
rect 7982 10852 7986 10908
rect 7922 10848 7986 10852
rect 8002 10908 8066 10912
rect 8002 10852 8006 10908
rect 8006 10852 8062 10908
rect 8062 10852 8066 10908
rect 8002 10848 8066 10852
rect 10862 10908 10926 10912
rect 10862 10852 10866 10908
rect 10866 10852 10922 10908
rect 10922 10852 10926 10908
rect 10862 10848 10926 10852
rect 10942 10908 11006 10912
rect 10942 10852 10946 10908
rect 10946 10852 11002 10908
rect 11002 10852 11006 10908
rect 10942 10848 11006 10852
rect 11022 10908 11086 10912
rect 11022 10852 11026 10908
rect 11026 10852 11082 10908
rect 11082 10852 11086 10908
rect 11022 10848 11086 10852
rect 11102 10908 11166 10912
rect 11102 10852 11106 10908
rect 11106 10852 11162 10908
rect 11162 10852 11166 10908
rect 11102 10848 11166 10852
rect 13962 10908 14026 10912
rect 13962 10852 13966 10908
rect 13966 10852 14022 10908
rect 14022 10852 14026 10908
rect 13962 10848 14026 10852
rect 14042 10908 14106 10912
rect 14042 10852 14046 10908
rect 14046 10852 14102 10908
rect 14102 10852 14106 10908
rect 14042 10848 14106 10852
rect 14122 10908 14186 10912
rect 14122 10852 14126 10908
rect 14126 10852 14182 10908
rect 14182 10852 14186 10908
rect 14122 10848 14186 10852
rect 14202 10908 14266 10912
rect 14202 10852 14206 10908
rect 14206 10852 14262 10908
rect 14262 10852 14266 10908
rect 14202 10848 14266 10852
rect 17062 10908 17126 10912
rect 17062 10852 17066 10908
rect 17066 10852 17122 10908
rect 17122 10852 17126 10908
rect 17062 10848 17126 10852
rect 17142 10908 17206 10912
rect 17142 10852 17146 10908
rect 17146 10852 17202 10908
rect 17202 10852 17206 10908
rect 17142 10848 17206 10852
rect 17222 10908 17286 10912
rect 17222 10852 17226 10908
rect 17226 10852 17282 10908
rect 17282 10852 17286 10908
rect 17222 10848 17286 10852
rect 17302 10908 17366 10912
rect 17302 10852 17306 10908
rect 17306 10852 17362 10908
rect 17362 10852 17366 10908
rect 17302 10848 17366 10852
rect 3112 10364 3176 10368
rect 3112 10308 3116 10364
rect 3116 10308 3172 10364
rect 3172 10308 3176 10364
rect 3112 10304 3176 10308
rect 3192 10364 3256 10368
rect 3192 10308 3196 10364
rect 3196 10308 3252 10364
rect 3252 10308 3256 10364
rect 3192 10304 3256 10308
rect 3272 10364 3336 10368
rect 3272 10308 3276 10364
rect 3276 10308 3332 10364
rect 3332 10308 3336 10364
rect 3272 10304 3336 10308
rect 3352 10364 3416 10368
rect 3352 10308 3356 10364
rect 3356 10308 3412 10364
rect 3412 10308 3416 10364
rect 3352 10304 3416 10308
rect 6212 10364 6276 10368
rect 6212 10308 6216 10364
rect 6216 10308 6272 10364
rect 6272 10308 6276 10364
rect 6212 10304 6276 10308
rect 6292 10364 6356 10368
rect 6292 10308 6296 10364
rect 6296 10308 6352 10364
rect 6352 10308 6356 10364
rect 6292 10304 6356 10308
rect 6372 10364 6436 10368
rect 6372 10308 6376 10364
rect 6376 10308 6432 10364
rect 6432 10308 6436 10364
rect 6372 10304 6436 10308
rect 6452 10364 6516 10368
rect 6452 10308 6456 10364
rect 6456 10308 6512 10364
rect 6512 10308 6516 10364
rect 6452 10304 6516 10308
rect 9312 10364 9376 10368
rect 9312 10308 9316 10364
rect 9316 10308 9372 10364
rect 9372 10308 9376 10364
rect 9312 10304 9376 10308
rect 9392 10364 9456 10368
rect 9392 10308 9396 10364
rect 9396 10308 9452 10364
rect 9452 10308 9456 10364
rect 9392 10304 9456 10308
rect 9472 10364 9536 10368
rect 9472 10308 9476 10364
rect 9476 10308 9532 10364
rect 9532 10308 9536 10364
rect 9472 10304 9536 10308
rect 9552 10364 9616 10368
rect 9552 10308 9556 10364
rect 9556 10308 9612 10364
rect 9612 10308 9616 10364
rect 9552 10304 9616 10308
rect 12412 10364 12476 10368
rect 12412 10308 12416 10364
rect 12416 10308 12472 10364
rect 12472 10308 12476 10364
rect 12412 10304 12476 10308
rect 12492 10364 12556 10368
rect 12492 10308 12496 10364
rect 12496 10308 12552 10364
rect 12552 10308 12556 10364
rect 12492 10304 12556 10308
rect 12572 10364 12636 10368
rect 12572 10308 12576 10364
rect 12576 10308 12632 10364
rect 12632 10308 12636 10364
rect 12572 10304 12636 10308
rect 12652 10364 12716 10368
rect 12652 10308 12656 10364
rect 12656 10308 12712 10364
rect 12712 10308 12716 10364
rect 12652 10304 12716 10308
rect 15512 10364 15576 10368
rect 15512 10308 15516 10364
rect 15516 10308 15572 10364
rect 15572 10308 15576 10364
rect 15512 10304 15576 10308
rect 15592 10364 15656 10368
rect 15592 10308 15596 10364
rect 15596 10308 15652 10364
rect 15652 10308 15656 10364
rect 15592 10304 15656 10308
rect 15672 10364 15736 10368
rect 15672 10308 15676 10364
rect 15676 10308 15732 10364
rect 15732 10308 15736 10364
rect 15672 10304 15736 10308
rect 15752 10364 15816 10368
rect 15752 10308 15756 10364
rect 15756 10308 15812 10364
rect 15812 10308 15816 10364
rect 15752 10304 15816 10308
rect 4662 9820 4726 9824
rect 4662 9764 4666 9820
rect 4666 9764 4722 9820
rect 4722 9764 4726 9820
rect 4662 9760 4726 9764
rect 4742 9820 4806 9824
rect 4742 9764 4746 9820
rect 4746 9764 4802 9820
rect 4802 9764 4806 9820
rect 4742 9760 4806 9764
rect 4822 9820 4886 9824
rect 4822 9764 4826 9820
rect 4826 9764 4882 9820
rect 4882 9764 4886 9820
rect 4822 9760 4886 9764
rect 4902 9820 4966 9824
rect 4902 9764 4906 9820
rect 4906 9764 4962 9820
rect 4962 9764 4966 9820
rect 4902 9760 4966 9764
rect 7762 9820 7826 9824
rect 7762 9764 7766 9820
rect 7766 9764 7822 9820
rect 7822 9764 7826 9820
rect 7762 9760 7826 9764
rect 7842 9820 7906 9824
rect 7842 9764 7846 9820
rect 7846 9764 7902 9820
rect 7902 9764 7906 9820
rect 7842 9760 7906 9764
rect 7922 9820 7986 9824
rect 7922 9764 7926 9820
rect 7926 9764 7982 9820
rect 7982 9764 7986 9820
rect 7922 9760 7986 9764
rect 8002 9820 8066 9824
rect 8002 9764 8006 9820
rect 8006 9764 8062 9820
rect 8062 9764 8066 9820
rect 8002 9760 8066 9764
rect 10862 9820 10926 9824
rect 10862 9764 10866 9820
rect 10866 9764 10922 9820
rect 10922 9764 10926 9820
rect 10862 9760 10926 9764
rect 10942 9820 11006 9824
rect 10942 9764 10946 9820
rect 10946 9764 11002 9820
rect 11002 9764 11006 9820
rect 10942 9760 11006 9764
rect 11022 9820 11086 9824
rect 11022 9764 11026 9820
rect 11026 9764 11082 9820
rect 11082 9764 11086 9820
rect 11022 9760 11086 9764
rect 11102 9820 11166 9824
rect 11102 9764 11106 9820
rect 11106 9764 11162 9820
rect 11162 9764 11166 9820
rect 11102 9760 11166 9764
rect 13962 9820 14026 9824
rect 13962 9764 13966 9820
rect 13966 9764 14022 9820
rect 14022 9764 14026 9820
rect 13962 9760 14026 9764
rect 14042 9820 14106 9824
rect 14042 9764 14046 9820
rect 14046 9764 14102 9820
rect 14102 9764 14106 9820
rect 14042 9760 14106 9764
rect 14122 9820 14186 9824
rect 14122 9764 14126 9820
rect 14126 9764 14182 9820
rect 14182 9764 14186 9820
rect 14122 9760 14186 9764
rect 14202 9820 14266 9824
rect 14202 9764 14206 9820
rect 14206 9764 14262 9820
rect 14262 9764 14266 9820
rect 14202 9760 14266 9764
rect 17062 9820 17126 9824
rect 17062 9764 17066 9820
rect 17066 9764 17122 9820
rect 17122 9764 17126 9820
rect 17062 9760 17126 9764
rect 17142 9820 17206 9824
rect 17142 9764 17146 9820
rect 17146 9764 17202 9820
rect 17202 9764 17206 9820
rect 17142 9760 17206 9764
rect 17222 9820 17286 9824
rect 17222 9764 17226 9820
rect 17226 9764 17282 9820
rect 17282 9764 17286 9820
rect 17222 9760 17286 9764
rect 17302 9820 17366 9824
rect 17302 9764 17306 9820
rect 17306 9764 17362 9820
rect 17362 9764 17366 9820
rect 17302 9760 17366 9764
rect 3112 9276 3176 9280
rect 3112 9220 3116 9276
rect 3116 9220 3172 9276
rect 3172 9220 3176 9276
rect 3112 9216 3176 9220
rect 3192 9276 3256 9280
rect 3192 9220 3196 9276
rect 3196 9220 3252 9276
rect 3252 9220 3256 9276
rect 3192 9216 3256 9220
rect 3272 9276 3336 9280
rect 3272 9220 3276 9276
rect 3276 9220 3332 9276
rect 3332 9220 3336 9276
rect 3272 9216 3336 9220
rect 3352 9276 3416 9280
rect 3352 9220 3356 9276
rect 3356 9220 3412 9276
rect 3412 9220 3416 9276
rect 3352 9216 3416 9220
rect 6212 9276 6276 9280
rect 6212 9220 6216 9276
rect 6216 9220 6272 9276
rect 6272 9220 6276 9276
rect 6212 9216 6276 9220
rect 6292 9276 6356 9280
rect 6292 9220 6296 9276
rect 6296 9220 6352 9276
rect 6352 9220 6356 9276
rect 6292 9216 6356 9220
rect 6372 9276 6436 9280
rect 6372 9220 6376 9276
rect 6376 9220 6432 9276
rect 6432 9220 6436 9276
rect 6372 9216 6436 9220
rect 6452 9276 6516 9280
rect 6452 9220 6456 9276
rect 6456 9220 6512 9276
rect 6512 9220 6516 9276
rect 6452 9216 6516 9220
rect 9312 9276 9376 9280
rect 9312 9220 9316 9276
rect 9316 9220 9372 9276
rect 9372 9220 9376 9276
rect 9312 9216 9376 9220
rect 9392 9276 9456 9280
rect 9392 9220 9396 9276
rect 9396 9220 9452 9276
rect 9452 9220 9456 9276
rect 9392 9216 9456 9220
rect 9472 9276 9536 9280
rect 9472 9220 9476 9276
rect 9476 9220 9532 9276
rect 9532 9220 9536 9276
rect 9472 9216 9536 9220
rect 9552 9276 9616 9280
rect 9552 9220 9556 9276
rect 9556 9220 9612 9276
rect 9612 9220 9616 9276
rect 9552 9216 9616 9220
rect 12412 9276 12476 9280
rect 12412 9220 12416 9276
rect 12416 9220 12472 9276
rect 12472 9220 12476 9276
rect 12412 9216 12476 9220
rect 12492 9276 12556 9280
rect 12492 9220 12496 9276
rect 12496 9220 12552 9276
rect 12552 9220 12556 9276
rect 12492 9216 12556 9220
rect 12572 9276 12636 9280
rect 12572 9220 12576 9276
rect 12576 9220 12632 9276
rect 12632 9220 12636 9276
rect 12572 9216 12636 9220
rect 12652 9276 12716 9280
rect 12652 9220 12656 9276
rect 12656 9220 12712 9276
rect 12712 9220 12716 9276
rect 12652 9216 12716 9220
rect 15512 9276 15576 9280
rect 15512 9220 15516 9276
rect 15516 9220 15572 9276
rect 15572 9220 15576 9276
rect 15512 9216 15576 9220
rect 15592 9276 15656 9280
rect 15592 9220 15596 9276
rect 15596 9220 15652 9276
rect 15652 9220 15656 9276
rect 15592 9216 15656 9220
rect 15672 9276 15736 9280
rect 15672 9220 15676 9276
rect 15676 9220 15732 9276
rect 15732 9220 15736 9276
rect 15672 9216 15736 9220
rect 15752 9276 15816 9280
rect 15752 9220 15756 9276
rect 15756 9220 15812 9276
rect 15812 9220 15816 9276
rect 15752 9216 15816 9220
rect 4662 8732 4726 8736
rect 4662 8676 4666 8732
rect 4666 8676 4722 8732
rect 4722 8676 4726 8732
rect 4662 8672 4726 8676
rect 4742 8732 4806 8736
rect 4742 8676 4746 8732
rect 4746 8676 4802 8732
rect 4802 8676 4806 8732
rect 4742 8672 4806 8676
rect 4822 8732 4886 8736
rect 4822 8676 4826 8732
rect 4826 8676 4882 8732
rect 4882 8676 4886 8732
rect 4822 8672 4886 8676
rect 4902 8732 4966 8736
rect 4902 8676 4906 8732
rect 4906 8676 4962 8732
rect 4962 8676 4966 8732
rect 4902 8672 4966 8676
rect 7762 8732 7826 8736
rect 7762 8676 7766 8732
rect 7766 8676 7822 8732
rect 7822 8676 7826 8732
rect 7762 8672 7826 8676
rect 7842 8732 7906 8736
rect 7842 8676 7846 8732
rect 7846 8676 7902 8732
rect 7902 8676 7906 8732
rect 7842 8672 7906 8676
rect 7922 8732 7986 8736
rect 7922 8676 7926 8732
rect 7926 8676 7982 8732
rect 7982 8676 7986 8732
rect 7922 8672 7986 8676
rect 8002 8732 8066 8736
rect 8002 8676 8006 8732
rect 8006 8676 8062 8732
rect 8062 8676 8066 8732
rect 8002 8672 8066 8676
rect 10862 8732 10926 8736
rect 10862 8676 10866 8732
rect 10866 8676 10922 8732
rect 10922 8676 10926 8732
rect 10862 8672 10926 8676
rect 10942 8732 11006 8736
rect 10942 8676 10946 8732
rect 10946 8676 11002 8732
rect 11002 8676 11006 8732
rect 10942 8672 11006 8676
rect 11022 8732 11086 8736
rect 11022 8676 11026 8732
rect 11026 8676 11082 8732
rect 11082 8676 11086 8732
rect 11022 8672 11086 8676
rect 11102 8732 11166 8736
rect 11102 8676 11106 8732
rect 11106 8676 11162 8732
rect 11162 8676 11166 8732
rect 11102 8672 11166 8676
rect 13962 8732 14026 8736
rect 13962 8676 13966 8732
rect 13966 8676 14022 8732
rect 14022 8676 14026 8732
rect 13962 8672 14026 8676
rect 14042 8732 14106 8736
rect 14042 8676 14046 8732
rect 14046 8676 14102 8732
rect 14102 8676 14106 8732
rect 14042 8672 14106 8676
rect 14122 8732 14186 8736
rect 14122 8676 14126 8732
rect 14126 8676 14182 8732
rect 14182 8676 14186 8732
rect 14122 8672 14186 8676
rect 14202 8732 14266 8736
rect 14202 8676 14206 8732
rect 14206 8676 14262 8732
rect 14262 8676 14266 8732
rect 14202 8672 14266 8676
rect 17062 8732 17126 8736
rect 17062 8676 17066 8732
rect 17066 8676 17122 8732
rect 17122 8676 17126 8732
rect 17062 8672 17126 8676
rect 17142 8732 17206 8736
rect 17142 8676 17146 8732
rect 17146 8676 17202 8732
rect 17202 8676 17206 8732
rect 17142 8672 17206 8676
rect 17222 8732 17286 8736
rect 17222 8676 17226 8732
rect 17226 8676 17282 8732
rect 17282 8676 17286 8732
rect 17222 8672 17286 8676
rect 17302 8732 17366 8736
rect 17302 8676 17306 8732
rect 17306 8676 17362 8732
rect 17362 8676 17366 8732
rect 17302 8672 17366 8676
rect 3112 8188 3176 8192
rect 3112 8132 3116 8188
rect 3116 8132 3172 8188
rect 3172 8132 3176 8188
rect 3112 8128 3176 8132
rect 3192 8188 3256 8192
rect 3192 8132 3196 8188
rect 3196 8132 3252 8188
rect 3252 8132 3256 8188
rect 3192 8128 3256 8132
rect 3272 8188 3336 8192
rect 3272 8132 3276 8188
rect 3276 8132 3332 8188
rect 3332 8132 3336 8188
rect 3272 8128 3336 8132
rect 3352 8188 3416 8192
rect 3352 8132 3356 8188
rect 3356 8132 3412 8188
rect 3412 8132 3416 8188
rect 3352 8128 3416 8132
rect 6212 8188 6276 8192
rect 6212 8132 6216 8188
rect 6216 8132 6272 8188
rect 6272 8132 6276 8188
rect 6212 8128 6276 8132
rect 6292 8188 6356 8192
rect 6292 8132 6296 8188
rect 6296 8132 6352 8188
rect 6352 8132 6356 8188
rect 6292 8128 6356 8132
rect 6372 8188 6436 8192
rect 6372 8132 6376 8188
rect 6376 8132 6432 8188
rect 6432 8132 6436 8188
rect 6372 8128 6436 8132
rect 6452 8188 6516 8192
rect 6452 8132 6456 8188
rect 6456 8132 6512 8188
rect 6512 8132 6516 8188
rect 6452 8128 6516 8132
rect 9312 8188 9376 8192
rect 9312 8132 9316 8188
rect 9316 8132 9372 8188
rect 9372 8132 9376 8188
rect 9312 8128 9376 8132
rect 9392 8188 9456 8192
rect 9392 8132 9396 8188
rect 9396 8132 9452 8188
rect 9452 8132 9456 8188
rect 9392 8128 9456 8132
rect 9472 8188 9536 8192
rect 9472 8132 9476 8188
rect 9476 8132 9532 8188
rect 9532 8132 9536 8188
rect 9472 8128 9536 8132
rect 9552 8188 9616 8192
rect 9552 8132 9556 8188
rect 9556 8132 9612 8188
rect 9612 8132 9616 8188
rect 9552 8128 9616 8132
rect 12412 8188 12476 8192
rect 12412 8132 12416 8188
rect 12416 8132 12472 8188
rect 12472 8132 12476 8188
rect 12412 8128 12476 8132
rect 12492 8188 12556 8192
rect 12492 8132 12496 8188
rect 12496 8132 12552 8188
rect 12552 8132 12556 8188
rect 12492 8128 12556 8132
rect 12572 8188 12636 8192
rect 12572 8132 12576 8188
rect 12576 8132 12632 8188
rect 12632 8132 12636 8188
rect 12572 8128 12636 8132
rect 12652 8188 12716 8192
rect 12652 8132 12656 8188
rect 12656 8132 12712 8188
rect 12712 8132 12716 8188
rect 12652 8128 12716 8132
rect 15512 8188 15576 8192
rect 15512 8132 15516 8188
rect 15516 8132 15572 8188
rect 15572 8132 15576 8188
rect 15512 8128 15576 8132
rect 15592 8188 15656 8192
rect 15592 8132 15596 8188
rect 15596 8132 15652 8188
rect 15652 8132 15656 8188
rect 15592 8128 15656 8132
rect 15672 8188 15736 8192
rect 15672 8132 15676 8188
rect 15676 8132 15732 8188
rect 15732 8132 15736 8188
rect 15672 8128 15736 8132
rect 15752 8188 15816 8192
rect 15752 8132 15756 8188
rect 15756 8132 15812 8188
rect 15812 8132 15816 8188
rect 15752 8128 15816 8132
rect 4662 7644 4726 7648
rect 4662 7588 4666 7644
rect 4666 7588 4722 7644
rect 4722 7588 4726 7644
rect 4662 7584 4726 7588
rect 4742 7644 4806 7648
rect 4742 7588 4746 7644
rect 4746 7588 4802 7644
rect 4802 7588 4806 7644
rect 4742 7584 4806 7588
rect 4822 7644 4886 7648
rect 4822 7588 4826 7644
rect 4826 7588 4882 7644
rect 4882 7588 4886 7644
rect 4822 7584 4886 7588
rect 4902 7644 4966 7648
rect 4902 7588 4906 7644
rect 4906 7588 4962 7644
rect 4962 7588 4966 7644
rect 4902 7584 4966 7588
rect 7762 7644 7826 7648
rect 7762 7588 7766 7644
rect 7766 7588 7822 7644
rect 7822 7588 7826 7644
rect 7762 7584 7826 7588
rect 7842 7644 7906 7648
rect 7842 7588 7846 7644
rect 7846 7588 7902 7644
rect 7902 7588 7906 7644
rect 7842 7584 7906 7588
rect 7922 7644 7986 7648
rect 7922 7588 7926 7644
rect 7926 7588 7982 7644
rect 7982 7588 7986 7644
rect 7922 7584 7986 7588
rect 8002 7644 8066 7648
rect 8002 7588 8006 7644
rect 8006 7588 8062 7644
rect 8062 7588 8066 7644
rect 8002 7584 8066 7588
rect 10862 7644 10926 7648
rect 10862 7588 10866 7644
rect 10866 7588 10922 7644
rect 10922 7588 10926 7644
rect 10862 7584 10926 7588
rect 10942 7644 11006 7648
rect 10942 7588 10946 7644
rect 10946 7588 11002 7644
rect 11002 7588 11006 7644
rect 10942 7584 11006 7588
rect 11022 7644 11086 7648
rect 11022 7588 11026 7644
rect 11026 7588 11082 7644
rect 11082 7588 11086 7644
rect 11022 7584 11086 7588
rect 11102 7644 11166 7648
rect 11102 7588 11106 7644
rect 11106 7588 11162 7644
rect 11162 7588 11166 7644
rect 11102 7584 11166 7588
rect 13962 7644 14026 7648
rect 13962 7588 13966 7644
rect 13966 7588 14022 7644
rect 14022 7588 14026 7644
rect 13962 7584 14026 7588
rect 14042 7644 14106 7648
rect 14042 7588 14046 7644
rect 14046 7588 14102 7644
rect 14102 7588 14106 7644
rect 14042 7584 14106 7588
rect 14122 7644 14186 7648
rect 14122 7588 14126 7644
rect 14126 7588 14182 7644
rect 14182 7588 14186 7644
rect 14122 7584 14186 7588
rect 14202 7644 14266 7648
rect 14202 7588 14206 7644
rect 14206 7588 14262 7644
rect 14262 7588 14266 7644
rect 14202 7584 14266 7588
rect 17062 7644 17126 7648
rect 17062 7588 17066 7644
rect 17066 7588 17122 7644
rect 17122 7588 17126 7644
rect 17062 7584 17126 7588
rect 17142 7644 17206 7648
rect 17142 7588 17146 7644
rect 17146 7588 17202 7644
rect 17202 7588 17206 7644
rect 17142 7584 17206 7588
rect 17222 7644 17286 7648
rect 17222 7588 17226 7644
rect 17226 7588 17282 7644
rect 17282 7588 17286 7644
rect 17222 7584 17286 7588
rect 17302 7644 17366 7648
rect 17302 7588 17306 7644
rect 17306 7588 17362 7644
rect 17362 7588 17366 7644
rect 17302 7584 17366 7588
rect 3112 7100 3176 7104
rect 3112 7044 3116 7100
rect 3116 7044 3172 7100
rect 3172 7044 3176 7100
rect 3112 7040 3176 7044
rect 3192 7100 3256 7104
rect 3192 7044 3196 7100
rect 3196 7044 3252 7100
rect 3252 7044 3256 7100
rect 3192 7040 3256 7044
rect 3272 7100 3336 7104
rect 3272 7044 3276 7100
rect 3276 7044 3332 7100
rect 3332 7044 3336 7100
rect 3272 7040 3336 7044
rect 3352 7100 3416 7104
rect 3352 7044 3356 7100
rect 3356 7044 3412 7100
rect 3412 7044 3416 7100
rect 3352 7040 3416 7044
rect 6212 7100 6276 7104
rect 6212 7044 6216 7100
rect 6216 7044 6272 7100
rect 6272 7044 6276 7100
rect 6212 7040 6276 7044
rect 6292 7100 6356 7104
rect 6292 7044 6296 7100
rect 6296 7044 6352 7100
rect 6352 7044 6356 7100
rect 6292 7040 6356 7044
rect 6372 7100 6436 7104
rect 6372 7044 6376 7100
rect 6376 7044 6432 7100
rect 6432 7044 6436 7100
rect 6372 7040 6436 7044
rect 6452 7100 6516 7104
rect 6452 7044 6456 7100
rect 6456 7044 6512 7100
rect 6512 7044 6516 7100
rect 6452 7040 6516 7044
rect 9312 7100 9376 7104
rect 9312 7044 9316 7100
rect 9316 7044 9372 7100
rect 9372 7044 9376 7100
rect 9312 7040 9376 7044
rect 9392 7100 9456 7104
rect 9392 7044 9396 7100
rect 9396 7044 9452 7100
rect 9452 7044 9456 7100
rect 9392 7040 9456 7044
rect 9472 7100 9536 7104
rect 9472 7044 9476 7100
rect 9476 7044 9532 7100
rect 9532 7044 9536 7100
rect 9472 7040 9536 7044
rect 9552 7100 9616 7104
rect 9552 7044 9556 7100
rect 9556 7044 9612 7100
rect 9612 7044 9616 7100
rect 9552 7040 9616 7044
rect 12412 7100 12476 7104
rect 12412 7044 12416 7100
rect 12416 7044 12472 7100
rect 12472 7044 12476 7100
rect 12412 7040 12476 7044
rect 12492 7100 12556 7104
rect 12492 7044 12496 7100
rect 12496 7044 12552 7100
rect 12552 7044 12556 7100
rect 12492 7040 12556 7044
rect 12572 7100 12636 7104
rect 12572 7044 12576 7100
rect 12576 7044 12632 7100
rect 12632 7044 12636 7100
rect 12572 7040 12636 7044
rect 12652 7100 12716 7104
rect 12652 7044 12656 7100
rect 12656 7044 12712 7100
rect 12712 7044 12716 7100
rect 12652 7040 12716 7044
rect 15512 7100 15576 7104
rect 15512 7044 15516 7100
rect 15516 7044 15572 7100
rect 15572 7044 15576 7100
rect 15512 7040 15576 7044
rect 15592 7100 15656 7104
rect 15592 7044 15596 7100
rect 15596 7044 15652 7100
rect 15652 7044 15656 7100
rect 15592 7040 15656 7044
rect 15672 7100 15736 7104
rect 15672 7044 15676 7100
rect 15676 7044 15732 7100
rect 15732 7044 15736 7100
rect 15672 7040 15736 7044
rect 15752 7100 15816 7104
rect 15752 7044 15756 7100
rect 15756 7044 15812 7100
rect 15812 7044 15816 7100
rect 15752 7040 15816 7044
rect 4662 6556 4726 6560
rect 4662 6500 4666 6556
rect 4666 6500 4722 6556
rect 4722 6500 4726 6556
rect 4662 6496 4726 6500
rect 4742 6556 4806 6560
rect 4742 6500 4746 6556
rect 4746 6500 4802 6556
rect 4802 6500 4806 6556
rect 4742 6496 4806 6500
rect 4822 6556 4886 6560
rect 4822 6500 4826 6556
rect 4826 6500 4882 6556
rect 4882 6500 4886 6556
rect 4822 6496 4886 6500
rect 4902 6556 4966 6560
rect 4902 6500 4906 6556
rect 4906 6500 4962 6556
rect 4962 6500 4966 6556
rect 4902 6496 4966 6500
rect 7762 6556 7826 6560
rect 7762 6500 7766 6556
rect 7766 6500 7822 6556
rect 7822 6500 7826 6556
rect 7762 6496 7826 6500
rect 7842 6556 7906 6560
rect 7842 6500 7846 6556
rect 7846 6500 7902 6556
rect 7902 6500 7906 6556
rect 7842 6496 7906 6500
rect 7922 6556 7986 6560
rect 7922 6500 7926 6556
rect 7926 6500 7982 6556
rect 7982 6500 7986 6556
rect 7922 6496 7986 6500
rect 8002 6556 8066 6560
rect 8002 6500 8006 6556
rect 8006 6500 8062 6556
rect 8062 6500 8066 6556
rect 8002 6496 8066 6500
rect 10862 6556 10926 6560
rect 10862 6500 10866 6556
rect 10866 6500 10922 6556
rect 10922 6500 10926 6556
rect 10862 6496 10926 6500
rect 10942 6556 11006 6560
rect 10942 6500 10946 6556
rect 10946 6500 11002 6556
rect 11002 6500 11006 6556
rect 10942 6496 11006 6500
rect 11022 6556 11086 6560
rect 11022 6500 11026 6556
rect 11026 6500 11082 6556
rect 11082 6500 11086 6556
rect 11022 6496 11086 6500
rect 11102 6556 11166 6560
rect 11102 6500 11106 6556
rect 11106 6500 11162 6556
rect 11162 6500 11166 6556
rect 11102 6496 11166 6500
rect 13962 6556 14026 6560
rect 13962 6500 13966 6556
rect 13966 6500 14022 6556
rect 14022 6500 14026 6556
rect 13962 6496 14026 6500
rect 14042 6556 14106 6560
rect 14042 6500 14046 6556
rect 14046 6500 14102 6556
rect 14102 6500 14106 6556
rect 14042 6496 14106 6500
rect 14122 6556 14186 6560
rect 14122 6500 14126 6556
rect 14126 6500 14182 6556
rect 14182 6500 14186 6556
rect 14122 6496 14186 6500
rect 14202 6556 14266 6560
rect 14202 6500 14206 6556
rect 14206 6500 14262 6556
rect 14262 6500 14266 6556
rect 14202 6496 14266 6500
rect 17062 6556 17126 6560
rect 17062 6500 17066 6556
rect 17066 6500 17122 6556
rect 17122 6500 17126 6556
rect 17062 6496 17126 6500
rect 17142 6556 17206 6560
rect 17142 6500 17146 6556
rect 17146 6500 17202 6556
rect 17202 6500 17206 6556
rect 17142 6496 17206 6500
rect 17222 6556 17286 6560
rect 17222 6500 17226 6556
rect 17226 6500 17282 6556
rect 17282 6500 17286 6556
rect 17222 6496 17286 6500
rect 17302 6556 17366 6560
rect 17302 6500 17306 6556
rect 17306 6500 17362 6556
rect 17362 6500 17366 6556
rect 17302 6496 17366 6500
rect 3112 6012 3176 6016
rect 3112 5956 3116 6012
rect 3116 5956 3172 6012
rect 3172 5956 3176 6012
rect 3112 5952 3176 5956
rect 3192 6012 3256 6016
rect 3192 5956 3196 6012
rect 3196 5956 3252 6012
rect 3252 5956 3256 6012
rect 3192 5952 3256 5956
rect 3272 6012 3336 6016
rect 3272 5956 3276 6012
rect 3276 5956 3332 6012
rect 3332 5956 3336 6012
rect 3272 5952 3336 5956
rect 3352 6012 3416 6016
rect 3352 5956 3356 6012
rect 3356 5956 3412 6012
rect 3412 5956 3416 6012
rect 3352 5952 3416 5956
rect 6212 6012 6276 6016
rect 6212 5956 6216 6012
rect 6216 5956 6272 6012
rect 6272 5956 6276 6012
rect 6212 5952 6276 5956
rect 6292 6012 6356 6016
rect 6292 5956 6296 6012
rect 6296 5956 6352 6012
rect 6352 5956 6356 6012
rect 6292 5952 6356 5956
rect 6372 6012 6436 6016
rect 6372 5956 6376 6012
rect 6376 5956 6432 6012
rect 6432 5956 6436 6012
rect 6372 5952 6436 5956
rect 6452 6012 6516 6016
rect 6452 5956 6456 6012
rect 6456 5956 6512 6012
rect 6512 5956 6516 6012
rect 6452 5952 6516 5956
rect 9312 6012 9376 6016
rect 9312 5956 9316 6012
rect 9316 5956 9372 6012
rect 9372 5956 9376 6012
rect 9312 5952 9376 5956
rect 9392 6012 9456 6016
rect 9392 5956 9396 6012
rect 9396 5956 9452 6012
rect 9452 5956 9456 6012
rect 9392 5952 9456 5956
rect 9472 6012 9536 6016
rect 9472 5956 9476 6012
rect 9476 5956 9532 6012
rect 9532 5956 9536 6012
rect 9472 5952 9536 5956
rect 9552 6012 9616 6016
rect 9552 5956 9556 6012
rect 9556 5956 9612 6012
rect 9612 5956 9616 6012
rect 9552 5952 9616 5956
rect 12412 6012 12476 6016
rect 12412 5956 12416 6012
rect 12416 5956 12472 6012
rect 12472 5956 12476 6012
rect 12412 5952 12476 5956
rect 12492 6012 12556 6016
rect 12492 5956 12496 6012
rect 12496 5956 12552 6012
rect 12552 5956 12556 6012
rect 12492 5952 12556 5956
rect 12572 6012 12636 6016
rect 12572 5956 12576 6012
rect 12576 5956 12632 6012
rect 12632 5956 12636 6012
rect 12572 5952 12636 5956
rect 12652 6012 12716 6016
rect 12652 5956 12656 6012
rect 12656 5956 12712 6012
rect 12712 5956 12716 6012
rect 12652 5952 12716 5956
rect 15512 6012 15576 6016
rect 15512 5956 15516 6012
rect 15516 5956 15572 6012
rect 15572 5956 15576 6012
rect 15512 5952 15576 5956
rect 15592 6012 15656 6016
rect 15592 5956 15596 6012
rect 15596 5956 15652 6012
rect 15652 5956 15656 6012
rect 15592 5952 15656 5956
rect 15672 6012 15736 6016
rect 15672 5956 15676 6012
rect 15676 5956 15732 6012
rect 15732 5956 15736 6012
rect 15672 5952 15736 5956
rect 15752 6012 15816 6016
rect 15752 5956 15756 6012
rect 15756 5956 15812 6012
rect 15812 5956 15816 6012
rect 15752 5952 15816 5956
rect 4662 5468 4726 5472
rect 4662 5412 4666 5468
rect 4666 5412 4722 5468
rect 4722 5412 4726 5468
rect 4662 5408 4726 5412
rect 4742 5468 4806 5472
rect 4742 5412 4746 5468
rect 4746 5412 4802 5468
rect 4802 5412 4806 5468
rect 4742 5408 4806 5412
rect 4822 5468 4886 5472
rect 4822 5412 4826 5468
rect 4826 5412 4882 5468
rect 4882 5412 4886 5468
rect 4822 5408 4886 5412
rect 4902 5468 4966 5472
rect 4902 5412 4906 5468
rect 4906 5412 4962 5468
rect 4962 5412 4966 5468
rect 4902 5408 4966 5412
rect 7762 5468 7826 5472
rect 7762 5412 7766 5468
rect 7766 5412 7822 5468
rect 7822 5412 7826 5468
rect 7762 5408 7826 5412
rect 7842 5468 7906 5472
rect 7842 5412 7846 5468
rect 7846 5412 7902 5468
rect 7902 5412 7906 5468
rect 7842 5408 7906 5412
rect 7922 5468 7986 5472
rect 7922 5412 7926 5468
rect 7926 5412 7982 5468
rect 7982 5412 7986 5468
rect 7922 5408 7986 5412
rect 8002 5468 8066 5472
rect 8002 5412 8006 5468
rect 8006 5412 8062 5468
rect 8062 5412 8066 5468
rect 8002 5408 8066 5412
rect 10862 5468 10926 5472
rect 10862 5412 10866 5468
rect 10866 5412 10922 5468
rect 10922 5412 10926 5468
rect 10862 5408 10926 5412
rect 10942 5468 11006 5472
rect 10942 5412 10946 5468
rect 10946 5412 11002 5468
rect 11002 5412 11006 5468
rect 10942 5408 11006 5412
rect 11022 5468 11086 5472
rect 11022 5412 11026 5468
rect 11026 5412 11082 5468
rect 11082 5412 11086 5468
rect 11022 5408 11086 5412
rect 11102 5468 11166 5472
rect 11102 5412 11106 5468
rect 11106 5412 11162 5468
rect 11162 5412 11166 5468
rect 11102 5408 11166 5412
rect 13962 5468 14026 5472
rect 13962 5412 13966 5468
rect 13966 5412 14022 5468
rect 14022 5412 14026 5468
rect 13962 5408 14026 5412
rect 14042 5468 14106 5472
rect 14042 5412 14046 5468
rect 14046 5412 14102 5468
rect 14102 5412 14106 5468
rect 14042 5408 14106 5412
rect 14122 5468 14186 5472
rect 14122 5412 14126 5468
rect 14126 5412 14182 5468
rect 14182 5412 14186 5468
rect 14122 5408 14186 5412
rect 14202 5468 14266 5472
rect 14202 5412 14206 5468
rect 14206 5412 14262 5468
rect 14262 5412 14266 5468
rect 14202 5408 14266 5412
rect 17062 5468 17126 5472
rect 17062 5412 17066 5468
rect 17066 5412 17122 5468
rect 17122 5412 17126 5468
rect 17062 5408 17126 5412
rect 17142 5468 17206 5472
rect 17142 5412 17146 5468
rect 17146 5412 17202 5468
rect 17202 5412 17206 5468
rect 17142 5408 17206 5412
rect 17222 5468 17286 5472
rect 17222 5412 17226 5468
rect 17226 5412 17282 5468
rect 17282 5412 17286 5468
rect 17222 5408 17286 5412
rect 17302 5468 17366 5472
rect 17302 5412 17306 5468
rect 17306 5412 17362 5468
rect 17362 5412 17366 5468
rect 17302 5408 17366 5412
rect 3112 4924 3176 4928
rect 3112 4868 3116 4924
rect 3116 4868 3172 4924
rect 3172 4868 3176 4924
rect 3112 4864 3176 4868
rect 3192 4924 3256 4928
rect 3192 4868 3196 4924
rect 3196 4868 3252 4924
rect 3252 4868 3256 4924
rect 3192 4864 3256 4868
rect 3272 4924 3336 4928
rect 3272 4868 3276 4924
rect 3276 4868 3332 4924
rect 3332 4868 3336 4924
rect 3272 4864 3336 4868
rect 3352 4924 3416 4928
rect 3352 4868 3356 4924
rect 3356 4868 3412 4924
rect 3412 4868 3416 4924
rect 3352 4864 3416 4868
rect 6212 4924 6276 4928
rect 6212 4868 6216 4924
rect 6216 4868 6272 4924
rect 6272 4868 6276 4924
rect 6212 4864 6276 4868
rect 6292 4924 6356 4928
rect 6292 4868 6296 4924
rect 6296 4868 6352 4924
rect 6352 4868 6356 4924
rect 6292 4864 6356 4868
rect 6372 4924 6436 4928
rect 6372 4868 6376 4924
rect 6376 4868 6432 4924
rect 6432 4868 6436 4924
rect 6372 4864 6436 4868
rect 6452 4924 6516 4928
rect 6452 4868 6456 4924
rect 6456 4868 6512 4924
rect 6512 4868 6516 4924
rect 6452 4864 6516 4868
rect 9312 4924 9376 4928
rect 9312 4868 9316 4924
rect 9316 4868 9372 4924
rect 9372 4868 9376 4924
rect 9312 4864 9376 4868
rect 9392 4924 9456 4928
rect 9392 4868 9396 4924
rect 9396 4868 9452 4924
rect 9452 4868 9456 4924
rect 9392 4864 9456 4868
rect 9472 4924 9536 4928
rect 9472 4868 9476 4924
rect 9476 4868 9532 4924
rect 9532 4868 9536 4924
rect 9472 4864 9536 4868
rect 9552 4924 9616 4928
rect 9552 4868 9556 4924
rect 9556 4868 9612 4924
rect 9612 4868 9616 4924
rect 9552 4864 9616 4868
rect 12412 4924 12476 4928
rect 12412 4868 12416 4924
rect 12416 4868 12472 4924
rect 12472 4868 12476 4924
rect 12412 4864 12476 4868
rect 12492 4924 12556 4928
rect 12492 4868 12496 4924
rect 12496 4868 12552 4924
rect 12552 4868 12556 4924
rect 12492 4864 12556 4868
rect 12572 4924 12636 4928
rect 12572 4868 12576 4924
rect 12576 4868 12632 4924
rect 12632 4868 12636 4924
rect 12572 4864 12636 4868
rect 12652 4924 12716 4928
rect 12652 4868 12656 4924
rect 12656 4868 12712 4924
rect 12712 4868 12716 4924
rect 12652 4864 12716 4868
rect 15512 4924 15576 4928
rect 15512 4868 15516 4924
rect 15516 4868 15572 4924
rect 15572 4868 15576 4924
rect 15512 4864 15576 4868
rect 15592 4924 15656 4928
rect 15592 4868 15596 4924
rect 15596 4868 15652 4924
rect 15652 4868 15656 4924
rect 15592 4864 15656 4868
rect 15672 4924 15736 4928
rect 15672 4868 15676 4924
rect 15676 4868 15732 4924
rect 15732 4868 15736 4924
rect 15672 4864 15736 4868
rect 15752 4924 15816 4928
rect 15752 4868 15756 4924
rect 15756 4868 15812 4924
rect 15812 4868 15816 4924
rect 15752 4864 15816 4868
rect 4662 4380 4726 4384
rect 4662 4324 4666 4380
rect 4666 4324 4722 4380
rect 4722 4324 4726 4380
rect 4662 4320 4726 4324
rect 4742 4380 4806 4384
rect 4742 4324 4746 4380
rect 4746 4324 4802 4380
rect 4802 4324 4806 4380
rect 4742 4320 4806 4324
rect 4822 4380 4886 4384
rect 4822 4324 4826 4380
rect 4826 4324 4882 4380
rect 4882 4324 4886 4380
rect 4822 4320 4886 4324
rect 4902 4380 4966 4384
rect 4902 4324 4906 4380
rect 4906 4324 4962 4380
rect 4962 4324 4966 4380
rect 4902 4320 4966 4324
rect 7762 4380 7826 4384
rect 7762 4324 7766 4380
rect 7766 4324 7822 4380
rect 7822 4324 7826 4380
rect 7762 4320 7826 4324
rect 7842 4380 7906 4384
rect 7842 4324 7846 4380
rect 7846 4324 7902 4380
rect 7902 4324 7906 4380
rect 7842 4320 7906 4324
rect 7922 4380 7986 4384
rect 7922 4324 7926 4380
rect 7926 4324 7982 4380
rect 7982 4324 7986 4380
rect 7922 4320 7986 4324
rect 8002 4380 8066 4384
rect 8002 4324 8006 4380
rect 8006 4324 8062 4380
rect 8062 4324 8066 4380
rect 8002 4320 8066 4324
rect 10862 4380 10926 4384
rect 10862 4324 10866 4380
rect 10866 4324 10922 4380
rect 10922 4324 10926 4380
rect 10862 4320 10926 4324
rect 10942 4380 11006 4384
rect 10942 4324 10946 4380
rect 10946 4324 11002 4380
rect 11002 4324 11006 4380
rect 10942 4320 11006 4324
rect 11022 4380 11086 4384
rect 11022 4324 11026 4380
rect 11026 4324 11082 4380
rect 11082 4324 11086 4380
rect 11022 4320 11086 4324
rect 11102 4380 11166 4384
rect 11102 4324 11106 4380
rect 11106 4324 11162 4380
rect 11162 4324 11166 4380
rect 11102 4320 11166 4324
rect 13962 4380 14026 4384
rect 13962 4324 13966 4380
rect 13966 4324 14022 4380
rect 14022 4324 14026 4380
rect 13962 4320 14026 4324
rect 14042 4380 14106 4384
rect 14042 4324 14046 4380
rect 14046 4324 14102 4380
rect 14102 4324 14106 4380
rect 14042 4320 14106 4324
rect 14122 4380 14186 4384
rect 14122 4324 14126 4380
rect 14126 4324 14182 4380
rect 14182 4324 14186 4380
rect 14122 4320 14186 4324
rect 14202 4380 14266 4384
rect 14202 4324 14206 4380
rect 14206 4324 14262 4380
rect 14262 4324 14266 4380
rect 14202 4320 14266 4324
rect 17062 4380 17126 4384
rect 17062 4324 17066 4380
rect 17066 4324 17122 4380
rect 17122 4324 17126 4380
rect 17062 4320 17126 4324
rect 17142 4380 17206 4384
rect 17142 4324 17146 4380
rect 17146 4324 17202 4380
rect 17202 4324 17206 4380
rect 17142 4320 17206 4324
rect 17222 4380 17286 4384
rect 17222 4324 17226 4380
rect 17226 4324 17282 4380
rect 17282 4324 17286 4380
rect 17222 4320 17286 4324
rect 17302 4380 17366 4384
rect 17302 4324 17306 4380
rect 17306 4324 17362 4380
rect 17362 4324 17366 4380
rect 17302 4320 17366 4324
rect 3112 3836 3176 3840
rect 3112 3780 3116 3836
rect 3116 3780 3172 3836
rect 3172 3780 3176 3836
rect 3112 3776 3176 3780
rect 3192 3836 3256 3840
rect 3192 3780 3196 3836
rect 3196 3780 3252 3836
rect 3252 3780 3256 3836
rect 3192 3776 3256 3780
rect 3272 3836 3336 3840
rect 3272 3780 3276 3836
rect 3276 3780 3332 3836
rect 3332 3780 3336 3836
rect 3272 3776 3336 3780
rect 3352 3836 3416 3840
rect 3352 3780 3356 3836
rect 3356 3780 3412 3836
rect 3412 3780 3416 3836
rect 3352 3776 3416 3780
rect 6212 3836 6276 3840
rect 6212 3780 6216 3836
rect 6216 3780 6272 3836
rect 6272 3780 6276 3836
rect 6212 3776 6276 3780
rect 6292 3836 6356 3840
rect 6292 3780 6296 3836
rect 6296 3780 6352 3836
rect 6352 3780 6356 3836
rect 6292 3776 6356 3780
rect 6372 3836 6436 3840
rect 6372 3780 6376 3836
rect 6376 3780 6432 3836
rect 6432 3780 6436 3836
rect 6372 3776 6436 3780
rect 6452 3836 6516 3840
rect 6452 3780 6456 3836
rect 6456 3780 6512 3836
rect 6512 3780 6516 3836
rect 6452 3776 6516 3780
rect 9312 3836 9376 3840
rect 9312 3780 9316 3836
rect 9316 3780 9372 3836
rect 9372 3780 9376 3836
rect 9312 3776 9376 3780
rect 9392 3836 9456 3840
rect 9392 3780 9396 3836
rect 9396 3780 9452 3836
rect 9452 3780 9456 3836
rect 9392 3776 9456 3780
rect 9472 3836 9536 3840
rect 9472 3780 9476 3836
rect 9476 3780 9532 3836
rect 9532 3780 9536 3836
rect 9472 3776 9536 3780
rect 9552 3836 9616 3840
rect 9552 3780 9556 3836
rect 9556 3780 9612 3836
rect 9612 3780 9616 3836
rect 9552 3776 9616 3780
rect 12412 3836 12476 3840
rect 12412 3780 12416 3836
rect 12416 3780 12472 3836
rect 12472 3780 12476 3836
rect 12412 3776 12476 3780
rect 12492 3836 12556 3840
rect 12492 3780 12496 3836
rect 12496 3780 12552 3836
rect 12552 3780 12556 3836
rect 12492 3776 12556 3780
rect 12572 3836 12636 3840
rect 12572 3780 12576 3836
rect 12576 3780 12632 3836
rect 12632 3780 12636 3836
rect 12572 3776 12636 3780
rect 12652 3836 12716 3840
rect 12652 3780 12656 3836
rect 12656 3780 12712 3836
rect 12712 3780 12716 3836
rect 12652 3776 12716 3780
rect 15512 3836 15576 3840
rect 15512 3780 15516 3836
rect 15516 3780 15572 3836
rect 15572 3780 15576 3836
rect 15512 3776 15576 3780
rect 15592 3836 15656 3840
rect 15592 3780 15596 3836
rect 15596 3780 15652 3836
rect 15652 3780 15656 3836
rect 15592 3776 15656 3780
rect 15672 3836 15736 3840
rect 15672 3780 15676 3836
rect 15676 3780 15732 3836
rect 15732 3780 15736 3836
rect 15672 3776 15736 3780
rect 15752 3836 15816 3840
rect 15752 3780 15756 3836
rect 15756 3780 15812 3836
rect 15812 3780 15816 3836
rect 15752 3776 15816 3780
rect 4662 3292 4726 3296
rect 4662 3236 4666 3292
rect 4666 3236 4722 3292
rect 4722 3236 4726 3292
rect 4662 3232 4726 3236
rect 4742 3292 4806 3296
rect 4742 3236 4746 3292
rect 4746 3236 4802 3292
rect 4802 3236 4806 3292
rect 4742 3232 4806 3236
rect 4822 3292 4886 3296
rect 4822 3236 4826 3292
rect 4826 3236 4882 3292
rect 4882 3236 4886 3292
rect 4822 3232 4886 3236
rect 4902 3292 4966 3296
rect 4902 3236 4906 3292
rect 4906 3236 4962 3292
rect 4962 3236 4966 3292
rect 4902 3232 4966 3236
rect 7762 3292 7826 3296
rect 7762 3236 7766 3292
rect 7766 3236 7822 3292
rect 7822 3236 7826 3292
rect 7762 3232 7826 3236
rect 7842 3292 7906 3296
rect 7842 3236 7846 3292
rect 7846 3236 7902 3292
rect 7902 3236 7906 3292
rect 7842 3232 7906 3236
rect 7922 3292 7986 3296
rect 7922 3236 7926 3292
rect 7926 3236 7982 3292
rect 7982 3236 7986 3292
rect 7922 3232 7986 3236
rect 8002 3292 8066 3296
rect 8002 3236 8006 3292
rect 8006 3236 8062 3292
rect 8062 3236 8066 3292
rect 8002 3232 8066 3236
rect 10862 3292 10926 3296
rect 10862 3236 10866 3292
rect 10866 3236 10922 3292
rect 10922 3236 10926 3292
rect 10862 3232 10926 3236
rect 10942 3292 11006 3296
rect 10942 3236 10946 3292
rect 10946 3236 11002 3292
rect 11002 3236 11006 3292
rect 10942 3232 11006 3236
rect 11022 3292 11086 3296
rect 11022 3236 11026 3292
rect 11026 3236 11082 3292
rect 11082 3236 11086 3292
rect 11022 3232 11086 3236
rect 11102 3292 11166 3296
rect 11102 3236 11106 3292
rect 11106 3236 11162 3292
rect 11162 3236 11166 3292
rect 11102 3232 11166 3236
rect 13962 3292 14026 3296
rect 13962 3236 13966 3292
rect 13966 3236 14022 3292
rect 14022 3236 14026 3292
rect 13962 3232 14026 3236
rect 14042 3292 14106 3296
rect 14042 3236 14046 3292
rect 14046 3236 14102 3292
rect 14102 3236 14106 3292
rect 14042 3232 14106 3236
rect 14122 3292 14186 3296
rect 14122 3236 14126 3292
rect 14126 3236 14182 3292
rect 14182 3236 14186 3292
rect 14122 3232 14186 3236
rect 14202 3292 14266 3296
rect 14202 3236 14206 3292
rect 14206 3236 14262 3292
rect 14262 3236 14266 3292
rect 14202 3232 14266 3236
rect 17062 3292 17126 3296
rect 17062 3236 17066 3292
rect 17066 3236 17122 3292
rect 17122 3236 17126 3292
rect 17062 3232 17126 3236
rect 17142 3292 17206 3296
rect 17142 3236 17146 3292
rect 17146 3236 17202 3292
rect 17202 3236 17206 3292
rect 17142 3232 17206 3236
rect 17222 3292 17286 3296
rect 17222 3236 17226 3292
rect 17226 3236 17282 3292
rect 17282 3236 17286 3292
rect 17222 3232 17286 3236
rect 17302 3292 17366 3296
rect 17302 3236 17306 3292
rect 17306 3236 17362 3292
rect 17362 3236 17366 3292
rect 17302 3232 17366 3236
rect 3112 2748 3176 2752
rect 3112 2692 3116 2748
rect 3116 2692 3172 2748
rect 3172 2692 3176 2748
rect 3112 2688 3176 2692
rect 3192 2748 3256 2752
rect 3192 2692 3196 2748
rect 3196 2692 3252 2748
rect 3252 2692 3256 2748
rect 3192 2688 3256 2692
rect 3272 2748 3336 2752
rect 3272 2692 3276 2748
rect 3276 2692 3332 2748
rect 3332 2692 3336 2748
rect 3272 2688 3336 2692
rect 3352 2748 3416 2752
rect 3352 2692 3356 2748
rect 3356 2692 3412 2748
rect 3412 2692 3416 2748
rect 3352 2688 3416 2692
rect 6212 2748 6276 2752
rect 6212 2692 6216 2748
rect 6216 2692 6272 2748
rect 6272 2692 6276 2748
rect 6212 2688 6276 2692
rect 6292 2748 6356 2752
rect 6292 2692 6296 2748
rect 6296 2692 6352 2748
rect 6352 2692 6356 2748
rect 6292 2688 6356 2692
rect 6372 2748 6436 2752
rect 6372 2692 6376 2748
rect 6376 2692 6432 2748
rect 6432 2692 6436 2748
rect 6372 2688 6436 2692
rect 6452 2748 6516 2752
rect 6452 2692 6456 2748
rect 6456 2692 6512 2748
rect 6512 2692 6516 2748
rect 6452 2688 6516 2692
rect 9312 2748 9376 2752
rect 9312 2692 9316 2748
rect 9316 2692 9372 2748
rect 9372 2692 9376 2748
rect 9312 2688 9376 2692
rect 9392 2748 9456 2752
rect 9392 2692 9396 2748
rect 9396 2692 9452 2748
rect 9452 2692 9456 2748
rect 9392 2688 9456 2692
rect 9472 2748 9536 2752
rect 9472 2692 9476 2748
rect 9476 2692 9532 2748
rect 9532 2692 9536 2748
rect 9472 2688 9536 2692
rect 9552 2748 9616 2752
rect 9552 2692 9556 2748
rect 9556 2692 9612 2748
rect 9612 2692 9616 2748
rect 9552 2688 9616 2692
rect 12412 2748 12476 2752
rect 12412 2692 12416 2748
rect 12416 2692 12472 2748
rect 12472 2692 12476 2748
rect 12412 2688 12476 2692
rect 12492 2748 12556 2752
rect 12492 2692 12496 2748
rect 12496 2692 12552 2748
rect 12552 2692 12556 2748
rect 12492 2688 12556 2692
rect 12572 2748 12636 2752
rect 12572 2692 12576 2748
rect 12576 2692 12632 2748
rect 12632 2692 12636 2748
rect 12572 2688 12636 2692
rect 12652 2748 12716 2752
rect 12652 2692 12656 2748
rect 12656 2692 12712 2748
rect 12712 2692 12716 2748
rect 12652 2688 12716 2692
rect 15512 2748 15576 2752
rect 15512 2692 15516 2748
rect 15516 2692 15572 2748
rect 15572 2692 15576 2748
rect 15512 2688 15576 2692
rect 15592 2748 15656 2752
rect 15592 2692 15596 2748
rect 15596 2692 15652 2748
rect 15652 2692 15656 2748
rect 15592 2688 15656 2692
rect 15672 2748 15736 2752
rect 15672 2692 15676 2748
rect 15676 2692 15732 2748
rect 15732 2692 15736 2748
rect 15672 2688 15736 2692
rect 15752 2748 15816 2752
rect 15752 2692 15756 2748
rect 15756 2692 15812 2748
rect 15812 2692 15816 2748
rect 15752 2688 15816 2692
rect 4662 2204 4726 2208
rect 4662 2148 4666 2204
rect 4666 2148 4722 2204
rect 4722 2148 4726 2204
rect 4662 2144 4726 2148
rect 4742 2204 4806 2208
rect 4742 2148 4746 2204
rect 4746 2148 4802 2204
rect 4802 2148 4806 2204
rect 4742 2144 4806 2148
rect 4822 2204 4886 2208
rect 4822 2148 4826 2204
rect 4826 2148 4882 2204
rect 4882 2148 4886 2204
rect 4822 2144 4886 2148
rect 4902 2204 4966 2208
rect 4902 2148 4906 2204
rect 4906 2148 4962 2204
rect 4962 2148 4966 2204
rect 4902 2144 4966 2148
rect 7762 2204 7826 2208
rect 7762 2148 7766 2204
rect 7766 2148 7822 2204
rect 7822 2148 7826 2204
rect 7762 2144 7826 2148
rect 7842 2204 7906 2208
rect 7842 2148 7846 2204
rect 7846 2148 7902 2204
rect 7902 2148 7906 2204
rect 7842 2144 7906 2148
rect 7922 2204 7986 2208
rect 7922 2148 7926 2204
rect 7926 2148 7982 2204
rect 7982 2148 7986 2204
rect 7922 2144 7986 2148
rect 8002 2204 8066 2208
rect 8002 2148 8006 2204
rect 8006 2148 8062 2204
rect 8062 2148 8066 2204
rect 8002 2144 8066 2148
rect 10862 2204 10926 2208
rect 10862 2148 10866 2204
rect 10866 2148 10922 2204
rect 10922 2148 10926 2204
rect 10862 2144 10926 2148
rect 10942 2204 11006 2208
rect 10942 2148 10946 2204
rect 10946 2148 11002 2204
rect 11002 2148 11006 2204
rect 10942 2144 11006 2148
rect 11022 2204 11086 2208
rect 11022 2148 11026 2204
rect 11026 2148 11082 2204
rect 11082 2148 11086 2204
rect 11022 2144 11086 2148
rect 11102 2204 11166 2208
rect 11102 2148 11106 2204
rect 11106 2148 11162 2204
rect 11162 2148 11166 2204
rect 11102 2144 11166 2148
rect 13962 2204 14026 2208
rect 13962 2148 13966 2204
rect 13966 2148 14022 2204
rect 14022 2148 14026 2204
rect 13962 2144 14026 2148
rect 14042 2204 14106 2208
rect 14042 2148 14046 2204
rect 14046 2148 14102 2204
rect 14102 2148 14106 2204
rect 14042 2144 14106 2148
rect 14122 2204 14186 2208
rect 14122 2148 14126 2204
rect 14126 2148 14182 2204
rect 14182 2148 14186 2204
rect 14122 2144 14186 2148
rect 14202 2204 14266 2208
rect 14202 2148 14206 2204
rect 14206 2148 14262 2204
rect 14262 2148 14266 2204
rect 14202 2144 14266 2148
rect 17062 2204 17126 2208
rect 17062 2148 17066 2204
rect 17066 2148 17122 2204
rect 17122 2148 17126 2204
rect 17062 2144 17126 2148
rect 17142 2204 17206 2208
rect 17142 2148 17146 2204
rect 17146 2148 17202 2204
rect 17202 2148 17206 2204
rect 17142 2144 17206 2148
rect 17222 2204 17286 2208
rect 17222 2148 17226 2204
rect 17226 2148 17282 2204
rect 17282 2148 17286 2204
rect 17222 2144 17286 2148
rect 17302 2204 17366 2208
rect 17302 2148 17306 2204
rect 17306 2148 17362 2204
rect 17362 2148 17366 2204
rect 17302 2144 17366 2148
rect 3112 1660 3176 1664
rect 3112 1604 3116 1660
rect 3116 1604 3172 1660
rect 3172 1604 3176 1660
rect 3112 1600 3176 1604
rect 3192 1660 3256 1664
rect 3192 1604 3196 1660
rect 3196 1604 3252 1660
rect 3252 1604 3256 1660
rect 3192 1600 3256 1604
rect 3272 1660 3336 1664
rect 3272 1604 3276 1660
rect 3276 1604 3332 1660
rect 3332 1604 3336 1660
rect 3272 1600 3336 1604
rect 3352 1660 3416 1664
rect 3352 1604 3356 1660
rect 3356 1604 3412 1660
rect 3412 1604 3416 1660
rect 3352 1600 3416 1604
rect 6212 1660 6276 1664
rect 6212 1604 6216 1660
rect 6216 1604 6272 1660
rect 6272 1604 6276 1660
rect 6212 1600 6276 1604
rect 6292 1660 6356 1664
rect 6292 1604 6296 1660
rect 6296 1604 6352 1660
rect 6352 1604 6356 1660
rect 6292 1600 6356 1604
rect 6372 1660 6436 1664
rect 6372 1604 6376 1660
rect 6376 1604 6432 1660
rect 6432 1604 6436 1660
rect 6372 1600 6436 1604
rect 6452 1660 6516 1664
rect 6452 1604 6456 1660
rect 6456 1604 6512 1660
rect 6512 1604 6516 1660
rect 6452 1600 6516 1604
rect 9312 1660 9376 1664
rect 9312 1604 9316 1660
rect 9316 1604 9372 1660
rect 9372 1604 9376 1660
rect 9312 1600 9376 1604
rect 9392 1660 9456 1664
rect 9392 1604 9396 1660
rect 9396 1604 9452 1660
rect 9452 1604 9456 1660
rect 9392 1600 9456 1604
rect 9472 1660 9536 1664
rect 9472 1604 9476 1660
rect 9476 1604 9532 1660
rect 9532 1604 9536 1660
rect 9472 1600 9536 1604
rect 9552 1660 9616 1664
rect 9552 1604 9556 1660
rect 9556 1604 9612 1660
rect 9612 1604 9616 1660
rect 9552 1600 9616 1604
rect 12412 1660 12476 1664
rect 12412 1604 12416 1660
rect 12416 1604 12472 1660
rect 12472 1604 12476 1660
rect 12412 1600 12476 1604
rect 12492 1660 12556 1664
rect 12492 1604 12496 1660
rect 12496 1604 12552 1660
rect 12552 1604 12556 1660
rect 12492 1600 12556 1604
rect 12572 1660 12636 1664
rect 12572 1604 12576 1660
rect 12576 1604 12632 1660
rect 12632 1604 12636 1660
rect 12572 1600 12636 1604
rect 12652 1660 12716 1664
rect 12652 1604 12656 1660
rect 12656 1604 12712 1660
rect 12712 1604 12716 1660
rect 12652 1600 12716 1604
rect 15512 1660 15576 1664
rect 15512 1604 15516 1660
rect 15516 1604 15572 1660
rect 15572 1604 15576 1660
rect 15512 1600 15576 1604
rect 15592 1660 15656 1664
rect 15592 1604 15596 1660
rect 15596 1604 15652 1660
rect 15652 1604 15656 1660
rect 15592 1600 15656 1604
rect 15672 1660 15736 1664
rect 15672 1604 15676 1660
rect 15676 1604 15732 1660
rect 15732 1604 15736 1660
rect 15672 1600 15736 1604
rect 15752 1660 15816 1664
rect 15752 1604 15756 1660
rect 15756 1604 15812 1660
rect 15812 1604 15816 1660
rect 15752 1600 15816 1604
rect 4662 1116 4726 1120
rect 4662 1060 4666 1116
rect 4666 1060 4722 1116
rect 4722 1060 4726 1116
rect 4662 1056 4726 1060
rect 4742 1116 4806 1120
rect 4742 1060 4746 1116
rect 4746 1060 4802 1116
rect 4802 1060 4806 1116
rect 4742 1056 4806 1060
rect 4822 1116 4886 1120
rect 4822 1060 4826 1116
rect 4826 1060 4882 1116
rect 4882 1060 4886 1116
rect 4822 1056 4886 1060
rect 4902 1116 4966 1120
rect 4902 1060 4906 1116
rect 4906 1060 4962 1116
rect 4962 1060 4966 1116
rect 4902 1056 4966 1060
rect 7762 1116 7826 1120
rect 7762 1060 7766 1116
rect 7766 1060 7822 1116
rect 7822 1060 7826 1116
rect 7762 1056 7826 1060
rect 7842 1116 7906 1120
rect 7842 1060 7846 1116
rect 7846 1060 7902 1116
rect 7902 1060 7906 1116
rect 7842 1056 7906 1060
rect 7922 1116 7986 1120
rect 7922 1060 7926 1116
rect 7926 1060 7982 1116
rect 7982 1060 7986 1116
rect 7922 1056 7986 1060
rect 8002 1116 8066 1120
rect 8002 1060 8006 1116
rect 8006 1060 8062 1116
rect 8062 1060 8066 1116
rect 8002 1056 8066 1060
rect 10862 1116 10926 1120
rect 10862 1060 10866 1116
rect 10866 1060 10922 1116
rect 10922 1060 10926 1116
rect 10862 1056 10926 1060
rect 10942 1116 11006 1120
rect 10942 1060 10946 1116
rect 10946 1060 11002 1116
rect 11002 1060 11006 1116
rect 10942 1056 11006 1060
rect 11022 1116 11086 1120
rect 11022 1060 11026 1116
rect 11026 1060 11082 1116
rect 11082 1060 11086 1116
rect 11022 1056 11086 1060
rect 11102 1116 11166 1120
rect 11102 1060 11106 1116
rect 11106 1060 11162 1116
rect 11162 1060 11166 1116
rect 11102 1056 11166 1060
rect 13962 1116 14026 1120
rect 13962 1060 13966 1116
rect 13966 1060 14022 1116
rect 14022 1060 14026 1116
rect 13962 1056 14026 1060
rect 14042 1116 14106 1120
rect 14042 1060 14046 1116
rect 14046 1060 14102 1116
rect 14102 1060 14106 1116
rect 14042 1056 14106 1060
rect 14122 1116 14186 1120
rect 14122 1060 14126 1116
rect 14126 1060 14182 1116
rect 14182 1060 14186 1116
rect 14122 1056 14186 1060
rect 14202 1116 14266 1120
rect 14202 1060 14206 1116
rect 14206 1060 14262 1116
rect 14262 1060 14266 1116
rect 14202 1056 14266 1060
rect 17062 1116 17126 1120
rect 17062 1060 17066 1116
rect 17066 1060 17122 1116
rect 17122 1060 17126 1116
rect 17062 1056 17126 1060
rect 17142 1116 17206 1120
rect 17142 1060 17146 1116
rect 17146 1060 17202 1116
rect 17202 1060 17206 1116
rect 17142 1056 17206 1060
rect 17222 1116 17286 1120
rect 17222 1060 17226 1116
rect 17226 1060 17282 1116
rect 17282 1060 17286 1116
rect 17222 1056 17286 1060
rect 17302 1116 17366 1120
rect 17302 1060 17306 1116
rect 17306 1060 17362 1116
rect 17362 1060 17366 1116
rect 17302 1056 17366 1060
rect 3112 572 3176 576
rect 3112 516 3116 572
rect 3116 516 3172 572
rect 3172 516 3176 572
rect 3112 512 3176 516
rect 3192 572 3256 576
rect 3192 516 3196 572
rect 3196 516 3252 572
rect 3252 516 3256 572
rect 3192 512 3256 516
rect 3272 572 3336 576
rect 3272 516 3276 572
rect 3276 516 3332 572
rect 3332 516 3336 572
rect 3272 512 3336 516
rect 3352 572 3416 576
rect 3352 516 3356 572
rect 3356 516 3412 572
rect 3412 516 3416 572
rect 3352 512 3416 516
rect 6212 572 6276 576
rect 6212 516 6216 572
rect 6216 516 6272 572
rect 6272 516 6276 572
rect 6212 512 6276 516
rect 6292 572 6356 576
rect 6292 516 6296 572
rect 6296 516 6352 572
rect 6352 516 6356 572
rect 6292 512 6356 516
rect 6372 572 6436 576
rect 6372 516 6376 572
rect 6376 516 6432 572
rect 6432 516 6436 572
rect 6372 512 6436 516
rect 6452 572 6516 576
rect 6452 516 6456 572
rect 6456 516 6512 572
rect 6512 516 6516 572
rect 6452 512 6516 516
rect 9312 572 9376 576
rect 9312 516 9316 572
rect 9316 516 9372 572
rect 9372 516 9376 572
rect 9312 512 9376 516
rect 9392 572 9456 576
rect 9392 516 9396 572
rect 9396 516 9452 572
rect 9452 516 9456 572
rect 9392 512 9456 516
rect 9472 572 9536 576
rect 9472 516 9476 572
rect 9476 516 9532 572
rect 9532 516 9536 572
rect 9472 512 9536 516
rect 9552 572 9616 576
rect 9552 516 9556 572
rect 9556 516 9612 572
rect 9612 516 9616 572
rect 9552 512 9616 516
rect 12412 572 12476 576
rect 12412 516 12416 572
rect 12416 516 12472 572
rect 12472 516 12476 572
rect 12412 512 12476 516
rect 12492 572 12556 576
rect 12492 516 12496 572
rect 12496 516 12552 572
rect 12552 516 12556 572
rect 12492 512 12556 516
rect 12572 572 12636 576
rect 12572 516 12576 572
rect 12576 516 12632 572
rect 12632 516 12636 572
rect 12572 512 12636 516
rect 12652 572 12716 576
rect 12652 516 12656 572
rect 12656 516 12712 572
rect 12712 516 12716 572
rect 12652 512 12716 516
rect 15512 572 15576 576
rect 15512 516 15516 572
rect 15516 516 15572 572
rect 15572 516 15576 572
rect 15512 512 15576 516
rect 15592 572 15656 576
rect 15592 516 15596 572
rect 15596 516 15652 572
rect 15652 516 15656 572
rect 15592 512 15656 516
rect 15672 572 15736 576
rect 15672 516 15676 572
rect 15676 516 15732 572
rect 15732 516 15736 572
rect 15672 512 15736 516
rect 15752 572 15816 576
rect 15752 516 15756 572
rect 15756 516 15812 572
rect 15812 516 15816 572
rect 15752 512 15816 516
rect 4662 28 4726 32
rect 4662 -28 4666 28
rect 4666 -28 4722 28
rect 4722 -28 4726 28
rect 4662 -32 4726 -28
rect 4742 28 4806 32
rect 4742 -28 4746 28
rect 4746 -28 4802 28
rect 4802 -28 4806 28
rect 4742 -32 4806 -28
rect 4822 28 4886 32
rect 4822 -28 4826 28
rect 4826 -28 4882 28
rect 4882 -28 4886 28
rect 4822 -32 4886 -28
rect 4902 28 4966 32
rect 4902 -28 4906 28
rect 4906 -28 4962 28
rect 4962 -28 4966 28
rect 4902 -32 4966 -28
rect 7762 28 7826 32
rect 7762 -28 7766 28
rect 7766 -28 7822 28
rect 7822 -28 7826 28
rect 7762 -32 7826 -28
rect 7842 28 7906 32
rect 7842 -28 7846 28
rect 7846 -28 7902 28
rect 7902 -28 7906 28
rect 7842 -32 7906 -28
rect 7922 28 7986 32
rect 7922 -28 7926 28
rect 7926 -28 7982 28
rect 7982 -28 7986 28
rect 7922 -32 7986 -28
rect 8002 28 8066 32
rect 8002 -28 8006 28
rect 8006 -28 8062 28
rect 8062 -28 8066 28
rect 8002 -32 8066 -28
rect 10862 28 10926 32
rect 10862 -28 10866 28
rect 10866 -28 10922 28
rect 10922 -28 10926 28
rect 10862 -32 10926 -28
rect 10942 28 11006 32
rect 10942 -28 10946 28
rect 10946 -28 11002 28
rect 11002 -28 11006 28
rect 10942 -32 11006 -28
rect 11022 28 11086 32
rect 11022 -28 11026 28
rect 11026 -28 11082 28
rect 11082 -28 11086 28
rect 11022 -32 11086 -28
rect 11102 28 11166 32
rect 11102 -28 11106 28
rect 11106 -28 11162 28
rect 11162 -28 11166 28
rect 11102 -32 11166 -28
rect 13962 28 14026 32
rect 13962 -28 13966 28
rect 13966 -28 14022 28
rect 14022 -28 14026 28
rect 13962 -32 14026 -28
rect 14042 28 14106 32
rect 14042 -28 14046 28
rect 14046 -28 14102 28
rect 14102 -28 14106 28
rect 14042 -32 14106 -28
rect 14122 28 14186 32
rect 14122 -28 14126 28
rect 14126 -28 14182 28
rect 14182 -28 14186 28
rect 14122 -32 14186 -28
rect 14202 28 14266 32
rect 14202 -28 14206 28
rect 14206 -28 14262 28
rect 14262 -28 14266 28
rect 14202 -32 14266 -28
rect 17062 28 17126 32
rect 17062 -28 17066 28
rect 17066 -28 17122 28
rect 17122 -28 17126 28
rect 17062 -32 17126 -28
rect 17142 28 17206 32
rect 17142 -28 17146 28
rect 17146 -28 17202 28
rect 17202 -28 17206 28
rect 17142 -32 17206 -28
rect 17222 28 17286 32
rect 17222 -28 17226 28
rect 17226 -28 17282 28
rect 17282 -28 17286 28
rect 17222 -32 17286 -28
rect 17302 28 17366 32
rect 17302 -28 17306 28
rect 17306 -28 17362 28
rect 17362 -28 17366 28
rect 17302 -32 17366 -28
<< metal4 >>
rect 3104 10368 3424 10928
rect 3104 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3272 10368
rect 3336 10304 3352 10368
rect 3416 10304 3424 10368
rect 3104 10160 3424 10304
rect 3104 9924 3146 10160
rect 3382 9924 3424 10160
rect 3104 9280 3424 9924
rect 3104 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3272 9280
rect 3336 9216 3352 9280
rect 3416 9216 3424 9280
rect 3104 8192 3424 9216
rect 3104 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3272 8192
rect 3336 8128 3352 8192
rect 3416 8128 3424 8192
rect 3104 7104 3424 8128
rect 3104 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3272 7104
rect 3336 7040 3352 7104
rect 3416 7040 3424 7104
rect 3104 6780 3424 7040
rect 3104 6544 3146 6780
rect 3382 6544 3424 6780
rect 3104 6016 3424 6544
rect 3104 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3272 6016
rect 3336 5952 3352 6016
rect 3416 5952 3424 6016
rect 3104 4928 3424 5952
rect 3104 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3272 4928
rect 3336 4864 3352 4928
rect 3416 4864 3424 4928
rect 3104 3840 3424 4864
rect 3104 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3272 3840
rect 3336 3776 3352 3840
rect 3416 3776 3424 3840
rect 3104 3400 3424 3776
rect 3104 3164 3146 3400
rect 3382 3164 3424 3400
rect 3104 2752 3424 3164
rect 3104 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3272 2752
rect 3336 2688 3352 2752
rect 3416 2688 3424 2752
rect 3104 1664 3424 2688
rect 3104 1600 3112 1664
rect 3176 1600 3192 1664
rect 3256 1600 3272 1664
rect 3336 1600 3352 1664
rect 3416 1600 3424 1664
rect 3104 576 3424 1600
rect 3104 512 3112 576
rect 3176 512 3192 576
rect 3256 512 3272 576
rect 3336 512 3352 576
rect 3416 512 3424 576
rect 3104 -48 3424 512
rect 4654 10912 4974 10928
rect 4654 10848 4662 10912
rect 4726 10848 4742 10912
rect 4806 10848 4822 10912
rect 4886 10848 4902 10912
rect 4966 10848 4974 10912
rect 4654 9824 4974 10848
rect 4654 9760 4662 9824
rect 4726 9760 4742 9824
rect 4806 9760 4822 9824
rect 4886 9760 4902 9824
rect 4966 9760 4974 9824
rect 4654 8736 4974 9760
rect 4654 8672 4662 8736
rect 4726 8672 4742 8736
rect 4806 8672 4822 8736
rect 4886 8672 4902 8736
rect 4966 8672 4974 8736
rect 4654 8470 4974 8672
rect 4654 8234 4696 8470
rect 4932 8234 4974 8470
rect 4654 7648 4974 8234
rect 4654 7584 4662 7648
rect 4726 7584 4742 7648
rect 4806 7584 4822 7648
rect 4886 7584 4902 7648
rect 4966 7584 4974 7648
rect 4654 6560 4974 7584
rect 4654 6496 4662 6560
rect 4726 6496 4742 6560
rect 4806 6496 4822 6560
rect 4886 6496 4902 6560
rect 4966 6496 4974 6560
rect 4654 5472 4974 6496
rect 4654 5408 4662 5472
rect 4726 5408 4742 5472
rect 4806 5408 4822 5472
rect 4886 5408 4902 5472
rect 4966 5408 4974 5472
rect 4654 5090 4974 5408
rect 4654 4854 4696 5090
rect 4932 4854 4974 5090
rect 4654 4384 4974 4854
rect 4654 4320 4662 4384
rect 4726 4320 4742 4384
rect 4806 4320 4822 4384
rect 4886 4320 4902 4384
rect 4966 4320 4974 4384
rect 4654 3296 4974 4320
rect 4654 3232 4662 3296
rect 4726 3232 4742 3296
rect 4806 3232 4822 3296
rect 4886 3232 4902 3296
rect 4966 3232 4974 3296
rect 4654 2208 4974 3232
rect 4654 2144 4662 2208
rect 4726 2144 4742 2208
rect 4806 2144 4822 2208
rect 4886 2144 4902 2208
rect 4966 2144 4974 2208
rect 4654 1120 4974 2144
rect 4654 1056 4662 1120
rect 4726 1056 4742 1120
rect 4806 1056 4822 1120
rect 4886 1056 4902 1120
rect 4966 1056 4974 1120
rect 4654 32 4974 1056
rect 4654 -32 4662 32
rect 4726 -32 4742 32
rect 4806 -32 4822 32
rect 4886 -32 4902 32
rect 4966 -32 4974 32
rect 4654 -48 4974 -32
rect 6204 10368 6524 10928
rect 6204 10304 6212 10368
rect 6276 10304 6292 10368
rect 6356 10304 6372 10368
rect 6436 10304 6452 10368
rect 6516 10304 6524 10368
rect 6204 10160 6524 10304
rect 6204 9924 6246 10160
rect 6482 9924 6524 10160
rect 6204 9280 6524 9924
rect 6204 9216 6212 9280
rect 6276 9216 6292 9280
rect 6356 9216 6372 9280
rect 6436 9216 6452 9280
rect 6516 9216 6524 9280
rect 6204 8192 6524 9216
rect 6204 8128 6212 8192
rect 6276 8128 6292 8192
rect 6356 8128 6372 8192
rect 6436 8128 6452 8192
rect 6516 8128 6524 8192
rect 6204 7104 6524 8128
rect 6204 7040 6212 7104
rect 6276 7040 6292 7104
rect 6356 7040 6372 7104
rect 6436 7040 6452 7104
rect 6516 7040 6524 7104
rect 6204 6780 6524 7040
rect 6204 6544 6246 6780
rect 6482 6544 6524 6780
rect 6204 6016 6524 6544
rect 6204 5952 6212 6016
rect 6276 5952 6292 6016
rect 6356 5952 6372 6016
rect 6436 5952 6452 6016
rect 6516 5952 6524 6016
rect 6204 4928 6524 5952
rect 6204 4864 6212 4928
rect 6276 4864 6292 4928
rect 6356 4864 6372 4928
rect 6436 4864 6452 4928
rect 6516 4864 6524 4928
rect 6204 3840 6524 4864
rect 6204 3776 6212 3840
rect 6276 3776 6292 3840
rect 6356 3776 6372 3840
rect 6436 3776 6452 3840
rect 6516 3776 6524 3840
rect 6204 3400 6524 3776
rect 6204 3164 6246 3400
rect 6482 3164 6524 3400
rect 6204 2752 6524 3164
rect 6204 2688 6212 2752
rect 6276 2688 6292 2752
rect 6356 2688 6372 2752
rect 6436 2688 6452 2752
rect 6516 2688 6524 2752
rect 6204 1664 6524 2688
rect 6204 1600 6212 1664
rect 6276 1600 6292 1664
rect 6356 1600 6372 1664
rect 6436 1600 6452 1664
rect 6516 1600 6524 1664
rect 6204 576 6524 1600
rect 6204 512 6212 576
rect 6276 512 6292 576
rect 6356 512 6372 576
rect 6436 512 6452 576
rect 6516 512 6524 576
rect 6204 -48 6524 512
rect 7754 10912 8074 10928
rect 7754 10848 7762 10912
rect 7826 10848 7842 10912
rect 7906 10848 7922 10912
rect 7986 10848 8002 10912
rect 8066 10848 8074 10912
rect 7754 9824 8074 10848
rect 7754 9760 7762 9824
rect 7826 9760 7842 9824
rect 7906 9760 7922 9824
rect 7986 9760 8002 9824
rect 8066 9760 8074 9824
rect 7754 8736 8074 9760
rect 7754 8672 7762 8736
rect 7826 8672 7842 8736
rect 7906 8672 7922 8736
rect 7986 8672 8002 8736
rect 8066 8672 8074 8736
rect 7754 8470 8074 8672
rect 7754 8234 7796 8470
rect 8032 8234 8074 8470
rect 7754 7648 8074 8234
rect 7754 7584 7762 7648
rect 7826 7584 7842 7648
rect 7906 7584 7922 7648
rect 7986 7584 8002 7648
rect 8066 7584 8074 7648
rect 7754 6560 8074 7584
rect 7754 6496 7762 6560
rect 7826 6496 7842 6560
rect 7906 6496 7922 6560
rect 7986 6496 8002 6560
rect 8066 6496 8074 6560
rect 7754 5472 8074 6496
rect 7754 5408 7762 5472
rect 7826 5408 7842 5472
rect 7906 5408 7922 5472
rect 7986 5408 8002 5472
rect 8066 5408 8074 5472
rect 7754 5090 8074 5408
rect 7754 4854 7796 5090
rect 8032 4854 8074 5090
rect 7754 4384 8074 4854
rect 7754 4320 7762 4384
rect 7826 4320 7842 4384
rect 7906 4320 7922 4384
rect 7986 4320 8002 4384
rect 8066 4320 8074 4384
rect 7754 3296 8074 4320
rect 7754 3232 7762 3296
rect 7826 3232 7842 3296
rect 7906 3232 7922 3296
rect 7986 3232 8002 3296
rect 8066 3232 8074 3296
rect 7754 2208 8074 3232
rect 7754 2144 7762 2208
rect 7826 2144 7842 2208
rect 7906 2144 7922 2208
rect 7986 2144 8002 2208
rect 8066 2144 8074 2208
rect 7754 1120 8074 2144
rect 7754 1056 7762 1120
rect 7826 1056 7842 1120
rect 7906 1056 7922 1120
rect 7986 1056 8002 1120
rect 8066 1056 8074 1120
rect 7754 32 8074 1056
rect 7754 -32 7762 32
rect 7826 -32 7842 32
rect 7906 -32 7922 32
rect 7986 -32 8002 32
rect 8066 -32 8074 32
rect 7754 -48 8074 -32
rect 9304 10368 9624 10928
rect 9304 10304 9312 10368
rect 9376 10304 9392 10368
rect 9456 10304 9472 10368
rect 9536 10304 9552 10368
rect 9616 10304 9624 10368
rect 9304 10160 9624 10304
rect 9304 9924 9346 10160
rect 9582 9924 9624 10160
rect 9304 9280 9624 9924
rect 9304 9216 9312 9280
rect 9376 9216 9392 9280
rect 9456 9216 9472 9280
rect 9536 9216 9552 9280
rect 9616 9216 9624 9280
rect 9304 8192 9624 9216
rect 9304 8128 9312 8192
rect 9376 8128 9392 8192
rect 9456 8128 9472 8192
rect 9536 8128 9552 8192
rect 9616 8128 9624 8192
rect 9304 7104 9624 8128
rect 9304 7040 9312 7104
rect 9376 7040 9392 7104
rect 9456 7040 9472 7104
rect 9536 7040 9552 7104
rect 9616 7040 9624 7104
rect 9304 6780 9624 7040
rect 9304 6544 9346 6780
rect 9582 6544 9624 6780
rect 9304 6016 9624 6544
rect 9304 5952 9312 6016
rect 9376 5952 9392 6016
rect 9456 5952 9472 6016
rect 9536 5952 9552 6016
rect 9616 5952 9624 6016
rect 9304 4928 9624 5952
rect 9304 4864 9312 4928
rect 9376 4864 9392 4928
rect 9456 4864 9472 4928
rect 9536 4864 9552 4928
rect 9616 4864 9624 4928
rect 9304 3840 9624 4864
rect 9304 3776 9312 3840
rect 9376 3776 9392 3840
rect 9456 3776 9472 3840
rect 9536 3776 9552 3840
rect 9616 3776 9624 3840
rect 9304 3400 9624 3776
rect 9304 3164 9346 3400
rect 9582 3164 9624 3400
rect 9304 2752 9624 3164
rect 9304 2688 9312 2752
rect 9376 2688 9392 2752
rect 9456 2688 9472 2752
rect 9536 2688 9552 2752
rect 9616 2688 9624 2752
rect 9304 1664 9624 2688
rect 9304 1600 9312 1664
rect 9376 1600 9392 1664
rect 9456 1600 9472 1664
rect 9536 1600 9552 1664
rect 9616 1600 9624 1664
rect 9304 576 9624 1600
rect 9304 512 9312 576
rect 9376 512 9392 576
rect 9456 512 9472 576
rect 9536 512 9552 576
rect 9616 512 9624 576
rect 9304 -48 9624 512
rect 10854 10912 11174 10928
rect 10854 10848 10862 10912
rect 10926 10848 10942 10912
rect 11006 10848 11022 10912
rect 11086 10848 11102 10912
rect 11166 10848 11174 10912
rect 10854 9824 11174 10848
rect 10854 9760 10862 9824
rect 10926 9760 10942 9824
rect 11006 9760 11022 9824
rect 11086 9760 11102 9824
rect 11166 9760 11174 9824
rect 10854 8736 11174 9760
rect 10854 8672 10862 8736
rect 10926 8672 10942 8736
rect 11006 8672 11022 8736
rect 11086 8672 11102 8736
rect 11166 8672 11174 8736
rect 10854 8470 11174 8672
rect 10854 8234 10896 8470
rect 11132 8234 11174 8470
rect 10854 7648 11174 8234
rect 10854 7584 10862 7648
rect 10926 7584 10942 7648
rect 11006 7584 11022 7648
rect 11086 7584 11102 7648
rect 11166 7584 11174 7648
rect 10854 6560 11174 7584
rect 10854 6496 10862 6560
rect 10926 6496 10942 6560
rect 11006 6496 11022 6560
rect 11086 6496 11102 6560
rect 11166 6496 11174 6560
rect 10854 5472 11174 6496
rect 10854 5408 10862 5472
rect 10926 5408 10942 5472
rect 11006 5408 11022 5472
rect 11086 5408 11102 5472
rect 11166 5408 11174 5472
rect 10854 5090 11174 5408
rect 10854 4854 10896 5090
rect 11132 4854 11174 5090
rect 10854 4384 11174 4854
rect 10854 4320 10862 4384
rect 10926 4320 10942 4384
rect 11006 4320 11022 4384
rect 11086 4320 11102 4384
rect 11166 4320 11174 4384
rect 10854 3296 11174 4320
rect 10854 3232 10862 3296
rect 10926 3232 10942 3296
rect 11006 3232 11022 3296
rect 11086 3232 11102 3296
rect 11166 3232 11174 3296
rect 10854 2208 11174 3232
rect 10854 2144 10862 2208
rect 10926 2144 10942 2208
rect 11006 2144 11022 2208
rect 11086 2144 11102 2208
rect 11166 2144 11174 2208
rect 10854 1120 11174 2144
rect 10854 1056 10862 1120
rect 10926 1056 10942 1120
rect 11006 1056 11022 1120
rect 11086 1056 11102 1120
rect 11166 1056 11174 1120
rect 10854 32 11174 1056
rect 10854 -32 10862 32
rect 10926 -32 10942 32
rect 11006 -32 11022 32
rect 11086 -32 11102 32
rect 11166 -32 11174 32
rect 10854 -48 11174 -32
rect 12404 10368 12724 10928
rect 12404 10304 12412 10368
rect 12476 10304 12492 10368
rect 12556 10304 12572 10368
rect 12636 10304 12652 10368
rect 12716 10304 12724 10368
rect 12404 10160 12724 10304
rect 12404 9924 12446 10160
rect 12682 9924 12724 10160
rect 12404 9280 12724 9924
rect 12404 9216 12412 9280
rect 12476 9216 12492 9280
rect 12556 9216 12572 9280
rect 12636 9216 12652 9280
rect 12716 9216 12724 9280
rect 12404 8192 12724 9216
rect 12404 8128 12412 8192
rect 12476 8128 12492 8192
rect 12556 8128 12572 8192
rect 12636 8128 12652 8192
rect 12716 8128 12724 8192
rect 12404 7104 12724 8128
rect 12404 7040 12412 7104
rect 12476 7040 12492 7104
rect 12556 7040 12572 7104
rect 12636 7040 12652 7104
rect 12716 7040 12724 7104
rect 12404 6780 12724 7040
rect 12404 6544 12446 6780
rect 12682 6544 12724 6780
rect 12404 6016 12724 6544
rect 12404 5952 12412 6016
rect 12476 5952 12492 6016
rect 12556 5952 12572 6016
rect 12636 5952 12652 6016
rect 12716 5952 12724 6016
rect 12404 4928 12724 5952
rect 12404 4864 12412 4928
rect 12476 4864 12492 4928
rect 12556 4864 12572 4928
rect 12636 4864 12652 4928
rect 12716 4864 12724 4928
rect 12404 3840 12724 4864
rect 12404 3776 12412 3840
rect 12476 3776 12492 3840
rect 12556 3776 12572 3840
rect 12636 3776 12652 3840
rect 12716 3776 12724 3840
rect 12404 3400 12724 3776
rect 12404 3164 12446 3400
rect 12682 3164 12724 3400
rect 12404 2752 12724 3164
rect 12404 2688 12412 2752
rect 12476 2688 12492 2752
rect 12556 2688 12572 2752
rect 12636 2688 12652 2752
rect 12716 2688 12724 2752
rect 12404 1664 12724 2688
rect 12404 1600 12412 1664
rect 12476 1600 12492 1664
rect 12556 1600 12572 1664
rect 12636 1600 12652 1664
rect 12716 1600 12724 1664
rect 12404 576 12724 1600
rect 12404 512 12412 576
rect 12476 512 12492 576
rect 12556 512 12572 576
rect 12636 512 12652 576
rect 12716 512 12724 576
rect 12404 -48 12724 512
rect 13954 10912 14274 10928
rect 13954 10848 13962 10912
rect 14026 10848 14042 10912
rect 14106 10848 14122 10912
rect 14186 10848 14202 10912
rect 14266 10848 14274 10912
rect 13954 9824 14274 10848
rect 13954 9760 13962 9824
rect 14026 9760 14042 9824
rect 14106 9760 14122 9824
rect 14186 9760 14202 9824
rect 14266 9760 14274 9824
rect 13954 8736 14274 9760
rect 13954 8672 13962 8736
rect 14026 8672 14042 8736
rect 14106 8672 14122 8736
rect 14186 8672 14202 8736
rect 14266 8672 14274 8736
rect 13954 8470 14274 8672
rect 13954 8234 13996 8470
rect 14232 8234 14274 8470
rect 13954 7648 14274 8234
rect 13954 7584 13962 7648
rect 14026 7584 14042 7648
rect 14106 7584 14122 7648
rect 14186 7584 14202 7648
rect 14266 7584 14274 7648
rect 13954 6560 14274 7584
rect 13954 6496 13962 6560
rect 14026 6496 14042 6560
rect 14106 6496 14122 6560
rect 14186 6496 14202 6560
rect 14266 6496 14274 6560
rect 13954 5472 14274 6496
rect 13954 5408 13962 5472
rect 14026 5408 14042 5472
rect 14106 5408 14122 5472
rect 14186 5408 14202 5472
rect 14266 5408 14274 5472
rect 13954 5090 14274 5408
rect 13954 4854 13996 5090
rect 14232 4854 14274 5090
rect 13954 4384 14274 4854
rect 13954 4320 13962 4384
rect 14026 4320 14042 4384
rect 14106 4320 14122 4384
rect 14186 4320 14202 4384
rect 14266 4320 14274 4384
rect 13954 3296 14274 4320
rect 13954 3232 13962 3296
rect 14026 3232 14042 3296
rect 14106 3232 14122 3296
rect 14186 3232 14202 3296
rect 14266 3232 14274 3296
rect 13954 2208 14274 3232
rect 13954 2144 13962 2208
rect 14026 2144 14042 2208
rect 14106 2144 14122 2208
rect 14186 2144 14202 2208
rect 14266 2144 14274 2208
rect 13954 1120 14274 2144
rect 13954 1056 13962 1120
rect 14026 1056 14042 1120
rect 14106 1056 14122 1120
rect 14186 1056 14202 1120
rect 14266 1056 14274 1120
rect 13954 32 14274 1056
rect 13954 -32 13962 32
rect 14026 -32 14042 32
rect 14106 -32 14122 32
rect 14186 -32 14202 32
rect 14266 -32 14274 32
rect 13954 -48 14274 -32
rect 15504 10368 15824 10928
rect 15504 10304 15512 10368
rect 15576 10304 15592 10368
rect 15656 10304 15672 10368
rect 15736 10304 15752 10368
rect 15816 10304 15824 10368
rect 15504 10160 15824 10304
rect 15504 9924 15546 10160
rect 15782 9924 15824 10160
rect 15504 9280 15824 9924
rect 15504 9216 15512 9280
rect 15576 9216 15592 9280
rect 15656 9216 15672 9280
rect 15736 9216 15752 9280
rect 15816 9216 15824 9280
rect 15504 8192 15824 9216
rect 15504 8128 15512 8192
rect 15576 8128 15592 8192
rect 15656 8128 15672 8192
rect 15736 8128 15752 8192
rect 15816 8128 15824 8192
rect 15504 7104 15824 8128
rect 15504 7040 15512 7104
rect 15576 7040 15592 7104
rect 15656 7040 15672 7104
rect 15736 7040 15752 7104
rect 15816 7040 15824 7104
rect 15504 6780 15824 7040
rect 15504 6544 15546 6780
rect 15782 6544 15824 6780
rect 15504 6016 15824 6544
rect 15504 5952 15512 6016
rect 15576 5952 15592 6016
rect 15656 5952 15672 6016
rect 15736 5952 15752 6016
rect 15816 5952 15824 6016
rect 15504 4928 15824 5952
rect 15504 4864 15512 4928
rect 15576 4864 15592 4928
rect 15656 4864 15672 4928
rect 15736 4864 15752 4928
rect 15816 4864 15824 4928
rect 15504 3840 15824 4864
rect 15504 3776 15512 3840
rect 15576 3776 15592 3840
rect 15656 3776 15672 3840
rect 15736 3776 15752 3840
rect 15816 3776 15824 3840
rect 15504 3400 15824 3776
rect 15504 3164 15546 3400
rect 15782 3164 15824 3400
rect 15504 2752 15824 3164
rect 15504 2688 15512 2752
rect 15576 2688 15592 2752
rect 15656 2688 15672 2752
rect 15736 2688 15752 2752
rect 15816 2688 15824 2752
rect 15504 1664 15824 2688
rect 15504 1600 15512 1664
rect 15576 1600 15592 1664
rect 15656 1600 15672 1664
rect 15736 1600 15752 1664
rect 15816 1600 15824 1664
rect 15504 576 15824 1600
rect 15504 512 15512 576
rect 15576 512 15592 576
rect 15656 512 15672 576
rect 15736 512 15752 576
rect 15816 512 15824 576
rect 15504 -48 15824 512
rect 17054 10912 17374 10928
rect 17054 10848 17062 10912
rect 17126 10848 17142 10912
rect 17206 10848 17222 10912
rect 17286 10848 17302 10912
rect 17366 10848 17374 10912
rect 17054 9824 17374 10848
rect 17054 9760 17062 9824
rect 17126 9760 17142 9824
rect 17206 9760 17222 9824
rect 17286 9760 17302 9824
rect 17366 9760 17374 9824
rect 17054 8736 17374 9760
rect 17054 8672 17062 8736
rect 17126 8672 17142 8736
rect 17206 8672 17222 8736
rect 17286 8672 17302 8736
rect 17366 8672 17374 8736
rect 17054 8470 17374 8672
rect 17054 8234 17096 8470
rect 17332 8234 17374 8470
rect 17054 7648 17374 8234
rect 17054 7584 17062 7648
rect 17126 7584 17142 7648
rect 17206 7584 17222 7648
rect 17286 7584 17302 7648
rect 17366 7584 17374 7648
rect 17054 6560 17374 7584
rect 17054 6496 17062 6560
rect 17126 6496 17142 6560
rect 17206 6496 17222 6560
rect 17286 6496 17302 6560
rect 17366 6496 17374 6560
rect 17054 5472 17374 6496
rect 17054 5408 17062 5472
rect 17126 5408 17142 5472
rect 17206 5408 17222 5472
rect 17286 5408 17302 5472
rect 17366 5408 17374 5472
rect 17054 5090 17374 5408
rect 17054 4854 17096 5090
rect 17332 4854 17374 5090
rect 17054 4384 17374 4854
rect 17054 4320 17062 4384
rect 17126 4320 17142 4384
rect 17206 4320 17222 4384
rect 17286 4320 17302 4384
rect 17366 4320 17374 4384
rect 17054 3296 17374 4320
rect 17054 3232 17062 3296
rect 17126 3232 17142 3296
rect 17206 3232 17222 3296
rect 17286 3232 17302 3296
rect 17366 3232 17374 3296
rect 17054 2208 17374 3232
rect 17054 2144 17062 2208
rect 17126 2144 17142 2208
rect 17206 2144 17222 2208
rect 17286 2144 17302 2208
rect 17366 2144 17374 2208
rect 17054 1120 17374 2144
rect 17054 1056 17062 1120
rect 17126 1056 17142 1120
rect 17206 1056 17222 1120
rect 17286 1056 17302 1120
rect 17366 1056 17374 1120
rect 17054 32 17374 1056
rect 17054 -32 17062 32
rect 17126 -32 17142 32
rect 17206 -32 17222 32
rect 17286 -32 17302 32
rect 17366 -32 17374 32
rect 17054 -48 17374 -32
<< via4 >>
rect 3146 9924 3382 10160
rect 3146 6544 3382 6780
rect 3146 3164 3382 3400
rect 4696 8234 4932 8470
rect 4696 4854 4932 5090
rect 6246 9924 6482 10160
rect 6246 6544 6482 6780
rect 6246 3164 6482 3400
rect 7796 8234 8032 8470
rect 7796 4854 8032 5090
rect 9346 9924 9582 10160
rect 9346 6544 9582 6780
rect 9346 3164 9582 3400
rect 10896 8234 11132 8470
rect 10896 4854 11132 5090
rect 12446 9924 12682 10160
rect 12446 6544 12682 6780
rect 12446 3164 12682 3400
rect 13996 8234 14232 8470
rect 13996 4854 14232 5090
rect 15546 9924 15782 10160
rect 15546 6544 15782 6780
rect 15546 3164 15782 3400
rect 17096 8234 17332 8470
rect 17096 4854 17332 5090
<< metal5 >>
rect 0 10160 18860 10202
rect 0 9924 3146 10160
rect 3382 9924 6246 10160
rect 6482 9924 9346 10160
rect 9582 9924 12446 10160
rect 12682 9924 15546 10160
rect 15782 9924 18860 10160
rect 0 9882 18860 9924
rect 0 8470 18860 8512
rect 0 8234 4696 8470
rect 4932 8234 7796 8470
rect 8032 8234 10896 8470
rect 11132 8234 13996 8470
rect 14232 8234 17096 8470
rect 17332 8234 18860 8470
rect 0 8192 18860 8234
rect 0 6780 18860 6822
rect 0 6544 3146 6780
rect 3382 6544 6246 6780
rect 6482 6544 9346 6780
rect 9582 6544 12446 6780
rect 12682 6544 15546 6780
rect 15782 6544 18860 6780
rect 0 6502 18860 6544
rect 0 5090 18860 5132
rect 0 4854 4696 5090
rect 4932 4854 7796 5090
rect 8032 4854 10896 5090
rect 11132 4854 13996 5090
rect 14232 4854 17096 5090
rect 17332 4854 18860 5090
rect 0 4812 18860 4854
rect 0 3400 18860 3442
rect 0 3164 3146 3400
rect 3382 3164 6246 3400
rect 6482 3164 9346 3400
rect 9582 3164 12446 3400
rect 12682 3164 15546 3400
rect 15782 3164 18860 3400
rect 0 3122 18860 3164
use sky130_fd_sc_hd__decap_8  FILLER_0_15 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 1380 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 2116 0 1 0
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 276 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1636915332
transform 1 0 1380 0 -1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1636915332
transform 1 0 276 0 -1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_0 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 0 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1636915332
transform 1 0 0 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _336_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 3312 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _334__6 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 2300 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 2576 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_36 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 3312 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_31 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 2852 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_27
timestamp 1636915332
transform 1 0 2484 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _335_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 4232 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _311_
timestamp 1636915332
transform -1 0 3956 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_46
timestamp 1636915332
transform 1 0 4232 0 -1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dfstp_1  _441_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 2668 0 1 0
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _382_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 5612 0 1 0
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _355_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 5244 0 -1 1088
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1636915332
transform 1 0 5152 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1636915332
transform 1 0 5152 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1636915332
transform 1 0 4968 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57
timestamp 1636915332
transform 1 0 5244 0 1 0
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 4600 0 1 0
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _381_
timestamp 1636915332
transform 1 0 5980 0 -1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_1_74
timestamp 1636915332
transform 1 0 6808 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_64
timestamp 1636915332
transform 1 0 5888 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_70
timestamp 1636915332
transform 1 0 6440 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1636915332
transform 1 0 7544 0 1 0
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_85
timestamp 1636915332
transform 1 0 7820 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1636915332
transform 1 0 7728 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_1  _289_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 9200 0 1 0
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _290_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 8832 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _402_
timestamp 1636915332
transform 1 0 9108 0 -1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__dfstp_1  _452_
timestamp 1636915332
transform 1 0 7176 0 -1 1088
box -38 -48 1970 592
use sky130_fd_sc_hd__nor2_1  _360_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 10304 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_108
timestamp 1636915332
transform 1 0 9936 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _401_
timestamp 1636915332
transform 1 0 10488 0 -1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _359_
timestamp 1636915332
transform 1 0 10396 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _275_
timestamp 1636915332
transform 1 0 11316 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1636915332
transform 1 0 10304 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1636915332
transform 1 0 10304 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_113
timestamp 1636915332
transform 1 0 10396 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_120
timestamp 1636915332
transform 1 0 11040 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_100
timestamp 1636915332
transform 1 0 9200 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_132
timestamp 1636915332
transform 1 0 12144 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_1_126
timestamp 1636915332
transform 1 0 11592 0 -1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1636915332
transform 1 0 12880 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_1  _291_
timestamp 1636915332
transform 1 0 12144 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _292_
timestamp 1636915332
transform 1 0 12512 0 -1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _405_
timestamp 1636915332
transform 1 0 13248 0 -1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__dfrtp_2  _451_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 12972 0 1 0
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_6  FILLER_0_162
timestamp 1636915332
transform 1 0 14904 0 1 0
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_169
timestamp 1636915332
transform 1 0 15548 0 1 0
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_157
timestamp 1636915332
transform 1 0 14444 0 -1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_165
timestamp 1636915332
transform 1 0 15180 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1636915332
transform 1 0 15456 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1636915332
transform 1 0 15456 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_1  _329_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 16100 0 -1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_2  _358_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 14444 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _325_
timestamp 1636915332
transform -1 0 17296 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_183
timestamp 1636915332
transform 1 0 16836 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_175
timestamp 1636915332
transform 1 0 16100 0 -1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__or2b_1  _324_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 18400 0 -1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _323_
timestamp 1636915332
transform -1 0 17848 0 -1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1636915332
transform 1 0 18032 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1636915332
transform 1 0 18124 0 1 0
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1636915332
transform 1 0 17940 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_191
timestamp 1636915332
transform 1 0 17572 0 1 0
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _415_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 16100 0 1 0
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_1_200
timestamp 1636915332
transform 1 0 18400 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1636915332
transform -1 0 18860 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1636915332
transform -1 0 18860 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input1 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 18308 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3
timestamp 1636915332
transform 1 0 276 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_7
timestamp 1636915332
transform 1 0 644 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1636915332
transform 1 0 0 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtn_1  _442_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 736 0 1 1088
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_2_29
timestamp 1636915332
transform 1 0 2668 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_34
timestamp 1636915332
transform 1 0 3128 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_45
timestamp 1636915332
transform 1 0 4140 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1636915332
transform 1 0 2576 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__nor3b_2  _308_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 5336 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _310_
timestamp 1636915332
transform -1 0 3864 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _312_
timestamp 1636915332
transform 1 0 3220 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _332_
timestamp 1636915332
transform -1 0 4140 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _333_
timestamp 1636915332
transform -1 0 3128 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _356_
timestamp 1636915332
transform -1 0 5612 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _407_
timestamp 1636915332
transform 1 0 5612 0 1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer9 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 6440 0 1 1088
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1636915332
transform 1 0 7084 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1636915332
transform 1 0 7636 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_85
timestamp 1636915332
transform 1 0 7820 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_91
timestamp 1636915332
transform 1 0 8372 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1636915332
transform 1 0 7728 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__a21bo_1  _288_
timestamp 1636915332
transform -1 0 9200 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_100
timestamp 1636915332
transform 1 0 9200 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_108
timestamp 1636915332
transform 1 0 9936 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_116
timestamp 1636915332
transform 1 0 10672 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _274_
timestamp 1636915332
transform 1 0 11224 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _276_
timestamp 1636915332
transform 1 0 10856 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _361_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 10028 0 1 1088
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_2_125
timestamp 1636915332
transform 1 0 11500 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_133
timestamp 1636915332
transform 1 0 12236 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1636915332
transform 1 0 12788 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_141
timestamp 1636915332
transform 1 0 12972 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1636915332
transform 1 0 12880 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _345_
timestamp 1636915332
transform -1 0 12788 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _404_
timestamp 1636915332
transform 1 0 13524 0 1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_2_156
timestamp 1636915332
transform 1 0 14352 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _443_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 16560 0 1 1088
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1636915332
transform 1 0 18032 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _374_
timestamp 1636915332
transform -1 0 18400 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _414_
timestamp 1636915332
transform 1 0 16560 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_2_200
timestamp 1636915332
transform 1 0 18400 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1636915332
transform -1 0 18860 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1636915332
transform 1 0 1380 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1636915332
transform 1 0 276 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1636915332
transform 1 0 0 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_27
timestamp 1636915332
transform 1 0 2484 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_35
timestamp 1636915332
transform 1 0 3220 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _337_
timestamp 1636915332
transform -1 0 3680 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _338_
timestamp 1636915332
transform -1 0 3956 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _386_
timestamp 1636915332
transform 1 0 3956 0 -1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_3_52
timestamp 1636915332
transform 1 0 4784 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_64
timestamp 1636915332
transform 1 0 5888 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_74
timestamp 1636915332
transform 1 0 6808 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1636915332
transform 1 0 5152 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__xor2_1  _357_
timestamp 1636915332
transform 1 0 5244 0 -1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _406_
timestamp 1636915332
transform 1 0 5980 0 -1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__dfrtp_1  _453_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 7360 0 -1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  FILLER_3_100
timestamp 1636915332
transform 1 0 9200 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_113
timestamp 1636915332
transform 1 0 10396 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_123
timestamp 1636915332
transform 1 0 11316 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1636915332
transform 1 0 10304 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _398_
timestamp 1636915332
transform 1 0 10488 0 -1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _399_
timestamp 1636915332
transform 1 0 9476 0 -1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_131
timestamp 1636915332
transform 1 0 12052 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_145
timestamp 1636915332
transform 1 0 13340 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__nand3b_1  _279_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 12788 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__o21bai_1  _284_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 13340 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_153
timestamp 1636915332
transform 1 0 14076 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_169
timestamp 1636915332
transform 1 0 15548 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1636915332
transform 1 0 15456 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_1  _278_
timestamp 1636915332
transform 1 0 14904 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _326_
timestamp 1636915332
transform -1 0 14444 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _327_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 14444 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__dfrtp_1  _427_
timestamp 1636915332
transform 1 0 15640 0 -1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_12  FILLER_3_190
timestamp 1636915332
transform 1 0 17480 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1636915332
transform -1 0 18860 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_3
timestamp 1636915332
transform 1 0 276 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_7
timestamp 1636915332
transform 1 0 644 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1636915332
transform 1 0 0 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtn_1  _440_
timestamp 1636915332
transform 1 0 736 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_4_29
timestamp 1636915332
transform 1 0 2668 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_37
timestamp 1636915332
transform 1 0 3404 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1636915332
transform 1 0 2576 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _331_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 4508 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _339_
timestamp 1636915332
transform -1 0 3404 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _385_
timestamp 1636915332
transform 1 0 4508 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_4_58
timestamp 1636915332
transform 1 0 5336 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_67
timestamp 1636915332
transform 1 0 6164 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _309_
timestamp 1636915332
transform 1 0 6532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__o21bai_1  _315_
timestamp 1636915332
transform -1 0 6164 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_75
timestamp 1636915332
transform 1 0 6900 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_79
timestamp 1636915332
transform 1 0 7268 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_85
timestamp 1636915332
transform 1 0 7820 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_97
timestamp 1636915332
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1636915332
transform 1 0 7728 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _281_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 7360 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _287_
timestamp 1636915332
transform -1 0 8924 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_112
timestamp 1636915332
transform 1 0 10304 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_124
timestamp 1636915332
transform 1 0 11408 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _307_
timestamp 1636915332
transform -1 0 10304 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_141
timestamp 1636915332
transform 1 0 12972 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_149
timestamp 1636915332
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1636915332
transform 1 0 12880 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _277_
timestamp 1636915332
transform 1 0 12604 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _285_
timestamp 1636915332
transform -1 0 12604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _349_
timestamp 1636915332
transform 1 0 11592 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_4_172
timestamp 1636915332
transform 1 0 15824 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  _328_
timestamp 1636915332
transform 1 0 15456 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _416_
timestamp 1636915332
transform -1 0 15456 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_4  _430_
timestamp 1636915332
transform -1 0 18032 0 1 2176
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_2  FILLER_4_197
timestamp 1636915332
transform 1 0 18124 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1636915332
transform 1 0 18032 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1636915332
transform -1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1636915332
transform 1 0 18308 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1636915332
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1636915332
transform 1 0 276 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1636915332
transform 1 0 0 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_27
timestamp 1636915332
transform 1 0 2484 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_31
timestamp 1636915332
transform 1 0 2852 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_41
timestamp 1636915332
transform 1 0 3772 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_49
timestamp 1636915332
transform 1 0 4508 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _294_
timestamp 1636915332
transform -1 0 3772 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _302_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 2944 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1636915332
transform 1 0 5060 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_57
timestamp 1636915332
transform 1 0 5244 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_68
timestamp 1636915332
transform 1 0 6256 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1636915332
transform 1 0 5152 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _280_
timestamp 1636915332
transform 1 0 4784 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _314_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 5980 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _330_
timestamp 1636915332
transform -1 0 6256 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_76
timestamp 1636915332
transform 1 0 6992 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_86
timestamp 1636915332
transform 1 0 7912 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _283_
timestamp 1636915332
transform 1 0 8004 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _286_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 7084 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _316_
timestamp 1636915332
transform -1 0 7912 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dfstp_1  _447_
timestamp 1636915332
transform 1 0 8372 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1636915332
transform 1 0 10304 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_1  _454_
timestamp 1636915332
transform 1 0 10396 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_5_134
timestamp 1636915332
transform 1 0 12328 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_144
timestamp 1636915332
transform 1 0 13248 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__and2b_2  _350_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 14076 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__o21bai_2  _351_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 13248 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_5_162
timestamp 1636915332
transform 1 0 14904 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_169
timestamp 1636915332
transform 1 0 15548 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1636915332
transform 1 0 15456 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _411_
timestamp 1636915332
transform 1 0 14076 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__dfstp_1  _428_
timestamp 1636915332
transform -1 0 17848 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer4
timestamp 1636915332
transform 1 0 17848 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_5_201
timestamp 1636915332
transform 1 0 18492 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1636915332
transform -1 0 18860 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_3
timestamp 1636915332
transform 1 0 276 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_7
timestamp 1636915332
transform 1 0 644 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1636915332
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1636915332
transform 1 0 276 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1636915332
transform 1 0 0 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1636915332
transform 1 0 0 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtn_1  _448_
timestamp 1636915332
transform 1 0 736 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_6_37
timestamp 1636915332
transform 1 0 3404 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_27
timestamp 1636915332
transform 1 0 2484 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1636915332
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1636915332
transform 1 0 2576 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__o21bai_1  _295_
timestamp 1636915332
transform 1 0 3588 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nand3b_1  _296_
timestamp 1636915332
transform -1 0 4692 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _303_
timestamp 1636915332
transform -1 0 3588 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _304_
timestamp 1636915332
transform -1 0 3404 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  rebuffer3 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 5060 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _313_
timestamp 1636915332
transform 1 0 4876 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2ai_1  _300_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 5244 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1636915332
transform 1 0 5152 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_57
timestamp 1636915332
transform 1 0 5244 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_51
timestamp 1636915332
transform 1 0 4692 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_55
timestamp 1636915332
transform 1 0 5060 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__dlymetal6s2s_1  rebuffer8
timestamp 1636915332
transform -1 0 6716 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _397_
timestamp 1636915332
transform 1 0 6256 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _293_
timestamp 1636915332
transform 1 0 5888 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_67
timestamp 1636915332
transform 1 0 6164 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _299_
timestamp 1636915332
transform 1 0 6716 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer11
timestamp 1636915332
transform 1 0 7084 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _306_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 7544 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1636915332
transform 1 0 7728 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_82
timestamp 1636915332
transform 1 0 7544 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_76
timestamp 1636915332
transform 1 0 6992 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer7
timestamp 1636915332
transform -1 0 9108 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _322_
timestamp 1636915332
transform -1 0 8096 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _321_
timestamp 1636915332
transform 1 0 8372 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_2  _282_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 8464 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_7_88
timestamp 1636915332
transform 1 0 8096 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _305__5
timestamp 1636915332
transform 1 0 9108 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _400_
timestamp 1636915332
transform 1 0 9200 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkinv_2  _362_
timestamp 1636915332
transform -1 0 9844 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_109
timestamp 1636915332
transform 1 0 10028 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_107
timestamp 1636915332
transform 1 0 9844 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_102
timestamp 1636915332
transform 1 0 9384 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _403_
timestamp 1636915332
transform 1 0 11224 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _363_
timestamp 1636915332
transform 1 0 10396 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _319_
timestamp 1636915332
transform 1 0 10396 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1636915332
transform 1 0 10304 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_120
timestamp 1636915332
transform 1 0 11040 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_132
timestamp 1636915332
transform 1 0 12144 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_141
timestamp 1636915332
transform 1 0 12972 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_149
timestamp 1636915332
transform 1 0 13708 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_140
timestamp 1636915332
transform 1 0 12880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1636915332
transform 1 0 12880 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__nand3b_1  _341_
timestamp 1636915332
transform 1 0 12328 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _342_
timestamp 1636915332
transform 1 0 13156 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _364_
timestamp 1636915332
transform 1 0 12052 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_171
timestamp 1636915332
transform 1 0 15732 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_150
timestamp 1636915332
transform 1 0 13800 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_7_159
timestamp 1636915332
transform 1 0 14628 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1636915332
transform 1 0 15364 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_169
timestamp 1636915332
transform 1 0 15548 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1636915332
transform 1 0 15456 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _348_
timestamp 1636915332
transform 1 0 14352 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_4  _431_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 15824 0 1 3264
box -38 -48 2246 592
use sky130_fd_sc_hd__dfstp_1  _439_
timestamp 1636915332
transform 1 0 13800 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_8  FILLER_7_179
timestamp 1636915332
transform 1 0 16468 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_187
timestamp 1636915332
transform 1 0 17204 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1636915332
transform 1 0 18032 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer5
timestamp 1636915332
transform -1 0 18584 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer6
timestamp 1636915332
transform -1 0 17940 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  split12
timestamp 1636915332
transform -1 0 16468 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  split2
timestamp 1636915332
transform -1 0 18492 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_201
timestamp 1636915332
transform 1 0 18492 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1636915332
transform -1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1636915332
transform -1 0 18860 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_15
timestamp 1636915332
transform 1 0 1380 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_23
timestamp 1636915332
transform 1 0 2116 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1636915332
transform 1 0 276 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1636915332
transform 1 0 0 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1636915332
transform 1 0 2576 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _301__4
timestamp 1636915332
transform 1 0 2300 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  _449_
timestamp 1636915332
transform 1 0 2668 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_2  FILLER_8_53
timestamp 1636915332
transform 1 0 4876 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _298_
timestamp 1636915332
transform -1 0 4876 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtn_1  _450_
timestamp 1636915332
transform -1 0 6900 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_8_75
timestamp 1636915332
transform 1 0 6900 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_80
timestamp 1636915332
transform 1 0 7360 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1636915332
transform 1 0 7728 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_2  _444_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 7820 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_pll_clk
timestamp 1636915332
transform -1 0 7360 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _445_
timestamp 1636915332
transform 1 0 9752 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_8_126
timestamp 1636915332
transform 1 0 11592 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1636915332
transform 1 0 12788 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1636915332
transform 1 0 12972 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1636915332
transform 1 0 12880 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__nor3_1  _317_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 12512 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _340_
timestamp 1636915332
transform 1 0 12512 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _424_
timestamp 1636915332
transform -1 0 15916 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _432_
timestamp 1636915332
transform -1 0 18032 0 1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_2  FILLER_8_197
timestamp 1636915332
transform 1 0 18124 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1636915332
transform 1 0 18032 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1636915332
transform -1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1636915332
transform 1 0 18308 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1636915332
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1636915332
transform 1 0 276 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1636915332
transform 1 0 0 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1636915332
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1636915332
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1636915332
transform 1 0 4692 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1636915332
transform 1 0 5060 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_57
timestamp 1636915332
transform 1 0 5244 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_61
timestamp 1636915332
transform 1 0 5612 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_65
timestamp 1636915332
transform 1 0 5980 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1636915332
transform 1 0 5152 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _297_
timestamp 1636915332
transform 1 0 5704 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_77
timestamp 1636915332
transform 1 0 7084 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_81
timestamp 1636915332
transform 1 0 7452 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_92
timestamp 1636915332
transform 1 0 8464 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _219_
timestamp 1636915332
transform 1 0 8924 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _221_
timestamp 1636915332
transform 1 0 8556 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _370_
timestamp 1636915332
transform -1 0 7820 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _371_
timestamp 1636915332
transform 1 0 7820 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_9_103
timestamp 1636915332
transform 1 0 9476 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_109
timestamp 1636915332
transform 1 0 10028 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_113
timestamp 1636915332
transform 1 0 10396 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_120
timestamp 1636915332
transform 1 0 11040 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1636915332
transform 1 0 10304 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _220_
timestamp 1636915332
transform 1 0 9200 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _320_
timestamp 1636915332
transform -1 0 10028 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_pll_clk
timestamp 1636915332
transform 1 0 10672 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _318_
timestamp 1636915332
transform 1 0 12144 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__dfrtp_1  _446_
timestamp 1636915332
transform -1 0 14628 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_9_159
timestamp 1636915332
transform 1 0 14628 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1636915332
transform 1 0 15364 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_169
timestamp 1636915332
transform 1 0 15548 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1636915332
transform 1 0 15456 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_181
timestamp 1636915332
transform 1 0 16652 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _429_
timestamp 1636915332
transform -1 0 18584 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1636915332
transform -1 0 18860 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_15
timestamp 1636915332
transform 1 0 1380 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_23
timestamp 1636915332
transform 1 0 2116 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1636915332
transform 1 0 276 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1636915332
transform 1 0 0 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1636915332
transform 1 0 2576 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _242__1
timestamp 1636915332
transform 1 0 2300 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  _461_
timestamp 1636915332
transform 1 0 2668 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_12  FILLER_10_50
timestamp 1636915332
transform 1 0 4600 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_62
timestamp 1636915332
transform 1 0 5704 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_1  _464_
timestamp 1636915332
transform 1 0 5796 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  FILLER_10_85
timestamp 1636915332
transform 1 0 7820 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1636915332
transform 1 0 7728 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_pll_clk OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 9936 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _463_
timestamp 1636915332
transform -1 0 11868 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_8  FILLER_10_129
timestamp 1636915332
transform 1 0 11868 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_137
timestamp 1636915332
transform 1 0 12604 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_144
timestamp 1636915332
transform 1 0 13248 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1636915332
transform 1 0 12880 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _205_
timestamp 1636915332
transform 1 0 12972 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_156
timestamp 1636915332
transform 1 0 14352 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__xor2_1  _377_
timestamp 1636915332
transform 1 0 14536 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__dfrtp_1  _470_
timestamp 1636915332
transform -1 0 17020 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_10_185
timestamp 1636915332
transform 1 0 17020 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_193
timestamp 1636915332
transform 1 0 17756 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1636915332
transform 1 0 18124 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1636915332
transform 1 0 18032 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1636915332
transform -1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1636915332
transform 1 0 18308 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_23
timestamp 1636915332
transform 1 0 2116 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1636915332
transform 1 0 0 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtn_1  _460_
timestamp 1636915332
transform 1 0 276 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_12  FILLER_11_29
timestamp 1636915332
transform 1 0 2668 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_41
timestamp 1636915332
transform 1 0 3772 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_47
timestamp 1636915332
transform 1 0 4324 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__a21bo_1  _229_
timestamp 1636915332
transform -1 0 5152 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _244_
timestamp 1636915332
transform 1 0 2300 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_70
timestamp 1636915332
transform 1 0 6440 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1636915332
transform 1 0 5152 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_1  _228_
timestamp 1636915332
transform 1 0 6072 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _230_
timestamp 1636915332
transform -1 0 6992 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _389_
timestamp 1636915332
transform 1 0 5244 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_11_76
timestamp 1636915332
transform 1 0 6992 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_84
timestamp 1636915332
transform 1 0 7728 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_96
timestamp 1636915332
transform 1 0 8832 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _388_
timestamp 1636915332
transform 1 0 8004 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1636915332
transform 1 0 10304 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_1  _232_
timestamp 1636915332
transform 1 0 9936 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _233_
timestamp 1636915332
transform 1 0 10396 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _379_
timestamp 1636915332
transform 1 0 11132 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_11_130
timestamp 1636915332
transform 1 0 11960 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _469_
timestamp 1636915332
transform 1 0 12236 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_11_164
timestamp 1636915332
transform 1 0 15088 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_169
timestamp 1636915332
transform 1 0 15548 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1636915332
transform 1 0 15456 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__xnor2_1  _373_
timestamp 1636915332
transform 1 0 14076 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _376_
timestamp 1636915332
transform 1 0 14720 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_177
timestamp 1636915332
transform 1 0 16284 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _207_
timestamp 1636915332
transform -1 0 16652 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  _468_
timestamp 1636915332
transform 1 0 16652 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1636915332
transform -1 0 18860 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_11
timestamp 1636915332
transform 1 0 1012 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_3
timestamp 1636915332
transform 1 0 276 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1636915332
transform 1 0 0 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _243_
timestamp 1636915332
transform 1 0 2024 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _245_
timestamp 1636915332
transform -1 0 2024 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_29
timestamp 1636915332
transform 1 0 2668 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_39
timestamp 1636915332
transform 1 0 3588 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_43
timestamp 1636915332
transform 1 0 3956 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1636915332
transform 1 0 2576 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _234_
timestamp 1636915332
transform 1 0 3312 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_1  _236_
timestamp 1636915332
transform 1 0 2760 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__dfrtp_1  _465_
timestamp 1636915332
transform 1 0 4048 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  FILLER_12_64
timestamp 1636915332
transform 1 0 5888 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _231_
timestamp 1636915332
transform -1 0 6900 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_85
timestamp 1636915332
transform 1 0 7820 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_96
timestamp 1636915332
transform 1 0 8832 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1636915332
transform 1 0 7728 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _391_
timestamp 1636915332
transform 1 0 8004 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _392_
timestamp 1636915332
transform 1 0 6900 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_12_102
timestamp 1636915332
transform 1 0 9384 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_106
timestamp 1636915332
transform 1 0 9752 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_114
timestamp 1636915332
transform 1 0 10488 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_1  _226_
timestamp 1636915332
transform -1 0 10488 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _347_
timestamp 1636915332
transform 1 0 9476 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _380_
timestamp 1636915332
transform 1 0 10764 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_12_130
timestamp 1636915332
transform 1 0 11960 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1636915332
transform 1 0 12696 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_141
timestamp 1636915332
transform 1 0 12972 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1636915332
transform 1 0 12880 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _204_
timestamp 1636915332
transform 1 0 13248 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkinv_2  _368_
timestamp 1636915332
transform 1 0 11592 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_153
timestamp 1636915332
transform 1 0 14076 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_171
timestamp 1636915332
transform 1 0 15732 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nor3b_1  _268_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 15180 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _410_
timestamp 1636915332
transform 1 0 14352 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_12_179
timestamp 1636915332
transform 1 0 16468 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1636915332
transform 1 0 17940 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_197
timestamp 1636915332
transform 1 0 18124 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1636915332
transform 1 0 18032 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _206_
timestamp 1636915332
transform 1 0 16744 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkinv_2  _372_
timestamp 1636915332
transform 1 0 17572 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1636915332
transform -1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1636915332
transform 1 0 18308 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_22
timestamp 1636915332
transform 1 0 2024 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1636915332
transform 1 0 276 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_23
timestamp 1636915332
transform 1 0 2116 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1636915332
transform 1 0 0 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1636915332
transform 1 0 0 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2ai_1  _241_
timestamp 1636915332
transform -1 0 2024 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__dfrtn_1  _462_
timestamp 1636915332
transform 1 0 276 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__nand2_1  _240_
timestamp 1636915332
transform 1 0 2300 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _238_
timestamp 1636915332
transform -1 0 2944 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_1  _237_
timestamp 1636915332
transform -1 0 3496 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _235_
timestamp 1636915332
transform -1 0 2852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1636915332
transform 1 0 2576 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_32
timestamp 1636915332
transform 1 0 2944 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1636915332
transform 1 0 2484 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_31
timestamp 1636915332
transform 1 0 2852 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  rebuffer10
timestamp 1636915332
transform 1 0 3864 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _254_
timestamp 1636915332
transform -1 0 3496 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _239_
timestamp 1636915332
transform -1 0 3772 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _216_
timestamp 1636915332
transform 1 0 3588 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_38
timestamp 1636915332
transform 1 0 3496 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_41
timestamp 1636915332
transform 1 0 3772 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o211ai_1  _255_
timestamp 1636915332
transform -1 0 4784 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_45
timestamp 1636915332
transform 1 0 4140 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_49
timestamp 1636915332
transform 1 0 4508 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_70
timestamp 1636915332
transform 1 0 6440 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1636915332
transform 1 0 5152 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_2  _215_
timestamp 1636915332
transform -1 0 6992 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _217_
timestamp 1636915332
transform 1 0 4692 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _224_
timestamp 1636915332
transform 1 0 5704 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _225_
timestamp 1636915332
transform 1 0 6072 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _247_
timestamp 1636915332
transform 1 0 4784 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_4  _390_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer2
timestamp 1636915332
transform 1 0 5060 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _369_
timestamp 1636915332
transform 1 0 7636 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _248_
timestamp 1636915332
transform -1 0 8096 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1636915332
transform 1 0 7728 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1636915332
transform 1 0 7544 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_82
timestamp 1636915332
transform 1 0 7544 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_76
timestamp 1636915332
transform 1 0 6992 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _212_
timestamp 1636915332
transform 1 0 8832 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__fill_2  FILLER_14_88
timestamp 1636915332
transform 1 0 8096 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_90
timestamp 1636915332
transform 1 0 8280 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _419_
timestamp 1636915332
transform -1 0 9752 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__nand3b_1  _223_
timestamp 1636915332
transform 1 0 9476 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _213_
timestamp 1636915332
transform 1 0 9752 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_13_109
timestamp 1636915332
transform 1 0 10028 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_101
timestamp 1636915332
transform 1 0 9292 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_1  _218_
timestamp 1636915332
transform 1 0 10304 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _214_
timestamp 1636915332
transform -1 0 11592 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _210_
timestamp 1636915332
transform -1 0 11224 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1636915332
transform 1 0 10304 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_113
timestamp 1636915332
transform 1 0 10396 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__dfstp_1  _466_
timestamp 1636915332
transform 1 0 10580 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_12  FILLER_13_139
timestamp 1636915332
transform 1 0 12788 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_130
timestamp 1636915332
transform 1 0 11960 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1636915332
transform 1 0 12788 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1636915332
transform 1 0 12880 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _222_
timestamp 1636915332
transform 1 0 12512 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _227_
timestamp 1636915332
transform -1 0 11960 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _353_
timestamp 1636915332
transform 1 0 12144 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2ai_2  _354_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__a21o_1  _271_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 14352 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_14_153
timestamp 1636915332
transform 1 0 14076 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_159
timestamp 1636915332
transform 1 0 14628 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_151
timestamp 1636915332
transform 1 0 13892 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _346_
timestamp 1636915332
transform -1 0 15180 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _272_
timestamp 1636915332
transform 1 0 14904 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _269_
timestamp 1636915332
transform -1 0 15548 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1636915332
transform 1 0 15456 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_169
timestamp 1636915332
transform 1 0 15548 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_165
timestamp 1636915332
transform 1 0 15180 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _436_
timestamp 1636915332
transform 1 0 15916 0 1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _433_
timestamp 1636915332
transform -1 0 17388 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_13_198
timestamp 1636915332
transform 1 0 18216 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_197
timestamp 1636915332
transform 1 0 18124 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1636915332
transform 1 0 18032 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _387_
timestamp 1636915332
transform 1 0 17388 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_14_201
timestamp 1636915332
transform 1 0 18492 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1636915332
transform -1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1636915332
transform -1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_15
timestamp 1636915332
transform 1 0 1380 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_23
timestamp 1636915332
transform 1 0 2116 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1636915332
transform 1 0 276 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1636915332
transform 1 0 0 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _265_
timestamp 1636915332
transform -1 0 2484 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_30
timestamp 1636915332
transform 1 0 2760 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_43
timestamp 1636915332
transform 1 0 3956 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o21bai_1  _256_
timestamp 1636915332
transform -1 0 4876 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _258_
timestamp 1636915332
transform 1 0 3680 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _266_
timestamp 1636915332
transform -1 0 2760 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _384_
timestamp 1636915332
transform 1 0 2852 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_15_53
timestamp 1636915332
transform 1 0 4876 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1636915332
transform 1 0 5152 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_1  _250_
timestamp 1636915332
transform 1 0 5244 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _257_
timestamp 1636915332
transform -1 0 5980 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dfstp_1  _459_
timestamp 1636915332
transform 1 0 6348 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_pll_clk90
timestamp 1636915332
transform -1 0 6348 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_90
timestamp 1636915332
transform 1 0 8280 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_pll_clk90
timestamp 1636915332
transform -1 0 10304 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1636915332
transform 1 0 10304 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _417_
timestamp 1636915332
transform 1 0 10396 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_15_133
timestamp 1636915332
transform 1 0 12236 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_141
timestamp 1636915332
transform 1 0 12972 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _413_
timestamp 1636915332
transform -1 0 14076 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_pll_clk90
timestamp 1636915332
transform 1 0 11868 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_153
timestamp 1636915332
transform 1 0 14076 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_159
timestamp 1636915332
transform 1 0 14628 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_164
timestamp 1636915332
transform 1 0 15088 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1636915332
transform 1 0 15548 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1636915332
transform 1 0 15456 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _270_
timestamp 1636915332
transform 1 0 14812 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _273_
timestamp 1636915332
transform -1 0 14628 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  _434_
timestamp 1636915332
transform -1 0 17664 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_6  FILLER_15_192
timestamp 1636915332
transform 1 0 17664 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_198
timestamp 1636915332
transform 1 0 18216 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1636915332
transform -1 0 18860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1636915332
transform 1 0 18308 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1636915332
transform 1 0 0 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _267_
timestamp 1636915332
transform -1 0 2484 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtn_1  _456_
timestamp 1636915332
transform 1 0 276 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1636915332
transform 1 0 2484 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1636915332
transform 1 0 2668 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1636915332
transform 1 0 2576 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _259_
timestamp 1636915332
transform 1 0 2852 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _383_
timestamp 1636915332
transform 1 0 3772 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_16_50
timestamp 1636915332
transform 1 0 4600 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_58
timestamp 1636915332
transform 1 0 5336 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_69
timestamp 1636915332
transform 1 0 6348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_73
timestamp 1636915332
transform 1 0 6716 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _246__2
timestamp 1636915332
transform -1 0 6716 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _409_
timestamp 1636915332
transform 1 0 5520 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_16_81
timestamp 1636915332
transform 1 0 7452 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1636915332
transform 1 0 7728 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _418_
timestamp 1636915332
transform 1 0 7820 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_16_101
timestamp 1636915332
transform 1 0 9292 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__or2b_1  _208_
timestamp 1636915332
transform 1 0 9384 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _412_
timestamp 1636915332
transform -1 0 10764 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__dfrtp_4  _467_
timestamp 1636915332
transform -1 0 12880 0 1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_4  FILLER_16_141
timestamp 1636915332
transform 1 0 12972 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_148
timestamp 1636915332
transform 1 0 13616 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1636915332
transform 1 0 12880 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _352_
timestamp 1636915332
transform -1 0 13616 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_4  _437_
timestamp 1636915332
transform 1 0 15824 0 1 8704
box -38 -48 2246 592
use sky130_fd_sc_hd__dfstp_1  _455_
timestamp 1636915332
transform -1 0 15824 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1636915332
transform 1 0 18032 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  split1
timestamp 1636915332
transform 1 0 18124 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_201
timestamp 1636915332
transform 1 0 18492 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1636915332
transform -1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_11
timestamp 1636915332
transform 1 0 1012 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_16
timestamp 1636915332
transform 1 0 1472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_20
timestamp 1636915332
transform 1 0 1840 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_3
timestamp 1636915332
transform 1 0 276 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1636915332
transform 1 0 0 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _260_
timestamp 1636915332
transform -1 0 1840 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _261_
timestamp 1636915332
transform -1 0 1472 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_35
timestamp 1636915332
transform 1 0 3220 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _263_
timestamp 1636915332
transform -1 0 3220 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _396_
timestamp 1636915332
transform 1 0 4324 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_17_57
timestamp 1636915332
transform 1 0 5244 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1636915332
transform 1 0 5152 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _395_
timestamp 1636915332
transform 1 0 5520 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _408_
timestamp 1636915332
transform 1 0 6348 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_17_78
timestamp 1636915332
transform 1 0 7176 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_90
timestamp 1636915332
transform 1 0 8280 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_1  _426_
timestamp 1636915332
transform -1 0 10304 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_17_113
timestamp 1636915332
transform 1 0 10396 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1636915332
transform 1 0 10304 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _425_
timestamp 1636915332
transform 1 0 10580 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  _393_
timestamp 1636915332
transform 1 0 12420 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__dfrtp_4  _438_
timestamp 1636915332
transform -1 0 15364 0 -1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1636915332
transform 1 0 15364 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_169
timestamp 1636915332
transform 1 0 15548 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1636915332
transform 1 0 15456 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_175
timestamp 1636915332
transform 1 0 16100 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_196
timestamp 1636915332
transform 1 0 18032 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__dfrtp_1  _435_
timestamp 1636915332
transform -1 0 18032 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1636915332
transform -1 0 18860 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1636915332
transform 1 0 0 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _251_
timestamp 1636915332
transform -1 0 2392 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtn_1  _458_
timestamp 1636915332
transform 1 0 276 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_18_26
timestamp 1636915332
transform 1 0 2392 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_43
timestamp 1636915332
transform 1 0 3956 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1636915332
transform 1 0 2576 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__nor3b_2  _249_
timestamp 1636915332
transform -1 0 5152 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _252_
timestamp 1636915332
transform -1 0 3956 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _253_
timestamp 1636915332
transform -1 0 3036 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _262__3
timestamp 1636915332
transform -1 0 3680 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _264_
timestamp 1636915332
transform -1 0 3404 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_56
timestamp 1636915332
transform 1 0 5152 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_68
timestamp 1636915332
transform 1 0 6256 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__xnor2_1  _365_
timestamp 1636915332
transform 1 0 5336 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _366_
timestamp 1636915332
transform 1 0 5980 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_80
timestamp 1636915332
transform 1 0 7360 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_94
timestamp 1636915332
transform 1 0 8648 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1636915332
transform 1 0 7728 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _211_
timestamp 1636915332
transform -1 0 9200 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _343_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 7820 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_18_100
timestamp 1636915332
transform 1 0 9200 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_124
timestamp 1636915332
transform 1 0 11408 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_ext_clk
timestamp 1636915332
transform 1 0 9568 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_18_128
timestamp 1636915332
transform 1 0 11776 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1636915332
transform 1 0 12236 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1636915332
transform 1 0 12788 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_145
timestamp 1636915332
transform 1 0 13340 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1636915332
transform 1 0 12880 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _378__13 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 13892 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_ext_clk
timestamp 1636915332
transform -1 0 12236 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 1636915332
transform -1 0 13340 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_151
timestamp 1636915332
transform 1 0 13892 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_159
timestamp 1636915332
transform 1 0 14628 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__dfstp_1  _422_
timestamp 1636915332
transform 1 0 14812 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_8  FILLER_18_182
timestamp 1636915332
transform 1 0 16744 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_190
timestamp 1636915332
transform 1 0 17480 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1636915332
transform 1 0 18124 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1636915332
transform 1 0 18032 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1636915332
transform 1 0 17756 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1636915332
transform -1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1636915332
transform 1 0 18308 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_11
timestamp 1636915332
transform 1 0 1012 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_3
timestamp 1636915332
transform 1 0 276 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1636915332
transform 1 0 0 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  input3 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 1104 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1636915332
transform 1 0 2576 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_1  _457_
timestamp 1636915332
transform 1 0 2668 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_6  FILLER_19_50
timestamp 1636915332
transform 1 0 4600 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_19_64
timestamp 1636915332
transform 1 0 5888 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_72
timestamp 1636915332
transform 1 0 6624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1636915332
transform 1 0 5152 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__xor2_1  _367_
timestamp 1636915332
transform 1 0 5244 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  output10
timestamp 1636915332
transform -1 0 6992 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_83
timestamp 1636915332
transform 1 0 7636 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1636915332
transform 1 0 7728 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _344_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 6992 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _420_
timestamp 1636915332
transform 1 0 7820 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_ext_clk
timestamp 1636915332
transform 1 0 7268 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_109
timestamp 1636915332
transform 1 0 10028 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_19_122
timestamp 1636915332
transform 1 0 11224 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1636915332
transform 1 0 10304 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__or2b_1  _209_
timestamp 1636915332
transform 1 0 10396 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold1 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 9292 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  output12
timestamp 1636915332
transform 1 0 10948 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_128
timestamp 1636915332
transform 1 0 11776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_138
timestamp 1636915332
transform 1 0 12696 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_141
timestamp 1636915332
transform 1 0 12972 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1636915332
transform 1 0 12880 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _394_
timestamp 1636915332
transform 1 0 11868 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__dfstp_1  _423_
timestamp 1636915332
transform 1 0 13248 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  FILLER_19_165
timestamp 1636915332
transform 1 0 15180 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_19_169
timestamp 1636915332
transform 1 0 15548 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1636915332
transform 1 0 15456 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1636915332
transform 1 0 18032 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _375_
timestamp 1636915332
transform 1 0 18124 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  _421_
timestamp 1636915332
transform 1 0 16100 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_2  FILLER_19_200
timestamp 1636915332
transform 1 0 18400 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1636915332
transform -1 0 18860 0 -1 10880
box -38 -48 314 592
<< labels >>
rlabel metal5 s 0 4812 18860 5132 6 VGND
port 0 nsew ground input
rlabel metal5 s 0 8192 18860 8512 6 VGND
port 0 nsew ground input
rlabel metal4 s 4654 -48 4974 10928 6 VGND
port 0 nsew ground input
rlabel metal4 s 7754 -48 8074 10928 6 VGND
port 0 nsew ground input
rlabel metal4 s 10854 -48 11174 10928 6 VGND
port 0 nsew ground input
rlabel metal4 s 13954 -48 14274 10928 6 VGND
port 0 nsew ground input
rlabel metal4 s 17054 -48 17374 10928 6 VGND
port 0 nsew ground input
rlabel metal5 s 0 3122 18860 3442 6 VPWR
port 1 nsew power input
rlabel metal5 s 0 6502 18860 6822 6 VPWR
port 1 nsew power input
rlabel metal5 s 0 9882 18860 10202 6 VPWR
port 1 nsew power input
rlabel metal4 s 3104 -48 3424 10928 6 VPWR
port 1 nsew power input
rlabel metal4 s 6204 -48 6524 10928 6 VPWR
port 1 nsew power input
rlabel metal4 s 9304 -48 9624 10928 6 VPWR
port 1 nsew power input
rlabel metal4 s 12404 -48 12724 10928 6 VPWR
port 1 nsew power input
rlabel metal4 s 15504 -48 15824 10928 6 VPWR
port 1 nsew power input
rlabel metal2 s 7102 11200 7158 12000 6 core_clk
port 2 nsew signal tristate
rlabel metal2 s 4250 11200 4306 12000 6 ext_clk
port 3 nsew signal input
rlabel metal3 s 19200 688 20000 808 6 ext_clk_sel
port 4 nsew signal input
rlabel metal3 s 19200 11160 20000 11280 6 ext_reset
port 5 nsew signal input
rlabel metal2 s 15658 11200 15714 12000 6 pll_clk
port 6 nsew signal input
rlabel metal2 s 18510 11200 18566 12000 6 pll_clk90
port 7 nsew signal input
rlabel metal2 s 1398 11200 1454 12000 6 resetb
port 8 nsew signal input
rlabel metal2 s 12806 11200 12862 12000 6 resetb_sync
port 9 nsew signal tristate
rlabel metal3 s 19200 6672 20000 6792 6 sel2[0]
port 10 nsew signal input
rlabel metal3 s 19200 8168 20000 8288 6 sel2[1]
port 11 nsew signal input
rlabel metal3 s 19200 9664 20000 9784 6 sel2[2]
port 12 nsew signal input
rlabel metal3 s 19200 2184 20000 2304 6 sel[0]
port 13 nsew signal input
rlabel metal3 s 19200 3680 20000 3800 6 sel[1]
port 14 nsew signal input
rlabel metal3 s 19200 5176 20000 5296 6 sel[2]
port 15 nsew signal input
rlabel metal2 s 9954 11200 10010 12000 6 user_clk
port 16 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 20000 12000
<< end >>
