VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ./mag/caravel_power_routing
  CLASS BLOCK ;
  FOREIGN ./mag/caravel_power_routing ;
  ORIGIN 0.000 0.000 ;
  SIZE 3588.000 BY 5188.000 ;
  PIN vccd_core
    PORT
      LAYER met3 ;
        RECT 197.280 390.755 229.220 413.720 ;
        RECT 197.280 341.280 229.220 364.500 ;
      LAYER via3 ;
        RECT 209.885 391.210 228.205 413.530 ;
        RECT 209.765 341.690 228.085 364.010 ;
      LAYER met4 ;
        RECT 220.930 1152.330 315.800 1167.330 ;
        RECT 448.500 1152.330 450.780 1170.320 ;
        RECT 468.500 1152.330 470.780 1170.320 ;
        RECT 548.500 1152.330 550.780 1170.320 ;
        RECT 568.500 1152.330 570.780 1170.320 ;
        RECT 665.300 1152.330 667.580 1167.320 ;
        RECT 740.550 1152.330 742.830 1167.320 ;
        RECT 815.800 1152.330 818.080 1167.320 ;
        RECT 891.050 1152.330 893.330 1167.320 ;
        RECT 966.300 1152.330 968.580 1167.320 ;
        RECT 1041.550 1152.330 1043.830 1167.320 ;
        RECT 1116.800 1152.330 1119.080 1167.320 ;
        RECT 1192.050 1152.330 1194.330 1167.320 ;
        RECT 1267.300 1152.330 1269.580 1167.320 ;
        RECT 1342.550 1152.330 1344.830 1167.320 ;
        RECT 1417.800 1152.330 1420.080 1167.320 ;
        RECT 1493.050 1152.330 1495.330 1167.320 ;
        RECT 1568.300 1152.330 1570.580 1167.320 ;
        RECT 1643.550 1152.330 1645.830 1167.320 ;
        RECT 1718.800 1152.330 1721.080 1167.320 ;
        RECT 1794.050 1152.330 1796.330 1167.320 ;
        RECT 1869.300 1152.330 1871.580 1167.320 ;
        RECT 1944.550 1152.330 1946.830 1167.320 ;
        RECT 2019.800 1152.330 2022.080 1167.320 ;
        RECT 2095.050 1152.330 2097.330 1167.320 ;
        RECT 2170.300 1152.330 2172.580 1167.320 ;
        RECT 2245.550 1152.330 2247.830 1167.320 ;
        RECT 2320.800 1152.330 2323.080 1167.320 ;
        RECT 2396.050 1152.330 2398.330 1167.320 ;
        RECT 2471.300 1152.330 2473.580 1167.320 ;
        RECT 2546.550 1152.330 2548.830 1167.320 ;
        RECT 2621.800 1152.330 2624.080 1167.320 ;
        RECT 2696.800 1152.330 2699.080 1167.320 ;
        RECT 2898.600 1152.330 2900.880 1170.320 ;
        RECT 2918.600 1152.330 2920.880 1170.320 ;
        RECT 220.990 1046.990 233.990 1152.330 ;
        RECT 2921.840 1047.520 2984.810 1062.520 ;
        RECT 3135.220 1047.640 3140.540 1062.300 ;
        RECT 3212.020 1047.640 3217.340 1062.300 ;
        RECT 3288.820 1047.640 3294.140 1062.300 ;
        RECT 220.990 1043.790 257.600 1046.990 ;
        RECT 220.990 996.990 233.990 1043.790 ;
        RECT 2983.210 1038.460 2984.810 1047.520 ;
        RECT 3136.810 1038.420 3138.410 1047.640 ;
        RECT 3213.610 1038.420 3215.210 1047.640 ;
        RECT 3290.410 1038.420 3292.010 1047.640 ;
        RECT 2922.480 997.300 2935.870 999.040 ;
        RECT 220.990 993.790 257.600 996.990 ;
        RECT 2922.480 995.700 2964.880 997.300 ;
        RECT 2922.480 994.620 2935.870 995.700 ;
        RECT 220.990 946.990 233.990 993.790 ;
        RECT 220.990 943.790 257.600 946.990 ;
        RECT 220.990 896.990 233.990 943.790 ;
        RECT 2922.480 919.100 2935.870 920.840 ;
        RECT 2922.480 917.500 2964.880 919.100 ;
        RECT 2922.480 916.420 2935.870 917.500 ;
        RECT 220.990 893.790 257.600 896.990 ;
        RECT 220.990 883.710 233.990 893.790 ;
        RECT 209.320 865.630 233.990 883.710 ;
        RECT 208.840 843.790 257.600 846.990 ;
        RECT 2922.480 840.900 2935.870 842.640 ;
        RECT 2922.480 839.300 2964.880 840.900 ;
        RECT 2922.480 838.220 2935.870 839.300 ;
        RECT 208.840 793.790 257.600 796.990 ;
        RECT 2922.480 762.700 2935.870 764.440 ;
        RECT 2922.480 761.100 2964.880 762.700 ;
        RECT 2922.480 760.020 2935.870 761.100 ;
        RECT 208.840 743.790 257.600 746.990 ;
        RECT 208.840 693.790 257.600 696.990 ;
        RECT 2922.480 684.500 2935.870 686.240 ;
        RECT 2922.480 682.900 2964.880 684.500 ;
        RECT 2922.480 681.820 2935.870 682.900 ;
        RECT 208.840 643.790 257.600 646.990 ;
        RECT 2922.480 600.300 2935.870 602.040 ;
        RECT 2959.660 600.300 2965.060 606.530 ;
        RECT 2922.480 598.700 2965.060 600.300 ;
        RECT 2922.480 597.620 2935.870 598.700 ;
        RECT 208.840 593.790 257.600 596.990 ;
        RECT 208.840 543.790 257.600 546.990 ;
        RECT 2922.480 528.100 2935.870 529.840 ;
        RECT 2922.480 526.500 2964.880 528.100 ;
        RECT 2922.480 525.420 2935.870 526.500 ;
        RECT 208.840 493.790 257.600 496.990 ;
        RECT 208.840 443.790 257.600 446.990 ;
        RECT 209.320 396.990 228.890 413.970 ;
        RECT 3161.770 404.620 3163.370 410.310 ;
        RECT 3201.770 405.080 3203.370 410.000 ;
        RECT 208.840 393.790 257.600 396.990 ;
        RECT 209.320 390.770 228.890 393.790 ;
        RECT 3160.360 390.990 3165.050 404.620 ;
        RECT 3200.490 390.670 3204.610 405.080 ;
        RECT 3141.590 369.140 3143.190 386.870 ;
        RECT 3157.090 369.140 3158.690 386.870 ;
        RECT 3172.590 369.140 3174.190 386.870 ;
        RECT 3188.090 369.140 3189.690 386.870 ;
        RECT 3203.590 369.140 3205.190 386.870 ;
        RECT 3219.090 369.140 3220.690 386.870 ;
        RECT 209.290 346.990 228.860 364.450 ;
        RECT 208.840 343.790 257.600 346.990 ;
        RECT 209.290 341.250 228.860 343.790 ;
        RECT 208.840 293.790 257.600 296.990 ;
        RECT 3141.570 262.550 3143.170 278.900 ;
        RECT 3157.070 262.550 3158.670 278.900 ;
        RECT 3172.570 262.550 3174.170 278.900 ;
        RECT 3188.070 262.550 3189.670 278.900 ;
        RECT 3203.570 262.550 3205.170 278.900 ;
        RECT 3219.070 262.550 3220.670 278.900 ;
        RECT 209.370 241.110 292.680 260.610 ;
        RECT 716.620 249.680 723.690 253.440 ;
        RECT 719.300 248.190 720.200 249.680 ;
        RECT 3306.350 234.955 3347.130 236.600 ;
      LAYER via4 ;
        RECT 282.770 1153.675 314.350 1166.055 ;
        RECT 448.900 1165.630 450.080 1166.810 ;
        RECT 448.900 1164.030 450.080 1165.210 ;
        RECT 448.900 1162.430 450.080 1163.610 ;
        RECT 448.900 1160.830 450.080 1162.010 ;
        RECT 448.900 1159.230 450.080 1160.410 ;
        RECT 448.900 1157.630 450.080 1158.810 ;
        RECT 448.900 1156.030 450.080 1157.210 ;
        RECT 448.900 1154.430 450.080 1155.610 ;
        RECT 448.900 1152.830 450.080 1154.010 ;
        RECT 468.900 1165.630 470.080 1166.810 ;
        RECT 468.900 1164.030 470.080 1165.210 ;
        RECT 468.900 1162.430 470.080 1163.610 ;
        RECT 468.900 1160.830 470.080 1162.010 ;
        RECT 468.900 1159.230 470.080 1160.410 ;
        RECT 468.900 1157.630 470.080 1158.810 ;
        RECT 468.900 1156.030 470.080 1157.210 ;
        RECT 468.900 1154.430 470.080 1155.610 ;
        RECT 468.900 1152.830 470.080 1154.010 ;
        RECT 548.900 1165.630 550.080 1166.810 ;
        RECT 548.900 1164.030 550.080 1165.210 ;
        RECT 548.900 1162.430 550.080 1163.610 ;
        RECT 548.900 1160.830 550.080 1162.010 ;
        RECT 548.900 1159.230 550.080 1160.410 ;
        RECT 548.900 1157.630 550.080 1158.810 ;
        RECT 548.900 1156.030 550.080 1157.210 ;
        RECT 548.900 1154.430 550.080 1155.610 ;
        RECT 548.900 1152.830 550.080 1154.010 ;
        RECT 568.900 1165.630 570.080 1166.810 ;
        RECT 568.900 1164.030 570.080 1165.210 ;
        RECT 568.900 1162.430 570.080 1163.610 ;
        RECT 568.900 1160.830 570.080 1162.010 ;
        RECT 568.900 1159.230 570.080 1160.410 ;
        RECT 568.900 1157.630 570.080 1158.810 ;
        RECT 568.900 1156.030 570.080 1157.210 ;
        RECT 568.900 1154.430 570.080 1155.610 ;
        RECT 568.900 1152.830 570.080 1154.010 ;
        RECT 665.700 1165.630 666.880 1166.810 ;
        RECT 665.700 1164.030 666.880 1165.210 ;
        RECT 665.700 1162.430 666.880 1163.610 ;
        RECT 665.700 1160.830 666.880 1162.010 ;
        RECT 665.700 1159.230 666.880 1160.410 ;
        RECT 665.700 1157.630 666.880 1158.810 ;
        RECT 665.700 1156.030 666.880 1157.210 ;
        RECT 665.700 1154.430 666.880 1155.610 ;
        RECT 665.700 1152.830 666.880 1154.010 ;
        RECT 740.950 1165.630 742.130 1166.810 ;
        RECT 740.950 1164.030 742.130 1165.210 ;
        RECT 740.950 1162.430 742.130 1163.610 ;
        RECT 740.950 1160.830 742.130 1162.010 ;
        RECT 740.950 1159.230 742.130 1160.410 ;
        RECT 740.950 1157.630 742.130 1158.810 ;
        RECT 740.950 1156.030 742.130 1157.210 ;
        RECT 740.950 1154.430 742.130 1155.610 ;
        RECT 740.950 1152.830 742.130 1154.010 ;
        RECT 816.200 1165.630 817.380 1166.810 ;
        RECT 816.200 1164.030 817.380 1165.210 ;
        RECT 816.200 1162.430 817.380 1163.610 ;
        RECT 816.200 1160.830 817.380 1162.010 ;
        RECT 816.200 1159.230 817.380 1160.410 ;
        RECT 816.200 1157.630 817.380 1158.810 ;
        RECT 816.200 1156.030 817.380 1157.210 ;
        RECT 816.200 1154.430 817.380 1155.610 ;
        RECT 816.200 1152.830 817.380 1154.010 ;
        RECT 891.450 1165.630 892.630 1166.810 ;
        RECT 891.450 1164.030 892.630 1165.210 ;
        RECT 891.450 1162.430 892.630 1163.610 ;
        RECT 891.450 1160.830 892.630 1162.010 ;
        RECT 891.450 1159.230 892.630 1160.410 ;
        RECT 891.450 1157.630 892.630 1158.810 ;
        RECT 891.450 1156.030 892.630 1157.210 ;
        RECT 891.450 1154.430 892.630 1155.610 ;
        RECT 891.450 1152.830 892.630 1154.010 ;
        RECT 966.700 1165.630 967.880 1166.810 ;
        RECT 966.700 1164.030 967.880 1165.210 ;
        RECT 966.700 1162.430 967.880 1163.610 ;
        RECT 966.700 1160.830 967.880 1162.010 ;
        RECT 966.700 1159.230 967.880 1160.410 ;
        RECT 966.700 1157.630 967.880 1158.810 ;
        RECT 966.700 1156.030 967.880 1157.210 ;
        RECT 966.700 1154.430 967.880 1155.610 ;
        RECT 966.700 1152.830 967.880 1154.010 ;
        RECT 1041.950 1165.630 1043.130 1166.810 ;
        RECT 1041.950 1164.030 1043.130 1165.210 ;
        RECT 1041.950 1162.430 1043.130 1163.610 ;
        RECT 1041.950 1160.830 1043.130 1162.010 ;
        RECT 1041.950 1159.230 1043.130 1160.410 ;
        RECT 1041.950 1157.630 1043.130 1158.810 ;
        RECT 1041.950 1156.030 1043.130 1157.210 ;
        RECT 1041.950 1154.430 1043.130 1155.610 ;
        RECT 1041.950 1152.830 1043.130 1154.010 ;
        RECT 1117.200 1165.630 1118.380 1166.810 ;
        RECT 1117.200 1164.030 1118.380 1165.210 ;
        RECT 1117.200 1162.430 1118.380 1163.610 ;
        RECT 1117.200 1160.830 1118.380 1162.010 ;
        RECT 1117.200 1159.230 1118.380 1160.410 ;
        RECT 1117.200 1157.630 1118.380 1158.810 ;
        RECT 1117.200 1156.030 1118.380 1157.210 ;
        RECT 1117.200 1154.430 1118.380 1155.610 ;
        RECT 1117.200 1152.830 1118.380 1154.010 ;
        RECT 1192.450 1165.630 1193.630 1166.810 ;
        RECT 1192.450 1164.030 1193.630 1165.210 ;
        RECT 1192.450 1162.430 1193.630 1163.610 ;
        RECT 1192.450 1160.830 1193.630 1162.010 ;
        RECT 1192.450 1159.230 1193.630 1160.410 ;
        RECT 1192.450 1157.630 1193.630 1158.810 ;
        RECT 1192.450 1156.030 1193.630 1157.210 ;
        RECT 1192.450 1154.430 1193.630 1155.610 ;
        RECT 1192.450 1152.830 1193.630 1154.010 ;
        RECT 1267.700 1165.630 1268.880 1166.810 ;
        RECT 1267.700 1164.030 1268.880 1165.210 ;
        RECT 1267.700 1162.430 1268.880 1163.610 ;
        RECT 1267.700 1160.830 1268.880 1162.010 ;
        RECT 1267.700 1159.230 1268.880 1160.410 ;
        RECT 1267.700 1157.630 1268.880 1158.810 ;
        RECT 1267.700 1156.030 1268.880 1157.210 ;
        RECT 1267.700 1154.430 1268.880 1155.610 ;
        RECT 1267.700 1152.830 1268.880 1154.010 ;
        RECT 1342.950 1165.630 1344.130 1166.810 ;
        RECT 1342.950 1164.030 1344.130 1165.210 ;
        RECT 1342.950 1162.430 1344.130 1163.610 ;
        RECT 1342.950 1160.830 1344.130 1162.010 ;
        RECT 1342.950 1159.230 1344.130 1160.410 ;
        RECT 1342.950 1157.630 1344.130 1158.810 ;
        RECT 1342.950 1156.030 1344.130 1157.210 ;
        RECT 1342.950 1154.430 1344.130 1155.610 ;
        RECT 1342.950 1152.830 1344.130 1154.010 ;
        RECT 1418.200 1165.630 1419.380 1166.810 ;
        RECT 1418.200 1164.030 1419.380 1165.210 ;
        RECT 1418.200 1162.430 1419.380 1163.610 ;
        RECT 1418.200 1160.830 1419.380 1162.010 ;
        RECT 1418.200 1159.230 1419.380 1160.410 ;
        RECT 1418.200 1157.630 1419.380 1158.810 ;
        RECT 1418.200 1156.030 1419.380 1157.210 ;
        RECT 1418.200 1154.430 1419.380 1155.610 ;
        RECT 1418.200 1152.830 1419.380 1154.010 ;
        RECT 1493.450 1165.630 1494.630 1166.810 ;
        RECT 1493.450 1164.030 1494.630 1165.210 ;
        RECT 1493.450 1162.430 1494.630 1163.610 ;
        RECT 1493.450 1160.830 1494.630 1162.010 ;
        RECT 1493.450 1159.230 1494.630 1160.410 ;
        RECT 1493.450 1157.630 1494.630 1158.810 ;
        RECT 1493.450 1156.030 1494.630 1157.210 ;
        RECT 1493.450 1154.430 1494.630 1155.610 ;
        RECT 1493.450 1152.830 1494.630 1154.010 ;
        RECT 1568.700 1165.630 1569.880 1166.810 ;
        RECT 1568.700 1164.030 1569.880 1165.210 ;
        RECT 1568.700 1162.430 1569.880 1163.610 ;
        RECT 1568.700 1160.830 1569.880 1162.010 ;
        RECT 1568.700 1159.230 1569.880 1160.410 ;
        RECT 1568.700 1157.630 1569.880 1158.810 ;
        RECT 1568.700 1156.030 1569.880 1157.210 ;
        RECT 1568.700 1154.430 1569.880 1155.610 ;
        RECT 1568.700 1152.830 1569.880 1154.010 ;
        RECT 1643.950 1165.630 1645.130 1166.810 ;
        RECT 1643.950 1164.030 1645.130 1165.210 ;
        RECT 1643.950 1162.430 1645.130 1163.610 ;
        RECT 1643.950 1160.830 1645.130 1162.010 ;
        RECT 1643.950 1159.230 1645.130 1160.410 ;
        RECT 1643.950 1157.630 1645.130 1158.810 ;
        RECT 1643.950 1156.030 1645.130 1157.210 ;
        RECT 1643.950 1154.430 1645.130 1155.610 ;
        RECT 1643.950 1152.830 1645.130 1154.010 ;
        RECT 1719.200 1165.630 1720.380 1166.810 ;
        RECT 1719.200 1164.030 1720.380 1165.210 ;
        RECT 1719.200 1162.430 1720.380 1163.610 ;
        RECT 1719.200 1160.830 1720.380 1162.010 ;
        RECT 1719.200 1159.230 1720.380 1160.410 ;
        RECT 1719.200 1157.630 1720.380 1158.810 ;
        RECT 1719.200 1156.030 1720.380 1157.210 ;
        RECT 1719.200 1154.430 1720.380 1155.610 ;
        RECT 1719.200 1152.830 1720.380 1154.010 ;
        RECT 1794.450 1165.630 1795.630 1166.810 ;
        RECT 1794.450 1164.030 1795.630 1165.210 ;
        RECT 1794.450 1162.430 1795.630 1163.610 ;
        RECT 1794.450 1160.830 1795.630 1162.010 ;
        RECT 1794.450 1159.230 1795.630 1160.410 ;
        RECT 1794.450 1157.630 1795.630 1158.810 ;
        RECT 1794.450 1156.030 1795.630 1157.210 ;
        RECT 1794.450 1154.430 1795.630 1155.610 ;
        RECT 1794.450 1152.830 1795.630 1154.010 ;
        RECT 1869.700 1165.630 1870.880 1166.810 ;
        RECT 1869.700 1164.030 1870.880 1165.210 ;
        RECT 1869.700 1162.430 1870.880 1163.610 ;
        RECT 1869.700 1160.830 1870.880 1162.010 ;
        RECT 1869.700 1159.230 1870.880 1160.410 ;
        RECT 1869.700 1157.630 1870.880 1158.810 ;
        RECT 1869.700 1156.030 1870.880 1157.210 ;
        RECT 1869.700 1154.430 1870.880 1155.610 ;
        RECT 1869.700 1152.830 1870.880 1154.010 ;
        RECT 1944.950 1165.630 1946.130 1166.810 ;
        RECT 1944.950 1164.030 1946.130 1165.210 ;
        RECT 1944.950 1162.430 1946.130 1163.610 ;
        RECT 1944.950 1160.830 1946.130 1162.010 ;
        RECT 1944.950 1159.230 1946.130 1160.410 ;
        RECT 1944.950 1157.630 1946.130 1158.810 ;
        RECT 1944.950 1156.030 1946.130 1157.210 ;
        RECT 1944.950 1154.430 1946.130 1155.610 ;
        RECT 1944.950 1152.830 1946.130 1154.010 ;
        RECT 2020.200 1165.630 2021.380 1166.810 ;
        RECT 2020.200 1164.030 2021.380 1165.210 ;
        RECT 2020.200 1162.430 2021.380 1163.610 ;
        RECT 2020.200 1160.830 2021.380 1162.010 ;
        RECT 2020.200 1159.230 2021.380 1160.410 ;
        RECT 2020.200 1157.630 2021.380 1158.810 ;
        RECT 2020.200 1156.030 2021.380 1157.210 ;
        RECT 2020.200 1154.430 2021.380 1155.610 ;
        RECT 2020.200 1152.830 2021.380 1154.010 ;
        RECT 2095.450 1165.630 2096.630 1166.810 ;
        RECT 2095.450 1164.030 2096.630 1165.210 ;
        RECT 2095.450 1162.430 2096.630 1163.610 ;
        RECT 2095.450 1160.830 2096.630 1162.010 ;
        RECT 2095.450 1159.230 2096.630 1160.410 ;
        RECT 2095.450 1157.630 2096.630 1158.810 ;
        RECT 2095.450 1156.030 2096.630 1157.210 ;
        RECT 2095.450 1154.430 2096.630 1155.610 ;
        RECT 2095.450 1152.830 2096.630 1154.010 ;
        RECT 2170.700 1165.630 2171.880 1166.810 ;
        RECT 2170.700 1164.030 2171.880 1165.210 ;
        RECT 2170.700 1162.430 2171.880 1163.610 ;
        RECT 2170.700 1160.830 2171.880 1162.010 ;
        RECT 2170.700 1159.230 2171.880 1160.410 ;
        RECT 2170.700 1157.630 2171.880 1158.810 ;
        RECT 2170.700 1156.030 2171.880 1157.210 ;
        RECT 2170.700 1154.430 2171.880 1155.610 ;
        RECT 2170.700 1152.830 2171.880 1154.010 ;
        RECT 2245.950 1165.630 2247.130 1166.810 ;
        RECT 2245.950 1164.030 2247.130 1165.210 ;
        RECT 2245.950 1162.430 2247.130 1163.610 ;
        RECT 2245.950 1160.830 2247.130 1162.010 ;
        RECT 2245.950 1159.230 2247.130 1160.410 ;
        RECT 2245.950 1157.630 2247.130 1158.810 ;
        RECT 2245.950 1156.030 2247.130 1157.210 ;
        RECT 2245.950 1154.430 2247.130 1155.610 ;
        RECT 2245.950 1152.830 2247.130 1154.010 ;
        RECT 2321.200 1165.630 2322.380 1166.810 ;
        RECT 2321.200 1164.030 2322.380 1165.210 ;
        RECT 2321.200 1162.430 2322.380 1163.610 ;
        RECT 2321.200 1160.830 2322.380 1162.010 ;
        RECT 2321.200 1159.230 2322.380 1160.410 ;
        RECT 2321.200 1157.630 2322.380 1158.810 ;
        RECT 2321.200 1156.030 2322.380 1157.210 ;
        RECT 2321.200 1154.430 2322.380 1155.610 ;
        RECT 2321.200 1152.830 2322.380 1154.010 ;
        RECT 2396.450 1165.630 2397.630 1166.810 ;
        RECT 2396.450 1164.030 2397.630 1165.210 ;
        RECT 2396.450 1162.430 2397.630 1163.610 ;
        RECT 2396.450 1160.830 2397.630 1162.010 ;
        RECT 2396.450 1159.230 2397.630 1160.410 ;
        RECT 2396.450 1157.630 2397.630 1158.810 ;
        RECT 2396.450 1156.030 2397.630 1157.210 ;
        RECT 2396.450 1154.430 2397.630 1155.610 ;
        RECT 2396.450 1152.830 2397.630 1154.010 ;
        RECT 2471.700 1165.630 2472.880 1166.810 ;
        RECT 2471.700 1164.030 2472.880 1165.210 ;
        RECT 2471.700 1162.430 2472.880 1163.610 ;
        RECT 2471.700 1160.830 2472.880 1162.010 ;
        RECT 2471.700 1159.230 2472.880 1160.410 ;
        RECT 2471.700 1157.630 2472.880 1158.810 ;
        RECT 2471.700 1156.030 2472.880 1157.210 ;
        RECT 2471.700 1154.430 2472.880 1155.610 ;
        RECT 2471.700 1152.830 2472.880 1154.010 ;
        RECT 2546.950 1165.630 2548.130 1166.810 ;
        RECT 2546.950 1164.030 2548.130 1165.210 ;
        RECT 2546.950 1162.430 2548.130 1163.610 ;
        RECT 2546.950 1160.830 2548.130 1162.010 ;
        RECT 2546.950 1159.230 2548.130 1160.410 ;
        RECT 2546.950 1157.630 2548.130 1158.810 ;
        RECT 2546.950 1156.030 2548.130 1157.210 ;
        RECT 2546.950 1154.430 2548.130 1155.610 ;
        RECT 2546.950 1152.830 2548.130 1154.010 ;
        RECT 2622.200 1165.630 2623.380 1166.810 ;
        RECT 2622.200 1164.030 2623.380 1165.210 ;
        RECT 2622.200 1162.430 2623.380 1163.610 ;
        RECT 2622.200 1160.830 2623.380 1162.010 ;
        RECT 2622.200 1159.230 2623.380 1160.410 ;
        RECT 2622.200 1157.630 2623.380 1158.810 ;
        RECT 2622.200 1156.030 2623.380 1157.210 ;
        RECT 2622.200 1154.430 2623.380 1155.610 ;
        RECT 2622.200 1152.830 2623.380 1154.010 ;
        RECT 2697.200 1165.630 2698.380 1166.810 ;
        RECT 2697.200 1164.030 2698.380 1165.210 ;
        RECT 2697.200 1162.430 2698.380 1163.610 ;
        RECT 2697.200 1160.830 2698.380 1162.010 ;
        RECT 2697.200 1159.230 2698.380 1160.410 ;
        RECT 2697.200 1157.630 2698.380 1158.810 ;
        RECT 2697.200 1156.030 2698.380 1157.210 ;
        RECT 2697.200 1154.430 2698.380 1155.610 ;
        RECT 2697.200 1152.830 2698.380 1154.010 ;
        RECT 2899.000 1165.630 2900.180 1166.810 ;
        RECT 2899.000 1164.030 2900.180 1165.210 ;
        RECT 2899.000 1162.430 2900.180 1163.610 ;
        RECT 2899.000 1160.830 2900.180 1162.010 ;
        RECT 2899.000 1159.230 2900.180 1160.410 ;
        RECT 2899.000 1157.630 2900.180 1158.810 ;
        RECT 2899.000 1156.030 2900.180 1157.210 ;
        RECT 2899.000 1154.430 2900.180 1155.610 ;
        RECT 2899.000 1152.830 2900.180 1154.010 ;
        RECT 2919.000 1165.630 2920.180 1166.810 ;
        RECT 2919.000 1164.030 2920.180 1165.210 ;
        RECT 2919.000 1162.430 2920.180 1163.610 ;
        RECT 2919.000 1160.830 2920.180 1162.010 ;
        RECT 2919.000 1159.230 2920.180 1160.410 ;
        RECT 2919.000 1157.630 2920.180 1158.810 ;
        RECT 2919.000 1156.030 2920.180 1157.210 ;
        RECT 2919.000 1154.430 2920.180 1155.610 ;
        RECT 2919.000 1152.830 2920.180 1154.010 ;
        RECT 2923.050 1048.975 2935.430 1061.355 ;
        RECT 2967.320 1048.975 2979.700 1061.355 ;
        RECT 3136.515 1048.790 3139.295 1061.170 ;
        RECT 3213.315 1048.790 3216.095 1061.170 ;
        RECT 3290.115 1048.790 3292.895 1061.170 ;
        RECT 256.155 1045.600 257.335 1046.780 ;
        RECT 256.155 1044.000 257.335 1045.180 ;
        RECT 256.155 995.600 257.335 996.780 ;
        RECT 256.155 994.000 257.335 995.180 ;
        RECT 2923.915 995.485 2934.695 998.265 ;
        RECT 2960.190 995.895 2961.370 997.075 ;
        RECT 2961.790 995.895 2962.970 997.075 ;
        RECT 2963.390 995.895 2964.570 997.075 ;
        RECT 256.155 945.600 257.335 946.780 ;
        RECT 256.155 944.000 257.335 945.180 ;
        RECT 2923.915 917.285 2934.695 920.065 ;
        RECT 2960.190 917.695 2961.370 918.875 ;
        RECT 2961.790 917.695 2962.970 918.875 ;
        RECT 2963.390 917.695 2964.570 918.875 ;
        RECT 256.155 895.600 257.335 896.780 ;
        RECT 256.155 894.000 257.335 895.180 ;
        RECT 210.435 868.545 227.615 882.525 ;
        RECT 212.465 844.850 213.645 846.030 ;
        RECT 214.065 844.850 215.245 846.030 ;
        RECT 215.665 844.850 216.845 846.030 ;
        RECT 217.265 844.850 218.445 846.030 ;
        RECT 218.865 844.850 220.045 846.030 ;
        RECT 220.465 844.850 221.645 846.030 ;
        RECT 222.065 844.850 223.245 846.030 ;
        RECT 223.665 844.850 224.845 846.030 ;
        RECT 225.265 844.850 226.445 846.030 ;
        RECT 256.155 845.600 257.335 846.780 ;
        RECT 256.155 844.000 257.335 845.180 ;
        RECT 2923.915 839.085 2934.695 841.865 ;
        RECT 2960.190 839.495 2961.370 840.675 ;
        RECT 2961.790 839.495 2962.970 840.675 ;
        RECT 2963.390 839.495 2964.570 840.675 ;
        RECT 212.465 794.850 213.645 796.030 ;
        RECT 214.065 794.850 215.245 796.030 ;
        RECT 215.665 794.850 216.845 796.030 ;
        RECT 217.265 794.850 218.445 796.030 ;
        RECT 218.865 794.850 220.045 796.030 ;
        RECT 220.465 794.850 221.645 796.030 ;
        RECT 222.065 794.850 223.245 796.030 ;
        RECT 223.665 794.850 224.845 796.030 ;
        RECT 225.265 794.850 226.445 796.030 ;
        RECT 256.155 795.600 257.335 796.780 ;
        RECT 256.155 794.000 257.335 795.180 ;
        RECT 2923.915 760.885 2934.695 763.665 ;
        RECT 2960.190 761.295 2961.370 762.475 ;
        RECT 2961.790 761.295 2962.970 762.475 ;
        RECT 2963.390 761.295 2964.570 762.475 ;
        RECT 212.465 744.850 213.645 746.030 ;
        RECT 214.065 744.850 215.245 746.030 ;
        RECT 215.665 744.850 216.845 746.030 ;
        RECT 217.265 744.850 218.445 746.030 ;
        RECT 218.865 744.850 220.045 746.030 ;
        RECT 220.465 744.850 221.645 746.030 ;
        RECT 222.065 744.850 223.245 746.030 ;
        RECT 223.665 744.850 224.845 746.030 ;
        RECT 225.265 744.850 226.445 746.030 ;
        RECT 256.155 745.600 257.335 746.780 ;
        RECT 256.155 744.000 257.335 745.180 ;
        RECT 212.465 694.850 213.645 696.030 ;
        RECT 214.065 694.850 215.245 696.030 ;
        RECT 215.665 694.850 216.845 696.030 ;
        RECT 217.265 694.850 218.445 696.030 ;
        RECT 218.865 694.850 220.045 696.030 ;
        RECT 220.465 694.850 221.645 696.030 ;
        RECT 222.065 694.850 223.245 696.030 ;
        RECT 223.665 694.850 224.845 696.030 ;
        RECT 225.265 694.850 226.445 696.030 ;
        RECT 256.155 695.600 257.335 696.780 ;
        RECT 256.155 694.000 257.335 695.180 ;
        RECT 2923.915 682.685 2934.695 685.465 ;
        RECT 2960.190 683.095 2961.370 684.275 ;
        RECT 2961.790 683.095 2962.970 684.275 ;
        RECT 2963.390 683.095 2964.570 684.275 ;
        RECT 212.465 644.850 213.645 646.030 ;
        RECT 214.065 644.850 215.245 646.030 ;
        RECT 215.665 644.850 216.845 646.030 ;
        RECT 217.265 644.850 218.445 646.030 ;
        RECT 218.865 644.850 220.045 646.030 ;
        RECT 220.465 644.850 221.645 646.030 ;
        RECT 222.065 644.850 223.245 646.030 ;
        RECT 223.665 644.850 224.845 646.030 ;
        RECT 225.265 644.850 226.445 646.030 ;
        RECT 256.155 645.600 257.335 646.780 ;
        RECT 256.155 644.000 257.335 645.180 ;
        RECT 2960.190 604.895 2961.370 606.075 ;
        RECT 2961.790 604.895 2962.970 606.075 ;
        RECT 2963.390 604.895 2964.570 606.075 ;
        RECT 2923.915 598.485 2934.695 601.265 ;
        RECT 212.465 594.850 213.645 596.030 ;
        RECT 214.065 594.850 215.245 596.030 ;
        RECT 215.665 594.850 216.845 596.030 ;
        RECT 217.265 594.850 218.445 596.030 ;
        RECT 218.865 594.850 220.045 596.030 ;
        RECT 220.465 594.850 221.645 596.030 ;
        RECT 222.065 594.850 223.245 596.030 ;
        RECT 223.665 594.850 224.845 596.030 ;
        RECT 225.265 594.850 226.445 596.030 ;
        RECT 256.155 595.600 257.335 596.780 ;
        RECT 256.155 594.000 257.335 595.180 ;
        RECT 212.465 544.850 213.645 546.030 ;
        RECT 214.065 544.850 215.245 546.030 ;
        RECT 215.665 544.850 216.845 546.030 ;
        RECT 217.265 544.850 218.445 546.030 ;
        RECT 218.865 544.850 220.045 546.030 ;
        RECT 220.465 544.850 221.645 546.030 ;
        RECT 222.065 544.850 223.245 546.030 ;
        RECT 223.665 544.850 224.845 546.030 ;
        RECT 225.265 544.850 226.445 546.030 ;
        RECT 256.155 545.600 257.335 546.780 ;
        RECT 256.155 544.000 257.335 545.180 ;
        RECT 2923.915 526.285 2934.695 529.065 ;
        RECT 2960.190 526.695 2961.370 527.875 ;
        RECT 2961.790 526.695 2962.970 527.875 ;
        RECT 2963.390 526.695 2964.570 527.875 ;
        RECT 212.465 494.850 213.645 496.030 ;
        RECT 214.065 494.850 215.245 496.030 ;
        RECT 215.665 494.850 216.845 496.030 ;
        RECT 217.265 494.850 218.445 496.030 ;
        RECT 218.865 494.850 220.045 496.030 ;
        RECT 220.465 494.850 221.645 496.030 ;
        RECT 222.065 494.850 223.245 496.030 ;
        RECT 223.665 494.850 224.845 496.030 ;
        RECT 225.265 494.850 226.445 496.030 ;
        RECT 256.155 495.600 257.335 496.780 ;
        RECT 256.155 494.000 257.335 495.180 ;
        RECT 212.465 444.850 213.645 446.030 ;
        RECT 214.065 444.850 215.245 446.030 ;
        RECT 215.665 444.850 216.845 446.030 ;
        RECT 217.265 444.850 218.445 446.030 ;
        RECT 218.865 444.850 220.045 446.030 ;
        RECT 220.465 444.850 221.645 446.030 ;
        RECT 222.065 444.850 223.245 446.030 ;
        RECT 223.665 444.850 224.845 446.030 ;
        RECT 225.265 444.850 226.445 446.030 ;
        RECT 256.155 445.600 257.335 446.780 ;
        RECT 256.155 444.000 257.335 445.180 ;
        RECT 210.455 391.380 227.635 413.360 ;
        RECT 256.155 395.600 257.335 396.780 ;
        RECT 256.155 394.000 257.335 395.180 ;
        RECT 3161.270 392.365 3164.050 403.145 ;
        RECT 3201.160 391.700 3203.940 404.080 ;
        RECT 3141.745 384.785 3142.925 385.965 ;
        RECT 3141.745 383.185 3142.925 384.365 ;
        RECT 3141.745 381.585 3142.925 382.765 ;
        RECT 3157.245 384.785 3158.425 385.965 ;
        RECT 3157.245 383.185 3158.425 384.365 ;
        RECT 3157.245 381.585 3158.425 382.765 ;
        RECT 3172.805 384.855 3173.985 386.035 ;
        RECT 3172.805 383.255 3173.985 384.435 ;
        RECT 3172.805 381.655 3173.985 382.835 ;
        RECT 3188.255 384.835 3189.435 386.015 ;
        RECT 3188.255 383.235 3189.435 384.415 ;
        RECT 3188.255 381.635 3189.435 382.815 ;
        RECT 3203.725 384.835 3204.905 386.015 ;
        RECT 3203.725 383.235 3204.905 384.415 ;
        RECT 3203.725 381.635 3204.905 382.815 ;
        RECT 3219.265 384.895 3220.445 386.075 ;
        RECT 3219.265 383.295 3220.445 384.475 ;
        RECT 3219.265 381.695 3220.445 382.875 ;
        RECT 210.335 341.860 227.515 363.840 ;
        RECT 256.155 345.600 257.335 346.780 ;
        RECT 256.155 344.000 257.335 345.180 ;
        RECT 212.465 294.750 213.645 295.930 ;
        RECT 214.065 294.750 215.245 295.930 ;
        RECT 215.665 294.750 216.845 295.930 ;
        RECT 217.265 294.750 218.445 295.930 ;
        RECT 218.865 294.750 220.045 295.930 ;
        RECT 220.465 294.750 221.645 295.930 ;
        RECT 222.065 294.750 223.245 295.930 ;
        RECT 223.665 294.750 224.845 295.930 ;
        RECT 225.265 294.750 226.445 295.930 ;
        RECT 256.155 295.600 257.335 296.780 ;
        RECT 256.155 294.000 257.335 295.180 ;
        RECT 3141.725 276.815 3142.905 277.995 ;
        RECT 3141.725 275.215 3142.905 276.395 ;
        RECT 3141.725 273.615 3142.905 274.795 ;
        RECT 3157.225 276.815 3158.405 277.995 ;
        RECT 3157.225 275.215 3158.405 276.395 ;
        RECT 3157.225 273.615 3158.405 274.795 ;
        RECT 3172.785 276.885 3173.965 278.065 ;
        RECT 3172.785 275.285 3173.965 276.465 ;
        RECT 3172.785 273.685 3173.965 274.865 ;
        RECT 3188.235 276.865 3189.415 278.045 ;
        RECT 3188.235 275.265 3189.415 276.445 ;
        RECT 3188.235 273.665 3189.415 274.845 ;
        RECT 3203.705 276.865 3204.885 278.045 ;
        RECT 3203.705 275.265 3204.885 276.445 ;
        RECT 3203.705 273.665 3204.885 274.845 ;
        RECT 3219.245 276.925 3220.425 278.105 ;
        RECT 3219.245 275.325 3220.425 276.505 ;
        RECT 3219.245 273.725 3220.425 274.905 ;
        RECT 210.400 242.390 227.580 259.570 ;
        RECT 273.250 242.220 290.430 259.400 ;
        RECT 717.115 250.180 723.095 252.960 ;
        RECT 3332.610 235.190 3333.790 236.370 ;
        RECT 3334.210 235.190 3335.390 236.370 ;
        RECT 3335.810 235.190 3336.990 236.370 ;
        RECT 3337.410 235.190 3338.590 236.370 ;
        RECT 3339.010 235.190 3340.190 236.370 ;
        RECT 3340.610 235.190 3341.790 236.370 ;
        RECT 3342.210 235.190 3343.390 236.370 ;
        RECT 3343.810 235.190 3344.990 236.370 ;
        RECT 3345.410 235.190 3346.590 236.370 ;
      LAYER met5 ;
        RECT 281.480 1152.330 2936.870 1167.330 ;
        RECT 255.920 1043.790 266.080 1046.990 ;
        RECT 2873.230 1043.790 2901.550 1046.990 ;
        RECT 2898.350 1037.390 2901.550 1043.790 ;
        RECT 2921.870 1037.390 2936.870 1152.330 ;
        RECT 3243.040 1129.360 3256.790 1130.960 ;
        RECT 3251.120 1110.960 3256.790 1129.360 ;
        RECT 3243.200 1109.360 3256.790 1110.960 ;
        RECT 3251.120 1062.520 3256.790 1109.360 ;
        RECT 2966.260 1047.520 3347.130 1062.520 ;
        RECT 2898.350 1034.210 2936.870 1037.390 ;
        RECT 2901.550 1034.190 2936.870 1034.210 ;
        RECT 2921.870 996.990 2936.870 1034.190 ;
        RECT 3332.130 997.300 3347.130 1047.520 ;
        RECT 255.920 993.790 266.080 996.990 ;
        RECT 2873.230 993.790 2936.870 996.990 ;
        RECT 2959.880 995.700 2967.970 997.300 ;
        RECT 3325.880 995.700 3347.130 997.300 ;
        RECT 2921.870 946.990 2936.870 993.790 ;
        RECT 255.920 943.790 266.080 946.990 ;
        RECT 2873.230 943.790 2936.870 946.990 ;
        RECT 2921.870 896.990 2936.870 943.790 ;
        RECT 3332.130 919.100 3347.130 995.700 ;
        RECT 2959.880 917.500 2967.970 919.100 ;
        RECT 3325.880 917.500 3347.130 919.100 ;
        RECT 255.920 893.790 266.080 896.990 ;
        RECT 2873.230 893.790 2936.870 896.990 ;
        RECT 208.840 240.370 228.840 884.370 ;
        RECT 2921.870 846.990 2936.870 893.790 ;
        RECT 255.920 843.790 266.080 846.990 ;
        RECT 2873.230 843.790 2936.870 846.990 ;
        RECT 2921.870 796.990 2936.870 843.790 ;
        RECT 3332.130 840.900 3347.130 917.500 ;
        RECT 2959.880 839.300 2967.970 840.900 ;
        RECT 3325.880 839.300 3347.130 840.900 ;
        RECT 255.920 793.790 266.080 796.990 ;
        RECT 2873.230 793.790 2936.870 796.990 ;
        RECT 2921.870 746.990 2936.870 793.790 ;
        RECT 3332.130 762.700 3347.130 839.300 ;
        RECT 2959.880 761.100 2967.970 762.700 ;
        RECT 3325.880 761.100 3347.130 762.700 ;
        RECT 255.920 743.790 266.080 746.990 ;
        RECT 2873.230 743.790 2936.870 746.990 ;
        RECT 2921.870 696.990 2936.870 743.790 ;
        RECT 255.920 693.790 266.080 696.990 ;
        RECT 2873.230 693.790 2936.870 696.990 ;
        RECT 2921.870 646.990 2936.870 693.790 ;
        RECT 3332.130 684.500 3347.130 761.100 ;
        RECT 2959.880 682.900 2967.970 684.500 ;
        RECT 3325.880 682.900 3347.130 684.500 ;
        RECT 255.920 643.790 266.080 646.990 ;
        RECT 2873.230 643.790 2936.870 646.990 ;
        RECT 2921.870 596.990 2936.870 643.790 ;
        RECT 3332.130 606.300 3347.130 682.900 ;
        RECT 2959.880 604.700 2967.970 606.300 ;
        RECT 3325.880 604.700 3347.130 606.300 ;
        RECT 255.920 593.790 266.080 596.990 ;
        RECT 2873.230 593.790 2936.870 596.990 ;
        RECT 2921.870 546.990 2936.870 593.790 ;
        RECT 255.920 543.790 266.080 546.990 ;
        RECT 2873.230 543.790 2936.870 546.990 ;
        RECT 2921.870 496.990 2936.870 543.790 ;
        RECT 3332.130 528.100 3347.130 604.700 ;
        RECT 2959.880 526.500 2967.970 528.100 ;
        RECT 3325.880 526.500 3347.130 528.100 ;
        RECT 255.920 493.790 266.080 496.990 ;
        RECT 2873.230 493.790 2936.870 496.990 ;
        RECT 2921.870 446.990 2936.870 493.790 ;
        RECT 3332.130 467.030 3347.130 526.500 ;
        RECT 3312.610 465.430 3347.130 467.030 ;
        RECT 3332.130 458.870 3347.130 465.430 ;
        RECT 3312.420 457.270 3347.130 458.870 ;
        RECT 3332.130 450.710 3347.130 457.270 ;
        RECT 3312.520 449.110 3347.130 450.710 ;
        RECT 255.920 443.790 266.080 446.990 ;
        RECT 2873.230 443.790 2936.870 446.990 ;
        RECT 2921.870 396.990 2936.870 443.790 ;
        RECT 3209.840 425.770 3232.720 427.370 ;
        RECT 3217.720 405.410 3232.720 425.770 ;
        RECT 3332.130 405.410 3347.130 449.110 ;
        RECT 255.920 393.790 266.080 396.990 ;
        RECT 2873.230 393.790 2936.870 396.990 ;
        RECT 2921.870 346.990 2936.870 393.790 ;
        RECT 3160.010 390.410 3347.130 405.410 ;
        RECT 3226.280 386.340 3235.420 390.410 ;
        RECT 3141.340 381.340 3235.420 386.340 ;
        RECT 3231.420 353.270 3235.420 381.340 ;
        RECT 3227.680 351.670 3235.420 353.270 ;
        RECT 255.920 343.790 266.080 346.990 ;
        RECT 2873.230 343.790 2936.870 346.990 ;
        RECT 2921.870 296.990 2936.870 343.790 ;
        RECT 3231.420 336.370 3235.420 351.670 ;
        RECT 3227.510 334.770 3235.420 336.370 ;
        RECT 3231.420 319.470 3235.420 334.770 ;
        RECT 3228.120 317.870 3235.420 319.470 ;
        RECT 3231.420 302.570 3235.420 317.870 ;
        RECT 3228.120 300.970 3235.420 302.570 ;
        RECT 255.920 293.790 266.080 296.990 ;
        RECT 2873.230 293.790 2936.870 296.990 ;
        RECT 2921.870 261.110 2936.870 293.790 ;
        RECT 3231.420 285.670 3235.420 300.970 ;
        RECT 3228.120 284.070 3235.420 285.670 ;
        RECT 3231.420 278.370 3235.420 284.070 ;
        RECT 3141.320 273.370 3235.420 278.370 ;
        RECT 271.870 241.110 2936.870 261.110 ;
        RECT 3332.130 234.890 3347.130 390.410 ;
    END
  END vccd_core
  PIN vssd_core
    PORT
      LAYER met1 ;
        RECT 3240.520 233.690 3248.350 235.940 ;
        RECT 3240.520 232.990 3250.800 233.690 ;
        RECT 3240.520 232.950 3248.350 232.990 ;
      LAYER via ;
        RECT 3240.945 233.370 3247.925 235.550 ;
      LAYER met2 ;
        RECT 3240.520 233.690 3248.350 235.940 ;
        RECT 3240.520 232.990 3250.800 233.690 ;
        RECT 3240.520 232.950 3248.350 232.990 ;
      LAYER via2 ;
        RECT 3240.895 233.320 3247.975 235.600 ;
      LAYER met3 ;
        RECT 3240.520 234.220 3248.350 235.940 ;
        RECT 1208.450 197.130 1230.245 233.430 ;
        RECT 1256.500 197.130 1278.510 233.430 ;
        RECT 3240.520 232.990 3250.790 234.220 ;
        RECT 3240.520 232.950 3248.350 232.990 ;
      LAYER via3 ;
        RECT 1208.755 214.285 1229.875 233.005 ;
        RECT 1257.015 214.355 1278.135 233.075 ;
        RECT 3240.875 233.300 3247.995 235.620 ;
      LAYER met4 ;
        RECT 238.930 1172.330 316.250 1187.330 ;
        RECT 702.220 1172.240 704.620 1187.370 ;
        RECT 777.620 1172.240 780.020 1187.370 ;
        RECT 852.870 1172.240 855.270 1187.370 ;
        RECT 927.920 1172.240 930.320 1187.370 ;
        RECT 1078.620 1172.240 1081.020 1187.370 ;
        RECT 1153.870 1172.240 1156.270 1187.370 ;
        RECT 1229.120 1172.240 1231.520 1187.370 ;
        RECT 1304.370 1172.240 1306.770 1187.370 ;
        RECT 1379.620 1172.240 1382.020 1187.370 ;
        RECT 1454.870 1172.240 1457.270 1187.370 ;
        RECT 1529.920 1172.240 1532.320 1187.370 ;
        RECT 1605.870 1172.240 1608.270 1187.370 ;
        RECT 1680.620 1172.240 1683.020 1187.370 ;
        RECT 1755.570 1172.240 1757.970 1187.370 ;
        RECT 1831.120 1172.240 1833.520 1187.370 ;
        RECT 1905.770 1172.240 1908.170 1187.370 ;
        RECT 1981.220 1172.240 1983.620 1187.370 ;
        RECT 2056.870 1172.240 2059.270 1187.370 ;
        RECT 2132.120 1172.240 2134.520 1187.370 ;
        RECT 2207.370 1172.240 2209.770 1187.370 ;
        RECT 2282.620 1172.240 2285.020 1187.370 ;
        RECT 2357.870 1172.240 2360.270 1187.370 ;
        RECT 2433.120 1172.240 2435.520 1187.370 ;
        RECT 2508.370 1172.240 2510.770 1187.370 ;
        RECT 2583.620 1172.240 2586.020 1187.370 ;
        RECT 2658.870 1172.240 2661.270 1187.370 ;
        RECT 2733.870 1172.240 2736.270 1187.370 ;
        RECT 2911.310 1039.310 2956.940 1042.510 ;
        RECT 2910.360 1005.310 2956.940 1008.510 ;
        RECT 2910.360 955.310 2956.940 958.510 ;
        RECT 2910.360 905.310 2956.940 908.510 ;
        RECT 2910.360 855.310 2956.940 858.510 ;
        RECT 2910.360 805.310 2956.940 808.510 ;
        RECT 2910.360 755.310 2956.940 758.510 ;
        RECT 2910.360 705.310 2956.940 708.510 ;
        RECT 2910.360 655.310 2956.940 658.510 ;
        RECT 2910.360 605.310 2956.940 608.510 ;
        RECT 2910.360 555.310 2956.940 558.510 ;
        RECT 2910.360 505.310 2956.940 508.510 ;
        RECT 2986.510 493.800 2988.110 511.580 ;
        RECT 3063.310 494.020 3064.910 511.190 ;
        RECT 3140.110 494.020 3141.710 511.190 ;
        RECT 3216.910 494.020 3218.510 511.190 ;
        RECT 3293.710 494.020 3295.310 510.650 ;
        RECT 2983.710 479.780 2990.760 493.800 ;
        RECT 3061.120 480.250 3067.710 494.020 ;
        RECT 3137.920 480.250 3144.510 494.020 ;
        RECT 3180.400 482.170 3184.970 493.790 ;
        RECT 3181.770 472.240 3183.370 482.170 ;
        RECT 3214.720 480.250 3225.000 494.020 ;
        RECT 3291.520 480.250 3297.965 494.020 ;
        RECT 3221.770 472.240 3223.370 480.250 ;
        RECT 2910.360 455.310 2956.940 458.510 ;
        RECT 2910.360 405.310 2956.940 408.510 ;
        RECT 3149.340 369.140 3150.940 386.870 ;
        RECT 3164.840 369.140 3166.440 386.870 ;
        RECT 3180.340 369.140 3181.940 386.870 ;
        RECT 3195.840 369.140 3197.440 386.870 ;
        RECT 3211.340 369.140 3212.940 386.870 ;
        RECT 3226.840 369.140 3228.440 386.870 ;
        RECT 2910.360 355.310 2956.940 358.510 ;
        RECT 2910.360 305.310 2956.940 308.510 ;
        RECT 3149.320 262.550 3150.920 278.900 ;
        RECT 3164.820 262.550 3166.420 278.900 ;
        RECT 3180.320 262.550 3181.920 278.900 ;
        RECT 3195.820 262.550 3197.420 278.900 ;
        RECT 3211.320 262.550 3212.920 278.900 ;
        RECT 3226.820 262.550 3228.420 278.900 ;
        RECT 712.800 226.980 713.700 236.280 ;
        RECT 708.880 226.970 714.330 226.980 ;
        RECT 706.880 220.650 714.330 226.970 ;
        RECT 1208.400 213.920 1230.280 233.460 ;
        RECT 1256.510 213.940 1278.500 233.420 ;
        RECT 3240.520 232.950 3248.350 235.940 ;
      LAYER via4 ;
        RECT 240.455 1173.695 252.835 1186.075 ;
        RECT 282.275 1173.725 315.455 1186.105 ;
        RECT 702.600 1185.625 703.780 1186.805 ;
        RECT 702.600 1184.025 703.780 1185.205 ;
        RECT 702.600 1182.425 703.780 1183.605 ;
        RECT 702.600 1180.825 703.780 1182.005 ;
        RECT 702.600 1179.225 703.780 1180.405 ;
        RECT 702.600 1177.625 703.780 1178.805 ;
        RECT 702.600 1176.025 703.780 1177.205 ;
        RECT 702.600 1174.425 703.780 1175.605 ;
        RECT 702.600 1172.825 703.780 1174.005 ;
        RECT 778.000 1185.625 779.180 1186.805 ;
        RECT 778.000 1184.025 779.180 1185.205 ;
        RECT 778.000 1182.425 779.180 1183.605 ;
        RECT 778.000 1180.825 779.180 1182.005 ;
        RECT 778.000 1179.225 779.180 1180.405 ;
        RECT 778.000 1177.625 779.180 1178.805 ;
        RECT 778.000 1176.025 779.180 1177.205 ;
        RECT 778.000 1174.425 779.180 1175.605 ;
        RECT 778.000 1172.825 779.180 1174.005 ;
        RECT 853.250 1185.625 854.430 1186.805 ;
        RECT 853.250 1184.025 854.430 1185.205 ;
        RECT 853.250 1182.425 854.430 1183.605 ;
        RECT 853.250 1180.825 854.430 1182.005 ;
        RECT 853.250 1179.225 854.430 1180.405 ;
        RECT 853.250 1177.625 854.430 1178.805 ;
        RECT 853.250 1176.025 854.430 1177.205 ;
        RECT 853.250 1174.425 854.430 1175.605 ;
        RECT 853.250 1172.825 854.430 1174.005 ;
        RECT 928.300 1185.625 929.480 1186.805 ;
        RECT 928.300 1184.025 929.480 1185.205 ;
        RECT 928.300 1182.425 929.480 1183.605 ;
        RECT 928.300 1180.825 929.480 1182.005 ;
        RECT 928.300 1179.225 929.480 1180.405 ;
        RECT 928.300 1177.625 929.480 1178.805 ;
        RECT 928.300 1176.025 929.480 1177.205 ;
        RECT 928.300 1174.425 929.480 1175.605 ;
        RECT 928.300 1172.825 929.480 1174.005 ;
        RECT 1079.000 1185.625 1080.180 1186.805 ;
        RECT 1079.000 1184.025 1080.180 1185.205 ;
        RECT 1079.000 1182.425 1080.180 1183.605 ;
        RECT 1079.000 1180.825 1080.180 1182.005 ;
        RECT 1079.000 1179.225 1080.180 1180.405 ;
        RECT 1079.000 1177.625 1080.180 1178.805 ;
        RECT 1079.000 1176.025 1080.180 1177.205 ;
        RECT 1079.000 1174.425 1080.180 1175.605 ;
        RECT 1079.000 1172.825 1080.180 1174.005 ;
        RECT 1154.250 1185.625 1155.430 1186.805 ;
        RECT 1154.250 1184.025 1155.430 1185.205 ;
        RECT 1154.250 1182.425 1155.430 1183.605 ;
        RECT 1154.250 1180.825 1155.430 1182.005 ;
        RECT 1154.250 1179.225 1155.430 1180.405 ;
        RECT 1154.250 1177.625 1155.430 1178.805 ;
        RECT 1154.250 1176.025 1155.430 1177.205 ;
        RECT 1154.250 1174.425 1155.430 1175.605 ;
        RECT 1154.250 1172.825 1155.430 1174.005 ;
        RECT 1229.500 1185.625 1230.680 1186.805 ;
        RECT 1229.500 1184.025 1230.680 1185.205 ;
        RECT 1229.500 1182.425 1230.680 1183.605 ;
        RECT 1229.500 1180.825 1230.680 1182.005 ;
        RECT 1229.500 1179.225 1230.680 1180.405 ;
        RECT 1229.500 1177.625 1230.680 1178.805 ;
        RECT 1229.500 1176.025 1230.680 1177.205 ;
        RECT 1229.500 1174.425 1230.680 1175.605 ;
        RECT 1229.500 1172.825 1230.680 1174.005 ;
        RECT 1304.750 1185.625 1305.930 1186.805 ;
        RECT 1304.750 1184.025 1305.930 1185.205 ;
        RECT 1304.750 1182.425 1305.930 1183.605 ;
        RECT 1304.750 1180.825 1305.930 1182.005 ;
        RECT 1304.750 1179.225 1305.930 1180.405 ;
        RECT 1304.750 1177.625 1305.930 1178.805 ;
        RECT 1304.750 1176.025 1305.930 1177.205 ;
        RECT 1304.750 1174.425 1305.930 1175.605 ;
        RECT 1304.750 1172.825 1305.930 1174.005 ;
        RECT 1380.000 1185.625 1381.180 1186.805 ;
        RECT 1380.000 1184.025 1381.180 1185.205 ;
        RECT 1380.000 1182.425 1381.180 1183.605 ;
        RECT 1380.000 1180.825 1381.180 1182.005 ;
        RECT 1380.000 1179.225 1381.180 1180.405 ;
        RECT 1380.000 1177.625 1381.180 1178.805 ;
        RECT 1380.000 1176.025 1381.180 1177.205 ;
        RECT 1380.000 1174.425 1381.180 1175.605 ;
        RECT 1380.000 1172.825 1381.180 1174.005 ;
        RECT 1455.250 1185.625 1456.430 1186.805 ;
        RECT 1455.250 1184.025 1456.430 1185.205 ;
        RECT 1455.250 1182.425 1456.430 1183.605 ;
        RECT 1455.250 1180.825 1456.430 1182.005 ;
        RECT 1455.250 1179.225 1456.430 1180.405 ;
        RECT 1455.250 1177.625 1456.430 1178.805 ;
        RECT 1455.250 1176.025 1456.430 1177.205 ;
        RECT 1455.250 1174.425 1456.430 1175.605 ;
        RECT 1455.250 1172.825 1456.430 1174.005 ;
        RECT 1530.300 1185.625 1531.480 1186.805 ;
        RECT 1530.300 1184.025 1531.480 1185.205 ;
        RECT 1530.300 1182.425 1531.480 1183.605 ;
        RECT 1530.300 1180.825 1531.480 1182.005 ;
        RECT 1530.300 1179.225 1531.480 1180.405 ;
        RECT 1530.300 1177.625 1531.480 1178.805 ;
        RECT 1530.300 1176.025 1531.480 1177.205 ;
        RECT 1530.300 1174.425 1531.480 1175.605 ;
        RECT 1530.300 1172.825 1531.480 1174.005 ;
        RECT 1606.250 1185.625 1607.430 1186.805 ;
        RECT 1606.250 1184.025 1607.430 1185.205 ;
        RECT 1606.250 1182.425 1607.430 1183.605 ;
        RECT 1606.250 1180.825 1607.430 1182.005 ;
        RECT 1606.250 1179.225 1607.430 1180.405 ;
        RECT 1606.250 1177.625 1607.430 1178.805 ;
        RECT 1606.250 1176.025 1607.430 1177.205 ;
        RECT 1606.250 1174.425 1607.430 1175.605 ;
        RECT 1606.250 1172.825 1607.430 1174.005 ;
        RECT 1681.000 1185.625 1682.180 1186.805 ;
        RECT 1681.000 1184.025 1682.180 1185.205 ;
        RECT 1681.000 1182.425 1682.180 1183.605 ;
        RECT 1681.000 1180.825 1682.180 1182.005 ;
        RECT 1681.000 1179.225 1682.180 1180.405 ;
        RECT 1681.000 1177.625 1682.180 1178.805 ;
        RECT 1681.000 1176.025 1682.180 1177.205 ;
        RECT 1681.000 1174.425 1682.180 1175.605 ;
        RECT 1681.000 1172.825 1682.180 1174.005 ;
        RECT 1755.950 1185.625 1757.130 1186.805 ;
        RECT 1755.950 1184.025 1757.130 1185.205 ;
        RECT 1755.950 1182.425 1757.130 1183.605 ;
        RECT 1755.950 1180.825 1757.130 1182.005 ;
        RECT 1755.950 1179.225 1757.130 1180.405 ;
        RECT 1755.950 1177.625 1757.130 1178.805 ;
        RECT 1755.950 1176.025 1757.130 1177.205 ;
        RECT 1755.950 1174.425 1757.130 1175.605 ;
        RECT 1755.950 1172.825 1757.130 1174.005 ;
        RECT 1831.500 1185.625 1832.680 1186.805 ;
        RECT 1831.500 1184.025 1832.680 1185.205 ;
        RECT 1831.500 1182.425 1832.680 1183.605 ;
        RECT 1831.500 1180.825 1832.680 1182.005 ;
        RECT 1831.500 1179.225 1832.680 1180.405 ;
        RECT 1831.500 1177.625 1832.680 1178.805 ;
        RECT 1831.500 1176.025 1832.680 1177.205 ;
        RECT 1831.500 1174.425 1832.680 1175.605 ;
        RECT 1831.500 1172.825 1832.680 1174.005 ;
        RECT 1906.150 1185.625 1907.330 1186.805 ;
        RECT 1906.150 1184.025 1907.330 1185.205 ;
        RECT 1906.150 1182.425 1907.330 1183.605 ;
        RECT 1906.150 1180.825 1907.330 1182.005 ;
        RECT 1906.150 1179.225 1907.330 1180.405 ;
        RECT 1906.150 1177.625 1907.330 1178.805 ;
        RECT 1906.150 1176.025 1907.330 1177.205 ;
        RECT 1906.150 1174.425 1907.330 1175.605 ;
        RECT 1906.150 1172.825 1907.330 1174.005 ;
        RECT 1981.600 1185.625 1982.780 1186.805 ;
        RECT 1981.600 1184.025 1982.780 1185.205 ;
        RECT 1981.600 1182.425 1982.780 1183.605 ;
        RECT 1981.600 1180.825 1982.780 1182.005 ;
        RECT 1981.600 1179.225 1982.780 1180.405 ;
        RECT 1981.600 1177.625 1982.780 1178.805 ;
        RECT 1981.600 1176.025 1982.780 1177.205 ;
        RECT 1981.600 1174.425 1982.780 1175.605 ;
        RECT 1981.600 1172.825 1982.780 1174.005 ;
        RECT 2057.250 1185.625 2058.430 1186.805 ;
        RECT 2057.250 1184.025 2058.430 1185.205 ;
        RECT 2057.250 1182.425 2058.430 1183.605 ;
        RECT 2057.250 1180.825 2058.430 1182.005 ;
        RECT 2057.250 1179.225 2058.430 1180.405 ;
        RECT 2057.250 1177.625 2058.430 1178.805 ;
        RECT 2057.250 1176.025 2058.430 1177.205 ;
        RECT 2057.250 1174.425 2058.430 1175.605 ;
        RECT 2057.250 1172.825 2058.430 1174.005 ;
        RECT 2132.500 1185.625 2133.680 1186.805 ;
        RECT 2132.500 1184.025 2133.680 1185.205 ;
        RECT 2132.500 1182.425 2133.680 1183.605 ;
        RECT 2132.500 1180.825 2133.680 1182.005 ;
        RECT 2132.500 1179.225 2133.680 1180.405 ;
        RECT 2132.500 1177.625 2133.680 1178.805 ;
        RECT 2132.500 1176.025 2133.680 1177.205 ;
        RECT 2132.500 1174.425 2133.680 1175.605 ;
        RECT 2132.500 1172.825 2133.680 1174.005 ;
        RECT 2207.750 1185.625 2208.930 1186.805 ;
        RECT 2207.750 1184.025 2208.930 1185.205 ;
        RECT 2207.750 1182.425 2208.930 1183.605 ;
        RECT 2207.750 1180.825 2208.930 1182.005 ;
        RECT 2207.750 1179.225 2208.930 1180.405 ;
        RECT 2207.750 1177.625 2208.930 1178.805 ;
        RECT 2207.750 1176.025 2208.930 1177.205 ;
        RECT 2207.750 1174.425 2208.930 1175.605 ;
        RECT 2207.750 1172.825 2208.930 1174.005 ;
        RECT 2283.000 1185.625 2284.180 1186.805 ;
        RECT 2283.000 1184.025 2284.180 1185.205 ;
        RECT 2283.000 1182.425 2284.180 1183.605 ;
        RECT 2283.000 1180.825 2284.180 1182.005 ;
        RECT 2283.000 1179.225 2284.180 1180.405 ;
        RECT 2283.000 1177.625 2284.180 1178.805 ;
        RECT 2283.000 1176.025 2284.180 1177.205 ;
        RECT 2283.000 1174.425 2284.180 1175.605 ;
        RECT 2283.000 1172.825 2284.180 1174.005 ;
        RECT 2358.250 1185.625 2359.430 1186.805 ;
        RECT 2358.250 1184.025 2359.430 1185.205 ;
        RECT 2358.250 1182.425 2359.430 1183.605 ;
        RECT 2358.250 1180.825 2359.430 1182.005 ;
        RECT 2358.250 1179.225 2359.430 1180.405 ;
        RECT 2358.250 1177.625 2359.430 1178.805 ;
        RECT 2358.250 1176.025 2359.430 1177.205 ;
        RECT 2358.250 1174.425 2359.430 1175.605 ;
        RECT 2358.250 1172.825 2359.430 1174.005 ;
        RECT 2433.500 1185.625 2434.680 1186.805 ;
        RECT 2433.500 1184.025 2434.680 1185.205 ;
        RECT 2433.500 1182.425 2434.680 1183.605 ;
        RECT 2433.500 1180.825 2434.680 1182.005 ;
        RECT 2433.500 1179.225 2434.680 1180.405 ;
        RECT 2433.500 1177.625 2434.680 1178.805 ;
        RECT 2433.500 1176.025 2434.680 1177.205 ;
        RECT 2433.500 1174.425 2434.680 1175.605 ;
        RECT 2433.500 1172.825 2434.680 1174.005 ;
        RECT 2508.750 1185.625 2509.930 1186.805 ;
        RECT 2508.750 1184.025 2509.930 1185.205 ;
        RECT 2508.750 1182.425 2509.930 1183.605 ;
        RECT 2508.750 1180.825 2509.930 1182.005 ;
        RECT 2508.750 1179.225 2509.930 1180.405 ;
        RECT 2508.750 1177.625 2509.930 1178.805 ;
        RECT 2508.750 1176.025 2509.930 1177.205 ;
        RECT 2508.750 1174.425 2509.930 1175.605 ;
        RECT 2508.750 1172.825 2509.930 1174.005 ;
        RECT 2584.000 1185.625 2585.180 1186.805 ;
        RECT 2584.000 1184.025 2585.180 1185.205 ;
        RECT 2584.000 1182.425 2585.180 1183.605 ;
        RECT 2584.000 1180.825 2585.180 1182.005 ;
        RECT 2584.000 1179.225 2585.180 1180.405 ;
        RECT 2584.000 1177.625 2585.180 1178.805 ;
        RECT 2584.000 1176.025 2585.180 1177.205 ;
        RECT 2584.000 1174.425 2585.180 1175.605 ;
        RECT 2584.000 1172.825 2585.180 1174.005 ;
        RECT 2659.250 1185.625 2660.430 1186.805 ;
        RECT 2659.250 1184.025 2660.430 1185.205 ;
        RECT 2659.250 1182.425 2660.430 1183.605 ;
        RECT 2659.250 1180.825 2660.430 1182.005 ;
        RECT 2659.250 1179.225 2660.430 1180.405 ;
        RECT 2659.250 1177.625 2660.430 1178.805 ;
        RECT 2659.250 1176.025 2660.430 1177.205 ;
        RECT 2659.250 1174.425 2660.430 1175.605 ;
        RECT 2659.250 1172.825 2660.430 1174.005 ;
        RECT 2734.250 1185.625 2735.430 1186.805 ;
        RECT 2734.250 1184.025 2735.430 1185.205 ;
        RECT 2734.250 1182.425 2735.430 1183.605 ;
        RECT 2734.250 1180.825 2735.430 1182.005 ;
        RECT 2734.250 1179.225 2735.430 1180.405 ;
        RECT 2734.250 1177.625 2735.430 1178.805 ;
        RECT 2734.250 1176.025 2735.430 1177.205 ;
        RECT 2734.250 1174.425 2735.430 1175.605 ;
        RECT 2734.250 1172.825 2735.430 1174.005 ;
        RECT 2912.000 1040.330 2913.180 1041.510 ;
        RECT 2913.600 1040.330 2914.780 1041.510 ;
        RECT 2915.200 1040.330 2916.380 1041.510 ;
        RECT 2916.800 1040.330 2917.980 1041.510 ;
        RECT 2942.465 1040.330 2943.645 1041.510 ;
        RECT 2944.065 1040.330 2945.245 1041.510 ;
        RECT 2945.665 1040.330 2946.845 1041.510 ;
        RECT 2947.265 1040.330 2948.445 1041.510 ;
        RECT 2948.865 1040.330 2950.045 1041.510 ;
        RECT 2950.465 1040.330 2951.645 1041.510 ;
        RECT 2952.065 1040.330 2953.245 1041.510 ;
        RECT 2953.665 1040.330 2954.845 1041.510 ;
        RECT 2955.265 1040.330 2956.445 1041.510 ;
        RECT 2911.020 1006.270 2912.200 1007.450 ;
        RECT 2912.620 1006.270 2913.800 1007.450 ;
        RECT 2942.465 1006.250 2943.645 1007.430 ;
        RECT 2944.065 1006.250 2945.245 1007.430 ;
        RECT 2945.665 1006.250 2946.845 1007.430 ;
        RECT 2947.265 1006.250 2948.445 1007.430 ;
        RECT 2948.865 1006.250 2950.045 1007.430 ;
        RECT 2950.465 1006.250 2951.645 1007.430 ;
        RECT 2952.065 1006.250 2953.245 1007.430 ;
        RECT 2953.665 1006.250 2954.845 1007.430 ;
        RECT 2955.265 1006.250 2956.445 1007.430 ;
        RECT 2911.020 956.270 2912.200 957.450 ;
        RECT 2912.620 956.270 2913.800 957.450 ;
        RECT 2942.465 956.250 2943.645 957.430 ;
        RECT 2944.065 956.250 2945.245 957.430 ;
        RECT 2945.665 956.250 2946.845 957.430 ;
        RECT 2947.265 956.250 2948.445 957.430 ;
        RECT 2948.865 956.250 2950.045 957.430 ;
        RECT 2950.465 956.250 2951.645 957.430 ;
        RECT 2952.065 956.250 2953.245 957.430 ;
        RECT 2953.665 956.250 2954.845 957.430 ;
        RECT 2955.265 956.250 2956.445 957.430 ;
        RECT 2911.020 906.270 2912.200 907.450 ;
        RECT 2912.620 906.270 2913.800 907.450 ;
        RECT 2942.465 906.250 2943.645 907.430 ;
        RECT 2944.065 906.250 2945.245 907.430 ;
        RECT 2945.665 906.250 2946.845 907.430 ;
        RECT 2947.265 906.250 2948.445 907.430 ;
        RECT 2948.865 906.250 2950.045 907.430 ;
        RECT 2950.465 906.250 2951.645 907.430 ;
        RECT 2952.065 906.250 2953.245 907.430 ;
        RECT 2953.665 906.250 2954.845 907.430 ;
        RECT 2955.265 906.250 2956.445 907.430 ;
        RECT 2911.020 856.270 2912.200 857.450 ;
        RECT 2912.620 856.270 2913.800 857.450 ;
        RECT 2942.465 856.250 2943.645 857.430 ;
        RECT 2944.065 856.250 2945.245 857.430 ;
        RECT 2945.665 856.250 2946.845 857.430 ;
        RECT 2947.265 856.250 2948.445 857.430 ;
        RECT 2948.865 856.250 2950.045 857.430 ;
        RECT 2950.465 856.250 2951.645 857.430 ;
        RECT 2952.065 856.250 2953.245 857.430 ;
        RECT 2953.665 856.250 2954.845 857.430 ;
        RECT 2955.265 856.250 2956.445 857.430 ;
        RECT 2911.020 806.270 2912.200 807.450 ;
        RECT 2912.620 806.270 2913.800 807.450 ;
        RECT 2942.465 806.250 2943.645 807.430 ;
        RECT 2944.065 806.250 2945.245 807.430 ;
        RECT 2945.665 806.250 2946.845 807.430 ;
        RECT 2947.265 806.250 2948.445 807.430 ;
        RECT 2948.865 806.250 2950.045 807.430 ;
        RECT 2950.465 806.250 2951.645 807.430 ;
        RECT 2952.065 806.250 2953.245 807.430 ;
        RECT 2953.665 806.250 2954.845 807.430 ;
        RECT 2955.265 806.250 2956.445 807.430 ;
        RECT 2911.020 756.270 2912.200 757.450 ;
        RECT 2912.620 756.270 2913.800 757.450 ;
        RECT 2942.465 756.250 2943.645 757.430 ;
        RECT 2944.065 756.250 2945.245 757.430 ;
        RECT 2945.665 756.250 2946.845 757.430 ;
        RECT 2947.265 756.250 2948.445 757.430 ;
        RECT 2948.865 756.250 2950.045 757.430 ;
        RECT 2950.465 756.250 2951.645 757.430 ;
        RECT 2952.065 756.250 2953.245 757.430 ;
        RECT 2953.665 756.250 2954.845 757.430 ;
        RECT 2955.265 756.250 2956.445 757.430 ;
        RECT 2911.020 706.270 2912.200 707.450 ;
        RECT 2912.620 706.270 2913.800 707.450 ;
        RECT 2942.465 706.250 2943.645 707.430 ;
        RECT 2944.065 706.250 2945.245 707.430 ;
        RECT 2945.665 706.250 2946.845 707.430 ;
        RECT 2947.265 706.250 2948.445 707.430 ;
        RECT 2948.865 706.250 2950.045 707.430 ;
        RECT 2950.465 706.250 2951.645 707.430 ;
        RECT 2952.065 706.250 2953.245 707.430 ;
        RECT 2953.665 706.250 2954.845 707.430 ;
        RECT 2955.265 706.250 2956.445 707.430 ;
        RECT 2911.020 656.270 2912.200 657.450 ;
        RECT 2912.620 656.270 2913.800 657.450 ;
        RECT 2942.465 656.250 2943.645 657.430 ;
        RECT 2944.065 656.250 2945.245 657.430 ;
        RECT 2945.665 656.250 2946.845 657.430 ;
        RECT 2947.265 656.250 2948.445 657.430 ;
        RECT 2948.865 656.250 2950.045 657.430 ;
        RECT 2950.465 656.250 2951.645 657.430 ;
        RECT 2952.065 656.250 2953.245 657.430 ;
        RECT 2953.665 656.250 2954.845 657.430 ;
        RECT 2955.265 656.250 2956.445 657.430 ;
        RECT 2911.020 606.270 2912.200 607.450 ;
        RECT 2912.620 606.270 2913.800 607.450 ;
        RECT 2942.465 606.250 2943.645 607.430 ;
        RECT 2944.065 606.250 2945.245 607.430 ;
        RECT 2945.665 606.250 2946.845 607.430 ;
        RECT 2947.265 606.250 2948.445 607.430 ;
        RECT 2948.865 606.250 2950.045 607.430 ;
        RECT 2950.465 606.250 2951.645 607.430 ;
        RECT 2952.065 606.250 2953.245 607.430 ;
        RECT 2953.665 606.250 2954.845 607.430 ;
        RECT 2955.265 606.250 2956.445 607.430 ;
        RECT 2911.020 556.270 2912.200 557.450 ;
        RECT 2912.620 556.270 2913.800 557.450 ;
        RECT 2942.465 556.250 2943.645 557.430 ;
        RECT 2944.065 556.250 2945.245 557.430 ;
        RECT 2945.665 556.250 2946.845 557.430 ;
        RECT 2947.265 556.250 2948.445 557.430 ;
        RECT 2948.865 556.250 2950.045 557.430 ;
        RECT 2950.465 556.250 2951.645 557.430 ;
        RECT 2952.065 556.250 2953.245 557.430 ;
        RECT 2953.665 556.250 2954.845 557.430 ;
        RECT 2955.265 556.250 2956.445 557.430 ;
        RECT 2911.020 506.270 2912.200 507.450 ;
        RECT 2912.620 506.270 2913.800 507.450 ;
        RECT 2942.465 506.250 2943.645 507.430 ;
        RECT 2944.065 506.250 2945.245 507.430 ;
        RECT 2945.665 506.250 2946.845 507.430 ;
        RECT 2947.265 506.250 2948.445 507.430 ;
        RECT 2948.865 506.250 2950.045 507.430 ;
        RECT 2950.465 506.250 2951.645 507.430 ;
        RECT 2952.065 506.250 2953.245 507.430 ;
        RECT 2953.665 506.250 2954.845 507.430 ;
        RECT 2955.265 506.250 2956.445 507.430 ;
        RECT 2985.060 480.635 2989.440 493.015 ;
        RECT 3062.315 480.945 3066.695 493.325 ;
        RECT 3139.115 480.945 3143.495 493.325 ;
        RECT 3181.295 483.425 3184.075 492.605 ;
        RECT 3215.915 480.945 3223.495 493.325 ;
        RECT 3292.715 480.945 3297.095 493.325 ;
        RECT 2911.020 456.270 2912.200 457.450 ;
        RECT 2912.620 456.270 2913.800 457.450 ;
        RECT 2942.465 456.250 2943.645 457.430 ;
        RECT 2944.065 456.250 2945.245 457.430 ;
        RECT 2945.665 456.250 2946.845 457.430 ;
        RECT 2947.265 456.250 2948.445 457.430 ;
        RECT 2948.865 456.250 2950.045 457.430 ;
        RECT 2950.465 456.250 2951.645 457.430 ;
        RECT 2952.065 456.250 2953.245 457.430 ;
        RECT 2953.665 456.250 2954.845 457.430 ;
        RECT 2955.265 456.250 2956.445 457.430 ;
        RECT 2911.020 406.270 2912.200 407.450 ;
        RECT 2912.620 406.270 2913.800 407.450 ;
        RECT 2942.465 406.250 2943.645 407.430 ;
        RECT 2944.065 406.250 2945.245 407.430 ;
        RECT 2945.665 406.250 2946.845 407.430 ;
        RECT 2947.265 406.250 2948.445 407.430 ;
        RECT 2948.865 406.250 2950.045 407.430 ;
        RECT 2950.465 406.250 2951.645 407.430 ;
        RECT 2952.065 406.250 2953.245 407.430 ;
        RECT 2953.665 406.250 2954.845 407.430 ;
        RECT 2955.265 406.250 2956.445 407.430 ;
        RECT 3149.505 377.775 3150.685 378.955 ;
        RECT 3149.505 376.175 3150.685 377.355 ;
        RECT 3149.505 374.575 3150.685 375.755 ;
        RECT 3165.005 377.775 3166.185 378.955 ;
        RECT 3165.005 376.175 3166.185 377.355 ;
        RECT 3165.005 374.575 3166.185 375.755 ;
        RECT 3180.475 377.795 3181.655 378.975 ;
        RECT 3180.475 376.195 3181.655 377.375 ;
        RECT 3180.475 374.595 3181.655 375.775 ;
        RECT 3196.015 377.815 3197.195 378.995 ;
        RECT 3196.015 376.215 3197.195 377.395 ;
        RECT 3196.015 374.615 3197.195 375.795 ;
        RECT 3211.535 377.775 3212.715 378.955 ;
        RECT 3211.535 376.175 3212.715 377.355 ;
        RECT 3211.535 374.575 3212.715 375.755 ;
        RECT 3227.045 377.905 3228.225 379.085 ;
        RECT 3227.045 376.305 3228.225 377.485 ;
        RECT 3227.045 374.705 3228.225 375.885 ;
        RECT 2911.020 356.270 2912.200 357.450 ;
        RECT 2912.620 356.270 2913.800 357.450 ;
        RECT 2942.465 356.250 2943.645 357.430 ;
        RECT 2944.065 356.250 2945.245 357.430 ;
        RECT 2945.665 356.250 2946.845 357.430 ;
        RECT 2947.265 356.250 2948.445 357.430 ;
        RECT 2948.865 356.250 2950.045 357.430 ;
        RECT 2950.465 356.250 2951.645 357.430 ;
        RECT 2952.065 356.250 2953.245 357.430 ;
        RECT 2953.665 356.250 2954.845 357.430 ;
        RECT 2955.265 356.250 2956.445 357.430 ;
        RECT 2911.020 306.270 2912.200 307.450 ;
        RECT 2912.620 306.270 2913.800 307.450 ;
        RECT 2942.465 306.250 2943.645 307.430 ;
        RECT 2944.065 306.250 2945.245 307.430 ;
        RECT 2945.665 306.250 2946.845 307.430 ;
        RECT 2947.265 306.250 2948.445 307.430 ;
        RECT 2948.865 306.250 2950.045 307.430 ;
        RECT 2950.465 306.250 2951.645 307.430 ;
        RECT 2952.065 306.250 2953.245 307.430 ;
        RECT 2953.665 306.250 2954.845 307.430 ;
        RECT 2955.265 306.250 2956.445 307.430 ;
        RECT 3149.485 269.805 3150.665 270.985 ;
        RECT 3149.485 268.205 3150.665 269.385 ;
        RECT 3149.485 266.605 3150.665 267.785 ;
        RECT 3164.985 269.805 3166.165 270.985 ;
        RECT 3164.985 268.205 3166.165 269.385 ;
        RECT 3164.985 266.605 3166.165 267.785 ;
        RECT 3180.455 269.825 3181.635 271.005 ;
        RECT 3180.455 268.225 3181.635 269.405 ;
        RECT 3180.455 266.625 3181.635 267.805 ;
        RECT 3195.995 269.845 3197.175 271.025 ;
        RECT 3195.995 268.245 3197.175 269.425 ;
        RECT 3195.995 266.645 3197.175 267.825 ;
        RECT 3211.515 269.805 3212.695 270.985 ;
        RECT 3211.515 268.205 3212.695 269.385 ;
        RECT 3211.515 266.605 3212.695 267.785 ;
        RECT 3227.025 269.935 3228.205 271.115 ;
        RECT 3227.025 268.335 3228.205 269.515 ;
        RECT 3227.025 266.735 3228.205 267.915 ;
        RECT 3241.445 233.870 3242.625 235.050 ;
        RECT 3243.045 233.870 3244.225 235.050 ;
        RECT 3244.645 233.870 3245.825 235.050 ;
        RECT 3246.245 233.870 3247.425 235.050 ;
        RECT 707.640 221.590 713.620 225.970 ;
        RECT 1209.125 214.255 1229.505 233.035 ;
        RECT 1257.385 214.325 1277.765 233.105 ;
      LAYER met5 ;
        RECT 239.180 1058.490 254.180 1188.060 ;
        RECT 281.440 1172.330 2956.950 1187.330 ;
        RECT 2941.950 1130.420 2956.950 1172.330 ;
        RECT 2941.950 1120.960 3201.830 1130.420 ;
        RECT 2941.950 1120.410 3209.990 1120.960 ;
        RECT 239.180 1055.290 266.160 1058.490 ;
        RECT 2873.230 1055.290 2914.550 1058.490 ;
        RECT 239.180 1008.490 254.180 1055.290 ;
        RECT 2911.350 1042.510 2914.550 1055.290 ;
        RECT 2911.350 1039.310 2918.710 1042.510 ;
        RECT 2941.950 1036.400 2956.950 1120.410 ;
        RECT 3197.330 1119.360 3209.990 1120.410 ;
        RECT 2941.950 1034.800 2967.970 1036.400 ;
        RECT 239.180 1005.290 266.160 1008.490 ;
        RECT 2873.230 1005.290 2914.550 1008.490 ;
        RECT 239.180 958.490 254.180 1005.290 ;
        RECT 239.180 955.290 266.160 958.490 ;
        RECT 2873.230 955.290 2914.550 958.490 ;
        RECT 2941.950 958.200 2956.950 1034.800 ;
        RECT 2941.950 956.600 2967.970 958.200 ;
        RECT 239.180 908.490 254.180 955.290 ;
        RECT 239.180 905.290 266.160 908.490 ;
        RECT 2873.230 905.290 2914.550 908.490 ;
        RECT 239.180 858.490 254.180 905.290 ;
        RECT 2941.950 880.000 2956.950 956.600 ;
        RECT 2941.950 878.400 2967.970 880.000 ;
        RECT 239.180 855.290 266.160 858.490 ;
        RECT 2873.230 855.290 2914.550 858.490 ;
        RECT 239.180 833.940 254.180 855.290 ;
        RECT 234.180 808.490 254.180 833.940 ;
        RECT 234.180 805.290 266.160 808.490 ;
        RECT 2873.230 805.290 2914.550 808.490 ;
        RECT 234.180 758.490 254.180 805.290 ;
        RECT 2941.950 801.800 2956.950 878.400 ;
        RECT 2941.950 800.200 2967.970 801.800 ;
        RECT 234.180 755.290 266.160 758.490 ;
        RECT 2873.230 755.290 2914.550 758.490 ;
        RECT 234.180 708.490 254.180 755.290 ;
        RECT 2941.950 723.600 2956.950 800.200 ;
        RECT 2941.950 722.000 2967.970 723.600 ;
        RECT 234.180 705.290 266.160 708.490 ;
        RECT 2873.230 705.290 2914.550 708.490 ;
        RECT 234.180 658.490 254.180 705.290 ;
        RECT 234.180 655.290 266.160 658.490 ;
        RECT 2873.230 655.290 2914.550 658.490 ;
        RECT 234.180 608.490 254.180 655.290 ;
        RECT 2941.950 645.400 2956.950 722.000 ;
        RECT 2941.950 643.800 2967.970 645.400 ;
        RECT 234.180 605.290 266.160 608.490 ;
        RECT 2873.230 605.290 2914.550 608.490 ;
        RECT 234.180 558.490 254.180 605.290 ;
        RECT 2941.950 567.200 2956.950 643.800 ;
        RECT 2941.950 565.600 2968.050 567.200 ;
        RECT 234.180 555.290 266.160 558.490 ;
        RECT 2873.230 555.290 2914.550 558.490 ;
        RECT 234.180 508.490 254.180 555.290 ;
        RECT 234.180 505.290 266.160 508.490 ;
        RECT 2873.230 505.290 2914.550 508.490 ;
        RECT 234.180 458.490 254.180 505.290 ;
        RECT 2941.950 494.780 2956.950 565.600 ;
        RECT 2941.950 479.780 3297.965 494.780 ;
        RECT 234.180 455.290 266.160 458.490 ;
        RECT 2873.230 455.290 2914.550 458.490 ;
        RECT 234.180 408.490 254.180 455.290 ;
        RECT 234.180 405.290 266.160 408.490 ;
        RECT 2873.230 405.290 2914.550 408.490 ;
        RECT 234.180 358.490 254.180 405.290 ;
        RECT 234.180 355.290 266.160 358.490 ;
        RECT 2873.230 355.290 2914.550 358.490 ;
        RECT 234.180 308.490 254.180 355.290 ;
        RECT 234.180 305.290 266.160 308.490 ;
        RECT 2873.230 305.290 2914.550 308.490 ;
        RECT 234.180 233.940 254.180 305.290 ;
        RECT 2941.950 235.940 2956.950 479.780 ;
        RECT 3124.120 447.370 3139.120 479.780 ;
        RECT 3254.970 462.950 3269.970 479.780 ;
        RECT 3254.970 461.350 3288.770 462.950 ;
        RECT 3254.970 454.790 3269.970 461.350 ;
        RECT 3254.970 453.190 3288.920 454.790 ;
        RECT 3254.970 452.610 3269.970 453.190 ;
        RECT 3124.120 445.770 3146.810 447.370 ;
        RECT 3124.120 445.060 3139.120 445.770 ;
        RECT 3128.090 379.340 3135.170 445.060 ;
        RECT 3128.090 374.340 3228.690 379.340 ;
        RECT 3128.090 361.720 3132.090 374.340 ;
        RECT 3128.090 360.120 3134.840 361.720 ;
        RECT 3128.090 344.820 3132.090 360.120 ;
        RECT 3128.090 343.220 3134.840 344.820 ;
        RECT 3128.090 327.920 3132.090 343.220 ;
        RECT 3128.090 326.320 3134.840 327.920 ;
        RECT 3128.090 311.020 3132.090 326.320 ;
        RECT 3128.090 309.420 3134.840 311.020 ;
        RECT 3128.090 294.120 3132.090 309.420 ;
        RECT 3128.090 292.520 3134.840 294.120 ;
        RECT 3128.090 271.370 3132.090 292.520 ;
        RECT 3128.070 266.370 3228.670 271.370 ;
        RECT 2941.950 233.940 3248.340 235.940 ;
        RECT 234.180 232.940 3248.340 233.940 ;
        RECT 234.180 213.940 2956.980 232.940 ;
    END
  END vssd_core
  PIN vccd2_core
    PORT
      LAYER met4 ;
        RECT 306.910 1342.690 310.010 1379.380 ;
        RECT 306.910 1339.590 326.260 1342.690 ;
        RECT 323.160 1207.330 326.260 1339.590 ;
        RECT 220.980 1192.330 326.260 1207.330 ;
        RECT 974.410 1192.330 976.070 1207.320 ;
        RECT 1025.010 1192.330 1026.670 1207.320 ;
        RECT 220.980 1172.330 234.010 1192.330 ;
        RECT 323.160 1192.000 326.260 1192.330 ;
        RECT 3262.690 1191.330 3265.790 1379.380 ;
      LAYER via4 ;
        RECT 222.040 1173.135 232.820 1206.315 ;
        RECT 282.830 1193.695 316.010 1206.075 ;
        RECT 324.065 1205.650 325.245 1206.830 ;
        RECT 324.065 1204.050 325.245 1205.230 ;
        RECT 324.065 1202.450 325.245 1203.630 ;
        RECT 324.065 1200.850 325.245 1202.030 ;
        RECT 324.065 1199.250 325.245 1200.430 ;
        RECT 324.065 1197.650 325.245 1198.830 ;
        RECT 324.065 1196.050 325.245 1197.230 ;
        RECT 324.065 1194.450 325.245 1195.630 ;
        RECT 324.065 1192.850 325.245 1194.030 ;
        RECT 974.650 1205.685 975.830 1206.865 ;
        RECT 974.650 1204.085 975.830 1205.265 ;
        RECT 974.650 1202.485 975.830 1203.665 ;
        RECT 974.650 1200.885 975.830 1202.065 ;
        RECT 974.650 1199.285 975.830 1200.465 ;
        RECT 974.650 1197.685 975.830 1198.865 ;
        RECT 974.650 1196.085 975.830 1197.265 ;
        RECT 974.650 1194.485 975.830 1195.665 ;
        RECT 974.650 1192.885 975.830 1194.065 ;
        RECT 1025.250 1205.685 1026.430 1206.865 ;
        RECT 1025.250 1204.085 1026.430 1205.265 ;
        RECT 1025.250 1202.485 1026.430 1203.665 ;
        RECT 1025.250 1200.885 1026.430 1202.065 ;
        RECT 1025.250 1199.285 1026.430 1200.465 ;
        RECT 1025.250 1197.685 1026.430 1198.865 ;
        RECT 1025.250 1196.085 1026.430 1197.265 ;
        RECT 1025.250 1194.485 1026.430 1195.665 ;
        RECT 1025.250 1192.885 1026.430 1194.065 ;
        RECT 3263.605 1205.675 3264.785 1206.855 ;
        RECT 3263.605 1204.075 3264.785 1205.255 ;
        RECT 3263.605 1202.475 3264.785 1203.655 ;
        RECT 3263.605 1200.875 3264.785 1202.055 ;
        RECT 3263.605 1199.275 3264.785 1200.455 ;
        RECT 3263.605 1197.675 3264.785 1198.855 ;
        RECT 3263.605 1196.075 3264.785 1197.255 ;
        RECT 3263.605 1194.475 3264.785 1195.655 ;
        RECT 3263.605 1192.875 3264.785 1194.055 ;
      LAYER met5 ;
        RECT 221.270 1172.660 233.590 1206.790 ;
        RECT 281.390 1192.330 3266.530 1207.330 ;
    END
  END vccd2_core
  PIN vssd2_core
    PORT
      LAYER met4 ;
        RECT 302.110 1337.890 305.210 1374.610 ;
        RECT 302.110 1334.790 321.460 1337.890 ;
        RECT 318.360 1227.330 321.460 1334.790 ;
        RECT 204.920 1212.330 321.460 1227.330 ;
        RECT 995.310 1212.330 996.970 1227.320 ;
        RECT 1045.610 1212.340 1047.270 1227.330 ;
        RECT 204.920 1191.330 218.060 1212.330 ;
        RECT 318.360 1211.790 321.460 1212.330 ;
        RECT 3267.490 1211.810 3270.590 1374.580 ;
      LAYER via4 ;
        RECT 206.100 1191.985 216.880 1226.765 ;
        RECT 282.755 1213.525 315.935 1225.905 ;
        RECT 319.315 1225.670 320.495 1226.850 ;
        RECT 319.315 1224.070 320.495 1225.250 ;
        RECT 319.315 1222.470 320.495 1223.650 ;
        RECT 319.315 1220.870 320.495 1222.050 ;
        RECT 319.315 1219.270 320.495 1220.450 ;
        RECT 319.315 1217.670 320.495 1218.850 ;
        RECT 319.315 1216.070 320.495 1217.250 ;
        RECT 319.315 1214.470 320.495 1215.650 ;
        RECT 319.315 1212.870 320.495 1214.050 ;
        RECT 995.550 1225.685 996.730 1226.865 ;
        RECT 995.550 1224.085 996.730 1225.265 ;
        RECT 995.550 1222.485 996.730 1223.665 ;
        RECT 995.550 1220.885 996.730 1222.065 ;
        RECT 995.550 1219.285 996.730 1220.465 ;
        RECT 995.550 1217.685 996.730 1218.865 ;
        RECT 995.550 1216.085 996.730 1217.265 ;
        RECT 995.550 1214.485 996.730 1215.665 ;
        RECT 995.550 1212.885 996.730 1214.065 ;
        RECT 1045.850 1225.695 1047.030 1226.875 ;
        RECT 1045.850 1224.095 1047.030 1225.275 ;
        RECT 1045.850 1222.495 1047.030 1223.675 ;
        RECT 1045.850 1220.895 1047.030 1222.075 ;
        RECT 1045.850 1219.295 1047.030 1220.475 ;
        RECT 1045.850 1217.695 1047.030 1218.875 ;
        RECT 1045.850 1216.095 1047.030 1217.275 ;
        RECT 1045.850 1214.495 1047.030 1215.675 ;
        RECT 1045.850 1212.895 1047.030 1214.075 ;
        RECT 3268.395 1225.685 3269.575 1226.865 ;
        RECT 3268.395 1224.085 3269.575 1225.265 ;
        RECT 3268.395 1222.485 3269.575 1223.665 ;
        RECT 3268.395 1220.885 3269.575 1222.065 ;
        RECT 3268.395 1219.285 3269.575 1220.465 ;
        RECT 3268.395 1217.685 3269.575 1218.865 ;
        RECT 3268.395 1216.085 3269.575 1217.265 ;
        RECT 3268.395 1214.485 3269.575 1215.665 ;
        RECT 3268.395 1212.885 3269.575 1214.065 ;
      LAYER met5 ;
        RECT 205.330 1191.810 217.650 1226.940 ;
        RECT 281.390 1212.330 3271.110 1227.330 ;
    END
  END vssd2_core
  PIN vdda2_core
    PORT
      LAYER met3 ;
        RECT 199.620 2465.390 261.460 2489.290 ;
        RECT 199.620 2415.495 261.460 2439.395 ;
      LAYER via3 ;
        RECT 251.980 2466.295 260.300 2488.615 ;
        RECT 251.920 2416.345 260.240 2438.665 ;
      LAYER met4 ;
        RECT 250.970 4943.680 282.170 4946.740 ;
        RECT 250.860 2465.420 260.980 2489.370 ;
        RECT 250.990 2415.470 261.110 2439.420 ;
        RECT 250.930 1363.190 260.990 1367.190 ;
        RECT 250.930 1360.130 282.030 1363.190 ;
        RECT 287.710 1323.490 290.810 1360.210 ;
        RECT 287.710 1320.390 307.060 1323.490 ;
        RECT 303.960 1287.330 307.060 1320.390 ;
        RECT 250.850 1272.330 307.060 1287.330 ;
        RECT 303.960 1272.110 307.060 1272.330 ;
        RECT 1922.930 1272.260 1928.540 1287.350 ;
        RECT 1998.430 1272.260 2004.040 1287.350 ;
        RECT 3281.890 1271.930 3284.990 1360.180 ;
      LAYER via4 ;
        RECT 251.400 4944.625 252.580 4945.805 ;
        RECT 253.000 4944.625 254.180 4945.805 ;
        RECT 254.600 4944.625 255.780 4945.805 ;
        RECT 256.200 4944.625 257.380 4945.805 ;
        RECT 257.800 4944.625 258.980 4945.805 ;
        RECT 259.400 4944.625 260.580 4945.805 ;
        RECT 279.165 4944.650 280.345 4945.830 ;
        RECT 280.765 4944.650 281.945 4945.830 ;
        RECT 252.350 2466.465 259.930 2488.445 ;
        RECT 252.290 2416.515 259.870 2438.495 ;
        RECT 251.365 1360.680 260.545 1366.660 ;
        RECT 279.010 1360.285 281.790 1363.065 ;
        RECT 252.355 1273.845 259.935 1286.225 ;
        RECT 282.820 1273.540 301.600 1285.920 ;
        RECT 304.900 1285.630 306.080 1286.810 ;
        RECT 304.900 1284.030 306.080 1285.210 ;
        RECT 304.900 1282.430 306.080 1283.610 ;
        RECT 304.900 1280.830 306.080 1282.010 ;
        RECT 304.900 1279.230 306.080 1280.410 ;
        RECT 304.900 1277.630 306.080 1278.810 ;
        RECT 304.900 1276.030 306.080 1277.210 ;
        RECT 304.900 1274.430 306.080 1275.610 ;
        RECT 304.900 1272.830 306.080 1274.010 ;
        RECT 1923.575 1272.850 1927.955 1286.830 ;
        RECT 1999.075 1272.850 2003.455 1286.830 ;
        RECT 3282.805 1285.595 3283.985 1286.775 ;
        RECT 3282.805 1283.995 3283.985 1285.175 ;
        RECT 3282.805 1282.395 3283.985 1283.575 ;
        RECT 3282.805 1280.795 3283.985 1281.975 ;
        RECT 3282.805 1279.195 3283.985 1280.375 ;
        RECT 3282.805 1277.595 3283.985 1278.775 ;
        RECT 3282.805 1275.995 3283.985 1277.175 ;
        RECT 3282.805 1274.395 3283.985 1275.575 ;
        RECT 3282.805 1272.795 3283.985 1273.975 ;
      LAYER met5 ;
        RECT 250.990 1272.490 260.990 4952.330 ;
        RECT 278.880 4943.640 287.760 4946.740 ;
        RECT 278.770 1360.120 287.730 1363.220 ;
        RECT 281.850 1272.330 3285.380 1287.330 ;
    END
  END vdda2_core
  PIN vssa2_core
    PORT
      LAYER met3 ;
        RECT 199.260 4188.390 250.010 4212.290 ;
        RECT 199.260 4138.495 250.010 4162.395 ;
      LAYER via3 ;
        RECT 239.645 4189.150 248.365 4211.470 ;
        RECT 239.645 4139.490 248.365 4161.810 ;
      LAYER met4 ;
        RECT 238.980 4948.460 282.910 4951.550 ;
        RECT 238.960 4188.290 249.110 4212.310 ;
        RECT 238.960 4138.510 249.110 4162.530 ;
        RECT 238.960 1355.410 283.080 1358.440 ;
        RECT 238.960 1355.290 286.010 1355.410 ;
        RECT 238.960 1351.290 249.010 1355.290 ;
        RECT 282.860 1307.330 286.010 1355.290 ;
        RECT 238.850 1292.330 297.350 1307.330 ;
        RECT 1959.720 1292.340 1964.230 1307.250 ;
        RECT 2035.320 1292.340 2039.830 1307.250 ;
        RECT 3286.690 1291.950 3289.790 1355.410 ;
      LAYER via4 ;
        RECT 239.370 4949.445 240.550 4950.625 ;
        RECT 240.970 4949.445 242.150 4950.625 ;
        RECT 242.570 4949.445 243.750 4950.625 ;
        RECT 244.170 4949.445 245.350 4950.625 ;
        RECT 245.770 4949.445 246.950 4950.625 ;
        RECT 247.370 4949.445 248.550 4950.625 ;
        RECT 279.145 4949.450 280.325 4950.630 ;
        RECT 280.745 4949.450 281.925 4950.630 ;
        RECT 240.215 4189.320 247.795 4211.300 ;
        RECT 240.215 4139.660 247.795 4161.640 ;
        RECT 239.395 1351.915 248.575 1357.895 ;
        RECT 279.280 1355.470 282.060 1358.250 ;
        RECT 240.355 1293.845 247.935 1306.225 ;
        RECT 282.775 1293.540 296.755 1305.920 ;
        RECT 1960.585 1293.565 1963.365 1305.945 ;
        RECT 2036.185 1293.565 2038.965 1305.945 ;
        RECT 3287.615 1305.685 3288.795 1306.865 ;
        RECT 3287.615 1304.085 3288.795 1305.265 ;
        RECT 3287.615 1302.485 3288.795 1303.665 ;
        RECT 3287.615 1300.885 3288.795 1302.065 ;
        RECT 3287.615 1299.285 3288.795 1300.465 ;
        RECT 3287.615 1297.685 3288.795 1298.865 ;
        RECT 3287.615 1296.085 3288.795 1297.265 ;
        RECT 3287.615 1294.485 3288.795 1295.665 ;
        RECT 3287.615 1292.885 3288.795 1294.065 ;
      LAYER met5 ;
        RECT 238.990 1292.420 248.990 4952.330 ;
        RECT 278.880 4948.440 282.980 4951.540 ;
        RECT 278.770 1355.320 282.950 1358.420 ;
        RECT 281.850 1292.330 3290.450 1307.330 ;
    END
  END vssa2_core
  PIN vssd1_core
    PORT
      LAYER met3 ;
        RECT 565.910 4977.510 571.910 5152.410 ;
        RECT 822.910 4977.510 828.910 5152.410 ;
        RECT 1079.910 4977.510 1085.910 5152.410 ;
        RECT 1336.910 4977.510 1342.910 5152.410 ;
        RECT 1594.910 4977.510 1600.910 5152.410 ;
        RECT 1846.910 4977.510 1852.910 5152.410 ;
        RECT 2183.910 4977.510 2189.910 5152.410 ;
        RECT 2568.910 4977.510 2574.910 5152.410 ;
        RECT 2825.910 4977.510 2831.910 5152.410 ;
        RECT 36.180 4740.910 283.050 4741.910 ;
        RECT 36.180 4735.910 314.720 4740.910 ;
        RECT 277.160 4734.910 314.720 4735.910 ;
        RECT 36.180 4106.910 314.720 4112.910 ;
        RECT 36.180 3890.910 314.720 3896.910 ;
        RECT 36.180 3674.910 314.720 3680.910 ;
        RECT 36.180 3458.910 314.720 3464.910 ;
        RECT 36.180 3242.910 314.720 3248.910 ;
        RECT 36.180 3026.910 314.720 3032.910 ;
        RECT 36.180 2810.910 314.720 2816.910 ;
        RECT 36.180 2172.910 314.720 2178.910 ;
        RECT 36.180 1956.910 314.720 1962.910 ;
        RECT 36.180 1740.910 314.720 1746.910 ;
        RECT 36.180 1524.910 314.720 1530.910 ;
        RECT 36.180 1308.910 269.080 1314.910 ;
        RECT 36.180 1092.910 269.080 1098.910 ;
      LAYER via3 ;
        RECT 566.165 5148.530 571.685 5151.650 ;
        RECT 566.335 4978.065 571.455 4983.185 ;
        RECT 823.165 5148.530 828.685 5151.650 ;
        RECT 823.335 4978.065 828.455 4983.185 ;
        RECT 1080.165 5148.530 1085.685 5151.650 ;
        RECT 1080.335 4978.065 1085.455 4983.185 ;
        RECT 1337.165 5148.530 1342.685 5151.650 ;
        RECT 1337.335 4978.065 1342.455 4983.185 ;
        RECT 1595.165 5148.530 1600.685 5151.650 ;
        RECT 1595.335 4978.065 1600.455 4983.185 ;
        RECT 1847.165 5148.530 1852.685 5151.650 ;
        RECT 1847.335 4978.065 1852.455 4983.185 ;
        RECT 2184.165 5148.530 2189.685 5151.650 ;
        RECT 2184.335 4978.065 2189.455 4983.185 ;
        RECT 2569.165 5148.530 2574.685 5151.650 ;
        RECT 2569.335 4978.065 2574.455 4983.185 ;
        RECT 2826.165 5148.530 2831.685 5151.650 ;
        RECT 2826.335 4978.065 2831.455 4983.185 ;
        RECT 36.940 4736.165 40.060 4741.685 ;
        RECT 263.405 4736.335 268.525 4741.455 ;
        RECT 312.055 4735.085 314.375 4740.605 ;
        RECT 36.940 4107.165 40.060 4112.685 ;
        RECT 263.405 4107.335 268.525 4112.455 ;
        RECT 312.055 4107.085 314.375 4112.605 ;
        RECT 36.940 3891.165 40.060 3896.685 ;
        RECT 263.405 3891.335 268.525 3896.455 ;
        RECT 312.055 3891.085 314.375 3896.605 ;
        RECT 36.940 3675.165 40.060 3680.685 ;
        RECT 263.405 3675.335 268.525 3680.455 ;
        RECT 312.055 3675.085 314.375 3680.605 ;
        RECT 36.940 3459.165 40.060 3464.685 ;
        RECT 263.405 3459.335 268.525 3464.455 ;
        RECT 312.055 3459.085 314.375 3464.605 ;
        RECT 36.940 3243.165 40.060 3248.685 ;
        RECT 263.405 3243.335 268.525 3248.455 ;
        RECT 312.055 3243.085 314.375 3248.605 ;
        RECT 36.940 3027.165 40.060 3032.685 ;
        RECT 263.405 3027.335 268.525 3032.455 ;
        RECT 312.055 3027.085 314.375 3032.605 ;
        RECT 36.940 2811.165 40.060 2816.685 ;
        RECT 263.405 2811.335 268.525 2816.455 ;
        RECT 312.055 2811.085 314.375 2816.605 ;
        RECT 36.940 2173.165 40.060 2178.685 ;
        RECT 263.405 2173.335 268.525 2178.455 ;
        RECT 312.055 2173.085 314.375 2178.605 ;
        RECT 36.940 1957.165 40.060 1962.685 ;
        RECT 263.405 1957.335 268.525 1962.455 ;
        RECT 312.055 1957.085 314.375 1962.605 ;
        RECT 36.940 1741.165 40.060 1746.685 ;
        RECT 263.405 1741.335 268.525 1746.455 ;
        RECT 312.055 1741.085 314.375 1746.605 ;
        RECT 36.940 1525.165 40.060 1530.685 ;
        RECT 263.405 1525.335 268.525 1530.455 ;
        RECT 312.055 1525.085 314.375 1530.605 ;
        RECT 36.940 1309.165 40.060 1314.685 ;
        RECT 263.405 1309.335 268.525 1314.455 ;
        RECT 36.940 1093.165 40.060 1098.685 ;
        RECT 263.405 1093.335 268.525 1098.455 ;
      LAYER met4 ;
        RECT 505.380 5148.060 572.210 5152.060 ;
        RECT 762.380 5148.060 829.210 5152.060 ;
        RECT 1019.380 5148.060 1086.210 5152.060 ;
        RECT 1276.380 5148.060 1343.210 5152.060 ;
        RECT 1534.380 5148.060 1601.210 5152.060 ;
        RECT 1786.380 5148.060 1853.210 5152.060 ;
        RECT 2123.380 5148.060 2190.210 5152.060 ;
        RECT 2508.380 5148.060 2575.210 5152.060 ;
        RECT 2765.380 5148.060 2832.210 5152.060 ;
        RECT 565.870 4977.660 571.940 4983.690 ;
        RECT 822.870 4977.660 828.940 4983.690 ;
        RECT 1079.870 4977.660 1085.940 4983.690 ;
        RECT 1336.870 4977.660 1342.940 4983.690 ;
        RECT 1594.870 4977.660 1600.940 4983.690 ;
        RECT 1846.870 4977.660 1852.940 4983.690 ;
        RECT 2183.870 4977.660 2189.940 4983.690 ;
        RECT 2568.870 4977.660 2574.940 4983.690 ;
        RECT 2825.870 4977.660 2831.940 4983.690 ;
        RECT 3354.080 4983.460 3367.130 4983.480 ;
        RECT 3354.040 4977.460 3383.270 4983.460 ;
        RECT 3354.080 4951.000 3367.130 4977.460 ;
        RECT 262.980 4919.640 282.020 4922.740 ;
        RECT 36.530 4675.380 40.530 4742.210 ;
        RECT 262.900 4735.870 268.930 4741.940 ;
        RECT 311.910 4735.070 314.520 4740.620 ;
        RECT 36.530 4046.380 40.530 4113.210 ;
        RECT 262.900 4106.870 268.930 4112.940 ;
        RECT 311.910 4107.070 314.520 4112.620 ;
        RECT 36.530 3830.380 40.530 3897.210 ;
        RECT 262.900 3890.870 268.930 3896.940 ;
        RECT 311.910 3891.070 314.520 3896.620 ;
        RECT 36.530 3614.380 40.530 3681.210 ;
        RECT 262.900 3674.870 268.930 3680.940 ;
        RECT 311.910 3675.070 314.520 3680.620 ;
        RECT 36.530 3398.380 40.530 3465.210 ;
        RECT 262.900 3458.870 268.930 3464.940 ;
        RECT 311.910 3459.070 314.520 3464.620 ;
        RECT 36.530 3182.380 40.530 3249.210 ;
        RECT 262.900 3242.870 268.930 3248.940 ;
        RECT 311.910 3243.070 314.520 3248.620 ;
        RECT 36.530 2966.380 40.530 3033.210 ;
        RECT 262.900 3026.870 268.930 3032.940 ;
        RECT 311.910 3027.070 314.520 3032.620 ;
        RECT 36.530 2750.380 40.530 2817.210 ;
        RECT 262.900 2810.870 268.930 2816.940 ;
        RECT 311.910 2811.070 314.520 2816.620 ;
        RECT 36.530 2112.380 40.530 2179.210 ;
        RECT 262.900 2172.870 268.930 2178.940 ;
        RECT 311.910 2173.070 314.520 2178.620 ;
        RECT 36.530 1896.380 40.530 1963.210 ;
        RECT 262.900 1956.870 268.930 1962.940 ;
        RECT 311.910 1957.070 314.520 1962.620 ;
        RECT 36.530 1680.380 40.530 1747.210 ;
        RECT 262.900 1740.870 268.930 1746.940 ;
        RECT 311.910 1741.070 314.520 1746.620 ;
        RECT 36.530 1464.380 40.530 1531.210 ;
        RECT 262.900 1524.870 268.930 1530.940 ;
        RECT 311.910 1525.070 314.520 1530.620 ;
        RECT 262.910 1387.230 269.000 1390.230 ;
        RECT 262.910 1384.110 282.080 1387.230 ;
        RECT 311.710 1347.490 314.810 1384.170 ;
        RECT 311.710 1344.390 331.060 1347.490 ;
        RECT 36.530 1248.380 40.530 1315.210 ;
        RECT 262.900 1308.870 268.930 1314.940 ;
        RECT 262.890 1252.330 316.460 1267.330 ;
        RECT 327.960 1251.930 331.060 1344.390 ;
        RECT 1383.610 1252.350 1386.300 1267.360 ;
        RECT 1458.610 1252.350 1461.300 1267.360 ;
        RECT 1533.810 1252.350 1536.500 1267.360 ;
        RECT 1609.410 1252.350 1612.100 1267.360 ;
        RECT 3257.890 1251.960 3260.990 1384.220 ;
        RECT 36.530 1032.380 40.530 1099.210 ;
        RECT 262.900 1092.870 268.930 1098.940 ;
      LAYER via4 ;
        RECT 505.795 5150.285 506.975 5151.465 ;
        RECT 522.710 5150.285 523.890 5151.465 ;
        RECT 539.590 5150.275 540.770 5151.455 ;
        RECT 505.795 5148.685 506.975 5149.865 ;
        RECT 522.710 5148.685 523.890 5149.865 ;
        RECT 539.590 5148.675 540.770 5149.855 ;
        RECT 762.795 5150.285 763.975 5151.465 ;
        RECT 779.710 5150.285 780.890 5151.465 ;
        RECT 796.590 5150.275 797.770 5151.455 ;
        RECT 762.795 5148.685 763.975 5149.865 ;
        RECT 779.710 5148.685 780.890 5149.865 ;
        RECT 796.590 5148.675 797.770 5149.855 ;
        RECT 1019.795 5150.285 1020.975 5151.465 ;
        RECT 1036.710 5150.285 1037.890 5151.465 ;
        RECT 1053.590 5150.275 1054.770 5151.455 ;
        RECT 1019.795 5148.685 1020.975 5149.865 ;
        RECT 1036.710 5148.685 1037.890 5149.865 ;
        RECT 1053.590 5148.675 1054.770 5149.855 ;
        RECT 1276.795 5150.285 1277.975 5151.465 ;
        RECT 1293.710 5150.285 1294.890 5151.465 ;
        RECT 1310.590 5150.275 1311.770 5151.455 ;
        RECT 1276.795 5148.685 1277.975 5149.865 ;
        RECT 1293.710 5148.685 1294.890 5149.865 ;
        RECT 1310.590 5148.675 1311.770 5149.855 ;
        RECT 1534.795 5150.285 1535.975 5151.465 ;
        RECT 1551.710 5150.285 1552.890 5151.465 ;
        RECT 1568.590 5150.275 1569.770 5151.455 ;
        RECT 1534.795 5148.685 1535.975 5149.865 ;
        RECT 1551.710 5148.685 1552.890 5149.865 ;
        RECT 1568.590 5148.675 1569.770 5149.855 ;
        RECT 1786.795 5150.285 1787.975 5151.465 ;
        RECT 1803.710 5150.285 1804.890 5151.465 ;
        RECT 1820.590 5150.275 1821.770 5151.455 ;
        RECT 1786.795 5148.685 1787.975 5149.865 ;
        RECT 1803.710 5148.685 1804.890 5149.865 ;
        RECT 1820.590 5148.675 1821.770 5149.855 ;
        RECT 2123.795 5150.285 2124.975 5151.465 ;
        RECT 2140.710 5150.285 2141.890 5151.465 ;
        RECT 2157.590 5150.275 2158.770 5151.455 ;
        RECT 2123.795 5148.685 2124.975 5149.865 ;
        RECT 2140.710 5148.685 2141.890 5149.865 ;
        RECT 2157.590 5148.675 2158.770 5149.855 ;
        RECT 2508.795 5150.285 2509.975 5151.465 ;
        RECT 2525.710 5150.285 2526.890 5151.465 ;
        RECT 2542.590 5150.275 2543.770 5151.455 ;
        RECT 2508.795 5148.685 2509.975 5149.865 ;
        RECT 2525.710 5148.685 2526.890 5149.865 ;
        RECT 2542.590 5148.675 2543.770 5149.855 ;
        RECT 2765.795 5150.285 2766.975 5151.465 ;
        RECT 2782.710 5150.285 2783.890 5151.465 ;
        RECT 2799.590 5150.275 2800.770 5151.455 ;
        RECT 2765.795 5148.685 2766.975 5149.865 ;
        RECT 2782.710 5148.685 2783.890 5149.865 ;
        RECT 2799.590 5148.675 2800.770 5149.855 ;
        RECT 566.705 4978.435 571.085 4982.815 ;
        RECT 823.705 4978.435 828.085 4982.815 ;
        RECT 1080.705 4978.435 1085.085 4982.815 ;
        RECT 1337.705 4978.435 1342.085 4982.815 ;
        RECT 1595.705 4978.435 1600.085 4982.815 ;
        RECT 1847.705 4978.435 1852.085 4982.815 ;
        RECT 2184.705 4978.435 2189.085 4982.815 ;
        RECT 2569.705 4978.435 2574.085 4982.815 ;
        RECT 2826.705 4978.435 2831.085 4982.815 ;
        RECT 3355.180 4978.340 3381.960 4982.720 ;
        RECT 3355.210 4951.820 3365.990 4962.600 ;
        RECT 263.795 4920.605 264.975 4921.785 ;
        RECT 265.395 4920.605 266.575 4921.785 ;
        RECT 266.995 4920.605 268.175 4921.785 ;
        RECT 279.055 4919.805 281.835 4922.585 ;
        RECT 263.775 4736.705 268.155 4741.085 ;
        RECT 37.135 4709.595 38.315 4710.775 ;
        RECT 38.735 4709.595 39.915 4710.775 ;
        RECT 37.140 4692.695 38.320 4693.875 ;
        RECT 38.740 4692.695 39.920 4693.875 ;
        RECT 37.125 4675.795 38.305 4676.975 ;
        RECT 38.725 4675.795 39.905 4676.975 ;
        RECT 263.775 4107.705 268.155 4112.085 ;
        RECT 37.135 4080.595 38.315 4081.775 ;
        RECT 38.735 4080.595 39.915 4081.775 ;
        RECT 37.140 4063.695 38.320 4064.875 ;
        RECT 38.740 4063.695 39.920 4064.875 ;
        RECT 37.125 4046.795 38.305 4047.975 ;
        RECT 38.725 4046.795 39.905 4047.975 ;
        RECT 263.775 3891.705 268.155 3896.085 ;
        RECT 37.135 3864.595 38.315 3865.775 ;
        RECT 38.735 3864.595 39.915 3865.775 ;
        RECT 37.140 3847.695 38.320 3848.875 ;
        RECT 38.740 3847.695 39.920 3848.875 ;
        RECT 37.125 3830.795 38.305 3831.975 ;
        RECT 38.725 3830.795 39.905 3831.975 ;
        RECT 263.775 3675.705 268.155 3680.085 ;
        RECT 37.135 3648.595 38.315 3649.775 ;
        RECT 38.735 3648.595 39.915 3649.775 ;
        RECT 37.140 3631.695 38.320 3632.875 ;
        RECT 38.740 3631.695 39.920 3632.875 ;
        RECT 37.125 3614.795 38.305 3615.975 ;
        RECT 38.725 3614.795 39.905 3615.975 ;
        RECT 263.775 3459.705 268.155 3464.085 ;
        RECT 37.135 3432.595 38.315 3433.775 ;
        RECT 38.735 3432.595 39.915 3433.775 ;
        RECT 37.140 3415.695 38.320 3416.875 ;
        RECT 38.740 3415.695 39.920 3416.875 ;
        RECT 37.125 3398.795 38.305 3399.975 ;
        RECT 38.725 3398.795 39.905 3399.975 ;
        RECT 263.775 3243.705 268.155 3248.085 ;
        RECT 37.135 3216.595 38.315 3217.775 ;
        RECT 38.735 3216.595 39.915 3217.775 ;
        RECT 37.140 3199.695 38.320 3200.875 ;
        RECT 38.740 3199.695 39.920 3200.875 ;
        RECT 37.125 3182.795 38.305 3183.975 ;
        RECT 38.725 3182.795 39.905 3183.975 ;
        RECT 263.775 3027.705 268.155 3032.085 ;
        RECT 37.135 3000.595 38.315 3001.775 ;
        RECT 38.735 3000.595 39.915 3001.775 ;
        RECT 37.140 2983.695 38.320 2984.875 ;
        RECT 38.740 2983.695 39.920 2984.875 ;
        RECT 37.125 2966.795 38.305 2967.975 ;
        RECT 38.725 2966.795 39.905 2967.975 ;
        RECT 263.775 2811.705 268.155 2816.085 ;
        RECT 37.135 2784.595 38.315 2785.775 ;
        RECT 38.735 2784.595 39.915 2785.775 ;
        RECT 37.140 2767.695 38.320 2768.875 ;
        RECT 38.740 2767.695 39.920 2768.875 ;
        RECT 37.125 2750.795 38.305 2751.975 ;
        RECT 38.725 2750.795 39.905 2751.975 ;
        RECT 263.775 2173.705 268.155 2178.085 ;
        RECT 37.135 2146.595 38.315 2147.775 ;
        RECT 38.735 2146.595 39.915 2147.775 ;
        RECT 37.140 2129.695 38.320 2130.875 ;
        RECT 38.740 2129.695 39.920 2130.875 ;
        RECT 37.125 2112.795 38.305 2113.975 ;
        RECT 38.725 2112.795 39.905 2113.975 ;
        RECT 263.775 1957.705 268.155 1962.085 ;
        RECT 37.135 1930.595 38.315 1931.775 ;
        RECT 38.735 1930.595 39.915 1931.775 ;
        RECT 37.140 1913.695 38.320 1914.875 ;
        RECT 38.740 1913.695 39.920 1914.875 ;
        RECT 37.125 1896.795 38.305 1897.975 ;
        RECT 38.725 1896.795 39.905 1897.975 ;
        RECT 263.775 1741.705 268.155 1746.085 ;
        RECT 37.135 1714.595 38.315 1715.775 ;
        RECT 38.735 1714.595 39.915 1715.775 ;
        RECT 37.140 1697.695 38.320 1698.875 ;
        RECT 38.740 1697.695 39.920 1698.875 ;
        RECT 37.125 1680.795 38.305 1681.975 ;
        RECT 38.725 1680.795 39.905 1681.975 ;
        RECT 263.775 1525.705 268.155 1530.085 ;
        RECT 37.135 1498.595 38.315 1499.775 ;
        RECT 38.735 1498.595 39.915 1499.775 ;
        RECT 37.140 1481.695 38.320 1482.875 ;
        RECT 38.740 1481.695 39.920 1482.875 ;
        RECT 37.125 1464.795 38.305 1465.975 ;
        RECT 38.725 1464.795 39.905 1465.975 ;
        RECT 263.765 1385.050 268.145 1389.430 ;
        RECT 279.030 1384.295 281.810 1387.075 ;
        RECT 263.775 1309.705 268.155 1314.085 ;
        RECT 37.135 1282.595 38.315 1283.775 ;
        RECT 38.735 1282.595 39.915 1283.775 ;
        RECT 37.140 1265.695 38.320 1266.875 ;
        RECT 38.740 1265.695 39.920 1266.875 ;
        RECT 263.810 1252.860 268.190 1266.840 ;
        RECT 281.160 1252.870 315.940 1266.850 ;
        RECT 328.875 1265.610 330.055 1266.790 ;
        RECT 328.875 1264.010 330.055 1265.190 ;
        RECT 328.875 1262.410 330.055 1263.590 ;
        RECT 328.875 1260.810 330.055 1261.990 ;
        RECT 328.875 1259.210 330.055 1260.390 ;
        RECT 328.875 1257.610 330.055 1258.790 ;
        RECT 328.875 1256.010 330.055 1257.190 ;
        RECT 328.875 1254.410 330.055 1255.590 ;
        RECT 328.875 1252.810 330.055 1253.990 ;
        RECT 1384.135 1265.700 1385.315 1266.880 ;
        RECT 1384.135 1264.100 1385.315 1265.280 ;
        RECT 1384.135 1262.500 1385.315 1263.680 ;
        RECT 1384.135 1260.900 1385.315 1262.080 ;
        RECT 1384.135 1259.300 1385.315 1260.480 ;
        RECT 1384.135 1257.700 1385.315 1258.880 ;
        RECT 1384.135 1256.100 1385.315 1257.280 ;
        RECT 1384.135 1254.500 1385.315 1255.680 ;
        RECT 1384.135 1252.900 1385.315 1254.080 ;
        RECT 1459.135 1265.700 1460.315 1266.880 ;
        RECT 1459.135 1264.100 1460.315 1265.280 ;
        RECT 1459.135 1262.500 1460.315 1263.680 ;
        RECT 1459.135 1260.900 1460.315 1262.080 ;
        RECT 1459.135 1259.300 1460.315 1260.480 ;
        RECT 1459.135 1257.700 1460.315 1258.880 ;
        RECT 1459.135 1256.100 1460.315 1257.280 ;
        RECT 1459.135 1254.500 1460.315 1255.680 ;
        RECT 1459.135 1252.900 1460.315 1254.080 ;
        RECT 1534.335 1265.700 1535.515 1266.880 ;
        RECT 1534.335 1264.100 1535.515 1265.280 ;
        RECT 1534.335 1262.500 1535.515 1263.680 ;
        RECT 1534.335 1260.900 1535.515 1262.080 ;
        RECT 1534.335 1259.300 1535.515 1260.480 ;
        RECT 1534.335 1257.700 1535.515 1258.880 ;
        RECT 1534.335 1256.100 1535.515 1257.280 ;
        RECT 1534.335 1254.500 1535.515 1255.680 ;
        RECT 1534.335 1252.900 1535.515 1254.080 ;
        RECT 1609.935 1265.700 1611.115 1266.880 ;
        RECT 1609.935 1264.100 1611.115 1265.280 ;
        RECT 1609.935 1262.500 1611.115 1263.680 ;
        RECT 1609.935 1260.900 1611.115 1262.080 ;
        RECT 1609.935 1259.300 1611.115 1260.480 ;
        RECT 1609.935 1257.700 1611.115 1258.880 ;
        RECT 1609.935 1256.100 1611.115 1257.280 ;
        RECT 1609.935 1254.500 1611.115 1255.680 ;
        RECT 1609.935 1252.900 1611.115 1254.080 ;
        RECT 3258.070 1252.805 3260.850 1266.785 ;
        RECT 37.125 1248.795 38.305 1249.975 ;
        RECT 38.725 1248.795 39.905 1249.975 ;
        RECT 263.775 1093.705 268.155 1098.085 ;
        RECT 37.135 1066.595 38.315 1067.775 ;
        RECT 38.735 1066.595 39.915 1067.775 ;
        RECT 37.140 1049.695 38.320 1050.875 ;
        RECT 38.740 1049.695 39.920 1050.875 ;
        RECT 37.125 1032.795 38.305 1033.975 ;
        RECT 38.725 1032.795 39.905 1033.975 ;
      LAYER met5 ;
        RECT 505.510 5147.980 507.260 5152.140 ;
        RECT 505.590 5145.520 507.190 5147.980 ;
        RECT 522.400 5147.940 524.130 5152.320 ;
        RECT 539.340 5147.970 541.070 5152.350 ;
        RECT 762.510 5147.980 764.260 5152.140 ;
        RECT 522.490 5145.680 524.090 5147.940 ;
        RECT 539.390 5145.680 540.990 5147.970 ;
        RECT 762.590 5145.520 764.190 5147.980 ;
        RECT 779.400 5147.940 781.130 5152.320 ;
        RECT 796.340 5147.970 798.070 5152.350 ;
        RECT 1019.510 5147.980 1021.260 5152.140 ;
        RECT 779.490 5145.680 781.090 5147.940 ;
        RECT 796.390 5145.680 797.990 5147.970 ;
        RECT 1019.590 5145.520 1021.190 5147.980 ;
        RECT 1036.400 5147.940 1038.130 5152.320 ;
        RECT 1053.340 5147.970 1055.070 5152.350 ;
        RECT 1276.510 5147.980 1278.260 5152.140 ;
        RECT 1036.490 5145.680 1038.090 5147.940 ;
        RECT 1053.390 5145.680 1054.990 5147.970 ;
        RECT 1276.590 5145.520 1278.190 5147.980 ;
        RECT 1293.400 5147.940 1295.130 5152.320 ;
        RECT 1310.340 5147.970 1312.070 5152.350 ;
        RECT 1534.510 5147.980 1536.260 5152.140 ;
        RECT 1293.490 5145.680 1295.090 5147.940 ;
        RECT 1310.390 5145.680 1311.990 5147.970 ;
        RECT 1534.590 5145.520 1536.190 5147.980 ;
        RECT 1551.400 5147.940 1553.130 5152.320 ;
        RECT 1568.340 5147.970 1570.070 5152.350 ;
        RECT 1786.510 5147.980 1788.260 5152.140 ;
        RECT 1551.490 5145.680 1553.090 5147.940 ;
        RECT 1568.390 5145.680 1569.990 5147.970 ;
        RECT 1786.590 5145.520 1788.190 5147.980 ;
        RECT 1803.400 5147.940 1805.130 5152.320 ;
        RECT 1820.340 5147.970 1822.070 5152.350 ;
        RECT 2123.510 5147.980 2125.260 5152.140 ;
        RECT 1803.490 5145.680 1805.090 5147.940 ;
        RECT 1820.390 5145.680 1821.990 5147.970 ;
        RECT 2123.590 5145.520 2125.190 5147.980 ;
        RECT 2140.400 5147.940 2142.130 5152.320 ;
        RECT 2157.340 5147.970 2159.070 5152.350 ;
        RECT 2508.510 5147.980 2510.260 5152.140 ;
        RECT 2140.490 5145.680 2142.090 5147.940 ;
        RECT 2157.390 5145.680 2158.990 5147.970 ;
        RECT 2508.590 5145.520 2510.190 5147.980 ;
        RECT 2525.400 5147.940 2527.130 5152.320 ;
        RECT 2542.340 5147.970 2544.070 5152.350 ;
        RECT 2765.510 5147.980 2767.260 5152.140 ;
        RECT 2525.490 5145.680 2527.090 5147.940 ;
        RECT 2542.390 5145.680 2543.990 5147.970 ;
        RECT 2765.590 5145.520 2767.190 5147.980 ;
        RECT 2782.400 5147.940 2784.130 5152.320 ;
        RECT 2799.340 5147.970 2801.070 5152.350 ;
        RECT 2782.490 5145.680 2784.090 5147.940 ;
        RECT 2799.390 5145.680 2800.990 5147.970 ;
        RECT 262.990 4977.510 3383.300 4983.510 ;
        RECT 36.395 4710.990 40.590 4711.095 ;
        RECT 36.300 4709.390 42.910 4710.990 ;
        RECT 36.395 4709.290 40.590 4709.390 ;
        RECT 36.485 4694.090 40.680 4694.205 ;
        RECT 36.330 4692.490 42.910 4694.090 ;
        RECT 36.485 4692.400 40.680 4692.490 ;
        RECT 36.385 4677.190 40.860 4677.265 ;
        RECT 36.385 4675.590 43.070 4677.190 ;
        RECT 36.385 4675.510 40.860 4675.590 ;
        RECT 36.395 4081.990 40.590 4082.095 ;
        RECT 36.300 4080.390 42.910 4081.990 ;
        RECT 36.395 4080.290 40.590 4080.390 ;
        RECT 36.485 4065.090 40.680 4065.205 ;
        RECT 36.330 4063.490 42.910 4065.090 ;
        RECT 36.485 4063.400 40.680 4063.490 ;
        RECT 36.385 4048.190 40.860 4048.265 ;
        RECT 36.385 4046.590 43.070 4048.190 ;
        RECT 36.385 4046.510 40.860 4046.590 ;
        RECT 36.395 3865.990 40.590 3866.095 ;
        RECT 36.300 3864.390 42.910 3865.990 ;
        RECT 36.395 3864.290 40.590 3864.390 ;
        RECT 36.485 3849.090 40.680 3849.205 ;
        RECT 36.330 3847.490 42.910 3849.090 ;
        RECT 36.485 3847.400 40.680 3847.490 ;
        RECT 36.385 3832.190 40.860 3832.265 ;
        RECT 36.385 3830.590 43.070 3832.190 ;
        RECT 36.385 3830.510 40.860 3830.590 ;
        RECT 36.395 3649.990 40.590 3650.095 ;
        RECT 36.300 3648.390 42.910 3649.990 ;
        RECT 36.395 3648.290 40.590 3648.390 ;
        RECT 36.485 3633.090 40.680 3633.205 ;
        RECT 36.330 3631.490 42.910 3633.090 ;
        RECT 36.485 3631.400 40.680 3631.490 ;
        RECT 36.385 3616.190 40.860 3616.265 ;
        RECT 36.385 3614.590 43.070 3616.190 ;
        RECT 36.385 3614.510 40.860 3614.590 ;
        RECT 36.395 3433.990 40.590 3434.095 ;
        RECT 36.300 3432.390 42.910 3433.990 ;
        RECT 36.395 3432.290 40.590 3432.390 ;
        RECT 36.485 3417.090 40.680 3417.205 ;
        RECT 36.330 3415.490 42.910 3417.090 ;
        RECT 36.485 3415.400 40.680 3415.490 ;
        RECT 36.385 3400.190 40.860 3400.265 ;
        RECT 36.385 3398.590 43.070 3400.190 ;
        RECT 36.385 3398.510 40.860 3398.590 ;
        RECT 36.395 3217.990 40.590 3218.095 ;
        RECT 36.300 3216.390 42.910 3217.990 ;
        RECT 36.395 3216.290 40.590 3216.390 ;
        RECT 36.485 3201.090 40.680 3201.205 ;
        RECT 36.330 3199.490 42.910 3201.090 ;
        RECT 36.485 3199.400 40.680 3199.490 ;
        RECT 36.385 3184.190 40.860 3184.265 ;
        RECT 36.385 3182.590 43.070 3184.190 ;
        RECT 36.385 3182.510 40.860 3182.590 ;
        RECT 36.395 3001.990 40.590 3002.095 ;
        RECT 36.300 3000.390 42.910 3001.990 ;
        RECT 36.395 3000.290 40.590 3000.390 ;
        RECT 36.485 2985.090 40.680 2985.205 ;
        RECT 36.330 2983.490 42.910 2985.090 ;
        RECT 36.485 2983.400 40.680 2983.490 ;
        RECT 36.385 2968.190 40.860 2968.265 ;
        RECT 36.385 2966.590 43.070 2968.190 ;
        RECT 36.385 2966.510 40.860 2966.590 ;
        RECT 36.395 2785.990 40.590 2786.095 ;
        RECT 36.300 2784.390 42.910 2785.990 ;
        RECT 36.395 2784.290 40.590 2784.390 ;
        RECT 36.485 2769.090 40.680 2769.205 ;
        RECT 36.330 2767.490 42.910 2769.090 ;
        RECT 36.485 2767.400 40.680 2767.490 ;
        RECT 36.385 2752.190 40.860 2752.265 ;
        RECT 36.385 2750.590 43.070 2752.190 ;
        RECT 36.385 2750.510 40.860 2750.590 ;
        RECT 36.395 2147.990 40.590 2148.095 ;
        RECT 36.300 2146.390 42.910 2147.990 ;
        RECT 36.395 2146.290 40.590 2146.390 ;
        RECT 36.485 2131.090 40.680 2131.205 ;
        RECT 36.330 2129.490 42.910 2131.090 ;
        RECT 36.485 2129.400 40.680 2129.490 ;
        RECT 36.385 2114.190 40.860 2114.265 ;
        RECT 36.385 2112.590 43.070 2114.190 ;
        RECT 36.385 2112.510 40.860 2112.590 ;
        RECT 36.395 1931.990 40.590 1932.095 ;
        RECT 36.300 1930.390 42.910 1931.990 ;
        RECT 36.395 1930.290 40.590 1930.390 ;
        RECT 36.485 1915.090 40.680 1915.205 ;
        RECT 36.330 1913.490 42.910 1915.090 ;
        RECT 36.485 1913.400 40.680 1913.490 ;
        RECT 36.385 1898.190 40.860 1898.265 ;
        RECT 36.385 1896.590 43.070 1898.190 ;
        RECT 36.385 1896.510 40.860 1896.590 ;
        RECT 36.395 1715.990 40.590 1716.095 ;
        RECT 36.300 1714.390 42.910 1715.990 ;
        RECT 36.395 1714.290 40.590 1714.390 ;
        RECT 36.485 1699.090 40.680 1699.205 ;
        RECT 36.330 1697.490 42.910 1699.090 ;
        RECT 36.485 1697.400 40.680 1697.490 ;
        RECT 36.385 1682.190 40.860 1682.265 ;
        RECT 36.385 1680.590 43.070 1682.190 ;
        RECT 36.385 1680.510 40.860 1680.590 ;
        RECT 36.395 1499.990 40.590 1500.095 ;
        RECT 36.300 1498.390 42.910 1499.990 ;
        RECT 36.395 1498.290 40.590 1498.390 ;
        RECT 36.485 1483.090 40.680 1483.205 ;
        RECT 36.330 1481.490 42.910 1483.090 ;
        RECT 36.485 1481.400 40.680 1481.490 ;
        RECT 36.385 1466.190 40.860 1466.265 ;
        RECT 36.385 1464.590 43.070 1466.190 ;
        RECT 36.385 1464.510 40.860 1464.590 ;
        RECT 36.395 1283.990 40.590 1284.095 ;
        RECT 36.300 1282.390 42.910 1283.990 ;
        RECT 36.395 1282.290 40.590 1282.390 ;
        RECT 36.485 1267.090 40.680 1267.205 ;
        RECT 36.330 1265.490 42.910 1267.090 ;
        RECT 36.485 1265.400 40.680 1265.490 ;
        RECT 36.385 1250.190 40.860 1250.265 ;
        RECT 36.385 1248.590 43.070 1250.190 ;
        RECT 36.385 1248.510 40.860 1248.590 ;
        RECT 262.990 1088.710 268.990 4977.510 ;
        RECT 3354.880 4951.770 3366.320 4962.650 ;
        RECT 278.880 4919.640 311.790 4922.740 ;
        RECT 278.770 1384.120 311.760 1387.220 ;
        RECT 280.630 1252.330 3354.930 1267.330 ;
        RECT 36.395 1067.990 40.590 1068.095 ;
        RECT 36.300 1066.390 42.910 1067.990 ;
        RECT 36.395 1066.290 40.590 1066.390 ;
        RECT 36.485 1051.090 40.680 1051.205 ;
        RECT 36.330 1049.490 42.910 1051.090 ;
        RECT 36.485 1049.400 40.680 1049.490 ;
        RECT 36.385 1034.190 40.860 1034.265 ;
        RECT 36.385 1032.590 43.070 1034.190 ;
        RECT 36.385 1032.510 40.860 1032.590 ;
    END
  END vssd1_core
  PIN vccd1_core
    PORT
      LAYER met3 ;
        RECT 573.910 4969.290 579.910 5158.480 ;
        RECT 830.910 4969.290 836.910 5158.480 ;
        RECT 1087.910 4969.290 1093.910 5158.480 ;
        RECT 1344.910 4969.290 1350.910 5158.480 ;
        RECT 1602.910 4969.290 1608.910 5158.480 ;
        RECT 1854.910 4969.290 1860.910 5158.480 ;
        RECT 2191.910 4969.290 2197.910 5158.480 ;
        RECT 2576.910 4969.290 2582.910 5158.480 ;
        RECT 2833.910 4969.290 2839.910 5158.480 ;
        RECT 30.110 4748.410 291.090 4749.910 ;
        RECT 30.110 4743.910 319.610 4748.410 ;
        RECT 285.190 4742.410 319.610 4743.910 ;
        RECT 30.110 4114.910 319.610 4120.910 ;
        RECT 280.390 3904.910 319.610 3910.910 ;
        RECT 30.110 3898.910 286.850 3904.910 ;
        RECT 30.110 3682.910 319.610 3688.910 ;
        RECT 30.110 3466.910 319.610 3472.910 ;
        RECT 30.110 3250.910 319.610 3256.910 ;
        RECT 30.110 3034.910 319.610 3040.910 ;
        RECT 30.110 2818.910 319.610 2824.910 ;
        RECT 30.110 2180.910 319.610 2186.910 ;
        RECT 30.110 1964.910 319.610 1970.910 ;
        RECT 279.840 1754.910 319.610 1758.910 ;
        RECT 30.110 1752.910 319.610 1754.910 ;
        RECT 30.110 1748.910 286.320 1752.910 ;
        RECT 30.110 1532.910 319.610 1538.910 ;
        RECT 30.110 1316.910 277.300 1322.910 ;
        RECT 30.110 1100.910 277.300 1106.910 ;
      LAYER via3 ;
        RECT 574.145 5154.520 579.665 5157.640 ;
        RECT 574.425 4970.095 579.545 4975.215 ;
        RECT 831.145 5154.520 836.665 5157.640 ;
        RECT 831.425 4970.095 836.545 4975.215 ;
        RECT 1088.145 5154.520 1093.665 5157.640 ;
        RECT 1088.425 4970.095 1093.545 4975.215 ;
        RECT 1345.145 5154.520 1350.665 5157.640 ;
        RECT 1345.425 4970.095 1350.545 4975.215 ;
        RECT 1603.145 5154.520 1608.665 5157.640 ;
        RECT 1603.425 4970.095 1608.545 4975.215 ;
        RECT 1855.145 5154.520 1860.665 5157.640 ;
        RECT 1855.425 4970.095 1860.545 4975.215 ;
        RECT 2192.145 5154.520 2197.665 5157.640 ;
        RECT 2192.425 4970.095 2197.545 4975.215 ;
        RECT 2577.145 5154.520 2582.665 5157.640 ;
        RECT 2577.425 4970.095 2582.545 4975.215 ;
        RECT 2834.145 5154.520 2839.665 5157.640 ;
        RECT 2834.425 4970.095 2839.545 4975.215 ;
        RECT 30.950 4744.145 34.070 4749.665 ;
        RECT 271.375 4744.425 276.495 4749.545 ;
        RECT 316.895 4742.625 319.215 4748.145 ;
        RECT 30.950 4115.145 34.070 4120.665 ;
        RECT 271.375 4115.425 276.495 4120.545 ;
        RECT 316.895 4115.125 319.215 4120.645 ;
        RECT 316.895 3905.125 319.215 3910.645 ;
        RECT 30.950 3899.145 34.070 3904.665 ;
        RECT 271.375 3899.425 276.495 3904.545 ;
        RECT 30.950 3683.145 34.070 3688.665 ;
        RECT 271.375 3683.425 276.495 3688.545 ;
        RECT 316.895 3683.125 319.215 3688.645 ;
        RECT 30.950 3467.145 34.070 3472.665 ;
        RECT 271.375 3467.425 276.495 3472.545 ;
        RECT 316.895 3467.125 319.215 3472.645 ;
        RECT 30.950 3251.145 34.070 3256.665 ;
        RECT 271.375 3251.425 276.495 3256.545 ;
        RECT 316.895 3251.125 319.215 3256.645 ;
        RECT 30.950 3035.145 34.070 3040.665 ;
        RECT 271.375 3035.425 276.495 3040.545 ;
        RECT 316.895 3035.125 319.215 3040.645 ;
        RECT 30.950 2819.145 34.070 2824.665 ;
        RECT 271.375 2819.425 276.495 2824.545 ;
        RECT 316.895 2819.125 319.215 2824.645 ;
        RECT 30.950 2181.145 34.070 2186.665 ;
        RECT 271.375 2181.425 276.495 2186.545 ;
        RECT 316.895 2181.125 319.215 2186.645 ;
        RECT 30.950 1965.145 34.070 1970.665 ;
        RECT 271.375 1965.425 276.495 1970.545 ;
        RECT 316.895 1965.125 319.215 1970.645 ;
        RECT 30.950 1749.145 34.070 1754.665 ;
        RECT 271.375 1749.425 276.495 1754.545 ;
        RECT 316.895 1753.125 319.215 1758.645 ;
        RECT 30.950 1533.145 34.070 1538.665 ;
        RECT 271.375 1533.425 276.495 1538.545 ;
        RECT 316.895 1533.125 319.215 1538.645 ;
        RECT 30.950 1317.145 34.070 1322.665 ;
        RECT 271.375 1317.425 276.495 1322.545 ;
        RECT 30.950 1101.145 34.070 1106.665 ;
        RECT 271.375 1101.425 276.495 1106.545 ;
      LAYER met4 ;
        RECT 496.730 5154.060 580.350 5158.060 ;
        RECT 753.730 5154.060 837.350 5158.060 ;
        RECT 1010.730 5154.060 1094.350 5158.060 ;
        RECT 1267.730 5154.060 1351.350 5158.060 ;
        RECT 1525.730 5154.060 1609.350 5158.060 ;
        RECT 1777.730 5154.060 1861.350 5158.060 ;
        RECT 2114.730 5154.060 2198.350 5158.060 ;
        RECT 2499.730 5154.060 2583.350 5158.060 ;
        RECT 2756.730 5154.060 2840.350 5158.060 ;
        RECT 573.870 4969.640 579.940 4975.670 ;
        RECT 830.870 4969.640 836.940 4975.670 ;
        RECT 1087.870 4969.640 1093.940 4975.670 ;
        RECT 1344.870 4969.640 1350.940 4975.670 ;
        RECT 1602.870 4969.640 1608.940 4975.670 ;
        RECT 1854.870 4969.640 1860.940 4975.670 ;
        RECT 2191.870 4969.640 2197.940 4975.670 ;
        RECT 2576.870 4969.640 2582.940 4975.670 ;
        RECT 2833.870 4969.640 2839.940 4975.670 ;
        RECT 30.530 4666.730 34.530 4750.350 ;
        RECT 270.920 4743.870 276.950 4749.940 ;
        RECT 316.750 4742.610 319.360 4748.160 ;
        RECT 30.530 4037.730 34.530 4121.350 ;
        RECT 270.920 4114.870 276.950 4120.940 ;
        RECT 316.750 4115.110 319.360 4120.660 ;
        RECT 30.530 3821.730 34.530 3905.350 ;
        RECT 316.750 3905.110 319.360 3910.660 ;
        RECT 270.920 3898.870 276.950 3904.940 ;
        RECT 30.530 3605.730 34.530 3689.350 ;
        RECT 270.920 3682.870 276.950 3688.940 ;
        RECT 316.750 3683.110 319.360 3688.660 ;
        RECT 30.530 3389.730 34.530 3473.350 ;
        RECT 270.920 3466.870 276.950 3472.940 ;
        RECT 316.750 3467.110 319.360 3472.660 ;
        RECT 30.530 3173.730 34.530 3257.350 ;
        RECT 270.920 3250.870 276.950 3256.940 ;
        RECT 316.750 3251.110 319.360 3256.660 ;
        RECT 30.530 2957.730 34.530 3041.350 ;
        RECT 270.920 3034.870 276.950 3040.940 ;
        RECT 316.750 3035.110 319.360 3040.660 ;
        RECT 30.530 2741.730 34.530 2825.350 ;
        RECT 270.920 2818.870 276.950 2824.940 ;
        RECT 316.750 2819.110 319.360 2824.660 ;
        RECT 30.530 2103.730 34.530 2187.350 ;
        RECT 270.920 2180.870 276.950 2186.940 ;
        RECT 316.750 2181.110 319.360 2186.660 ;
        RECT 30.530 1887.730 34.530 1971.350 ;
        RECT 270.920 1964.870 276.950 1970.940 ;
        RECT 316.750 1965.110 319.360 1970.660 ;
        RECT 30.530 1671.730 34.530 1755.350 ;
        RECT 270.920 1748.870 276.950 1754.940 ;
        RECT 316.750 1753.110 319.360 1758.660 ;
        RECT 30.530 1455.730 34.530 1539.350 ;
        RECT 270.920 1532.870 276.950 1538.940 ;
        RECT 316.750 1533.110 319.360 1538.660 ;
        RECT 316.510 1352.290 319.610 1388.960 ;
        RECT 316.510 1349.190 335.860 1352.290 ;
        RECT 30.530 1239.730 34.530 1323.350 ;
        RECT 270.920 1316.870 276.950 1322.940 ;
        RECT 332.760 1231.740 335.860 1349.190 ;
        RECT 1346.820 1232.340 1349.060 1246.620 ;
        RECT 1421.770 1232.340 1424.010 1246.620 ;
        RECT 1496.770 1232.340 1499.010 1246.620 ;
        RECT 1573.070 1232.340 1575.310 1246.620 ;
        RECT 3253.090 1231.480 3256.190 1388.990 ;
        RECT 3334.450 1232.330 3383.350 1247.380 ;
        RECT 30.530 1023.730 34.530 1107.350 ;
        RECT 270.920 1100.870 276.950 1106.940 ;
      LAYER via4 ;
        RECT 497.355 5156.255 498.535 5157.435 ;
        RECT 514.290 5156.275 515.470 5157.455 ;
        RECT 531.140 5156.265 532.320 5157.445 ;
        RECT 497.355 5154.655 498.535 5155.835 ;
        RECT 514.290 5154.675 515.470 5155.855 ;
        RECT 531.140 5154.665 532.320 5155.845 ;
        RECT 754.355 5156.255 755.535 5157.435 ;
        RECT 771.290 5156.275 772.470 5157.455 ;
        RECT 788.140 5156.265 789.320 5157.445 ;
        RECT 754.355 5154.655 755.535 5155.835 ;
        RECT 771.290 5154.675 772.470 5155.855 ;
        RECT 788.140 5154.665 789.320 5155.845 ;
        RECT 1011.355 5156.255 1012.535 5157.435 ;
        RECT 1028.290 5156.275 1029.470 5157.455 ;
        RECT 1045.140 5156.265 1046.320 5157.445 ;
        RECT 1011.355 5154.655 1012.535 5155.835 ;
        RECT 1028.290 5154.675 1029.470 5155.855 ;
        RECT 1045.140 5154.665 1046.320 5155.845 ;
        RECT 1268.355 5156.255 1269.535 5157.435 ;
        RECT 1285.290 5156.275 1286.470 5157.455 ;
        RECT 1302.140 5156.265 1303.320 5157.445 ;
        RECT 1268.355 5154.655 1269.535 5155.835 ;
        RECT 1285.290 5154.675 1286.470 5155.855 ;
        RECT 1302.140 5154.665 1303.320 5155.845 ;
        RECT 1526.355 5156.255 1527.535 5157.435 ;
        RECT 1543.290 5156.275 1544.470 5157.455 ;
        RECT 1560.140 5156.265 1561.320 5157.445 ;
        RECT 1526.355 5154.655 1527.535 5155.835 ;
        RECT 1543.290 5154.675 1544.470 5155.855 ;
        RECT 1560.140 5154.665 1561.320 5155.845 ;
        RECT 1778.355 5156.255 1779.535 5157.435 ;
        RECT 1795.290 5156.275 1796.470 5157.455 ;
        RECT 1812.140 5156.265 1813.320 5157.445 ;
        RECT 1778.355 5154.655 1779.535 5155.835 ;
        RECT 1795.290 5154.675 1796.470 5155.855 ;
        RECT 1812.140 5154.665 1813.320 5155.845 ;
        RECT 2115.355 5156.255 2116.535 5157.435 ;
        RECT 2132.290 5156.275 2133.470 5157.455 ;
        RECT 2149.140 5156.265 2150.320 5157.445 ;
        RECT 2115.355 5154.655 2116.535 5155.835 ;
        RECT 2132.290 5154.675 2133.470 5155.855 ;
        RECT 2149.140 5154.665 2150.320 5155.845 ;
        RECT 2500.355 5156.255 2501.535 5157.435 ;
        RECT 2517.290 5156.275 2518.470 5157.455 ;
        RECT 2534.140 5156.265 2535.320 5157.445 ;
        RECT 2500.355 5154.655 2501.535 5155.835 ;
        RECT 2517.290 5154.675 2518.470 5155.855 ;
        RECT 2534.140 5154.665 2535.320 5155.845 ;
        RECT 2757.355 5156.255 2758.535 5157.435 ;
        RECT 2774.290 5156.275 2775.470 5157.455 ;
        RECT 2791.140 5156.265 2792.320 5157.445 ;
        RECT 2757.355 5154.655 2758.535 5155.835 ;
        RECT 2774.290 5154.675 2775.470 5155.855 ;
        RECT 2791.140 5154.665 2792.320 5155.845 ;
        RECT 574.795 4970.465 579.175 4974.845 ;
        RECT 831.795 4970.465 836.175 4974.845 ;
        RECT 1088.795 4970.465 1093.175 4974.845 ;
        RECT 1345.795 4970.465 1350.175 4974.845 ;
        RECT 1603.795 4970.465 1608.175 4974.845 ;
        RECT 1855.795 4970.465 1860.175 4974.845 ;
        RECT 2192.795 4970.465 2197.175 4974.845 ;
        RECT 2577.795 4970.465 2582.175 4974.845 ;
        RECT 2834.795 4970.465 2839.175 4974.845 ;
        RECT 271.745 4744.795 276.125 4749.175 ;
        RECT 31.120 4701.135 32.300 4702.315 ;
        RECT 32.720 4701.135 33.900 4702.315 ;
        RECT 31.150 4684.305 32.330 4685.485 ;
        RECT 32.750 4684.305 33.930 4685.485 ;
        RECT 31.155 4667.355 32.335 4668.535 ;
        RECT 32.755 4667.355 33.935 4668.535 ;
        RECT 271.745 4115.795 276.125 4120.175 ;
        RECT 31.120 4072.135 32.300 4073.315 ;
        RECT 32.720 4072.135 33.900 4073.315 ;
        RECT 31.150 4055.305 32.330 4056.485 ;
        RECT 32.750 4055.305 33.930 4056.485 ;
        RECT 31.155 4038.355 32.335 4039.535 ;
        RECT 32.755 4038.355 33.935 4039.535 ;
        RECT 271.745 3899.795 276.125 3904.175 ;
        RECT 31.120 3856.135 32.300 3857.315 ;
        RECT 32.720 3856.135 33.900 3857.315 ;
        RECT 31.150 3839.305 32.330 3840.485 ;
        RECT 32.750 3839.305 33.930 3840.485 ;
        RECT 31.155 3822.355 32.335 3823.535 ;
        RECT 32.755 3822.355 33.935 3823.535 ;
        RECT 271.745 3683.795 276.125 3688.175 ;
        RECT 31.120 3640.135 32.300 3641.315 ;
        RECT 32.720 3640.135 33.900 3641.315 ;
        RECT 31.150 3623.305 32.330 3624.485 ;
        RECT 32.750 3623.305 33.930 3624.485 ;
        RECT 31.155 3606.355 32.335 3607.535 ;
        RECT 32.755 3606.355 33.935 3607.535 ;
        RECT 271.745 3467.795 276.125 3472.175 ;
        RECT 31.120 3424.135 32.300 3425.315 ;
        RECT 32.720 3424.135 33.900 3425.315 ;
        RECT 31.150 3407.305 32.330 3408.485 ;
        RECT 32.750 3407.305 33.930 3408.485 ;
        RECT 31.155 3390.355 32.335 3391.535 ;
        RECT 32.755 3390.355 33.935 3391.535 ;
        RECT 271.745 3251.795 276.125 3256.175 ;
        RECT 31.120 3208.135 32.300 3209.315 ;
        RECT 32.720 3208.135 33.900 3209.315 ;
        RECT 31.150 3191.305 32.330 3192.485 ;
        RECT 32.750 3191.305 33.930 3192.485 ;
        RECT 31.155 3174.355 32.335 3175.535 ;
        RECT 32.755 3174.355 33.935 3175.535 ;
        RECT 271.745 3035.795 276.125 3040.175 ;
        RECT 31.120 2992.135 32.300 2993.315 ;
        RECT 32.720 2992.135 33.900 2993.315 ;
        RECT 31.150 2975.305 32.330 2976.485 ;
        RECT 32.750 2975.305 33.930 2976.485 ;
        RECT 31.155 2958.355 32.335 2959.535 ;
        RECT 32.755 2958.355 33.935 2959.535 ;
        RECT 271.745 2819.795 276.125 2824.175 ;
        RECT 31.120 2776.135 32.300 2777.315 ;
        RECT 32.720 2776.135 33.900 2777.315 ;
        RECT 31.150 2759.305 32.330 2760.485 ;
        RECT 32.750 2759.305 33.930 2760.485 ;
        RECT 31.155 2742.355 32.335 2743.535 ;
        RECT 32.755 2742.355 33.935 2743.535 ;
        RECT 271.745 2181.795 276.125 2186.175 ;
        RECT 31.120 2138.135 32.300 2139.315 ;
        RECT 32.720 2138.135 33.900 2139.315 ;
        RECT 31.150 2121.305 32.330 2122.485 ;
        RECT 32.750 2121.305 33.930 2122.485 ;
        RECT 31.155 2104.355 32.335 2105.535 ;
        RECT 32.755 2104.355 33.935 2105.535 ;
        RECT 271.745 1965.795 276.125 1970.175 ;
        RECT 31.120 1922.135 32.300 1923.315 ;
        RECT 32.720 1922.135 33.900 1923.315 ;
        RECT 31.150 1905.305 32.330 1906.485 ;
        RECT 32.750 1905.305 33.930 1906.485 ;
        RECT 31.155 1888.355 32.335 1889.535 ;
        RECT 32.755 1888.355 33.935 1889.535 ;
        RECT 271.745 1749.795 276.125 1754.175 ;
        RECT 31.120 1706.135 32.300 1707.315 ;
        RECT 32.720 1706.135 33.900 1707.315 ;
        RECT 31.150 1689.305 32.330 1690.485 ;
        RECT 32.750 1689.305 33.930 1690.485 ;
        RECT 31.155 1672.355 32.335 1673.535 ;
        RECT 32.755 1672.355 33.935 1673.535 ;
        RECT 271.745 1533.795 276.125 1538.175 ;
        RECT 31.120 1490.135 32.300 1491.315 ;
        RECT 32.720 1490.135 33.900 1491.315 ;
        RECT 31.150 1473.305 32.330 1474.485 ;
        RECT 32.750 1473.305 33.930 1474.485 ;
        RECT 31.155 1456.355 32.335 1457.535 ;
        RECT 32.755 1456.355 33.935 1457.535 ;
        RECT 271.745 1317.795 276.125 1322.175 ;
        RECT 31.120 1274.135 32.300 1275.315 ;
        RECT 32.720 1274.135 33.900 1275.315 ;
        RECT 31.150 1257.305 32.330 1258.485 ;
        RECT 32.750 1257.305 33.930 1258.485 ;
        RECT 31.155 1240.355 32.335 1241.535 ;
        RECT 32.755 1240.355 33.935 1241.535 ;
        RECT 333.695 1245.670 334.875 1246.850 ;
        RECT 333.695 1244.070 334.875 1245.250 ;
        RECT 333.695 1242.470 334.875 1243.650 ;
        RECT 333.695 1240.870 334.875 1242.050 ;
        RECT 333.695 1239.270 334.875 1240.450 ;
        RECT 333.695 1237.670 334.875 1238.850 ;
        RECT 333.695 1236.070 334.875 1237.250 ;
        RECT 333.695 1234.470 334.875 1235.650 ;
        RECT 333.695 1232.870 334.875 1234.050 ;
        RECT 1347.350 1244.705 1348.530 1245.885 ;
        RECT 1347.350 1243.105 1348.530 1244.285 ;
        RECT 1347.350 1241.505 1348.530 1242.685 ;
        RECT 1347.350 1239.905 1348.530 1241.085 ;
        RECT 1347.350 1238.305 1348.530 1239.485 ;
        RECT 1347.350 1236.705 1348.530 1237.885 ;
        RECT 1347.350 1235.105 1348.530 1236.285 ;
        RECT 1347.350 1233.505 1348.530 1234.685 ;
        RECT 1422.300 1244.705 1423.480 1245.885 ;
        RECT 1422.300 1243.105 1423.480 1244.285 ;
        RECT 1422.300 1241.505 1423.480 1242.685 ;
        RECT 1422.300 1239.905 1423.480 1241.085 ;
        RECT 1422.300 1238.305 1423.480 1239.485 ;
        RECT 1422.300 1236.705 1423.480 1237.885 ;
        RECT 1422.300 1235.105 1423.480 1236.285 ;
        RECT 1422.300 1233.505 1423.480 1234.685 ;
        RECT 1497.300 1244.705 1498.480 1245.885 ;
        RECT 1497.300 1243.105 1498.480 1244.285 ;
        RECT 1497.300 1241.505 1498.480 1242.685 ;
        RECT 1497.300 1239.905 1498.480 1241.085 ;
        RECT 1497.300 1238.305 1498.480 1239.485 ;
        RECT 1497.300 1236.705 1498.480 1237.885 ;
        RECT 1497.300 1235.105 1498.480 1236.285 ;
        RECT 1497.300 1233.505 1498.480 1234.685 ;
        RECT 1573.600 1244.705 1574.780 1245.885 ;
        RECT 1573.600 1243.105 1574.780 1244.285 ;
        RECT 1573.600 1241.505 1574.780 1242.685 ;
        RECT 1573.600 1239.905 1574.780 1241.085 ;
        RECT 1573.600 1238.305 1574.780 1239.485 ;
        RECT 1573.600 1236.705 1574.780 1237.885 ;
        RECT 1573.600 1235.105 1574.780 1236.285 ;
        RECT 1573.600 1233.505 1574.780 1234.685 ;
        RECT 3253.240 1232.895 3256.020 1246.875 ;
        RECT 3335.560 1233.685 3347.940 1246.065 ;
        RECT 3371.130 1233.590 3381.910 1245.970 ;
        RECT 271.745 1101.795 276.125 1106.175 ;
        RECT 31.120 1058.135 32.300 1059.315 ;
        RECT 32.720 1058.135 33.900 1059.315 ;
        RECT 31.150 1041.305 32.330 1042.485 ;
        RECT 32.750 1041.305 33.930 1042.485 ;
        RECT 31.155 1024.355 32.335 1025.535 ;
        RECT 32.755 1024.355 33.935 1025.535 ;
      LAYER met5 ;
        RECT 497.060 5153.970 498.810 5158.130 ;
        RECT 514.010 5154.010 515.740 5158.390 ;
        RECT 497.140 5145.520 498.740 5153.970 ;
        RECT 514.040 5145.680 515.640 5154.010 ;
        RECT 530.830 5153.990 532.560 5158.370 ;
        RECT 530.940 5145.680 532.540 5153.990 ;
        RECT 754.060 5153.970 755.810 5158.130 ;
        RECT 771.010 5154.010 772.740 5158.390 ;
        RECT 754.140 5145.520 755.740 5153.970 ;
        RECT 771.040 5145.680 772.640 5154.010 ;
        RECT 787.830 5153.990 789.560 5158.370 ;
        RECT 787.940 5145.680 789.540 5153.990 ;
        RECT 1011.060 5153.970 1012.810 5158.130 ;
        RECT 1028.010 5154.010 1029.740 5158.390 ;
        RECT 1011.140 5145.520 1012.740 5153.970 ;
        RECT 1028.040 5145.680 1029.640 5154.010 ;
        RECT 1044.830 5153.990 1046.560 5158.370 ;
        RECT 1044.940 5145.680 1046.540 5153.990 ;
        RECT 1268.060 5153.970 1269.810 5158.130 ;
        RECT 1285.010 5154.010 1286.740 5158.390 ;
        RECT 1268.140 5145.520 1269.740 5153.970 ;
        RECT 1285.040 5145.680 1286.640 5154.010 ;
        RECT 1301.830 5153.990 1303.560 5158.370 ;
        RECT 1301.940 5145.680 1303.540 5153.990 ;
        RECT 1526.060 5153.970 1527.810 5158.130 ;
        RECT 1543.010 5154.010 1544.740 5158.390 ;
        RECT 1526.140 5145.520 1527.740 5153.970 ;
        RECT 1543.040 5145.680 1544.640 5154.010 ;
        RECT 1559.830 5153.990 1561.560 5158.370 ;
        RECT 1559.940 5145.680 1561.540 5153.990 ;
        RECT 1778.060 5153.970 1779.810 5158.130 ;
        RECT 1795.010 5154.010 1796.740 5158.390 ;
        RECT 1778.140 5145.520 1779.740 5153.970 ;
        RECT 1795.040 5145.680 1796.640 5154.010 ;
        RECT 1811.830 5153.990 1813.560 5158.370 ;
        RECT 1811.940 5145.680 1813.540 5153.990 ;
        RECT 2115.060 5153.970 2116.810 5158.130 ;
        RECT 2132.010 5154.010 2133.740 5158.390 ;
        RECT 2115.140 5145.520 2116.740 5153.970 ;
        RECT 2132.040 5145.680 2133.640 5154.010 ;
        RECT 2148.830 5153.990 2150.560 5158.370 ;
        RECT 2148.940 5145.680 2150.540 5153.990 ;
        RECT 2500.060 5153.970 2501.810 5158.130 ;
        RECT 2517.010 5154.010 2518.740 5158.390 ;
        RECT 2500.140 5145.520 2501.740 5153.970 ;
        RECT 2517.040 5145.680 2518.640 5154.010 ;
        RECT 2533.830 5153.990 2535.560 5158.370 ;
        RECT 2533.940 5145.680 2535.540 5153.990 ;
        RECT 2757.060 5153.970 2758.810 5158.130 ;
        RECT 2774.010 5154.010 2775.740 5158.390 ;
        RECT 2757.140 5145.520 2758.740 5153.970 ;
        RECT 2774.040 5145.680 2775.640 5154.010 ;
        RECT 2790.830 5153.990 2792.560 5158.370 ;
        RECT 2790.940 5145.680 2792.540 5153.990 ;
        RECT 270.990 4969.510 3383.100 4975.510 ;
        RECT 270.990 4917.940 276.990 4969.510 ;
        RECT 3370.100 4963.480 3383.100 4969.510 ;
        RECT 270.990 4914.840 316.580 4917.940 ;
        RECT 30.440 4702.540 34.635 4702.700 ;
        RECT 30.240 4700.940 42.910 4702.540 ;
        RECT 30.440 4700.895 34.635 4700.940 ;
        RECT 30.170 4685.640 34.645 4685.770 ;
        RECT 30.170 4684.040 42.910 4685.640 ;
        RECT 30.170 4684.030 34.645 4684.040 ;
        RECT 30.425 4668.740 34.900 4668.850 ;
        RECT 30.425 4667.140 43.070 4668.740 ;
        RECT 30.425 4667.040 34.900 4667.140 ;
        RECT 30.440 4073.540 34.635 4073.700 ;
        RECT 30.240 4071.940 42.910 4073.540 ;
        RECT 30.440 4071.895 34.635 4071.940 ;
        RECT 30.170 4056.640 34.645 4056.770 ;
        RECT 30.170 4055.040 42.910 4056.640 ;
        RECT 30.170 4055.030 34.645 4055.040 ;
        RECT 30.425 4039.740 34.900 4039.850 ;
        RECT 30.425 4038.140 43.070 4039.740 ;
        RECT 30.425 4038.040 34.900 4038.140 ;
        RECT 30.440 3857.540 34.635 3857.700 ;
        RECT 30.240 3855.940 42.910 3857.540 ;
        RECT 30.440 3855.895 34.635 3855.940 ;
        RECT 30.170 3840.640 34.645 3840.770 ;
        RECT 30.170 3839.040 42.910 3840.640 ;
        RECT 30.170 3839.030 34.645 3839.040 ;
        RECT 30.425 3823.740 34.900 3823.850 ;
        RECT 30.425 3822.140 43.070 3823.740 ;
        RECT 30.425 3822.040 34.900 3822.140 ;
        RECT 30.440 3641.540 34.635 3641.700 ;
        RECT 30.240 3639.940 42.910 3641.540 ;
        RECT 30.440 3639.895 34.635 3639.940 ;
        RECT 30.170 3624.640 34.645 3624.770 ;
        RECT 30.170 3623.040 42.910 3624.640 ;
        RECT 30.170 3623.030 34.645 3623.040 ;
        RECT 30.425 3607.740 34.900 3607.850 ;
        RECT 30.425 3606.140 43.070 3607.740 ;
        RECT 30.425 3606.040 34.900 3606.140 ;
        RECT 30.440 3425.540 34.635 3425.700 ;
        RECT 30.240 3423.940 42.910 3425.540 ;
        RECT 30.440 3423.895 34.635 3423.940 ;
        RECT 30.170 3408.640 34.645 3408.770 ;
        RECT 30.170 3407.040 42.910 3408.640 ;
        RECT 30.170 3407.030 34.645 3407.040 ;
        RECT 30.425 3391.740 34.900 3391.850 ;
        RECT 30.425 3390.140 43.070 3391.740 ;
        RECT 30.425 3390.040 34.900 3390.140 ;
        RECT 30.440 3209.540 34.635 3209.700 ;
        RECT 30.240 3207.940 42.910 3209.540 ;
        RECT 30.440 3207.895 34.635 3207.940 ;
        RECT 30.170 3192.640 34.645 3192.770 ;
        RECT 30.170 3191.040 42.910 3192.640 ;
        RECT 30.170 3191.030 34.645 3191.040 ;
        RECT 30.425 3175.740 34.900 3175.850 ;
        RECT 30.425 3174.140 43.070 3175.740 ;
        RECT 30.425 3174.040 34.900 3174.140 ;
        RECT 30.440 2993.540 34.635 2993.700 ;
        RECT 30.240 2991.940 42.910 2993.540 ;
        RECT 30.440 2991.895 34.635 2991.940 ;
        RECT 30.170 2976.640 34.645 2976.770 ;
        RECT 30.170 2975.040 42.910 2976.640 ;
        RECT 30.170 2975.030 34.645 2975.040 ;
        RECT 30.425 2959.740 34.900 2959.850 ;
        RECT 30.425 2958.140 43.070 2959.740 ;
        RECT 30.425 2958.040 34.900 2958.140 ;
        RECT 30.440 2777.540 34.635 2777.700 ;
        RECT 30.240 2775.940 42.910 2777.540 ;
        RECT 30.440 2775.895 34.635 2775.940 ;
        RECT 30.170 2760.640 34.645 2760.770 ;
        RECT 30.170 2759.040 42.910 2760.640 ;
        RECT 30.170 2759.030 34.645 2759.040 ;
        RECT 30.425 2743.740 34.900 2743.850 ;
        RECT 30.425 2742.140 43.070 2743.740 ;
        RECT 30.425 2742.040 34.900 2742.140 ;
        RECT 30.440 2139.540 34.635 2139.700 ;
        RECT 30.240 2137.940 42.910 2139.540 ;
        RECT 30.440 2137.895 34.635 2137.940 ;
        RECT 30.170 2122.640 34.645 2122.770 ;
        RECT 30.170 2121.040 42.910 2122.640 ;
        RECT 30.170 2121.030 34.645 2121.040 ;
        RECT 30.425 2105.740 34.900 2105.850 ;
        RECT 30.425 2104.140 43.070 2105.740 ;
        RECT 30.425 2104.040 34.900 2104.140 ;
        RECT 30.440 1923.540 34.635 1923.700 ;
        RECT 30.240 1921.940 42.910 1923.540 ;
        RECT 30.440 1921.895 34.635 1921.940 ;
        RECT 30.170 1906.640 34.645 1906.770 ;
        RECT 30.170 1905.040 42.910 1906.640 ;
        RECT 30.170 1905.030 34.645 1905.040 ;
        RECT 30.425 1889.740 34.900 1889.850 ;
        RECT 30.425 1888.140 43.070 1889.740 ;
        RECT 30.425 1888.040 34.900 1888.140 ;
        RECT 30.440 1707.540 34.635 1707.700 ;
        RECT 30.240 1705.940 42.910 1707.540 ;
        RECT 30.440 1705.895 34.635 1705.940 ;
        RECT 30.170 1690.640 34.645 1690.770 ;
        RECT 30.170 1689.040 42.910 1690.640 ;
        RECT 30.170 1689.030 34.645 1689.040 ;
        RECT 30.425 1673.740 34.900 1673.850 ;
        RECT 30.425 1672.140 43.070 1673.740 ;
        RECT 30.425 1672.040 34.900 1672.140 ;
        RECT 30.440 1491.540 34.635 1491.700 ;
        RECT 30.240 1489.940 42.910 1491.540 ;
        RECT 30.440 1489.895 34.635 1489.940 ;
        RECT 30.170 1474.640 34.645 1474.770 ;
        RECT 30.170 1473.040 42.910 1474.640 ;
        RECT 30.170 1473.030 34.645 1473.040 ;
        RECT 30.425 1457.740 34.900 1457.850 ;
        RECT 30.425 1456.140 43.070 1457.740 ;
        RECT 30.425 1456.040 34.900 1456.140 ;
        RECT 270.990 1392.020 276.990 4914.840 ;
        RECT 270.990 1388.920 316.560 1392.020 ;
        RECT 30.440 1275.540 34.635 1275.700 ;
        RECT 30.240 1273.940 42.910 1275.540 ;
        RECT 30.440 1273.895 34.635 1273.940 ;
        RECT 30.170 1258.640 34.645 1258.770 ;
        RECT 30.170 1257.040 42.910 1258.640 ;
        RECT 30.170 1257.030 34.645 1257.040 ;
        RECT 270.990 1247.330 276.990 1388.920 ;
        RECT 30.425 1241.740 34.900 1241.850 ;
        RECT 30.425 1240.140 43.070 1241.740 ;
        RECT 30.425 1240.040 34.900 1240.140 ;
        RECT 270.990 1232.330 3349.450 1247.330 ;
        RECT 3370.780 1233.080 3382.260 1246.480 ;
        RECT 270.990 1096.710 276.990 1232.330 ;
        RECT 30.440 1059.540 34.635 1059.700 ;
        RECT 30.240 1057.940 42.910 1059.540 ;
        RECT 30.440 1057.895 34.635 1057.940 ;
        RECT 30.170 1042.640 34.645 1042.770 ;
        RECT 30.170 1041.040 42.910 1042.640 ;
        RECT 30.170 1041.030 34.645 1041.040 ;
        RECT 30.425 1025.740 34.900 1025.850 ;
        RECT 30.425 1024.140 43.070 1025.740 ;
        RECT 30.425 1024.040 34.900 1024.140 ;
    END
  END vccd1_core
  PIN vssa1_core
    PORT
      LAYER met3 ;
        RECT 2878.500 4975.160 2902.395 4988.390 ;
        RECT 2928.390 4975.160 2952.290 4988.390 ;
        RECT 3319.570 2128.740 3388.560 2152.505 ;
        RECT 3319.570 2127.810 3335.550 2128.740 ;
        RECT 3319.570 2078.710 3388.560 2102.610 ;
      LAYER via3 ;
        RECT 2879.070 4975.715 2901.790 4985.235 ;
        RECT 2928.920 4975.745 2951.640 4985.265 ;
        RECT 3320.725 2128.425 3332.645 2151.945 ;
        RECT 3320.640 2079.435 3332.560 2102.155 ;
      LAYER met4 ;
        RECT 2878.400 4953.940 2902.390 4985.650 ;
        RECT 2928.350 4954.010 2952.340 4985.720 ;
        RECT 3320.040 2127.860 3333.060 2152.450 ;
        RECT 3320.090 2078.800 3333.170 2102.620 ;
        RECT 292.510 1332.040 295.610 1364.960 ;
        RECT 1953.860 1332.370 1957.790 1347.350 ;
        RECT 2029.110 1332.370 2033.040 1347.350 ;
        RECT 1956.870 1311.040 1957.770 1332.370 ;
        RECT 2032.120 1311.040 2033.020 1332.370 ;
        RECT 3277.090 1331.930 3280.190 1365.020 ;
      LAYER via4 ;
        RECT 2879.375 4955.105 2901.355 4965.885 ;
        RECT 2929.355 4955.175 2951.335 4965.955 ;
        RECT 3321.295 2129.195 3332.075 2151.175 ;
        RECT 3321.210 2079.805 3331.990 2101.785 ;
        RECT 293.445 1345.640 294.625 1346.820 ;
        RECT 293.445 1344.040 294.625 1345.220 ;
        RECT 293.445 1342.440 294.625 1343.620 ;
        RECT 293.445 1340.840 294.625 1342.020 ;
        RECT 293.445 1339.240 294.625 1340.420 ;
        RECT 293.445 1337.640 294.625 1338.820 ;
        RECT 293.445 1336.040 294.625 1337.220 ;
        RECT 293.445 1334.440 294.625 1335.620 ;
        RECT 293.445 1332.840 294.625 1334.020 ;
        RECT 1954.455 1332.825 1957.235 1346.805 ;
        RECT 2029.705 1332.825 2032.485 1346.805 ;
        RECT 3278.035 1345.625 3279.215 1346.805 ;
        RECT 3278.035 1344.025 3279.215 1345.205 ;
        RECT 3278.035 1342.425 3279.215 1343.605 ;
        RECT 3278.035 1340.825 3279.215 1342.005 ;
        RECT 3278.035 1339.225 3279.215 1340.405 ;
        RECT 3278.035 1337.625 3279.215 1338.805 ;
        RECT 3278.035 1336.025 3279.215 1337.205 ;
        RECT 3278.035 1334.425 3279.215 1335.605 ;
        RECT 3278.035 1332.825 3279.215 1334.005 ;
      LAYER met5 ;
        RECT 2878.200 4953.980 3333.100 4966.980 ;
        RECT 3320.100 4941.940 3333.100 4953.980 ;
        RECT 3280.190 4938.840 3333.100 4941.940 ;
        RECT 3320.100 1368.020 3333.100 4938.840 ;
        RECT 3280.130 1364.920 3333.100 1368.020 ;
        RECT 3320.100 1347.330 3333.100 1364.920 ;
        RECT 291.940 1332.330 3333.100 1347.330 ;
    END
  END vssa1_core
  PIN vdda1_core
    PORT
      LAYER met3 ;
        RECT 3335.860 4142.605 3389.090 4166.505 ;
        RECT 3335.860 4092.710 3389.090 4116.610 ;
        RECT 3335.310 2569.605 3388.500 2593.505 ;
        RECT 3335.310 2519.710 3388.500 2543.610 ;
      LAYER via3 ;
        RECT 3336.580 4143.230 3348.500 4165.950 ;
        RECT 3336.510 4093.260 3348.430 4115.980 ;
        RECT 3336.845 2570.435 3348.365 2592.755 ;
        RECT 3336.915 2520.485 3348.435 2542.805 ;
      LAYER met4 ;
        RECT 3291.900 4934.060 3349.130 4937.180 ;
        RECT 3336.010 4142.600 3349.010 4166.550 ;
        RECT 3336.070 4092.730 3349.070 4116.680 ;
        RECT 3336.030 2569.600 3349.070 2593.480 ;
        RECT 3336.090 2519.750 3349.130 2543.630 ;
        RECT 297.310 1333.090 300.410 1369.760 ;
        RECT 297.310 1329.990 316.660 1333.090 ;
        RECT 313.560 1312.010 316.660 1329.990 ;
        RECT 1919.970 1327.310 1920.870 1327.380 ;
        RECT 1995.220 1327.310 1996.120 1327.380 ;
        RECT 1916.830 1314.270 1920.870 1327.310 ;
        RECT 1992.080 1314.270 1996.120 1327.310 ;
        RECT 1919.970 1311.220 1920.870 1314.270 ;
        RECT 1995.220 1311.220 1996.120 1314.270 ;
        RECT 3272.290 1311.810 3275.390 1369.780 ;
        RECT 3294.750 1369.690 3349.060 1372.870 ;
        RECT 3336.080 1365.690 3349.060 1369.690 ;
      LAYER via4 ;
        RECT 3292.885 4935.030 3294.065 4936.210 ;
        RECT 3294.485 4935.030 3295.665 4936.210 ;
        RECT 3296.085 4935.030 3297.265 4936.210 ;
        RECT 3297.685 4935.030 3298.865 4936.210 ;
        RECT 3299.285 4935.030 3300.465 4936.210 ;
        RECT 3300.885 4935.030 3302.065 4936.210 ;
        RECT 3302.485 4935.030 3303.665 4936.210 ;
        RECT 3304.085 4935.030 3305.265 4936.210 ;
        RECT 3305.685 4935.030 3306.865 4936.210 ;
        RECT 3307.285 4935.030 3308.465 4936.210 ;
        RECT 3308.885 4935.030 3310.065 4936.210 ;
        RECT 3310.485 4935.030 3311.665 4936.210 ;
        RECT 3312.085 4935.030 3313.265 4936.210 ;
        RECT 3313.685 4935.030 3314.865 4936.210 ;
        RECT 3336.405 4935.055 3337.585 4936.235 ;
        RECT 3338.005 4935.055 3339.185 4936.235 ;
        RECT 3339.605 4935.055 3340.785 4936.235 ;
        RECT 3341.205 4935.055 3342.385 4936.235 ;
        RECT 3342.805 4935.055 3343.985 4936.235 ;
        RECT 3344.405 4935.055 3345.585 4936.235 ;
        RECT 3346.005 4935.055 3347.185 4936.235 ;
        RECT 3347.605 4935.055 3348.785 4936.235 ;
        RECT 3337.150 4143.600 3347.930 4165.580 ;
        RECT 3337.080 4093.630 3347.860 4115.610 ;
        RECT 3337.215 2570.605 3347.995 2592.585 ;
        RECT 3337.285 2520.655 3348.065 2542.635 ;
        RECT 3295.925 1370.645 3297.105 1371.825 ;
        RECT 3297.525 1370.645 3298.705 1371.825 ;
        RECT 3299.125 1370.645 3300.305 1371.825 ;
        RECT 3300.725 1370.645 3301.905 1371.825 ;
        RECT 3302.325 1370.645 3303.505 1371.825 ;
        RECT 3303.925 1370.645 3305.105 1371.825 ;
        RECT 3305.525 1370.645 3306.705 1371.825 ;
        RECT 3307.125 1370.645 3308.305 1371.825 ;
        RECT 3308.725 1370.645 3309.905 1371.825 ;
        RECT 3310.325 1370.645 3311.505 1371.825 ;
        RECT 3311.925 1370.645 3313.105 1371.825 ;
        RECT 3313.525 1370.645 3314.705 1371.825 ;
        RECT 314.485 1325.620 315.665 1326.800 ;
        RECT 314.485 1324.020 315.665 1325.200 ;
        RECT 314.485 1322.420 315.665 1323.600 ;
        RECT 314.485 1320.820 315.665 1322.000 ;
        RECT 314.485 1319.220 315.665 1320.400 ;
        RECT 314.485 1317.620 315.665 1318.800 ;
        RECT 314.485 1316.020 315.665 1317.200 ;
        RECT 314.485 1314.420 315.665 1315.600 ;
        RECT 1917.435 1315.260 1920.215 1326.040 ;
        RECT 1992.685 1315.260 1995.465 1326.040 ;
        RECT 314.485 1312.820 315.665 1314.000 ;
        RECT 3337.240 1366.280 3348.020 1372.260 ;
        RECT 3273.245 1325.615 3274.425 1326.795 ;
        RECT 3273.245 1324.015 3274.425 1325.195 ;
        RECT 3273.245 1322.415 3274.425 1323.595 ;
        RECT 3273.245 1320.815 3274.425 1321.995 ;
        RECT 3273.245 1319.215 3274.425 1320.395 ;
        RECT 3273.245 1317.615 3274.425 1318.795 ;
        RECT 3273.245 1316.015 3274.425 1317.195 ;
        RECT 3273.245 1314.415 3274.425 1315.595 ;
        RECT 3273.245 1312.815 3274.425 1313.995 ;
      LAYER met5 ;
        RECT 3275.390 4934.040 3315.890 4937.140 ;
        RECT 3275.300 1369.720 3315.790 1372.820 ;
        RECT 3336.100 1327.330 3349.100 4937.830 ;
        RECT 312.670 1312.330 3349.100 1327.330 ;
    END
  END vdda1_core
  OBS
      LAYER met2 ;
        RECT 2208.095 203.885 2209.960 211.885 ;
        RECT 2208.015 202.820 2210.045 203.885 ;
      LAYER via2 ;
        RECT 2208.285 203.020 2209.765 203.700 ;
      LAYER met3 ;
        RECT 549.500 4996.630 555.500 5093.480 ;
        RECT 557.500 5029.580 563.500 5099.450 ;
        RECT 806.500 4996.630 812.500 5093.480 ;
        RECT 814.500 5029.580 820.500 5099.450 ;
        RECT 842.905 4986.595 844.770 5034.235 ;
        RECT 848.895 4985.700 850.745 5001.540 ;
        RECT 1063.500 4996.630 1069.500 5093.480 ;
        RECT 1071.500 5029.580 1077.500 5099.450 ;
        RECT 1320.500 4996.630 1326.500 5093.480 ;
        RECT 1328.500 5029.580 1334.500 5099.450 ;
        RECT 1578.500 4996.630 1584.500 5093.480 ;
        RECT 1586.500 5029.580 1592.500 5099.450 ;
        RECT 1830.500 4996.630 1836.500 5093.480 ;
        RECT 1838.500 5029.580 1844.500 5099.450 ;
        RECT 2085.090 4986.595 2086.955 5034.235 ;
        RECT 2091.080 4985.695 2092.930 5001.535 ;
        RECT 2167.500 4996.630 2173.500 5093.480 ;
        RECT 2175.500 5029.580 2181.500 5099.450 ;
        RECT 2552.500 4996.630 2558.500 5093.480 ;
        RECT 2560.500 5029.580 2566.500 5099.450 ;
        RECT 2809.500 4996.630 2815.500 5093.480 ;
        RECT 2817.500 5029.580 2823.500 5099.450 ;
        RECT 3318.140 4986.595 3320.005 5034.235 ;
        RECT 3324.130 4985.695 3325.980 5001.535 ;
        RECT 220.990 4759.620 309.980 4765.620 ;
        RECT 204.920 4751.620 305.160 4757.620 ;
        RECT 89.140 4727.500 158.310 4733.500 ;
        RECT 3253.080 4725.910 3559.020 4731.910 ;
        RECT 95.110 4719.500 191.260 4725.500 ;
        RECT 3257.900 4717.910 3552.950 4723.910 ;
        RECT 3429.570 4709.500 3499.990 4715.500 ;
        RECT 3396.620 4701.500 3494.020 4707.500 ;
        RECT 3253.080 4499.910 3379.150 4505.910 ;
        RECT 3257.900 4491.910 3363.380 4497.910 ;
        RECT 153.765 4446.875 202.365 4448.740 ;
        RECT 186.465 4440.905 202.345 4442.755 ;
        RECT 3253.080 4274.910 3376.320 4280.910 ;
        RECT 3257.900 4266.910 3363.540 4272.910 ;
        RECT 220.990 4130.620 309.980 4136.620 ;
        RECT 204.920 4122.620 305.160 4128.620 ;
        RECT 89.140 4098.500 158.310 4104.500 ;
        RECT 95.110 4090.500 191.260 4096.500 ;
        RECT 220.990 3922.620 309.980 3928.620 ;
        RECT 204.920 3914.620 305.160 3920.620 ;
        RECT 89.140 3882.500 158.310 3888.500 ;
        RECT 95.110 3874.500 191.260 3880.500 ;
        RECT 3253.080 3833.910 3559.070 3839.910 ;
        RECT 3257.900 3825.910 3553.000 3831.910 ;
        RECT 3429.620 3817.500 3500.040 3823.500 ;
        RECT 3396.670 3809.500 3494.070 3815.500 ;
        RECT 220.990 3698.620 309.980 3704.620 ;
        RECT 204.920 3690.620 305.160 3696.620 ;
        RECT 89.140 3666.500 158.310 3672.500 ;
        RECT 95.110 3658.500 191.260 3664.500 ;
        RECT 3386.595 3622.445 3434.235 3624.310 ;
        RECT 3385.695 3616.470 3401.535 3618.320 ;
        RECT 3253.080 3608.910 3559.070 3614.910 ;
        RECT 3257.900 3600.910 3553.000 3606.910 ;
        RECT 3429.620 3592.500 3500.040 3598.500 ;
        RECT 3396.670 3584.500 3494.070 3590.500 ;
        RECT 220.990 3482.620 309.980 3488.620 ;
        RECT 204.920 3474.620 305.160 3480.620 ;
        RECT 89.140 3450.500 158.310 3456.500 ;
        RECT 95.110 3442.500 191.260 3448.500 ;
        RECT 3253.080 3382.910 3559.070 3388.910 ;
        RECT 3257.900 3374.910 3553.000 3380.910 ;
        RECT 3429.620 3366.500 3500.040 3372.500 ;
        RECT 3396.670 3358.500 3494.070 3364.500 ;
        RECT 220.990 3266.620 309.980 3272.620 ;
        RECT 204.920 3258.620 305.160 3264.620 ;
        RECT 89.140 3234.500 158.310 3240.500 ;
        RECT 95.110 3226.500 191.260 3232.500 ;
        RECT 3253.080 3157.910 3559.070 3163.910 ;
        RECT 3296.550 3149.910 3553.000 3155.910 ;
        RECT 3257.900 3143.910 3303.000 3149.910 ;
        RECT 3429.620 3141.500 3500.040 3147.500 ;
        RECT 3396.670 3133.500 3494.070 3139.500 ;
        RECT 220.990 3055.920 309.980 3061.920 ;
        RECT 204.920 3047.920 305.160 3053.920 ;
        RECT 153.865 3024.500 202.150 3024.870 ;
        RECT 89.140 3023.005 202.150 3024.500 ;
        RECT 89.140 3018.500 158.310 3023.005 ;
        RECT 188.000 3017.035 201.990 3018.885 ;
        RECT 188.000 3016.500 191.260 3017.035 ;
        RECT 95.110 3010.500 191.260 3016.500 ;
        RECT 3253.080 2931.910 3559.070 2937.910 ;
        RECT 3257.900 2923.910 3553.000 2929.910 ;
        RECT 3429.620 2915.500 3500.040 2921.500 ;
        RECT 3396.670 2907.500 3494.070 2913.500 ;
        RECT 220.990 2834.620 309.980 2840.620 ;
        RECT 204.920 2826.620 305.160 2832.620 ;
        RECT 89.140 2802.500 158.310 2808.500 ;
        RECT 95.110 2794.500 191.260 2800.500 ;
        RECT 3253.080 2706.910 3559.070 2712.910 ;
        RECT 3257.900 2698.910 3553.000 2704.910 ;
        RECT 3429.620 2690.500 3500.040 2696.500 ;
        RECT 3396.670 2682.500 3494.070 2688.500 ;
        RECT 3253.080 2492.910 3298.790 2495.910 ;
        RECT 3253.080 2489.910 3559.070 2492.910 ;
        RECT 3292.840 2486.910 3559.070 2489.910 ;
        RECT 3257.900 2478.910 3553.000 2484.910 ;
        RECT 3429.620 2470.500 3500.040 2476.500 ;
        RECT 3396.670 2462.500 3494.070 2468.500 ;
        RECT 3386.595 2240.440 3434.235 2242.305 ;
        RECT 3385.695 2234.465 3401.535 2236.315 ;
        RECT 220.990 2196.620 309.980 2202.620 ;
        RECT 204.920 2188.620 305.160 2194.620 ;
        RECT 89.140 2164.500 158.310 2170.500 ;
        RECT 95.110 2156.500 191.260 2162.500 ;
        RECT 3253.080 2045.910 3559.070 2051.910 ;
        RECT 3257.900 2037.910 3553.000 2043.910 ;
        RECT 3429.620 2029.500 3500.040 2035.500 ;
        RECT 3396.670 2021.500 3494.070 2027.500 ;
        RECT 220.990 1980.620 309.980 1986.620 ;
        RECT 204.920 1972.620 305.160 1978.620 ;
        RECT 89.140 1948.500 158.310 1954.500 ;
        RECT 95.110 1940.500 191.260 1946.500 ;
        RECT 3253.080 1826.910 3328.320 1832.910 ;
        RECT 3322.320 1825.910 3328.320 1826.910 ;
        RECT 3322.320 1819.910 3559.070 1825.910 ;
        RECT 3257.900 1811.910 3553.000 1817.910 ;
        RECT 3429.620 1803.500 3500.040 1809.500 ;
        RECT 3396.670 1795.500 3494.070 1801.500 ;
        RECT 220.990 1769.620 309.980 1775.620 ;
        RECT 204.920 1761.620 305.160 1767.620 ;
        RECT 89.140 1736.615 158.310 1738.500 ;
        RECT 89.140 1734.750 202.545 1736.615 ;
        RECT 89.140 1732.500 158.310 1734.750 ;
        RECT 186.465 1730.500 203.595 1730.630 ;
        RECT 95.110 1728.780 203.595 1730.500 ;
        RECT 95.110 1724.500 191.260 1728.780 ;
        RECT 3253.080 1594.910 3559.070 1600.910 ;
        RECT 3257.900 1586.910 3553.000 1592.910 ;
        RECT 3429.620 1578.500 3500.040 1584.500 ;
        RECT 3396.670 1570.500 3494.070 1576.500 ;
        RECT 220.990 1548.620 309.980 1554.620 ;
        RECT 204.920 1540.620 305.160 1546.620 ;
        RECT 89.140 1516.500 158.310 1522.500 ;
        RECT 95.110 1508.500 191.260 1514.500 ;
        RECT 3376.380 1369.910 3559.070 1375.910 ;
        RECT 3358.100 1361.910 3553.000 1367.910 ;
        RECT 3429.620 1353.500 3500.040 1359.500 ;
        RECT 3396.670 1345.500 3494.070 1351.500 ;
        RECT 89.140 1300.500 158.310 1306.500 ;
        RECT 95.110 1292.500 191.260 1298.500 ;
        RECT 3376.380 1143.910 3559.070 1149.910 ;
        RECT 3358.100 1135.910 3553.000 1141.910 ;
        RECT 3429.620 1127.500 3500.040 1133.500 ;
        RECT 3396.670 1119.500 3494.070 1125.500 ;
        RECT 89.140 1084.500 158.310 1090.500 ;
        RECT 95.110 1076.500 191.260 1082.500 ;
        RECT 3376.380 918.910 3559.070 924.910 ;
        RECT 3358.100 910.910 3553.000 916.910 ;
        RECT 3429.620 902.500 3500.040 908.500 ;
        RECT 3396.670 894.500 3494.070 900.500 ;
        RECT 3376.380 692.910 3559.070 698.910 ;
        RECT 3358.100 684.910 3553.000 690.910 ;
        RECT 3429.620 676.500 3500.040 682.500 ;
        RECT 3396.670 668.500 3494.070 674.500 ;
        RECT 730.965 209.380 732.815 211.400 ;
        RECT 736.940 209.835 746.570 210.455 ;
        RECT 2202.265 209.980 2202.585 210.300 ;
        RECT 2202.665 209.980 2202.985 210.300 ;
        RECT 2203.065 209.980 2203.385 210.300 ;
        RECT 2203.465 209.980 2203.785 210.300 ;
        RECT 643.050 169.500 647.340 208.000 ;
        RECT 730.965 207.390 740.895 209.380 ;
        RECT 650.710 175.570 655.000 204.610 ;
        RECT 738.975 186.505 740.900 203.515 ;
        RECT 2130.090 154.030 2131.995 203.810 ;
        RECT 2135.095 186.700 2137.000 205.790 ;
        RECT 2208.015 202.820 2210.045 203.885 ;
        RECT 2281.685 186.700 2283.590 203.810 ;
        RECT 2286.695 154.030 2288.600 203.810 ;
        RECT 3209.770 169.600 3218.470 220.130 ;
        RECT 3267.310 179.040 3284.550 225.780 ;
      LAYER via3 ;
        RECT 557.750 5095.525 563.270 5099.045 ;
        RECT 549.760 5089.505 555.280 5093.025 ;
        RECT 814.750 5095.525 820.270 5099.045 ;
        RECT 557.905 5030.145 563.025 5033.665 ;
        RECT 806.760 5089.505 812.280 5093.025 ;
        RECT 550.050 4997.435 555.170 5000.955 ;
        RECT 1071.750 5095.525 1077.270 5099.045 ;
        RECT 1063.760 5089.505 1069.280 5093.025 ;
        RECT 814.905 5030.145 820.025 5033.665 ;
        RECT 843.255 5029.885 844.375 5033.405 ;
        RECT 807.050 4997.435 812.170 5000.955 ;
        RECT 849.235 4997.440 850.355 5000.960 ;
        RECT 1328.750 5095.525 1334.270 5099.045 ;
        RECT 1071.905 5030.145 1077.025 5033.665 ;
        RECT 1320.760 5089.505 1326.280 5093.025 ;
        RECT 1064.050 4997.435 1069.170 5000.955 ;
        RECT 1586.750 5095.525 1592.270 5099.045 ;
        RECT 1328.905 5030.145 1334.025 5033.665 ;
        RECT 1578.760 5089.505 1584.280 5093.025 ;
        RECT 1321.050 4997.435 1326.170 5000.955 ;
        RECT 1838.750 5095.525 1844.270 5099.045 ;
        RECT 1586.905 5030.145 1592.025 5033.665 ;
        RECT 1830.760 5089.505 1836.280 5093.025 ;
        RECT 1579.050 4997.435 1584.170 5000.955 ;
        RECT 2175.750 5095.525 2181.270 5099.045 ;
        RECT 2167.760 5089.505 2173.280 5093.025 ;
        RECT 1838.905 5030.145 1844.025 5033.665 ;
        RECT 2085.440 5029.885 2086.560 5033.405 ;
        RECT 1831.050 4997.435 1836.170 5000.955 ;
        RECT 2091.420 4997.435 2092.540 5000.955 ;
        RECT 2560.750 5095.525 2566.270 5099.045 ;
        RECT 2175.905 5030.145 2181.025 5033.665 ;
        RECT 2552.760 5089.505 2558.280 5093.025 ;
        RECT 2168.050 4997.435 2173.170 5000.955 ;
        RECT 2817.750 5095.525 2823.270 5099.045 ;
        RECT 2560.905 5030.145 2566.025 5033.665 ;
        RECT 2809.760 5089.505 2815.280 5093.025 ;
        RECT 2553.050 4997.435 2558.170 5000.955 ;
        RECT 2817.905 5030.145 2823.025 5033.665 ;
        RECT 3318.490 5029.885 3319.610 5033.405 ;
        RECT 2810.050 4997.435 2815.170 5000.955 ;
        RECT 3324.470 4997.435 3325.590 5000.955 ;
        RECT 221.570 4759.955 233.490 4765.075 ;
        RECT 307.305 4759.840 309.625 4765.360 ;
        RECT 205.520 4752.045 217.440 4757.165 ;
        RECT 302.485 4751.880 304.805 4757.400 ;
        RECT 89.545 4727.750 93.065 4733.270 ;
        RECT 154.225 4727.905 157.745 4733.025 ;
        RECT 3253.280 4726.165 3256.000 4731.685 ;
        RECT 3377.135 4726.425 3382.255 4731.545 ;
        RECT 3555.060 4726.145 3558.180 4731.665 ;
        RECT 95.565 4719.760 99.085 4725.280 ;
        RECT 186.935 4720.050 190.455 4725.170 ;
        RECT 3258.070 4718.145 3260.790 4723.665 ;
        RECT 3358.605 4718.335 3363.725 4723.455 ;
        RECT 3549.070 4718.165 3552.190 4723.685 ;
        RECT 3430.135 4709.905 3433.655 4715.025 ;
        RECT 3496.065 4709.750 3499.585 4715.270 ;
        RECT 3397.425 4702.050 3400.945 4707.170 ;
        RECT 3490.045 4701.760 3493.565 4707.280 ;
        RECT 3253.280 4500.165 3256.000 4505.685 ;
        RECT 3373.825 4500.405 3378.545 4505.525 ;
        RECT 3258.070 4492.145 3260.790 4497.665 ;
        RECT 3357.845 4492.365 3362.965 4497.485 ;
        RECT 154.235 4447.440 157.755 4448.560 ;
        RECT 186.935 4441.455 190.455 4442.575 ;
        RECT 3253.280 4275.165 3256.000 4280.685 ;
        RECT 3370.680 4275.360 3375.800 4280.480 ;
        RECT 3258.070 4267.145 3260.790 4272.665 ;
        RECT 3357.960 4267.350 3363.080 4272.470 ;
        RECT 221.570 4130.955 233.490 4136.075 ;
        RECT 307.305 4130.840 309.625 4136.360 ;
        RECT 205.520 4123.045 217.440 4128.165 ;
        RECT 302.485 4122.880 304.805 4128.400 ;
        RECT 89.545 4098.750 93.065 4104.270 ;
        RECT 154.225 4098.905 157.745 4104.025 ;
        RECT 95.565 4090.760 99.085 4096.280 ;
        RECT 186.935 4091.050 190.455 4096.170 ;
        RECT 221.570 3922.955 233.490 3928.075 ;
        RECT 307.305 3922.840 309.625 3928.360 ;
        RECT 205.520 3915.045 217.440 3920.165 ;
        RECT 302.485 3914.880 304.805 3920.400 ;
        RECT 89.545 3882.750 93.065 3888.270 ;
        RECT 154.225 3882.905 157.745 3888.025 ;
        RECT 95.565 3874.760 99.085 3880.280 ;
        RECT 186.935 3875.050 190.455 3880.170 ;
        RECT 3253.280 3834.165 3256.000 3839.685 ;
        RECT 3377.185 3834.425 3382.305 3839.545 ;
        RECT 3555.110 3834.145 3558.230 3839.665 ;
        RECT 3258.070 3826.145 3260.790 3831.665 ;
        RECT 3358.655 3826.335 3363.775 3831.455 ;
        RECT 3549.120 3826.165 3552.240 3831.685 ;
        RECT 3430.185 3817.905 3433.705 3823.025 ;
        RECT 3496.115 3817.750 3499.635 3823.270 ;
        RECT 3397.475 3810.050 3400.995 3815.170 ;
        RECT 3490.095 3809.760 3493.615 3815.280 ;
        RECT 221.570 3698.955 233.490 3704.075 ;
        RECT 307.305 3698.840 309.625 3704.360 ;
        RECT 205.520 3691.045 217.440 3696.165 ;
        RECT 302.485 3690.880 304.805 3696.400 ;
        RECT 89.545 3666.750 93.065 3672.270 ;
        RECT 154.225 3666.905 157.745 3672.025 ;
        RECT 95.565 3658.760 99.085 3664.280 ;
        RECT 186.935 3659.050 190.455 3664.170 ;
        RECT 3429.885 3622.840 3433.405 3623.960 ;
        RECT 3397.435 3616.860 3400.955 3617.980 ;
        RECT 3253.280 3609.165 3256.000 3614.685 ;
        RECT 3377.185 3609.425 3382.305 3614.545 ;
        RECT 3555.110 3609.145 3558.230 3614.665 ;
        RECT 3258.070 3601.145 3260.790 3606.665 ;
        RECT 3358.655 3601.335 3363.775 3606.455 ;
        RECT 3549.120 3601.165 3552.240 3606.685 ;
        RECT 3430.185 3592.905 3433.705 3598.025 ;
        RECT 3496.115 3592.750 3499.635 3598.270 ;
        RECT 3397.475 3585.050 3400.995 3590.170 ;
        RECT 3490.095 3584.760 3493.615 3590.280 ;
        RECT 221.570 3482.955 233.490 3488.075 ;
        RECT 307.305 3482.840 309.625 3488.360 ;
        RECT 205.520 3475.045 217.440 3480.165 ;
        RECT 302.485 3474.880 304.805 3480.400 ;
        RECT 89.545 3450.750 93.065 3456.270 ;
        RECT 154.225 3450.905 157.745 3456.025 ;
        RECT 95.565 3442.760 99.085 3448.280 ;
        RECT 186.935 3443.050 190.455 3448.170 ;
        RECT 3253.280 3383.165 3256.000 3388.685 ;
        RECT 3377.185 3383.425 3382.305 3388.545 ;
        RECT 3555.110 3383.145 3558.230 3388.665 ;
        RECT 3258.070 3375.145 3260.790 3380.665 ;
        RECT 3358.655 3375.335 3363.775 3380.455 ;
        RECT 3549.120 3375.165 3552.240 3380.685 ;
        RECT 3430.185 3366.905 3433.705 3372.025 ;
        RECT 3496.115 3366.750 3499.635 3372.270 ;
        RECT 3397.475 3359.050 3400.995 3364.170 ;
        RECT 3490.095 3358.760 3493.615 3364.280 ;
        RECT 221.570 3266.955 233.490 3272.075 ;
        RECT 307.305 3266.840 309.625 3272.360 ;
        RECT 205.520 3259.045 217.440 3264.165 ;
        RECT 302.485 3258.880 304.805 3264.400 ;
        RECT 89.545 3234.750 93.065 3240.270 ;
        RECT 154.225 3234.905 157.745 3240.025 ;
        RECT 95.565 3226.760 99.085 3232.280 ;
        RECT 186.935 3227.050 190.455 3232.170 ;
        RECT 3253.280 3158.165 3256.000 3163.685 ;
        RECT 3377.185 3158.425 3382.305 3163.545 ;
        RECT 3555.110 3158.145 3558.230 3163.665 ;
        RECT 3358.655 3150.335 3363.775 3155.455 ;
        RECT 3549.120 3150.165 3552.240 3155.685 ;
        RECT 3258.070 3144.145 3260.790 3149.665 ;
        RECT 3430.185 3141.905 3433.705 3147.025 ;
        RECT 3496.115 3141.750 3499.635 3147.270 ;
        RECT 3397.475 3134.050 3400.995 3139.170 ;
        RECT 3490.095 3133.760 3493.615 3139.280 ;
        RECT 221.570 3056.255 233.490 3061.375 ;
        RECT 307.305 3056.140 309.625 3061.660 ;
        RECT 205.520 3048.345 217.440 3053.465 ;
        RECT 302.485 3048.180 304.805 3053.700 ;
        RECT 89.545 3018.750 93.065 3024.270 ;
        RECT 154.225 3018.905 157.745 3024.025 ;
        RECT 95.565 3010.760 99.085 3016.280 ;
        RECT 186.935 3011.050 190.455 3016.170 ;
        RECT 3253.280 2932.165 3256.000 2937.685 ;
        RECT 3377.185 2932.425 3382.305 2937.545 ;
        RECT 3555.110 2932.145 3558.230 2937.665 ;
        RECT 3258.070 2924.145 3260.790 2929.665 ;
        RECT 3358.655 2924.335 3363.775 2929.455 ;
        RECT 3549.120 2924.165 3552.240 2929.685 ;
        RECT 3430.185 2915.905 3433.705 2921.025 ;
        RECT 3496.115 2915.750 3499.635 2921.270 ;
        RECT 3397.475 2908.050 3400.995 2913.170 ;
        RECT 3490.095 2907.760 3493.615 2913.280 ;
        RECT 221.570 2834.955 233.490 2840.075 ;
        RECT 307.305 2834.840 309.625 2840.360 ;
        RECT 205.520 2827.045 217.440 2832.165 ;
        RECT 302.485 2826.880 304.805 2832.400 ;
        RECT 89.545 2802.750 93.065 2808.270 ;
        RECT 154.225 2802.905 157.745 2808.025 ;
        RECT 95.565 2794.760 99.085 2800.280 ;
        RECT 186.935 2795.050 190.455 2800.170 ;
        RECT 3253.280 2707.165 3256.000 2712.685 ;
        RECT 3377.185 2707.425 3382.305 2712.545 ;
        RECT 3555.110 2707.145 3558.230 2712.665 ;
        RECT 3258.070 2699.145 3260.790 2704.665 ;
        RECT 3358.655 2699.335 3363.775 2704.455 ;
        RECT 3549.120 2699.165 3552.240 2704.685 ;
        RECT 3430.185 2690.905 3433.705 2696.025 ;
        RECT 3496.115 2690.750 3499.635 2696.270 ;
        RECT 3397.475 2683.050 3400.995 2688.170 ;
        RECT 3490.095 2682.760 3493.615 2688.280 ;
        RECT 3253.280 2490.165 3256.000 2495.685 ;
        RECT 3377.185 2487.425 3382.305 2492.545 ;
        RECT 3555.110 2487.145 3558.230 2492.665 ;
        RECT 3258.070 2479.145 3260.790 2484.665 ;
        RECT 3358.655 2479.335 3363.775 2484.455 ;
        RECT 3549.120 2479.165 3552.240 2484.685 ;
        RECT 3430.185 2470.905 3433.705 2476.025 ;
        RECT 3496.115 2470.750 3499.635 2476.270 ;
        RECT 3397.475 2463.050 3400.995 2468.170 ;
        RECT 3490.095 2462.760 3493.615 2468.280 ;
        RECT 3429.885 2240.835 3433.405 2241.955 ;
        RECT 3397.435 2234.855 3400.955 2235.975 ;
        RECT 221.570 2196.955 233.490 2202.075 ;
        RECT 307.305 2196.840 309.625 2202.360 ;
        RECT 205.520 2189.045 217.440 2194.165 ;
        RECT 302.485 2188.880 304.805 2194.400 ;
        RECT 89.545 2164.750 93.065 2170.270 ;
        RECT 154.225 2164.905 157.745 2170.025 ;
        RECT 95.565 2156.760 99.085 2162.280 ;
        RECT 186.935 2157.050 190.455 2162.170 ;
        RECT 3253.280 2046.165 3256.000 2051.685 ;
        RECT 3377.185 2046.425 3382.305 2051.545 ;
        RECT 3555.110 2046.145 3558.230 2051.665 ;
        RECT 3258.070 2038.145 3260.790 2043.665 ;
        RECT 3358.655 2038.335 3363.775 2043.455 ;
        RECT 3549.120 2038.165 3552.240 2043.685 ;
        RECT 3430.185 2029.905 3433.705 2035.025 ;
        RECT 3496.115 2029.750 3499.635 2035.270 ;
        RECT 3397.475 2022.050 3400.995 2027.170 ;
        RECT 3490.095 2021.760 3493.615 2027.280 ;
        RECT 221.570 1980.955 233.490 1986.075 ;
        RECT 307.305 1980.840 309.625 1986.360 ;
        RECT 205.520 1973.045 217.440 1978.165 ;
        RECT 302.485 1972.880 304.805 1978.400 ;
        RECT 89.545 1948.750 93.065 1954.270 ;
        RECT 154.225 1948.905 157.745 1954.025 ;
        RECT 95.565 1940.760 99.085 1946.280 ;
        RECT 186.935 1941.050 190.455 1946.170 ;
        RECT 3253.280 1827.165 3256.000 1832.685 ;
        RECT 3377.185 1820.425 3382.305 1825.545 ;
        RECT 3555.110 1820.145 3558.230 1825.665 ;
        RECT 3258.070 1812.145 3260.790 1817.665 ;
        RECT 3358.655 1812.335 3363.775 1817.455 ;
        RECT 3549.120 1812.165 3552.240 1817.685 ;
        RECT 3430.185 1803.905 3433.705 1809.025 ;
        RECT 3496.115 1803.750 3499.635 1809.270 ;
        RECT 3397.475 1796.050 3400.995 1801.170 ;
        RECT 3490.095 1795.760 3493.615 1801.280 ;
        RECT 221.570 1769.955 233.490 1775.075 ;
        RECT 307.305 1769.840 309.625 1775.360 ;
        RECT 205.520 1762.045 217.440 1767.165 ;
        RECT 302.485 1761.880 304.805 1767.400 ;
        RECT 89.545 1732.750 93.065 1738.270 ;
        RECT 154.225 1732.905 157.745 1738.025 ;
        RECT 95.565 1724.760 99.085 1730.280 ;
        RECT 186.935 1725.050 190.455 1730.170 ;
        RECT 3253.280 1595.165 3256.000 1600.685 ;
        RECT 3377.185 1595.425 3382.305 1600.545 ;
        RECT 3555.110 1595.145 3558.230 1600.665 ;
        RECT 3258.070 1587.145 3260.790 1592.665 ;
        RECT 3358.655 1587.335 3363.775 1592.455 ;
        RECT 3549.120 1587.165 3552.240 1592.685 ;
        RECT 3430.185 1578.905 3433.705 1584.025 ;
        RECT 3496.115 1578.750 3499.635 1584.270 ;
        RECT 3397.475 1571.050 3400.995 1576.170 ;
        RECT 3490.095 1570.760 3493.615 1576.280 ;
        RECT 221.570 1548.955 233.490 1554.075 ;
        RECT 307.305 1548.840 309.625 1554.360 ;
        RECT 205.520 1541.045 217.440 1546.165 ;
        RECT 302.485 1540.880 304.805 1546.400 ;
        RECT 89.545 1516.750 93.065 1522.270 ;
        RECT 154.225 1516.905 157.745 1522.025 ;
        RECT 95.565 1508.760 99.085 1514.280 ;
        RECT 186.935 1509.050 190.455 1514.170 ;
        RECT 3377.185 1370.425 3382.305 1375.545 ;
        RECT 3555.110 1370.145 3558.230 1375.665 ;
        RECT 3358.655 1362.335 3363.775 1367.455 ;
        RECT 3549.120 1362.165 3552.240 1367.685 ;
        RECT 3430.185 1353.905 3433.705 1359.025 ;
        RECT 3496.115 1353.750 3499.635 1359.270 ;
        RECT 3397.475 1346.050 3400.995 1351.170 ;
        RECT 3490.095 1345.760 3493.615 1351.280 ;
        RECT 89.545 1300.750 93.065 1306.270 ;
        RECT 154.225 1300.905 157.745 1306.025 ;
        RECT 95.565 1292.760 99.085 1298.280 ;
        RECT 186.935 1293.050 190.455 1298.170 ;
        RECT 3377.185 1144.425 3382.305 1149.545 ;
        RECT 3555.110 1144.145 3558.230 1149.665 ;
        RECT 3358.655 1136.335 3363.775 1141.455 ;
        RECT 3549.120 1136.165 3552.240 1141.685 ;
        RECT 3430.185 1127.905 3433.705 1133.025 ;
        RECT 3496.115 1127.750 3499.635 1133.270 ;
        RECT 3397.475 1120.050 3400.995 1125.170 ;
        RECT 3490.095 1119.760 3493.615 1125.280 ;
        RECT 89.545 1084.750 93.065 1090.270 ;
        RECT 154.225 1084.905 157.745 1090.025 ;
        RECT 95.565 1076.760 99.085 1082.280 ;
        RECT 186.935 1077.050 190.455 1082.170 ;
        RECT 3377.185 919.425 3382.305 924.545 ;
        RECT 3555.110 919.145 3558.230 924.665 ;
        RECT 3358.655 911.335 3363.775 916.455 ;
        RECT 3549.120 911.165 3552.240 916.685 ;
        RECT 3430.185 902.905 3433.705 908.025 ;
        RECT 3496.115 902.750 3499.635 908.270 ;
        RECT 3397.475 895.050 3400.995 900.170 ;
        RECT 3490.095 894.760 3493.615 900.280 ;
        RECT 3377.185 693.425 3382.305 698.545 ;
        RECT 3555.110 693.145 3558.230 698.665 ;
        RECT 3358.655 685.335 3363.775 690.455 ;
        RECT 3549.120 685.165 3552.240 690.685 ;
        RECT 3430.185 676.905 3433.705 682.025 ;
        RECT 3496.115 676.750 3499.635 682.270 ;
        RECT 3397.475 669.050 3400.995 674.170 ;
        RECT 3490.095 668.760 3493.615 674.280 ;
        RECT 3209.975 211.105 3218.295 219.825 ;
        RECT 745.760 210.055 746.080 210.375 ;
        RECT 746.160 210.055 746.480 210.375 ;
        RECT 643.235 206.790 647.155 207.910 ;
        RECT 739.180 207.640 740.700 209.160 ;
        RECT 2135.295 204.980 2136.815 205.700 ;
        RECT 650.895 203.000 654.815 204.120 ;
        RECT 739.170 200.545 740.690 203.265 ;
        RECT 739.180 186.850 740.700 190.770 ;
        RECT 2130.290 203.000 2131.810 203.720 ;
        RECT 650.910 175.945 654.830 179.865 ;
        RECT 643.260 169.905 647.180 173.825 ;
        RECT 2208.265 203.000 2209.785 203.720 ;
        RECT 2135.285 187.050 2136.805 190.570 ;
        RECT 2281.885 200.080 2283.405 203.600 ;
        RECT 2281.885 187.050 2283.405 190.570 ;
        RECT 2286.890 200.080 2288.410 203.600 ;
        RECT 2130.280 154.380 2131.800 157.900 ;
        RECT 3267.915 213.190 3283.835 225.110 ;
        RECT 3210.190 170.110 3218.110 173.630 ;
        RECT 2286.890 154.380 2288.410 157.900 ;
      LAYER met4 ;
        RECT 500.110 5095.240 563.550 5099.240 ;
        RECT 757.110 5095.240 820.550 5099.240 ;
        RECT 1014.110 5095.240 1077.550 5099.240 ;
        RECT 1271.110 5095.240 1334.550 5099.240 ;
        RECT 1529.110 5095.240 1592.550 5099.240 ;
        RECT 1781.110 5095.240 1844.550 5099.240 ;
        RECT 2118.110 5095.240 2181.550 5099.240 ;
        RECT 2503.110 5095.240 2566.550 5099.240 ;
        RECT 2760.110 5095.240 2823.550 5099.240 ;
        RECT 491.740 5089.240 556.660 5093.240 ;
        RECT 748.740 5089.240 813.660 5093.240 ;
        RECT 1005.740 5089.240 1070.660 5093.240 ;
        RECT 1262.740 5089.240 1327.660 5093.240 ;
        RECT 1520.740 5089.240 1585.660 5093.240 ;
        RECT 1772.740 5089.240 1837.660 5093.240 ;
        RECT 2109.740 5089.240 2174.660 5093.240 ;
        RECT 2494.740 5089.240 2559.660 5093.240 ;
        RECT 2751.740 5089.240 2816.660 5093.240 ;
        RECT 557.770 5030.020 563.160 5033.790 ;
        RECT 814.770 5030.020 820.160 5033.790 ;
        RECT 843.255 5029.885 844.375 5033.405 ;
        RECT 1071.770 5030.020 1077.160 5033.790 ;
        RECT 1328.770 5030.020 1334.160 5033.790 ;
        RECT 1586.770 5030.020 1592.160 5033.790 ;
        RECT 1838.770 5030.020 1844.160 5033.790 ;
        RECT 2085.440 5029.885 2086.560 5033.405 ;
        RECT 2175.770 5030.020 2181.160 5033.790 ;
        RECT 2560.770 5030.020 2566.160 5033.790 ;
        RECT 2817.770 5030.020 2823.160 5033.790 ;
        RECT 3318.490 5029.885 3319.610 5033.405 ;
        RECT 549.900 4997.290 555.320 5001.100 ;
        RECT 806.900 4997.290 812.320 5001.100 ;
        RECT 849.235 4997.440 850.355 5000.960 ;
        RECT 1063.900 4997.290 1069.320 5001.100 ;
        RECT 1320.900 4997.290 1326.320 5001.100 ;
        RECT 1578.900 4997.290 1584.320 5001.100 ;
        RECT 1830.900 4997.290 1836.320 5001.100 ;
        RECT 2091.420 4997.435 2092.540 5000.955 ;
        RECT 2167.900 4997.290 2173.320 5001.100 ;
        RECT 2552.900 4997.290 2558.320 5001.100 ;
        RECT 2809.900 4997.290 2815.320 5001.100 ;
        RECT 3324.470 4997.435 3325.590 5000.955 ;
        RECT 204.965 4929.270 282.070 4932.340 ;
        RECT 221.000 4924.370 282.200 4927.630 ;
        RECT 3291.580 4919.640 3367.150 4922.850 ;
        RECT 3291.440 4914.800 3383.120 4918.010 ;
        RECT 221.000 4759.610 233.960 4765.630 ;
        RECT 307.120 4759.800 309.810 4765.400 ;
        RECT 204.970 4751.630 217.940 4757.610 ;
        RECT 302.300 4751.840 304.990 4757.440 ;
        RECT 89.350 4670.110 93.350 4733.550 ;
        RECT 154.100 4727.770 157.870 4733.160 ;
        RECT 95.350 4661.740 99.350 4726.660 ;
        RECT 3253.270 4726.120 3256.010 4731.730 ;
        RECT 3376.680 4725.870 3382.710 4731.940 ;
        RECT 186.790 4719.900 190.600 4725.320 ;
        RECT 3258.010 4718.060 3260.850 4723.750 ;
        RECT 3358.200 4717.870 3364.230 4723.940 ;
        RECT 3430.010 4709.770 3433.780 4715.160 ;
        RECT 3397.280 4701.900 3401.090 4707.320 ;
        RECT 3489.780 4643.740 3493.780 4708.660 ;
        RECT 3495.780 4652.110 3499.780 4715.550 ;
        RECT 3548.600 4657.380 3552.600 4724.210 ;
        RECT 3554.600 4648.730 3558.600 4732.350 ;
        RECT 3253.270 4500.120 3256.010 4505.730 ;
        RECT 3373.150 4499.910 3379.150 4505.910 ;
        RECT 3258.010 4492.060 3260.850 4497.750 ;
        RECT 3357.380 4491.910 3363.380 4497.910 ;
        RECT 154.235 4447.440 157.755 4448.560 ;
        RECT 186.935 4441.455 190.455 4442.575 ;
        RECT 3253.270 4275.120 3256.010 4280.730 ;
        RECT 3370.270 4274.910 3376.270 4280.910 ;
        RECT 3258.010 4267.060 3260.850 4272.750 ;
        RECT 3357.540 4266.910 3363.540 4272.910 ;
        RECT 221.000 4130.610 233.960 4136.630 ;
        RECT 307.120 4130.800 309.810 4136.400 ;
        RECT 204.970 4122.630 217.940 4128.610 ;
        RECT 302.300 4122.840 304.990 4128.440 ;
        RECT 89.350 4041.110 93.350 4104.550 ;
        RECT 154.100 4098.770 157.870 4104.160 ;
        RECT 95.350 4032.740 99.350 4097.660 ;
        RECT 186.790 4090.900 190.600 4096.320 ;
        RECT 221.000 3922.610 233.960 3928.630 ;
        RECT 307.120 3922.800 309.810 3928.400 ;
        RECT 204.970 3914.630 217.940 3920.610 ;
        RECT 302.300 3914.840 304.990 3920.440 ;
        RECT 89.350 3825.110 93.350 3888.550 ;
        RECT 154.100 3882.770 157.870 3888.160 ;
        RECT 95.350 3816.740 99.350 3881.660 ;
        RECT 186.790 3874.900 190.600 3880.320 ;
        RECT 3253.270 3834.120 3256.010 3839.730 ;
        RECT 3376.730 3833.870 3382.760 3839.940 ;
        RECT 3258.010 3826.060 3260.850 3831.750 ;
        RECT 3358.250 3825.870 3364.280 3831.940 ;
        RECT 3430.060 3817.770 3433.830 3823.160 ;
        RECT 3397.330 3809.900 3401.140 3815.320 ;
        RECT 3489.830 3751.740 3493.830 3816.660 ;
        RECT 3495.830 3760.110 3499.830 3823.550 ;
        RECT 3548.650 3765.380 3552.650 3832.210 ;
        RECT 3554.650 3756.730 3558.650 3840.350 ;
        RECT 221.000 3698.610 233.960 3704.630 ;
        RECT 307.120 3698.800 309.810 3704.400 ;
        RECT 204.970 3690.630 217.940 3696.610 ;
        RECT 302.300 3690.840 304.990 3696.440 ;
        RECT 89.350 3609.110 93.350 3672.550 ;
        RECT 154.100 3666.770 157.870 3672.160 ;
        RECT 95.350 3600.740 99.350 3665.660 ;
        RECT 186.790 3658.900 190.600 3664.320 ;
        RECT 3429.885 3622.840 3433.405 3623.960 ;
        RECT 3397.435 3616.860 3400.955 3617.980 ;
        RECT 3253.270 3609.120 3256.010 3614.730 ;
        RECT 3376.730 3608.870 3382.760 3614.940 ;
        RECT 3258.010 3601.060 3260.850 3606.750 ;
        RECT 3358.250 3600.870 3364.280 3606.940 ;
        RECT 3430.060 3592.770 3433.830 3598.160 ;
        RECT 3397.330 3584.900 3401.140 3590.320 ;
        RECT 3489.830 3526.740 3493.830 3591.660 ;
        RECT 3495.830 3535.110 3499.830 3598.550 ;
        RECT 3548.650 3540.380 3552.650 3607.210 ;
        RECT 3554.650 3531.730 3558.650 3615.350 ;
        RECT 221.000 3482.610 233.960 3488.630 ;
        RECT 307.120 3482.800 309.810 3488.400 ;
        RECT 204.970 3474.630 217.940 3480.610 ;
        RECT 302.300 3474.840 304.990 3480.440 ;
        RECT 89.350 3393.110 93.350 3456.550 ;
        RECT 154.100 3450.770 157.870 3456.160 ;
        RECT 95.350 3384.740 99.350 3449.660 ;
        RECT 186.790 3442.900 190.600 3448.320 ;
        RECT 3253.270 3383.120 3256.010 3388.730 ;
        RECT 3376.730 3382.870 3382.760 3388.940 ;
        RECT 3258.010 3375.060 3260.850 3380.750 ;
        RECT 3358.250 3374.870 3364.280 3380.940 ;
        RECT 3430.060 3366.770 3433.830 3372.160 ;
        RECT 3397.330 3358.900 3401.140 3364.320 ;
        RECT 3489.830 3300.740 3493.830 3365.660 ;
        RECT 3495.830 3309.110 3499.830 3372.550 ;
        RECT 3548.650 3314.380 3552.650 3381.210 ;
        RECT 3554.650 3305.730 3558.650 3389.350 ;
        RECT 221.000 3266.610 233.960 3272.630 ;
        RECT 307.120 3266.800 309.810 3272.400 ;
        RECT 204.970 3258.630 217.940 3264.610 ;
        RECT 302.300 3258.840 304.990 3264.440 ;
        RECT 89.350 3177.110 93.350 3240.550 ;
        RECT 154.100 3234.770 157.870 3240.160 ;
        RECT 95.350 3168.740 99.350 3233.660 ;
        RECT 186.790 3226.900 190.600 3232.320 ;
        RECT 3253.270 3158.120 3256.010 3163.730 ;
        RECT 3376.730 3157.870 3382.760 3163.940 ;
        RECT 3358.250 3149.870 3364.280 3155.940 ;
        RECT 3258.010 3144.060 3260.850 3149.750 ;
        RECT 3430.060 3141.770 3433.830 3147.160 ;
        RECT 3397.330 3133.900 3401.140 3139.320 ;
        RECT 3489.830 3075.740 3493.830 3140.660 ;
        RECT 3495.830 3084.110 3499.830 3147.550 ;
        RECT 3548.650 3089.380 3552.650 3156.210 ;
        RECT 3554.650 3080.730 3558.650 3164.350 ;
        RECT 221.000 3055.910 233.960 3061.930 ;
        RECT 307.120 3056.100 309.810 3061.700 ;
        RECT 204.970 3047.930 217.940 3053.910 ;
        RECT 302.300 3048.140 304.990 3053.740 ;
        RECT 89.350 2961.110 93.350 3024.550 ;
        RECT 154.100 3018.770 157.870 3024.160 ;
        RECT 95.350 2952.740 99.350 3017.660 ;
        RECT 186.790 3010.900 190.600 3016.320 ;
        RECT 3253.270 2932.120 3256.010 2937.730 ;
        RECT 3376.730 2931.870 3382.760 2937.940 ;
        RECT 3258.010 2924.060 3260.850 2929.750 ;
        RECT 3358.250 2923.870 3364.280 2929.940 ;
        RECT 3430.060 2915.770 3433.830 2921.160 ;
        RECT 3397.330 2907.900 3401.140 2913.320 ;
        RECT 3489.830 2849.740 3493.830 2914.660 ;
        RECT 3495.830 2858.110 3499.830 2921.550 ;
        RECT 3548.650 2863.380 3552.650 2930.210 ;
        RECT 3554.650 2854.730 3558.650 2938.350 ;
        RECT 221.000 2834.610 233.960 2840.630 ;
        RECT 307.120 2834.800 309.810 2840.400 ;
        RECT 204.970 2826.630 217.940 2832.610 ;
        RECT 302.300 2826.840 304.990 2832.440 ;
        RECT 89.350 2745.110 93.350 2808.550 ;
        RECT 154.100 2802.770 157.870 2808.160 ;
        RECT 95.350 2736.740 99.350 2801.660 ;
        RECT 186.790 2794.900 190.600 2800.320 ;
        RECT 3253.270 2707.120 3256.010 2712.730 ;
        RECT 3376.730 2706.870 3382.760 2712.940 ;
        RECT 3258.010 2699.060 3260.850 2704.750 ;
        RECT 3358.250 2698.870 3364.280 2704.940 ;
        RECT 3430.060 2690.770 3433.830 2696.160 ;
        RECT 3397.330 2682.900 3401.140 2688.320 ;
        RECT 3489.830 2624.740 3493.830 2689.660 ;
        RECT 3495.830 2633.110 3499.830 2696.550 ;
        RECT 3548.650 2638.380 3552.650 2705.210 ;
        RECT 3554.650 2629.730 3558.650 2713.350 ;
        RECT 3253.270 2490.120 3256.010 2495.730 ;
        RECT 3376.730 2486.870 3382.760 2492.940 ;
        RECT 3258.010 2479.060 3260.850 2484.750 ;
        RECT 3358.250 2478.870 3364.280 2484.940 ;
        RECT 3430.060 2470.770 3433.830 2476.160 ;
        RECT 3397.330 2462.900 3401.140 2468.320 ;
        RECT 3489.830 2404.740 3493.830 2469.660 ;
        RECT 3495.830 2413.110 3499.830 2476.550 ;
        RECT 3548.650 2418.380 3552.650 2485.210 ;
        RECT 3554.650 2409.730 3558.650 2493.350 ;
        RECT 3429.885 2240.835 3433.405 2241.955 ;
        RECT 3397.435 2234.855 3400.955 2235.975 ;
        RECT 221.000 2196.610 233.960 2202.630 ;
        RECT 307.120 2196.800 309.810 2202.400 ;
        RECT 204.970 2188.630 217.940 2194.610 ;
        RECT 302.300 2188.840 304.990 2194.440 ;
        RECT 89.350 2107.110 93.350 2170.550 ;
        RECT 154.100 2164.770 157.870 2170.160 ;
        RECT 95.350 2098.740 99.350 2163.660 ;
        RECT 186.790 2156.900 190.600 2162.320 ;
        RECT 3253.270 2046.120 3256.010 2051.730 ;
        RECT 3376.730 2045.870 3382.760 2051.940 ;
        RECT 3258.010 2038.060 3260.850 2043.750 ;
        RECT 3358.250 2037.870 3364.280 2043.940 ;
        RECT 3430.060 2029.770 3433.830 2035.160 ;
        RECT 3397.330 2021.900 3401.140 2027.320 ;
        RECT 221.000 1980.610 233.960 1986.630 ;
        RECT 307.120 1980.800 309.810 1986.400 ;
        RECT 204.970 1972.630 217.940 1978.610 ;
        RECT 302.300 1972.840 304.990 1978.440 ;
        RECT 3489.830 1963.740 3493.830 2028.660 ;
        RECT 3495.830 1972.110 3499.830 2035.550 ;
        RECT 3548.650 1977.380 3552.650 2044.210 ;
        RECT 3554.650 1968.730 3558.650 2052.350 ;
        RECT 89.350 1891.110 93.350 1954.550 ;
        RECT 154.100 1948.770 157.870 1954.160 ;
        RECT 95.350 1882.740 99.350 1947.660 ;
        RECT 186.790 1940.900 190.600 1946.320 ;
        RECT 3253.270 1827.120 3256.010 1832.730 ;
        RECT 3376.730 1819.870 3382.760 1825.940 ;
        RECT 3258.010 1812.060 3260.850 1817.750 ;
        RECT 3358.250 1811.870 3364.280 1817.940 ;
        RECT 3430.060 1803.770 3433.830 1809.160 ;
        RECT 3397.330 1795.900 3401.140 1801.320 ;
        RECT 221.000 1769.610 233.960 1775.630 ;
        RECT 307.120 1769.800 309.810 1775.400 ;
        RECT 204.970 1761.630 217.940 1767.610 ;
        RECT 302.300 1761.840 304.990 1767.440 ;
        RECT 89.350 1675.110 93.350 1738.550 ;
        RECT 154.100 1732.770 157.870 1738.160 ;
        RECT 3489.830 1737.740 3493.830 1802.660 ;
        RECT 3495.830 1746.110 3499.830 1809.550 ;
        RECT 3548.650 1751.380 3552.650 1818.210 ;
        RECT 3554.650 1742.730 3558.650 1826.350 ;
        RECT 95.350 1666.740 99.350 1731.660 ;
        RECT 186.790 1724.900 190.600 1730.320 ;
        RECT 3253.270 1595.120 3256.010 1600.730 ;
        RECT 3376.730 1594.870 3382.760 1600.940 ;
        RECT 3258.010 1587.060 3260.850 1592.750 ;
        RECT 3358.250 1586.870 3364.280 1592.940 ;
        RECT 3430.060 1578.770 3433.830 1584.160 ;
        RECT 3397.330 1570.900 3401.140 1576.320 ;
        RECT 221.000 1548.610 233.960 1554.630 ;
        RECT 307.120 1548.800 309.810 1554.400 ;
        RECT 204.970 1540.630 217.940 1546.610 ;
        RECT 302.300 1540.840 304.990 1546.440 ;
        RECT 89.350 1459.110 93.350 1522.550 ;
        RECT 154.100 1516.770 157.870 1522.160 ;
        RECT 95.350 1450.740 99.350 1515.660 ;
        RECT 186.790 1508.900 190.600 1514.320 ;
        RECT 3489.830 1512.740 3493.830 1577.660 ;
        RECT 3495.830 1521.110 3499.830 1584.550 ;
        RECT 3548.650 1526.380 3552.650 1593.210 ;
        RECT 3554.650 1517.730 3558.650 1601.350 ;
        RECT 3294.410 1388.870 3383.140 1392.030 ;
        RECT 220.975 1382.420 234.010 1386.420 ;
        RECT 3294.280 1384.080 3367.250 1387.280 ;
        RECT 220.975 1379.290 282.160 1382.420 ;
        RECT 3354.090 1380.080 3367.250 1384.080 ;
        RECT 3370.080 1383.870 3383.140 1388.870 ;
        RECT 213.730 1374.530 282.240 1377.660 ;
        RECT 213.730 1346.390 218.050 1374.530 ;
        RECT 3376.730 1369.870 3382.760 1375.940 ;
        RECT 3358.250 1361.870 3364.280 1367.940 ;
        RECT 3430.060 1353.770 3433.830 1359.160 ;
        RECT 3397.330 1345.900 3401.140 1351.320 ;
        RECT 89.350 1243.110 93.350 1306.550 ;
        RECT 154.100 1300.770 157.870 1306.160 ;
        RECT 95.350 1234.740 99.350 1299.660 ;
        RECT 186.790 1292.900 190.600 1298.320 ;
        RECT 3489.830 1287.740 3493.830 1352.660 ;
        RECT 3495.830 1296.110 3499.830 1359.550 ;
        RECT 3548.650 1301.380 3552.650 1368.210 ;
        RECT 3554.650 1292.730 3558.650 1376.350 ;
        RECT 3376.730 1143.870 3382.760 1149.940 ;
        RECT 3358.250 1135.870 3364.280 1141.940 ;
        RECT 3430.060 1127.770 3433.830 1133.160 ;
        RECT 3397.330 1119.900 3401.140 1125.320 ;
        RECT 89.350 1027.110 93.350 1090.550 ;
        RECT 154.100 1084.770 157.870 1090.160 ;
        RECT 95.350 1018.740 99.350 1083.660 ;
        RECT 186.790 1076.900 190.600 1082.320 ;
        RECT 3489.830 1061.740 3493.830 1126.660 ;
        RECT 3495.830 1070.110 3499.830 1133.550 ;
        RECT 3548.650 1075.380 3552.650 1142.210 ;
        RECT 3554.650 1066.730 3558.650 1150.350 ;
        RECT 3376.730 918.870 3382.760 924.940 ;
        RECT 3358.250 910.870 3364.280 916.940 ;
        RECT 3430.060 902.770 3433.830 908.160 ;
        RECT 3397.330 894.900 3401.140 900.320 ;
        RECT 3489.830 836.740 3493.830 901.660 ;
        RECT 3495.830 845.110 3499.830 908.550 ;
        RECT 3548.650 850.380 3552.650 917.210 ;
        RECT 3554.650 841.730 3558.650 925.350 ;
        RECT 3376.730 692.870 3382.760 698.940 ;
        RECT 3358.250 684.870 3364.280 690.940 ;
        RECT 3430.060 676.770 3433.830 682.160 ;
        RECT 3397.330 668.900 3401.140 674.320 ;
        RECT 3489.830 610.740 3493.830 675.660 ;
        RECT 3495.830 619.110 3499.830 682.550 ;
        RECT 3548.650 624.380 3552.650 691.210 ;
        RECT 3554.650 615.730 3558.650 699.350 ;
        RECT 2281.685 243.200 2299.120 245.200 ;
        RECT 717.200 208.000 718.100 236.480 ;
        RECT 643.050 206.310 647.340 208.000 ;
        RECT 716.450 206.310 718.230 208.000 ;
        RECT 723.700 204.610 724.600 236.700 ;
        RECT 745.670 209.380 746.570 210.455 ;
        RECT 650.710 202.910 655.000 204.610 ;
        RECT 722.950 202.910 724.725 204.610 ;
        RECT 738.970 200.290 740.895 209.380 ;
        RECT 2202.120 205.790 2203.970 210.390 ;
        RECT 2135.095 204.890 2203.970 205.790 ;
        RECT 2208.015 203.810 2210.045 203.885 ;
        RECT 2130.090 202.910 2210.045 203.810 ;
        RECT 2208.015 202.820 2210.045 202.910 ;
        RECT 2281.685 199.890 2283.590 243.200 ;
        RECT 2302.000 241.200 2303.600 245.200 ;
        RECT 2286.695 239.200 2303.600 241.200 ;
        RECT 2286.695 199.890 2288.600 239.200 ;
        RECT 3209.680 238.135 3251.010 240.135 ;
        RECT 3209.680 210.820 3218.590 238.135 ;
        RECT 3267.160 212.440 3284.560 235.270 ;
        RECT 739.085 186.710 740.800 190.915 ;
        RECT 2135.225 186.860 2136.865 190.765 ;
        RECT 2281.825 186.860 2283.465 190.765 ;
        RECT 650.860 175.830 654.880 179.980 ;
        RECT 643.210 169.790 647.230 173.940 ;
        RECT 3210.130 169.940 3218.170 173.800 ;
        RECT 2130.220 154.190 2131.860 158.095 ;
        RECT 2286.830 154.190 2288.470 158.095 ;
      LAYER via4 ;
        RECT 500.540 5097.460 501.720 5098.640 ;
        RECT 517.450 5097.470 518.630 5098.650 ;
        RECT 534.360 5097.440 535.540 5098.620 ;
        RECT 558.395 5097.460 559.575 5098.640 ;
        RECT 500.540 5095.860 501.720 5097.040 ;
        RECT 517.450 5095.870 518.630 5097.050 ;
        RECT 534.360 5095.840 535.540 5097.020 ;
        RECT 558.395 5095.860 559.575 5097.040 ;
        RECT 757.540 5097.460 758.720 5098.640 ;
        RECT 774.450 5097.470 775.630 5098.650 ;
        RECT 791.360 5097.440 792.540 5098.620 ;
        RECT 815.395 5097.460 816.575 5098.640 ;
        RECT 757.540 5095.860 758.720 5097.040 ;
        RECT 774.450 5095.870 775.630 5097.050 ;
        RECT 791.360 5095.840 792.540 5097.020 ;
        RECT 815.395 5095.860 816.575 5097.040 ;
        RECT 1014.540 5097.460 1015.720 5098.640 ;
        RECT 1031.450 5097.470 1032.630 5098.650 ;
        RECT 1048.360 5097.440 1049.540 5098.620 ;
        RECT 1072.395 5097.460 1073.575 5098.640 ;
        RECT 1014.540 5095.860 1015.720 5097.040 ;
        RECT 1031.450 5095.870 1032.630 5097.050 ;
        RECT 1048.360 5095.840 1049.540 5097.020 ;
        RECT 1072.395 5095.860 1073.575 5097.040 ;
        RECT 1271.540 5097.460 1272.720 5098.640 ;
        RECT 1288.450 5097.470 1289.630 5098.650 ;
        RECT 1305.360 5097.440 1306.540 5098.620 ;
        RECT 1329.395 5097.460 1330.575 5098.640 ;
        RECT 1271.540 5095.860 1272.720 5097.040 ;
        RECT 1288.450 5095.870 1289.630 5097.050 ;
        RECT 1305.360 5095.840 1306.540 5097.020 ;
        RECT 1329.395 5095.860 1330.575 5097.040 ;
        RECT 1529.540 5097.460 1530.720 5098.640 ;
        RECT 1546.450 5097.470 1547.630 5098.650 ;
        RECT 1563.360 5097.440 1564.540 5098.620 ;
        RECT 1587.395 5097.460 1588.575 5098.640 ;
        RECT 1529.540 5095.860 1530.720 5097.040 ;
        RECT 1546.450 5095.870 1547.630 5097.050 ;
        RECT 1563.360 5095.840 1564.540 5097.020 ;
        RECT 1587.395 5095.860 1588.575 5097.040 ;
        RECT 1781.540 5097.460 1782.720 5098.640 ;
        RECT 1798.450 5097.470 1799.630 5098.650 ;
        RECT 1815.360 5097.440 1816.540 5098.620 ;
        RECT 1839.395 5097.460 1840.575 5098.640 ;
        RECT 1781.540 5095.860 1782.720 5097.040 ;
        RECT 1798.450 5095.870 1799.630 5097.050 ;
        RECT 1815.360 5095.840 1816.540 5097.020 ;
        RECT 1839.395 5095.860 1840.575 5097.040 ;
        RECT 2118.540 5097.460 2119.720 5098.640 ;
        RECT 2135.450 5097.470 2136.630 5098.650 ;
        RECT 2152.360 5097.440 2153.540 5098.620 ;
        RECT 2176.395 5097.460 2177.575 5098.640 ;
        RECT 2118.540 5095.860 2119.720 5097.040 ;
        RECT 2135.450 5095.870 2136.630 5097.050 ;
        RECT 2152.360 5095.840 2153.540 5097.020 ;
        RECT 2176.395 5095.860 2177.575 5097.040 ;
        RECT 2503.540 5097.460 2504.720 5098.640 ;
        RECT 2520.450 5097.470 2521.630 5098.650 ;
        RECT 2537.360 5097.440 2538.540 5098.620 ;
        RECT 2561.395 5097.460 2562.575 5098.640 ;
        RECT 2503.540 5095.860 2504.720 5097.040 ;
        RECT 2520.450 5095.870 2521.630 5097.050 ;
        RECT 2537.360 5095.840 2538.540 5097.020 ;
        RECT 2561.395 5095.860 2562.575 5097.040 ;
        RECT 2760.540 5097.460 2761.720 5098.640 ;
        RECT 2777.450 5097.470 2778.630 5098.650 ;
        RECT 2794.360 5097.440 2795.540 5098.620 ;
        RECT 2818.395 5097.460 2819.575 5098.640 ;
        RECT 2760.540 5095.860 2761.720 5097.040 ;
        RECT 2777.450 5095.870 2778.630 5097.050 ;
        RECT 2794.360 5095.840 2795.540 5097.020 ;
        RECT 2818.395 5095.860 2819.575 5097.040 ;
        RECT 492.110 5091.440 493.290 5092.620 ;
        RECT 509.010 5091.440 510.190 5092.620 ;
        RECT 525.910 5091.460 527.090 5092.640 ;
        RECT 554.875 5091.460 556.055 5092.640 ;
        RECT 492.110 5089.840 493.290 5091.020 ;
        RECT 509.010 5089.840 510.190 5091.020 ;
        RECT 525.910 5089.860 527.090 5091.040 ;
        RECT 554.875 5089.860 556.055 5091.040 ;
        RECT 749.110 5091.440 750.290 5092.620 ;
        RECT 766.010 5091.440 767.190 5092.620 ;
        RECT 782.910 5091.460 784.090 5092.640 ;
        RECT 811.875 5091.460 813.055 5092.640 ;
        RECT 749.110 5089.840 750.290 5091.020 ;
        RECT 766.010 5089.840 767.190 5091.020 ;
        RECT 782.910 5089.860 784.090 5091.040 ;
        RECT 811.875 5089.860 813.055 5091.040 ;
        RECT 1006.110 5091.440 1007.290 5092.620 ;
        RECT 1023.010 5091.440 1024.190 5092.620 ;
        RECT 1039.910 5091.460 1041.090 5092.640 ;
        RECT 1068.875 5091.460 1070.055 5092.640 ;
        RECT 1006.110 5089.840 1007.290 5091.020 ;
        RECT 1023.010 5089.840 1024.190 5091.020 ;
        RECT 1039.910 5089.860 1041.090 5091.040 ;
        RECT 1068.875 5089.860 1070.055 5091.040 ;
        RECT 1263.110 5091.440 1264.290 5092.620 ;
        RECT 1280.010 5091.440 1281.190 5092.620 ;
        RECT 1296.910 5091.460 1298.090 5092.640 ;
        RECT 1325.875 5091.460 1327.055 5092.640 ;
        RECT 1263.110 5089.840 1264.290 5091.020 ;
        RECT 1280.010 5089.840 1281.190 5091.020 ;
        RECT 1296.910 5089.860 1298.090 5091.040 ;
        RECT 1325.875 5089.860 1327.055 5091.040 ;
        RECT 1521.110 5091.440 1522.290 5092.620 ;
        RECT 1538.010 5091.440 1539.190 5092.620 ;
        RECT 1554.910 5091.460 1556.090 5092.640 ;
        RECT 1583.875 5091.460 1585.055 5092.640 ;
        RECT 1521.110 5089.840 1522.290 5091.020 ;
        RECT 1538.010 5089.840 1539.190 5091.020 ;
        RECT 1554.910 5089.860 1556.090 5091.040 ;
        RECT 1583.875 5089.860 1585.055 5091.040 ;
        RECT 1773.110 5091.440 1774.290 5092.620 ;
        RECT 1790.010 5091.440 1791.190 5092.620 ;
        RECT 1806.910 5091.460 1808.090 5092.640 ;
        RECT 1835.875 5091.460 1837.055 5092.640 ;
        RECT 1773.110 5089.840 1774.290 5091.020 ;
        RECT 1790.010 5089.840 1791.190 5091.020 ;
        RECT 1806.910 5089.860 1808.090 5091.040 ;
        RECT 1835.875 5089.860 1837.055 5091.040 ;
        RECT 2110.110 5091.440 2111.290 5092.620 ;
        RECT 2127.010 5091.440 2128.190 5092.620 ;
        RECT 2143.910 5091.460 2145.090 5092.640 ;
        RECT 2172.875 5091.460 2174.055 5092.640 ;
        RECT 2110.110 5089.840 2111.290 5091.020 ;
        RECT 2127.010 5089.840 2128.190 5091.020 ;
        RECT 2143.910 5089.860 2145.090 5091.040 ;
        RECT 2172.875 5089.860 2174.055 5091.040 ;
        RECT 2495.110 5091.440 2496.290 5092.620 ;
        RECT 2512.010 5091.440 2513.190 5092.620 ;
        RECT 2528.910 5091.460 2530.090 5092.640 ;
        RECT 2557.875 5091.460 2559.055 5092.640 ;
        RECT 2495.110 5089.840 2496.290 5091.020 ;
        RECT 2512.010 5089.840 2513.190 5091.020 ;
        RECT 2528.910 5089.860 2530.090 5091.040 ;
        RECT 2557.875 5089.860 2559.055 5091.040 ;
        RECT 2752.110 5091.440 2753.290 5092.620 ;
        RECT 2769.010 5091.440 2770.190 5092.620 ;
        RECT 2785.910 5091.460 2787.090 5092.640 ;
        RECT 2814.875 5091.460 2816.055 5092.640 ;
        RECT 2752.110 5089.840 2753.290 5091.020 ;
        RECT 2769.010 5089.840 2770.190 5091.020 ;
        RECT 2785.910 5089.860 2787.090 5091.040 ;
        RECT 2814.875 5089.860 2816.055 5091.040 ;
        RECT 205.330 4929.425 217.710 4932.205 ;
        RECT 279.065 4930.215 280.245 4931.395 ;
        RECT 280.665 4930.215 281.845 4931.395 ;
        RECT 221.345 4924.650 233.725 4927.430 ;
        RECT 279.140 4924.595 281.920 4927.375 ;
        RECT 3291.955 4920.600 3293.135 4921.780 ;
        RECT 3293.555 4920.600 3294.735 4921.780 ;
        RECT 3295.155 4920.600 3296.335 4921.780 ;
        RECT 3296.755 4920.600 3297.935 4921.780 ;
        RECT 3298.355 4920.600 3299.535 4921.780 ;
        RECT 3299.955 4920.600 3301.135 4921.780 ;
        RECT 3301.555 4920.600 3302.735 4921.780 ;
        RECT 3303.155 4920.600 3304.335 4921.780 ;
        RECT 3304.755 4920.600 3305.935 4921.780 ;
        RECT 3306.355 4920.600 3307.535 4921.780 ;
        RECT 3307.955 4920.600 3309.135 4921.780 ;
        RECT 3309.555 4920.600 3310.735 4921.780 ;
        RECT 3311.155 4920.600 3312.335 4921.780 ;
        RECT 3312.755 4920.600 3313.935 4921.780 ;
        RECT 3314.355 4920.600 3315.535 4921.780 ;
        RECT 3354.415 4919.825 3366.795 4922.605 ;
        RECT 3291.865 4915.820 3293.045 4917.000 ;
        RECT 3293.465 4915.820 3294.645 4917.000 ;
        RECT 3295.065 4915.820 3296.245 4917.000 ;
        RECT 3296.665 4915.820 3297.845 4917.000 ;
        RECT 3298.265 4915.820 3299.445 4917.000 ;
        RECT 3299.865 4915.820 3301.045 4917.000 ;
        RECT 3301.465 4915.820 3302.645 4917.000 ;
        RECT 3303.065 4915.820 3304.245 4917.000 ;
        RECT 3304.665 4915.820 3305.845 4917.000 ;
        RECT 3306.265 4915.820 3307.445 4917.000 ;
        RECT 3307.865 4915.820 3309.045 4917.000 ;
        RECT 3309.465 4915.820 3310.645 4917.000 ;
        RECT 3311.065 4915.820 3312.245 4917.000 ;
        RECT 3312.665 4915.820 3313.845 4917.000 ;
        RECT 3314.265 4915.820 3315.445 4917.000 ;
        RECT 3370.405 4915.015 3382.785 4917.795 ;
        RECT 222.140 4760.325 232.920 4764.705 ;
        RECT 206.090 4752.415 216.870 4756.795 ;
        RECT 89.950 4728.395 91.130 4729.575 ;
        RECT 91.550 4728.395 92.730 4729.575 ;
        RECT 89.970 4704.360 91.150 4705.540 ;
        RECT 91.570 4704.360 92.750 4705.540 ;
        RECT 89.940 4687.450 91.120 4688.630 ;
        RECT 91.540 4687.450 92.720 4688.630 ;
        RECT 89.950 4670.540 91.130 4671.720 ;
        RECT 91.550 4670.540 92.730 4671.720 ;
        RECT 3377.505 4726.795 3381.885 4731.175 ;
        RECT 95.950 4724.875 97.130 4726.055 ;
        RECT 97.550 4724.875 98.730 4726.055 ;
        RECT 3358.975 4718.705 3363.355 4723.085 ;
        RECT 3496.400 4710.395 3497.580 4711.575 ;
        RECT 3498.000 4710.395 3499.180 4711.575 ;
        RECT 3490.400 4706.875 3491.580 4708.055 ;
        RECT 3492.000 4706.875 3493.180 4708.055 ;
        RECT 95.950 4695.910 97.130 4697.090 ;
        RECT 97.550 4695.910 98.730 4697.090 ;
        RECT 95.970 4679.010 97.150 4680.190 ;
        RECT 97.570 4679.010 98.750 4680.190 ;
        RECT 95.970 4662.110 97.150 4663.290 ;
        RECT 97.570 4662.110 98.750 4663.290 ;
        RECT 3490.400 4677.910 3491.580 4679.090 ;
        RECT 3492.000 4677.910 3493.180 4679.090 ;
        RECT 3490.380 4661.010 3491.560 4662.190 ;
        RECT 3491.980 4661.010 3493.160 4662.190 ;
        RECT 3496.380 4686.360 3497.560 4687.540 ;
        RECT 3497.980 4686.360 3499.160 4687.540 ;
        RECT 3496.410 4669.450 3497.590 4670.630 ;
        RECT 3498.010 4669.450 3499.190 4670.630 ;
        RECT 3549.205 4691.585 3550.385 4692.765 ;
        RECT 3550.805 4691.585 3551.985 4692.765 ;
        RECT 3549.215 4674.665 3550.395 4675.845 ;
        RECT 3550.815 4674.665 3551.995 4675.845 ;
        RECT 3549.225 4657.795 3550.405 4658.975 ;
        RECT 3550.825 4657.795 3552.005 4658.975 ;
        RECT 3555.215 4683.105 3556.395 4684.285 ;
        RECT 3556.815 4683.105 3557.995 4684.285 ;
        RECT 3555.185 4666.305 3556.365 4667.485 ;
        RECT 3556.785 4666.305 3557.965 4667.485 ;
        RECT 3496.400 4652.540 3497.580 4653.720 ;
        RECT 3498.000 4652.540 3499.180 4653.720 ;
        RECT 3555.195 4649.355 3556.375 4650.535 ;
        RECT 3556.795 4649.355 3557.975 4650.535 ;
        RECT 3490.380 4644.110 3491.560 4645.290 ;
        RECT 3491.980 4644.110 3493.160 4645.290 ;
        RECT 3373.995 4500.775 3378.375 4505.155 ;
        RECT 3358.215 4492.735 3362.595 4497.115 ;
        RECT 3371.050 4275.730 3375.430 4280.110 ;
        RECT 3358.330 4267.720 3362.710 4272.100 ;
        RECT 222.140 4131.325 232.920 4135.705 ;
        RECT 206.090 4123.415 216.870 4127.795 ;
        RECT 89.950 4099.395 91.130 4100.575 ;
        RECT 91.550 4099.395 92.730 4100.575 ;
        RECT 89.970 4075.360 91.150 4076.540 ;
        RECT 91.570 4075.360 92.750 4076.540 ;
        RECT 89.940 4058.450 91.120 4059.630 ;
        RECT 91.540 4058.450 92.720 4059.630 ;
        RECT 89.950 4041.540 91.130 4042.720 ;
        RECT 91.550 4041.540 92.730 4042.720 ;
        RECT 95.950 4095.875 97.130 4097.055 ;
        RECT 97.550 4095.875 98.730 4097.055 ;
        RECT 95.950 4066.910 97.130 4068.090 ;
        RECT 97.550 4066.910 98.730 4068.090 ;
        RECT 95.970 4050.010 97.150 4051.190 ;
        RECT 97.570 4050.010 98.750 4051.190 ;
        RECT 95.970 4033.110 97.150 4034.290 ;
        RECT 97.570 4033.110 98.750 4034.290 ;
        RECT 222.140 3923.325 232.920 3927.705 ;
        RECT 206.090 3915.415 216.870 3919.795 ;
        RECT 89.950 3883.395 91.130 3884.575 ;
        RECT 91.550 3883.395 92.730 3884.575 ;
        RECT 89.970 3859.360 91.150 3860.540 ;
        RECT 91.570 3859.360 92.750 3860.540 ;
        RECT 89.940 3842.450 91.120 3843.630 ;
        RECT 91.540 3842.450 92.720 3843.630 ;
        RECT 89.950 3825.540 91.130 3826.720 ;
        RECT 91.550 3825.540 92.730 3826.720 ;
        RECT 95.950 3879.875 97.130 3881.055 ;
        RECT 97.550 3879.875 98.730 3881.055 ;
        RECT 95.950 3850.910 97.130 3852.090 ;
        RECT 97.550 3850.910 98.730 3852.090 ;
        RECT 95.970 3834.010 97.150 3835.190 ;
        RECT 97.570 3834.010 98.750 3835.190 ;
        RECT 3377.555 3834.795 3381.935 3839.175 ;
        RECT 3359.025 3826.705 3363.405 3831.085 ;
        RECT 95.970 3817.110 97.150 3818.290 ;
        RECT 97.570 3817.110 98.750 3818.290 ;
        RECT 3496.450 3818.395 3497.630 3819.575 ;
        RECT 3498.050 3818.395 3499.230 3819.575 ;
        RECT 3490.450 3814.875 3491.630 3816.055 ;
        RECT 3492.050 3814.875 3493.230 3816.055 ;
        RECT 3490.450 3785.910 3491.630 3787.090 ;
        RECT 3492.050 3785.910 3493.230 3787.090 ;
        RECT 3490.430 3769.010 3491.610 3770.190 ;
        RECT 3492.030 3769.010 3493.210 3770.190 ;
        RECT 3496.430 3794.360 3497.610 3795.540 ;
        RECT 3498.030 3794.360 3499.210 3795.540 ;
        RECT 3496.460 3777.450 3497.640 3778.630 ;
        RECT 3498.060 3777.450 3499.240 3778.630 ;
        RECT 3549.255 3799.585 3550.435 3800.765 ;
        RECT 3550.855 3799.585 3552.035 3800.765 ;
        RECT 3549.265 3782.665 3550.445 3783.845 ;
        RECT 3550.865 3782.665 3552.045 3783.845 ;
        RECT 3549.275 3765.795 3550.455 3766.975 ;
        RECT 3550.875 3765.795 3552.055 3766.975 ;
        RECT 3555.265 3791.105 3556.445 3792.285 ;
        RECT 3556.865 3791.105 3558.045 3792.285 ;
        RECT 3555.235 3774.305 3556.415 3775.485 ;
        RECT 3556.835 3774.305 3558.015 3775.485 ;
        RECT 3496.450 3760.540 3497.630 3761.720 ;
        RECT 3498.050 3760.540 3499.230 3761.720 ;
        RECT 3555.245 3757.355 3556.425 3758.535 ;
        RECT 3556.845 3757.355 3558.025 3758.535 ;
        RECT 3490.430 3752.110 3491.610 3753.290 ;
        RECT 3492.030 3752.110 3493.210 3753.290 ;
        RECT 222.140 3699.325 232.920 3703.705 ;
        RECT 206.090 3691.415 216.870 3695.795 ;
        RECT 89.950 3667.395 91.130 3668.575 ;
        RECT 91.550 3667.395 92.730 3668.575 ;
        RECT 89.970 3643.360 91.150 3644.540 ;
        RECT 91.570 3643.360 92.750 3644.540 ;
        RECT 89.940 3626.450 91.120 3627.630 ;
        RECT 91.540 3626.450 92.720 3627.630 ;
        RECT 89.950 3609.540 91.130 3610.720 ;
        RECT 91.550 3609.540 92.730 3610.720 ;
        RECT 95.950 3663.875 97.130 3665.055 ;
        RECT 97.550 3663.875 98.730 3665.055 ;
        RECT 95.950 3634.910 97.130 3636.090 ;
        RECT 97.550 3634.910 98.730 3636.090 ;
        RECT 95.970 3618.010 97.150 3619.190 ;
        RECT 97.570 3618.010 98.750 3619.190 ;
        RECT 3377.555 3609.795 3381.935 3614.175 ;
        RECT 95.970 3601.110 97.150 3602.290 ;
        RECT 97.570 3601.110 98.750 3602.290 ;
        RECT 3359.025 3601.705 3363.405 3606.085 ;
        RECT 3496.450 3593.395 3497.630 3594.575 ;
        RECT 3498.050 3593.395 3499.230 3594.575 ;
        RECT 3490.450 3589.875 3491.630 3591.055 ;
        RECT 3492.050 3589.875 3493.230 3591.055 ;
        RECT 3490.450 3560.910 3491.630 3562.090 ;
        RECT 3492.050 3560.910 3493.230 3562.090 ;
        RECT 3490.430 3544.010 3491.610 3545.190 ;
        RECT 3492.030 3544.010 3493.210 3545.190 ;
        RECT 3496.430 3569.360 3497.610 3570.540 ;
        RECT 3498.030 3569.360 3499.210 3570.540 ;
        RECT 3496.460 3552.450 3497.640 3553.630 ;
        RECT 3498.060 3552.450 3499.240 3553.630 ;
        RECT 3549.255 3574.585 3550.435 3575.765 ;
        RECT 3550.855 3574.585 3552.035 3575.765 ;
        RECT 3549.265 3557.665 3550.445 3558.845 ;
        RECT 3550.865 3557.665 3552.045 3558.845 ;
        RECT 3549.275 3540.795 3550.455 3541.975 ;
        RECT 3550.875 3540.795 3552.055 3541.975 ;
        RECT 3555.265 3566.105 3556.445 3567.285 ;
        RECT 3556.865 3566.105 3558.045 3567.285 ;
        RECT 3555.235 3549.305 3556.415 3550.485 ;
        RECT 3556.835 3549.305 3558.015 3550.485 ;
        RECT 3496.450 3535.540 3497.630 3536.720 ;
        RECT 3498.050 3535.540 3499.230 3536.720 ;
        RECT 3555.245 3532.355 3556.425 3533.535 ;
        RECT 3556.845 3532.355 3558.025 3533.535 ;
        RECT 3490.430 3527.110 3491.610 3528.290 ;
        RECT 3492.030 3527.110 3493.210 3528.290 ;
        RECT 222.140 3483.325 232.920 3487.705 ;
        RECT 206.090 3475.415 216.870 3479.795 ;
        RECT 89.950 3451.395 91.130 3452.575 ;
        RECT 91.550 3451.395 92.730 3452.575 ;
        RECT 89.970 3427.360 91.150 3428.540 ;
        RECT 91.570 3427.360 92.750 3428.540 ;
        RECT 89.940 3410.450 91.120 3411.630 ;
        RECT 91.540 3410.450 92.720 3411.630 ;
        RECT 89.950 3393.540 91.130 3394.720 ;
        RECT 91.550 3393.540 92.730 3394.720 ;
        RECT 95.950 3447.875 97.130 3449.055 ;
        RECT 97.550 3447.875 98.730 3449.055 ;
        RECT 95.950 3418.910 97.130 3420.090 ;
        RECT 97.550 3418.910 98.730 3420.090 ;
        RECT 95.970 3402.010 97.150 3403.190 ;
        RECT 97.570 3402.010 98.750 3403.190 ;
        RECT 95.970 3385.110 97.150 3386.290 ;
        RECT 97.570 3385.110 98.750 3386.290 ;
        RECT 3377.555 3383.795 3381.935 3388.175 ;
        RECT 3359.025 3375.705 3363.405 3380.085 ;
        RECT 3496.450 3367.395 3497.630 3368.575 ;
        RECT 3498.050 3367.395 3499.230 3368.575 ;
        RECT 3490.450 3363.875 3491.630 3365.055 ;
        RECT 3492.050 3363.875 3493.230 3365.055 ;
        RECT 3490.450 3334.910 3491.630 3336.090 ;
        RECT 3492.050 3334.910 3493.230 3336.090 ;
        RECT 3490.430 3318.010 3491.610 3319.190 ;
        RECT 3492.030 3318.010 3493.210 3319.190 ;
        RECT 3496.430 3343.360 3497.610 3344.540 ;
        RECT 3498.030 3343.360 3499.210 3344.540 ;
        RECT 3496.460 3326.450 3497.640 3327.630 ;
        RECT 3498.060 3326.450 3499.240 3327.630 ;
        RECT 3549.255 3348.585 3550.435 3349.765 ;
        RECT 3550.855 3348.585 3552.035 3349.765 ;
        RECT 3549.265 3331.665 3550.445 3332.845 ;
        RECT 3550.865 3331.665 3552.045 3332.845 ;
        RECT 3549.275 3314.795 3550.455 3315.975 ;
        RECT 3550.875 3314.795 3552.055 3315.975 ;
        RECT 3555.265 3340.105 3556.445 3341.285 ;
        RECT 3556.865 3340.105 3558.045 3341.285 ;
        RECT 3555.235 3323.305 3556.415 3324.485 ;
        RECT 3556.835 3323.305 3558.015 3324.485 ;
        RECT 3496.450 3309.540 3497.630 3310.720 ;
        RECT 3498.050 3309.540 3499.230 3310.720 ;
        RECT 3555.245 3306.355 3556.425 3307.535 ;
        RECT 3556.845 3306.355 3558.025 3307.535 ;
        RECT 3490.430 3301.110 3491.610 3302.290 ;
        RECT 3492.030 3301.110 3493.210 3302.290 ;
        RECT 222.140 3267.325 232.920 3271.705 ;
        RECT 206.090 3259.415 216.870 3263.795 ;
        RECT 89.950 3235.395 91.130 3236.575 ;
        RECT 91.550 3235.395 92.730 3236.575 ;
        RECT 89.970 3211.360 91.150 3212.540 ;
        RECT 91.570 3211.360 92.750 3212.540 ;
        RECT 89.940 3194.450 91.120 3195.630 ;
        RECT 91.540 3194.450 92.720 3195.630 ;
        RECT 89.950 3177.540 91.130 3178.720 ;
        RECT 91.550 3177.540 92.730 3178.720 ;
        RECT 95.950 3231.875 97.130 3233.055 ;
        RECT 97.550 3231.875 98.730 3233.055 ;
        RECT 95.950 3202.910 97.130 3204.090 ;
        RECT 97.550 3202.910 98.730 3204.090 ;
        RECT 95.970 3186.010 97.150 3187.190 ;
        RECT 97.570 3186.010 98.750 3187.190 ;
        RECT 95.970 3169.110 97.150 3170.290 ;
        RECT 97.570 3169.110 98.750 3170.290 ;
        RECT 3377.555 3158.795 3381.935 3163.175 ;
        RECT 3359.025 3150.705 3363.405 3155.085 ;
        RECT 3496.450 3142.395 3497.630 3143.575 ;
        RECT 3498.050 3142.395 3499.230 3143.575 ;
        RECT 3490.450 3138.875 3491.630 3140.055 ;
        RECT 3492.050 3138.875 3493.230 3140.055 ;
        RECT 3490.450 3109.910 3491.630 3111.090 ;
        RECT 3492.050 3109.910 3493.230 3111.090 ;
        RECT 3490.430 3093.010 3491.610 3094.190 ;
        RECT 3492.030 3093.010 3493.210 3094.190 ;
        RECT 3496.430 3118.360 3497.610 3119.540 ;
        RECT 3498.030 3118.360 3499.210 3119.540 ;
        RECT 3496.460 3101.450 3497.640 3102.630 ;
        RECT 3498.060 3101.450 3499.240 3102.630 ;
        RECT 3549.255 3123.585 3550.435 3124.765 ;
        RECT 3550.855 3123.585 3552.035 3124.765 ;
        RECT 3549.265 3106.665 3550.445 3107.845 ;
        RECT 3550.865 3106.665 3552.045 3107.845 ;
        RECT 3549.275 3089.795 3550.455 3090.975 ;
        RECT 3550.875 3089.795 3552.055 3090.975 ;
        RECT 3555.265 3115.105 3556.445 3116.285 ;
        RECT 3556.865 3115.105 3558.045 3116.285 ;
        RECT 3555.235 3098.305 3556.415 3099.485 ;
        RECT 3556.835 3098.305 3558.015 3099.485 ;
        RECT 3496.450 3084.540 3497.630 3085.720 ;
        RECT 3498.050 3084.540 3499.230 3085.720 ;
        RECT 3555.245 3081.355 3556.425 3082.535 ;
        RECT 3556.845 3081.355 3558.025 3082.535 ;
        RECT 3490.430 3076.110 3491.610 3077.290 ;
        RECT 3492.030 3076.110 3493.210 3077.290 ;
        RECT 222.140 3056.625 232.920 3061.005 ;
        RECT 206.090 3048.715 216.870 3053.095 ;
        RECT 89.950 3019.395 91.130 3020.575 ;
        RECT 91.550 3019.395 92.730 3020.575 ;
        RECT 89.970 2995.360 91.150 2996.540 ;
        RECT 91.570 2995.360 92.750 2996.540 ;
        RECT 89.940 2978.450 91.120 2979.630 ;
        RECT 91.540 2978.450 92.720 2979.630 ;
        RECT 89.950 2961.540 91.130 2962.720 ;
        RECT 91.550 2961.540 92.730 2962.720 ;
        RECT 95.950 3015.875 97.130 3017.055 ;
        RECT 97.550 3015.875 98.730 3017.055 ;
        RECT 95.950 2986.910 97.130 2988.090 ;
        RECT 97.550 2986.910 98.730 2988.090 ;
        RECT 95.970 2970.010 97.150 2971.190 ;
        RECT 97.570 2970.010 98.750 2971.190 ;
        RECT 95.970 2953.110 97.150 2954.290 ;
        RECT 97.570 2953.110 98.750 2954.290 ;
        RECT 3377.555 2932.795 3381.935 2937.175 ;
        RECT 3359.025 2924.705 3363.405 2929.085 ;
        RECT 3496.450 2916.395 3497.630 2917.575 ;
        RECT 3498.050 2916.395 3499.230 2917.575 ;
        RECT 3490.450 2912.875 3491.630 2914.055 ;
        RECT 3492.050 2912.875 3493.230 2914.055 ;
        RECT 3490.450 2883.910 3491.630 2885.090 ;
        RECT 3492.050 2883.910 3493.230 2885.090 ;
        RECT 3490.430 2867.010 3491.610 2868.190 ;
        RECT 3492.030 2867.010 3493.210 2868.190 ;
        RECT 3496.430 2892.360 3497.610 2893.540 ;
        RECT 3498.030 2892.360 3499.210 2893.540 ;
        RECT 3496.460 2875.450 3497.640 2876.630 ;
        RECT 3498.060 2875.450 3499.240 2876.630 ;
        RECT 3549.255 2897.585 3550.435 2898.765 ;
        RECT 3550.855 2897.585 3552.035 2898.765 ;
        RECT 3549.265 2880.665 3550.445 2881.845 ;
        RECT 3550.865 2880.665 3552.045 2881.845 ;
        RECT 3549.275 2863.795 3550.455 2864.975 ;
        RECT 3550.875 2863.795 3552.055 2864.975 ;
        RECT 3555.265 2889.105 3556.445 2890.285 ;
        RECT 3556.865 2889.105 3558.045 2890.285 ;
        RECT 3555.235 2872.305 3556.415 2873.485 ;
        RECT 3556.835 2872.305 3558.015 2873.485 ;
        RECT 3496.450 2858.540 3497.630 2859.720 ;
        RECT 3498.050 2858.540 3499.230 2859.720 ;
        RECT 3555.245 2855.355 3556.425 2856.535 ;
        RECT 3556.845 2855.355 3558.025 2856.535 ;
        RECT 3490.430 2850.110 3491.610 2851.290 ;
        RECT 3492.030 2850.110 3493.210 2851.290 ;
        RECT 222.140 2835.325 232.920 2839.705 ;
        RECT 206.090 2827.415 216.870 2831.795 ;
        RECT 89.950 2803.395 91.130 2804.575 ;
        RECT 91.550 2803.395 92.730 2804.575 ;
        RECT 89.970 2779.360 91.150 2780.540 ;
        RECT 91.570 2779.360 92.750 2780.540 ;
        RECT 89.940 2762.450 91.120 2763.630 ;
        RECT 91.540 2762.450 92.720 2763.630 ;
        RECT 89.950 2745.540 91.130 2746.720 ;
        RECT 91.550 2745.540 92.730 2746.720 ;
        RECT 95.950 2799.875 97.130 2801.055 ;
        RECT 97.550 2799.875 98.730 2801.055 ;
        RECT 95.950 2770.910 97.130 2772.090 ;
        RECT 97.550 2770.910 98.730 2772.090 ;
        RECT 95.970 2754.010 97.150 2755.190 ;
        RECT 97.570 2754.010 98.750 2755.190 ;
        RECT 95.970 2737.110 97.150 2738.290 ;
        RECT 97.570 2737.110 98.750 2738.290 ;
        RECT 3377.555 2707.795 3381.935 2712.175 ;
        RECT 3359.025 2699.705 3363.405 2704.085 ;
        RECT 3496.450 2691.395 3497.630 2692.575 ;
        RECT 3498.050 2691.395 3499.230 2692.575 ;
        RECT 3490.450 2687.875 3491.630 2689.055 ;
        RECT 3492.050 2687.875 3493.230 2689.055 ;
        RECT 3490.450 2658.910 3491.630 2660.090 ;
        RECT 3492.050 2658.910 3493.230 2660.090 ;
        RECT 3490.430 2642.010 3491.610 2643.190 ;
        RECT 3492.030 2642.010 3493.210 2643.190 ;
        RECT 3496.430 2667.360 3497.610 2668.540 ;
        RECT 3498.030 2667.360 3499.210 2668.540 ;
        RECT 3496.460 2650.450 3497.640 2651.630 ;
        RECT 3498.060 2650.450 3499.240 2651.630 ;
        RECT 3549.255 2672.585 3550.435 2673.765 ;
        RECT 3550.855 2672.585 3552.035 2673.765 ;
        RECT 3549.265 2655.665 3550.445 2656.845 ;
        RECT 3550.865 2655.665 3552.045 2656.845 ;
        RECT 3549.275 2638.795 3550.455 2639.975 ;
        RECT 3550.875 2638.795 3552.055 2639.975 ;
        RECT 3555.265 2664.105 3556.445 2665.285 ;
        RECT 3556.865 2664.105 3558.045 2665.285 ;
        RECT 3555.235 2647.305 3556.415 2648.485 ;
        RECT 3556.835 2647.305 3558.015 2648.485 ;
        RECT 3496.450 2633.540 3497.630 2634.720 ;
        RECT 3498.050 2633.540 3499.230 2634.720 ;
        RECT 3555.245 2630.355 3556.425 2631.535 ;
        RECT 3556.845 2630.355 3558.025 2631.535 ;
        RECT 3490.430 2625.110 3491.610 2626.290 ;
        RECT 3492.030 2625.110 3493.210 2626.290 ;
        RECT 3377.555 2487.795 3381.935 2492.175 ;
        RECT 3359.025 2479.705 3363.405 2484.085 ;
        RECT 3496.450 2471.395 3497.630 2472.575 ;
        RECT 3498.050 2471.395 3499.230 2472.575 ;
        RECT 3490.450 2467.875 3491.630 2469.055 ;
        RECT 3492.050 2467.875 3493.230 2469.055 ;
        RECT 3490.450 2438.910 3491.630 2440.090 ;
        RECT 3492.050 2438.910 3493.230 2440.090 ;
        RECT 3490.430 2422.010 3491.610 2423.190 ;
        RECT 3492.030 2422.010 3493.210 2423.190 ;
        RECT 3496.430 2447.360 3497.610 2448.540 ;
        RECT 3498.030 2447.360 3499.210 2448.540 ;
        RECT 3496.460 2430.450 3497.640 2431.630 ;
        RECT 3498.060 2430.450 3499.240 2431.630 ;
        RECT 3549.255 2452.585 3550.435 2453.765 ;
        RECT 3550.855 2452.585 3552.035 2453.765 ;
        RECT 3549.265 2435.665 3550.445 2436.845 ;
        RECT 3550.865 2435.665 3552.045 2436.845 ;
        RECT 3549.275 2418.795 3550.455 2419.975 ;
        RECT 3550.875 2418.795 3552.055 2419.975 ;
        RECT 3555.265 2444.105 3556.445 2445.285 ;
        RECT 3556.865 2444.105 3558.045 2445.285 ;
        RECT 3555.235 2427.305 3556.415 2428.485 ;
        RECT 3556.835 2427.305 3558.015 2428.485 ;
        RECT 3496.450 2413.540 3497.630 2414.720 ;
        RECT 3498.050 2413.540 3499.230 2414.720 ;
        RECT 3555.245 2410.355 3556.425 2411.535 ;
        RECT 3556.845 2410.355 3558.025 2411.535 ;
        RECT 3490.430 2405.110 3491.610 2406.290 ;
        RECT 3492.030 2405.110 3493.210 2406.290 ;
        RECT 222.140 2197.325 232.920 2201.705 ;
        RECT 206.090 2189.415 216.870 2193.795 ;
        RECT 89.950 2165.395 91.130 2166.575 ;
        RECT 91.550 2165.395 92.730 2166.575 ;
        RECT 89.970 2141.360 91.150 2142.540 ;
        RECT 91.570 2141.360 92.750 2142.540 ;
        RECT 89.940 2124.450 91.120 2125.630 ;
        RECT 91.540 2124.450 92.720 2125.630 ;
        RECT 89.950 2107.540 91.130 2108.720 ;
        RECT 91.550 2107.540 92.730 2108.720 ;
        RECT 95.950 2161.875 97.130 2163.055 ;
        RECT 97.550 2161.875 98.730 2163.055 ;
        RECT 95.950 2132.910 97.130 2134.090 ;
        RECT 97.550 2132.910 98.730 2134.090 ;
        RECT 95.970 2116.010 97.150 2117.190 ;
        RECT 97.570 2116.010 98.750 2117.190 ;
        RECT 95.970 2099.110 97.150 2100.290 ;
        RECT 97.570 2099.110 98.750 2100.290 ;
        RECT 3377.555 2046.795 3381.935 2051.175 ;
        RECT 3359.025 2038.705 3363.405 2043.085 ;
        RECT 3496.450 2030.395 3497.630 2031.575 ;
        RECT 3498.050 2030.395 3499.230 2031.575 ;
        RECT 3490.450 2026.875 3491.630 2028.055 ;
        RECT 3492.050 2026.875 3493.230 2028.055 ;
        RECT 3490.450 1997.910 3491.630 1999.090 ;
        RECT 3492.050 1997.910 3493.230 1999.090 ;
        RECT 222.140 1981.325 232.920 1985.705 ;
        RECT 3490.430 1981.010 3491.610 1982.190 ;
        RECT 3492.030 1981.010 3493.210 1982.190 ;
        RECT 206.090 1973.415 216.870 1977.795 ;
        RECT 3496.430 2006.360 3497.610 2007.540 ;
        RECT 3498.030 2006.360 3499.210 2007.540 ;
        RECT 3496.460 1989.450 3497.640 1990.630 ;
        RECT 3498.060 1989.450 3499.240 1990.630 ;
        RECT 3549.255 2011.585 3550.435 2012.765 ;
        RECT 3550.855 2011.585 3552.035 2012.765 ;
        RECT 3549.265 1994.665 3550.445 1995.845 ;
        RECT 3550.865 1994.665 3552.045 1995.845 ;
        RECT 3549.275 1977.795 3550.455 1978.975 ;
        RECT 3550.875 1977.795 3552.055 1978.975 ;
        RECT 3555.265 2003.105 3556.445 2004.285 ;
        RECT 3556.865 2003.105 3558.045 2004.285 ;
        RECT 3555.235 1986.305 3556.415 1987.485 ;
        RECT 3556.835 1986.305 3558.015 1987.485 ;
        RECT 3496.450 1972.540 3497.630 1973.720 ;
        RECT 3498.050 1972.540 3499.230 1973.720 ;
        RECT 3555.245 1969.355 3556.425 1970.535 ;
        RECT 3556.845 1969.355 3558.025 1970.535 ;
        RECT 3490.430 1964.110 3491.610 1965.290 ;
        RECT 3492.030 1964.110 3493.210 1965.290 ;
        RECT 89.950 1949.395 91.130 1950.575 ;
        RECT 91.550 1949.395 92.730 1950.575 ;
        RECT 89.970 1925.360 91.150 1926.540 ;
        RECT 91.570 1925.360 92.750 1926.540 ;
        RECT 89.940 1908.450 91.120 1909.630 ;
        RECT 91.540 1908.450 92.720 1909.630 ;
        RECT 89.950 1891.540 91.130 1892.720 ;
        RECT 91.550 1891.540 92.730 1892.720 ;
        RECT 95.950 1945.875 97.130 1947.055 ;
        RECT 97.550 1945.875 98.730 1947.055 ;
        RECT 95.950 1916.910 97.130 1918.090 ;
        RECT 97.550 1916.910 98.730 1918.090 ;
        RECT 95.970 1900.010 97.150 1901.190 ;
        RECT 97.570 1900.010 98.750 1901.190 ;
        RECT 95.970 1883.110 97.150 1884.290 ;
        RECT 97.570 1883.110 98.750 1884.290 ;
        RECT 3377.555 1820.795 3381.935 1825.175 ;
        RECT 3359.025 1812.705 3363.405 1817.085 ;
        RECT 3496.450 1804.395 3497.630 1805.575 ;
        RECT 3498.050 1804.395 3499.230 1805.575 ;
        RECT 3490.450 1800.875 3491.630 1802.055 ;
        RECT 3492.050 1800.875 3493.230 1802.055 ;
        RECT 222.140 1770.325 232.920 1774.705 ;
        RECT 3490.450 1771.910 3491.630 1773.090 ;
        RECT 3492.050 1771.910 3493.230 1773.090 ;
        RECT 206.090 1762.415 216.870 1766.795 ;
        RECT 3490.430 1755.010 3491.610 1756.190 ;
        RECT 3492.030 1755.010 3493.210 1756.190 ;
        RECT 3496.430 1780.360 3497.610 1781.540 ;
        RECT 3498.030 1780.360 3499.210 1781.540 ;
        RECT 3496.460 1763.450 3497.640 1764.630 ;
        RECT 3498.060 1763.450 3499.240 1764.630 ;
        RECT 3549.255 1785.585 3550.435 1786.765 ;
        RECT 3550.855 1785.585 3552.035 1786.765 ;
        RECT 3549.265 1768.665 3550.445 1769.845 ;
        RECT 3550.865 1768.665 3552.045 1769.845 ;
        RECT 3549.275 1751.795 3550.455 1752.975 ;
        RECT 3550.875 1751.795 3552.055 1752.975 ;
        RECT 3555.265 1777.105 3556.445 1778.285 ;
        RECT 3556.865 1777.105 3558.045 1778.285 ;
        RECT 3555.235 1760.305 3556.415 1761.485 ;
        RECT 3556.835 1760.305 3558.015 1761.485 ;
        RECT 3496.450 1746.540 3497.630 1747.720 ;
        RECT 3498.050 1746.540 3499.230 1747.720 ;
        RECT 3555.245 1743.355 3556.425 1744.535 ;
        RECT 3556.845 1743.355 3558.025 1744.535 ;
        RECT 89.950 1733.395 91.130 1734.575 ;
        RECT 91.550 1733.395 92.730 1734.575 ;
        RECT 3490.430 1738.110 3491.610 1739.290 ;
        RECT 3492.030 1738.110 3493.210 1739.290 ;
        RECT 89.970 1709.360 91.150 1710.540 ;
        RECT 91.570 1709.360 92.750 1710.540 ;
        RECT 89.940 1692.450 91.120 1693.630 ;
        RECT 91.540 1692.450 92.720 1693.630 ;
        RECT 89.950 1675.540 91.130 1676.720 ;
        RECT 91.550 1675.540 92.730 1676.720 ;
        RECT 95.950 1729.875 97.130 1731.055 ;
        RECT 97.550 1729.875 98.730 1731.055 ;
        RECT 95.950 1700.910 97.130 1702.090 ;
        RECT 97.550 1700.910 98.730 1702.090 ;
        RECT 95.970 1684.010 97.150 1685.190 ;
        RECT 97.570 1684.010 98.750 1685.190 ;
        RECT 95.970 1667.110 97.150 1668.290 ;
        RECT 97.570 1667.110 98.750 1668.290 ;
        RECT 3377.555 1595.795 3381.935 1600.175 ;
        RECT 3359.025 1587.705 3363.405 1592.085 ;
        RECT 3496.450 1579.395 3497.630 1580.575 ;
        RECT 3498.050 1579.395 3499.230 1580.575 ;
        RECT 3490.450 1575.875 3491.630 1577.055 ;
        RECT 3492.050 1575.875 3493.230 1577.055 ;
        RECT 222.140 1549.325 232.920 1553.705 ;
        RECT 3490.450 1546.910 3491.630 1548.090 ;
        RECT 3492.050 1546.910 3493.230 1548.090 ;
        RECT 206.090 1541.415 216.870 1545.795 ;
        RECT 3490.430 1530.010 3491.610 1531.190 ;
        RECT 3492.030 1530.010 3493.210 1531.190 ;
        RECT 89.950 1517.395 91.130 1518.575 ;
        RECT 91.550 1517.395 92.730 1518.575 ;
        RECT 89.970 1493.360 91.150 1494.540 ;
        RECT 91.570 1493.360 92.750 1494.540 ;
        RECT 89.940 1476.450 91.120 1477.630 ;
        RECT 91.540 1476.450 92.720 1477.630 ;
        RECT 89.950 1459.540 91.130 1460.720 ;
        RECT 91.550 1459.540 92.730 1460.720 ;
        RECT 95.950 1513.875 97.130 1515.055 ;
        RECT 97.550 1513.875 98.730 1515.055 ;
        RECT 3496.430 1555.360 3497.610 1556.540 ;
        RECT 3498.030 1555.360 3499.210 1556.540 ;
        RECT 3496.460 1538.450 3497.640 1539.630 ;
        RECT 3498.060 1538.450 3499.240 1539.630 ;
        RECT 3549.255 1560.585 3550.435 1561.765 ;
        RECT 3550.855 1560.585 3552.035 1561.765 ;
        RECT 3549.265 1543.665 3550.445 1544.845 ;
        RECT 3550.865 1543.665 3552.045 1544.845 ;
        RECT 3549.275 1526.795 3550.455 1527.975 ;
        RECT 3550.875 1526.795 3552.055 1527.975 ;
        RECT 3555.265 1552.105 3556.445 1553.285 ;
        RECT 3556.865 1552.105 3558.045 1553.285 ;
        RECT 3555.235 1535.305 3556.415 1536.485 ;
        RECT 3556.835 1535.305 3558.015 1536.485 ;
        RECT 3496.450 1521.540 3497.630 1522.720 ;
        RECT 3498.050 1521.540 3499.230 1522.720 ;
        RECT 3555.245 1518.355 3556.425 1519.535 ;
        RECT 3556.845 1518.355 3558.025 1519.535 ;
        RECT 3490.430 1513.110 3491.610 1514.290 ;
        RECT 3492.030 1513.110 3493.210 1514.290 ;
        RECT 95.950 1484.910 97.130 1486.090 ;
        RECT 97.550 1484.910 98.730 1486.090 ;
        RECT 95.970 1468.010 97.150 1469.190 ;
        RECT 97.570 1468.010 98.750 1469.190 ;
        RECT 95.970 1451.110 97.150 1452.290 ;
        RECT 97.570 1451.110 98.750 1452.290 ;
        RECT 3294.920 1389.875 3296.100 1391.055 ;
        RECT 3296.520 1389.875 3297.700 1391.055 ;
        RECT 3298.120 1389.875 3299.300 1391.055 ;
        RECT 3299.720 1389.875 3300.900 1391.055 ;
        RECT 3301.320 1389.875 3302.500 1391.055 ;
        RECT 3302.920 1389.875 3304.100 1391.055 ;
        RECT 3304.520 1389.875 3305.700 1391.055 ;
        RECT 3306.120 1389.875 3307.300 1391.055 ;
        RECT 3307.720 1389.875 3308.900 1391.055 ;
        RECT 3309.320 1389.875 3310.500 1391.055 ;
        RECT 3310.920 1389.875 3312.100 1391.055 ;
        RECT 3312.520 1389.875 3313.700 1391.055 ;
        RECT 3314.120 1389.875 3315.300 1391.055 ;
        RECT 221.285 1379.885 233.665 1385.865 ;
        RECT 3294.825 1385.150 3296.005 1386.330 ;
        RECT 3296.425 1385.150 3297.605 1386.330 ;
        RECT 3298.025 1385.150 3299.205 1386.330 ;
        RECT 3299.625 1385.150 3300.805 1386.330 ;
        RECT 3301.225 1385.150 3302.405 1386.330 ;
        RECT 3302.825 1385.150 3304.005 1386.330 ;
        RECT 3304.425 1385.150 3305.605 1386.330 ;
        RECT 3306.025 1385.150 3307.205 1386.330 ;
        RECT 3307.625 1385.150 3308.805 1386.330 ;
        RECT 3309.225 1385.150 3310.405 1386.330 ;
        RECT 3310.825 1385.150 3312.005 1386.330 ;
        RECT 3312.425 1385.150 3313.605 1386.330 ;
        RECT 3314.025 1385.150 3315.205 1386.330 ;
        RECT 279.080 1380.260 280.260 1381.440 ;
        RECT 280.680 1380.260 281.860 1381.440 ;
        RECT 3354.430 1380.720 3366.810 1386.700 ;
        RECT 3370.430 1384.150 3382.810 1391.730 ;
        RECT 214.505 1347.100 217.285 1377.080 ;
        RECT 279.120 1375.490 280.300 1376.670 ;
        RECT 280.720 1375.490 281.900 1376.670 ;
        RECT 3377.555 1370.795 3381.935 1375.175 ;
        RECT 3359.025 1362.705 3363.405 1367.085 ;
        RECT 3496.450 1354.395 3497.630 1355.575 ;
        RECT 3498.050 1354.395 3499.230 1355.575 ;
        RECT 3490.450 1350.875 3491.630 1352.055 ;
        RECT 3492.050 1350.875 3493.230 1352.055 ;
        RECT 3490.450 1321.910 3491.630 1323.090 ;
        RECT 3492.050 1321.910 3493.230 1323.090 ;
        RECT 89.950 1301.395 91.130 1302.575 ;
        RECT 91.550 1301.395 92.730 1302.575 ;
        RECT 3490.430 1305.010 3491.610 1306.190 ;
        RECT 3492.030 1305.010 3493.210 1306.190 ;
        RECT 89.970 1277.360 91.150 1278.540 ;
        RECT 91.570 1277.360 92.750 1278.540 ;
        RECT 89.940 1260.450 91.120 1261.630 ;
        RECT 91.540 1260.450 92.720 1261.630 ;
        RECT 89.950 1243.540 91.130 1244.720 ;
        RECT 91.550 1243.540 92.730 1244.720 ;
        RECT 95.950 1297.875 97.130 1299.055 ;
        RECT 97.550 1297.875 98.730 1299.055 ;
        RECT 3496.430 1330.360 3497.610 1331.540 ;
        RECT 3498.030 1330.360 3499.210 1331.540 ;
        RECT 3496.460 1313.450 3497.640 1314.630 ;
        RECT 3498.060 1313.450 3499.240 1314.630 ;
        RECT 3549.255 1335.585 3550.435 1336.765 ;
        RECT 3550.855 1335.585 3552.035 1336.765 ;
        RECT 3549.265 1318.665 3550.445 1319.845 ;
        RECT 3550.865 1318.665 3552.045 1319.845 ;
        RECT 3549.275 1301.795 3550.455 1302.975 ;
        RECT 3550.875 1301.795 3552.055 1302.975 ;
        RECT 3555.265 1327.105 3556.445 1328.285 ;
        RECT 3556.865 1327.105 3558.045 1328.285 ;
        RECT 3555.235 1310.305 3556.415 1311.485 ;
        RECT 3556.835 1310.305 3558.015 1311.485 ;
        RECT 3496.450 1296.540 3497.630 1297.720 ;
        RECT 3498.050 1296.540 3499.230 1297.720 ;
        RECT 3555.245 1293.355 3556.425 1294.535 ;
        RECT 3556.845 1293.355 3558.025 1294.535 ;
        RECT 3490.430 1288.110 3491.610 1289.290 ;
        RECT 3492.030 1288.110 3493.210 1289.290 ;
        RECT 95.950 1268.910 97.130 1270.090 ;
        RECT 97.550 1268.910 98.730 1270.090 ;
        RECT 95.970 1252.010 97.150 1253.190 ;
        RECT 97.570 1252.010 98.750 1253.190 ;
        RECT 95.970 1235.110 97.150 1236.290 ;
        RECT 97.570 1235.110 98.750 1236.290 ;
        RECT 3377.555 1144.795 3381.935 1149.175 ;
        RECT 3359.025 1136.705 3363.405 1141.085 ;
        RECT 3496.450 1128.395 3497.630 1129.575 ;
        RECT 3498.050 1128.395 3499.230 1129.575 ;
        RECT 3490.450 1124.875 3491.630 1126.055 ;
        RECT 3492.050 1124.875 3493.230 1126.055 ;
        RECT 3490.450 1095.910 3491.630 1097.090 ;
        RECT 3492.050 1095.910 3493.230 1097.090 ;
        RECT 89.950 1085.395 91.130 1086.575 ;
        RECT 91.550 1085.395 92.730 1086.575 ;
        RECT 89.970 1061.360 91.150 1062.540 ;
        RECT 91.570 1061.360 92.750 1062.540 ;
        RECT 89.940 1044.450 91.120 1045.630 ;
        RECT 91.540 1044.450 92.720 1045.630 ;
        RECT 89.950 1027.540 91.130 1028.720 ;
        RECT 91.550 1027.540 92.730 1028.720 ;
        RECT 95.950 1081.875 97.130 1083.055 ;
        RECT 97.550 1081.875 98.730 1083.055 ;
        RECT 3490.430 1079.010 3491.610 1080.190 ;
        RECT 3492.030 1079.010 3493.210 1080.190 ;
        RECT 3496.430 1104.360 3497.610 1105.540 ;
        RECT 3498.030 1104.360 3499.210 1105.540 ;
        RECT 3496.460 1087.450 3497.640 1088.630 ;
        RECT 3498.060 1087.450 3499.240 1088.630 ;
        RECT 3549.255 1109.585 3550.435 1110.765 ;
        RECT 3550.855 1109.585 3552.035 1110.765 ;
        RECT 3549.265 1092.665 3550.445 1093.845 ;
        RECT 3550.865 1092.665 3552.045 1093.845 ;
        RECT 3549.275 1075.795 3550.455 1076.975 ;
        RECT 3550.875 1075.795 3552.055 1076.975 ;
        RECT 3555.265 1101.105 3556.445 1102.285 ;
        RECT 3556.865 1101.105 3558.045 1102.285 ;
        RECT 3555.235 1084.305 3556.415 1085.485 ;
        RECT 3556.835 1084.305 3558.015 1085.485 ;
        RECT 3496.450 1070.540 3497.630 1071.720 ;
        RECT 3498.050 1070.540 3499.230 1071.720 ;
        RECT 3555.245 1067.355 3556.425 1068.535 ;
        RECT 3556.845 1067.355 3558.025 1068.535 ;
        RECT 3490.430 1062.110 3491.610 1063.290 ;
        RECT 3492.030 1062.110 3493.210 1063.290 ;
        RECT 95.950 1052.910 97.130 1054.090 ;
        RECT 97.550 1052.910 98.730 1054.090 ;
        RECT 95.970 1036.010 97.150 1037.190 ;
        RECT 97.570 1036.010 98.750 1037.190 ;
        RECT 95.970 1019.110 97.150 1020.290 ;
        RECT 97.570 1019.110 98.750 1020.290 ;
        RECT 3377.555 919.795 3381.935 924.175 ;
        RECT 3359.025 911.705 3363.405 916.085 ;
        RECT 3496.450 903.395 3497.630 904.575 ;
        RECT 3498.050 903.395 3499.230 904.575 ;
        RECT 3490.450 899.875 3491.630 901.055 ;
        RECT 3492.050 899.875 3493.230 901.055 ;
        RECT 3490.450 870.910 3491.630 872.090 ;
        RECT 3492.050 870.910 3493.230 872.090 ;
        RECT 3490.430 854.010 3491.610 855.190 ;
        RECT 3492.030 854.010 3493.210 855.190 ;
        RECT 3496.430 879.360 3497.610 880.540 ;
        RECT 3498.030 879.360 3499.210 880.540 ;
        RECT 3496.460 862.450 3497.640 863.630 ;
        RECT 3498.060 862.450 3499.240 863.630 ;
        RECT 3549.255 884.585 3550.435 885.765 ;
        RECT 3550.855 884.585 3552.035 885.765 ;
        RECT 3549.265 867.665 3550.445 868.845 ;
        RECT 3550.865 867.665 3552.045 868.845 ;
        RECT 3549.275 850.795 3550.455 851.975 ;
        RECT 3550.875 850.795 3552.055 851.975 ;
        RECT 3555.265 876.105 3556.445 877.285 ;
        RECT 3556.865 876.105 3558.045 877.285 ;
        RECT 3555.235 859.305 3556.415 860.485 ;
        RECT 3556.835 859.305 3558.015 860.485 ;
        RECT 3496.450 845.540 3497.630 846.720 ;
        RECT 3498.050 845.540 3499.230 846.720 ;
        RECT 3555.245 842.355 3556.425 843.535 ;
        RECT 3556.845 842.355 3558.025 843.535 ;
        RECT 3490.430 837.110 3491.610 838.290 ;
        RECT 3492.030 837.110 3493.210 838.290 ;
        RECT 3377.555 693.795 3381.935 698.175 ;
        RECT 3359.025 685.705 3363.405 690.085 ;
        RECT 3496.450 677.395 3497.630 678.575 ;
        RECT 3498.050 677.395 3499.230 678.575 ;
        RECT 3490.450 673.875 3491.630 675.055 ;
        RECT 3492.050 673.875 3493.230 675.055 ;
        RECT 3490.450 644.910 3491.630 646.090 ;
        RECT 3492.050 644.910 3493.230 646.090 ;
        RECT 3490.430 628.010 3491.610 629.190 ;
        RECT 3492.030 628.010 3493.210 629.190 ;
        RECT 3496.430 653.360 3497.610 654.540 ;
        RECT 3498.030 653.360 3499.210 654.540 ;
        RECT 3496.460 636.450 3497.640 637.630 ;
        RECT 3498.060 636.450 3499.240 637.630 ;
        RECT 3549.255 658.585 3550.435 659.765 ;
        RECT 3550.855 658.585 3552.035 659.765 ;
        RECT 3549.265 641.665 3550.445 642.845 ;
        RECT 3550.865 641.665 3552.045 642.845 ;
        RECT 3549.275 624.795 3550.455 625.975 ;
        RECT 3550.875 624.795 3552.055 625.975 ;
        RECT 3555.265 650.105 3556.445 651.285 ;
        RECT 3556.865 650.105 3558.045 651.285 ;
        RECT 3555.235 633.305 3556.415 634.485 ;
        RECT 3556.835 633.305 3558.015 634.485 ;
        RECT 3496.450 619.540 3497.630 620.720 ;
        RECT 3498.050 619.540 3499.230 620.720 ;
        RECT 3555.245 616.355 3556.425 617.535 ;
        RECT 3556.845 616.355 3558.025 617.535 ;
        RECT 3490.430 611.110 3491.610 612.290 ;
        RECT 3492.030 611.110 3493.210 612.290 ;
        RECT 643.800 206.700 644.980 207.880 ;
        RECT 645.405 206.700 646.585 207.880 ;
        RECT 716.920 206.700 718.100 207.880 ;
        RECT 651.460 203.310 652.640 204.490 ;
        RECT 653.065 203.310 654.245 204.490 ;
        RECT 723.420 203.310 724.600 204.490 ;
      LAYER met5 ;
        RECT 491.900 5093.460 493.500 5101.470 ;
        RECT 500.350 5099.450 501.950 5101.470 ;
        RECT 500.280 5095.070 502.010 5099.450 ;
        RECT 508.800 5093.470 510.400 5101.470 ;
        RECT 517.250 5099.530 518.850 5101.470 ;
        RECT 517.140 5095.150 518.900 5099.530 ;
        RECT 525.700 5093.480 527.300 5101.470 ;
        RECT 534.150 5099.390 535.750 5101.470 ;
        RECT 534.110 5095.010 535.840 5099.390 ;
        RECT 491.840 5089.080 493.570 5093.460 ;
        RECT 508.740 5089.090 510.470 5093.470 ;
        RECT 525.620 5089.100 527.350 5093.480 ;
        RECT 554.650 5093.350 556.250 5117.040 ;
        RECT 558.150 5099.610 559.750 5117.040 ;
        RECT 558.130 5095.230 559.860 5099.610 ;
        RECT 748.900 5093.460 750.500 5101.470 ;
        RECT 757.350 5099.450 758.950 5101.470 ;
        RECT 757.280 5095.070 759.010 5099.450 ;
        RECT 765.800 5093.470 767.400 5101.470 ;
        RECT 774.250 5099.530 775.850 5101.470 ;
        RECT 774.140 5095.150 775.900 5099.530 ;
        RECT 782.700 5093.480 784.300 5101.470 ;
        RECT 791.150 5099.390 792.750 5101.470 ;
        RECT 791.110 5095.010 792.840 5099.390 ;
        RECT 525.700 5089.090 527.300 5089.100 ;
        RECT 554.620 5088.970 556.350 5093.350 ;
        RECT 748.840 5089.080 750.570 5093.460 ;
        RECT 765.740 5089.090 767.470 5093.470 ;
        RECT 782.620 5089.100 784.350 5093.480 ;
        RECT 811.650 5093.350 813.250 5117.040 ;
        RECT 815.150 5099.610 816.750 5117.040 ;
        RECT 815.130 5095.230 816.860 5099.610 ;
        RECT 1005.900 5093.460 1007.500 5101.470 ;
        RECT 1014.350 5099.450 1015.950 5101.470 ;
        RECT 1014.280 5095.070 1016.010 5099.450 ;
        RECT 1022.800 5093.470 1024.400 5101.470 ;
        RECT 1031.250 5099.530 1032.850 5101.470 ;
        RECT 1031.140 5095.150 1032.900 5099.530 ;
        RECT 1039.700 5093.480 1041.300 5101.470 ;
        RECT 1048.150 5099.390 1049.750 5101.470 ;
        RECT 1048.110 5095.010 1049.840 5099.390 ;
        RECT 782.700 5089.090 784.300 5089.100 ;
        RECT 811.620 5088.970 813.350 5093.350 ;
        RECT 1005.840 5089.080 1007.570 5093.460 ;
        RECT 1022.740 5089.090 1024.470 5093.470 ;
        RECT 1039.620 5089.100 1041.350 5093.480 ;
        RECT 1068.650 5093.350 1070.250 5117.040 ;
        RECT 1072.150 5099.610 1073.750 5117.040 ;
        RECT 1072.130 5095.230 1073.860 5099.610 ;
        RECT 1262.900 5093.460 1264.500 5101.470 ;
        RECT 1271.350 5099.450 1272.950 5101.470 ;
        RECT 1271.280 5095.070 1273.010 5099.450 ;
        RECT 1279.800 5093.470 1281.400 5101.470 ;
        RECT 1288.250 5099.530 1289.850 5101.470 ;
        RECT 1288.140 5095.150 1289.900 5099.530 ;
        RECT 1296.700 5093.480 1298.300 5101.470 ;
        RECT 1305.150 5099.390 1306.750 5101.470 ;
        RECT 1305.110 5095.010 1306.840 5099.390 ;
        RECT 1039.700 5089.090 1041.300 5089.100 ;
        RECT 1068.620 5088.970 1070.350 5093.350 ;
        RECT 1262.840 5089.080 1264.570 5093.460 ;
        RECT 1279.740 5089.090 1281.470 5093.470 ;
        RECT 1296.620 5089.100 1298.350 5093.480 ;
        RECT 1325.650 5093.350 1327.250 5117.040 ;
        RECT 1329.150 5099.610 1330.750 5117.040 ;
        RECT 1329.130 5095.230 1330.860 5099.610 ;
        RECT 1520.900 5093.460 1522.500 5101.470 ;
        RECT 1529.350 5099.450 1530.950 5101.470 ;
        RECT 1529.280 5095.070 1531.010 5099.450 ;
        RECT 1537.800 5093.470 1539.400 5101.470 ;
        RECT 1546.250 5099.530 1547.850 5101.470 ;
        RECT 1546.140 5095.150 1547.900 5099.530 ;
        RECT 1554.700 5093.480 1556.300 5101.470 ;
        RECT 1563.150 5099.390 1564.750 5101.470 ;
        RECT 1563.110 5095.010 1564.840 5099.390 ;
        RECT 1296.700 5089.090 1298.300 5089.100 ;
        RECT 1325.620 5088.970 1327.350 5093.350 ;
        RECT 1520.840 5089.080 1522.570 5093.460 ;
        RECT 1537.740 5089.090 1539.470 5093.470 ;
        RECT 1554.620 5089.100 1556.350 5093.480 ;
        RECT 1583.650 5093.350 1585.250 5117.040 ;
        RECT 1587.150 5099.610 1588.750 5117.040 ;
        RECT 1587.130 5095.230 1588.860 5099.610 ;
        RECT 1772.900 5093.460 1774.500 5101.470 ;
        RECT 1781.350 5099.450 1782.950 5101.470 ;
        RECT 1781.280 5095.070 1783.010 5099.450 ;
        RECT 1789.800 5093.470 1791.400 5101.470 ;
        RECT 1798.250 5099.530 1799.850 5101.470 ;
        RECT 1798.140 5095.150 1799.900 5099.530 ;
        RECT 1806.700 5093.480 1808.300 5101.470 ;
        RECT 1815.150 5099.390 1816.750 5101.470 ;
        RECT 1815.110 5095.010 1816.840 5099.390 ;
        RECT 1554.700 5089.090 1556.300 5089.100 ;
        RECT 1583.620 5088.970 1585.350 5093.350 ;
        RECT 1772.840 5089.080 1774.570 5093.460 ;
        RECT 1789.740 5089.090 1791.470 5093.470 ;
        RECT 1806.620 5089.100 1808.350 5093.480 ;
        RECT 1835.650 5093.350 1837.250 5117.040 ;
        RECT 1839.150 5099.610 1840.750 5117.040 ;
        RECT 1839.130 5095.230 1840.860 5099.610 ;
        RECT 2109.900 5093.460 2111.500 5101.470 ;
        RECT 2118.350 5099.450 2119.950 5101.470 ;
        RECT 2118.280 5095.070 2120.010 5099.450 ;
        RECT 2126.800 5093.470 2128.400 5101.470 ;
        RECT 2135.250 5099.530 2136.850 5101.470 ;
        RECT 2135.140 5095.150 2136.900 5099.530 ;
        RECT 2143.700 5093.480 2145.300 5101.470 ;
        RECT 2152.150 5099.390 2153.750 5101.470 ;
        RECT 2152.110 5095.010 2153.840 5099.390 ;
        RECT 1806.700 5089.090 1808.300 5089.100 ;
        RECT 1835.620 5088.970 1837.350 5093.350 ;
        RECT 2109.840 5089.080 2111.570 5093.460 ;
        RECT 2126.740 5089.090 2128.470 5093.470 ;
        RECT 2143.620 5089.100 2145.350 5093.480 ;
        RECT 2172.650 5093.350 2174.250 5117.040 ;
        RECT 2176.150 5099.610 2177.750 5117.040 ;
        RECT 2176.130 5095.230 2177.860 5099.610 ;
        RECT 2494.900 5093.460 2496.500 5101.470 ;
        RECT 2503.350 5099.450 2504.950 5101.470 ;
        RECT 2503.280 5095.070 2505.010 5099.450 ;
        RECT 2511.800 5093.470 2513.400 5101.470 ;
        RECT 2520.250 5099.530 2521.850 5101.470 ;
        RECT 2520.140 5095.150 2521.900 5099.530 ;
        RECT 2528.700 5093.480 2530.300 5101.470 ;
        RECT 2537.150 5099.390 2538.750 5101.470 ;
        RECT 2537.110 5095.010 2538.840 5099.390 ;
        RECT 2143.700 5089.090 2145.300 5089.100 ;
        RECT 2172.620 5088.970 2174.350 5093.350 ;
        RECT 2494.840 5089.080 2496.570 5093.460 ;
        RECT 2511.740 5089.090 2513.470 5093.470 ;
        RECT 2528.620 5089.100 2530.350 5093.480 ;
        RECT 2557.650 5093.350 2559.250 5117.040 ;
        RECT 2561.150 5099.610 2562.750 5117.040 ;
        RECT 2561.130 5095.230 2562.860 5099.610 ;
        RECT 2751.900 5093.460 2753.500 5101.470 ;
        RECT 2760.350 5099.450 2761.950 5101.470 ;
        RECT 2760.280 5095.070 2762.010 5099.450 ;
        RECT 2768.800 5093.470 2770.400 5101.470 ;
        RECT 2777.250 5099.530 2778.850 5101.470 ;
        RECT 2777.140 5095.150 2778.900 5099.530 ;
        RECT 2785.700 5093.480 2787.300 5101.470 ;
        RECT 2794.150 5099.390 2795.750 5101.470 ;
        RECT 2794.110 5095.010 2795.840 5099.390 ;
        RECT 2528.700 5089.090 2530.300 5089.100 ;
        RECT 2557.620 5088.970 2559.350 5093.350 ;
        RECT 2751.840 5089.080 2753.570 5093.460 ;
        RECT 2768.740 5089.090 2770.470 5093.470 ;
        RECT 2785.620 5089.100 2787.350 5093.480 ;
        RECT 2814.650 5093.350 2816.250 5117.040 ;
        RECT 2818.150 5099.610 2819.750 5117.040 ;
        RECT 2818.130 5095.230 2819.860 5099.610 ;
        RECT 2785.700 5089.090 2787.300 5089.100 ;
        RECT 2814.620 5088.970 2816.350 5093.350 ;
        RECT 205.170 4929.390 217.870 4932.240 ;
        RECT 278.880 4929.240 302.180 4932.340 ;
        RECT 221.210 4924.590 233.860 4927.490 ;
        RECT 278.880 4924.440 306.990 4927.540 ;
        RECT 3260.900 4919.640 3315.890 4922.740 ;
        RECT 3354.290 4919.750 3366.920 4922.680 ;
        RECT 3256.140 4914.840 3315.890 4917.940 ;
        RECT 3370.280 4914.940 3382.910 4917.870 ;
        RECT 221.390 4759.880 233.670 4765.150 ;
        RECT 205.340 4751.970 217.620 4757.240 ;
        RECT 89.230 4729.780 93.425 4729.895 ;
        RECT 71.550 4728.180 93.425 4729.780 ;
        RECT 89.230 4728.090 93.425 4728.180 ;
        RECT 95.260 4726.280 99.455 4726.350 ;
        RECT 71.550 4724.680 99.610 4726.280 ;
        RECT 3376.990 4726.240 3382.400 4731.730 ;
        RECT 95.260 4724.545 99.455 4724.680 ;
        RECT 3358.460 4718.150 3363.870 4723.640 ;
        RECT 3495.740 4711.780 3499.870 4711.840 ;
        RECT 3495.740 4710.180 3517.580 4711.780 ;
        RECT 3495.740 4710.125 3499.870 4710.180 ;
        RECT 3489.685 4708.280 3493.815 4708.355 ;
        RECT 3489.520 4706.680 3517.580 4708.280 ;
        RECT 3489.685 4706.640 3493.815 4706.680 ;
        RECT 89.245 4705.750 93.455 4705.840 ;
        RECT 87.120 4704.150 93.540 4705.750 ;
        RECT 89.245 4704.040 93.455 4704.150 ;
        RECT 95.280 4697.300 99.490 4697.365 ;
        RECT 87.120 4695.700 99.500 4697.300 ;
        RECT 95.280 4695.620 99.490 4695.700 ;
        RECT 3548.530 4692.990 3552.715 4693.075 ;
        RECT 3546.220 4691.390 3552.830 4692.990 ;
        RECT 3548.530 4691.300 3552.715 4691.390 ;
        RECT 89.285 4688.850 93.495 4688.890 ;
        RECT 87.120 4687.250 93.495 4688.850 ;
        RECT 89.285 4687.145 93.495 4687.250 ;
        RECT 3495.580 4687.750 3499.905 4687.850 ;
        RECT 3495.580 4686.150 3502.010 4687.750 ;
        RECT 3495.580 4686.080 3499.905 4686.150 ;
        RECT 3554.535 4684.540 3558.720 4684.620 ;
        RECT 3546.220 4682.940 3558.890 4684.540 ;
        RECT 3554.535 4682.845 3558.720 4682.940 ;
        RECT 95.265 4680.400 99.475 4680.475 ;
        RECT 87.120 4678.800 99.500 4680.400 ;
        RECT 3489.595 4679.300 3493.920 4679.360 ;
        RECT 95.265 4678.730 99.475 4678.800 ;
        RECT 3489.595 4677.700 3502.010 4679.300 ;
        RECT 3489.595 4677.590 3493.920 4677.700 ;
        RECT 3548.505 4676.090 3552.690 4676.205 ;
        RECT 3546.220 4674.490 3552.800 4676.090 ;
        RECT 3548.505 4674.430 3552.690 4674.490 ;
        RECT 89.265 4671.950 93.475 4672.025 ;
        RECT 87.120 4670.350 93.510 4671.950 ;
        RECT 3495.695 4670.850 3500.020 4670.935 ;
        RECT 89.265 4670.280 93.475 4670.350 ;
        RECT 3495.695 4669.250 3502.010 4670.850 ;
        RECT 3495.695 4669.165 3500.020 4669.250 ;
        RECT 3554.480 4667.640 3558.890 4667.750 ;
        RECT 3546.220 4666.140 3558.890 4667.640 ;
        RECT 3546.220 4666.060 3558.885 4666.140 ;
        RECT 3546.220 4666.040 3558.880 4666.060 ;
        RECT 95.310 4663.500 99.520 4663.575 ;
        RECT 87.120 4661.900 99.520 4663.500 ;
        RECT 95.310 4661.830 99.520 4661.900 ;
        RECT 3489.600 4662.400 3493.925 4662.460 ;
        RECT 3489.600 4660.800 3502.010 4662.400 ;
        RECT 3489.600 4660.690 3493.925 4660.800 ;
        RECT 3548.510 4659.190 3552.690 4659.280 ;
        RECT 3546.060 4657.590 3552.690 4659.190 ;
        RECT 3548.510 4657.480 3552.690 4657.590 ;
        RECT 3495.600 4653.950 3499.925 4654.055 ;
        RECT 3495.600 4652.350 3502.010 4653.950 ;
        RECT 3495.600 4652.285 3499.925 4652.350 ;
        RECT 3554.475 4650.740 3558.660 4650.820 ;
        RECT 3546.060 4649.140 3558.660 4650.740 ;
        RECT 3554.475 4649.045 3558.660 4649.140 ;
        RECT 3489.630 4645.500 3493.955 4645.600 ;
        RECT 3489.630 4643.900 3502.010 4645.500 ;
        RECT 3489.630 4643.830 3493.955 4643.900 ;
        RECT 3373.670 4500.370 3378.700 4505.560 ;
        RECT 3357.830 4492.330 3362.980 4497.520 ;
        RECT 3370.580 4275.260 3375.900 4280.580 ;
        RECT 3357.850 4267.210 3363.190 4272.610 ;
        RECT 221.390 4130.880 233.670 4136.150 ;
        RECT 205.340 4122.970 217.620 4128.240 ;
        RECT 89.230 4100.780 93.425 4100.895 ;
        RECT 71.550 4099.180 93.425 4100.780 ;
        RECT 89.230 4099.090 93.425 4099.180 ;
        RECT 95.260 4097.280 99.455 4097.350 ;
        RECT 71.550 4095.680 99.610 4097.280 ;
        RECT 95.260 4095.545 99.455 4095.680 ;
        RECT 89.245 4076.750 93.455 4076.840 ;
        RECT 87.120 4075.150 93.540 4076.750 ;
        RECT 89.245 4075.040 93.455 4075.150 ;
        RECT 95.280 4068.300 99.490 4068.365 ;
        RECT 87.120 4066.700 99.500 4068.300 ;
        RECT 95.280 4066.620 99.490 4066.700 ;
        RECT 89.285 4059.850 93.495 4059.890 ;
        RECT 87.120 4058.250 93.495 4059.850 ;
        RECT 89.285 4058.145 93.495 4058.250 ;
        RECT 95.265 4051.400 99.475 4051.475 ;
        RECT 87.120 4049.800 99.500 4051.400 ;
        RECT 95.265 4049.730 99.475 4049.800 ;
        RECT 89.265 4042.950 93.475 4043.025 ;
        RECT 87.120 4041.350 93.510 4042.950 ;
        RECT 89.265 4041.280 93.475 4041.350 ;
        RECT 95.310 4034.500 99.520 4034.575 ;
        RECT 87.120 4032.900 99.520 4034.500 ;
        RECT 95.310 4032.830 99.520 4032.900 ;
        RECT 221.390 3922.880 233.670 3928.150 ;
        RECT 205.340 3914.970 217.620 3920.240 ;
        RECT 89.230 3884.780 93.425 3884.895 ;
        RECT 71.550 3883.180 93.425 3884.780 ;
        RECT 89.230 3883.090 93.425 3883.180 ;
        RECT 95.260 3881.280 99.455 3881.350 ;
        RECT 71.550 3879.680 99.610 3881.280 ;
        RECT 95.260 3879.545 99.455 3879.680 ;
        RECT 89.245 3860.750 93.455 3860.840 ;
        RECT 87.120 3859.150 93.540 3860.750 ;
        RECT 89.245 3859.040 93.455 3859.150 ;
        RECT 95.280 3852.300 99.490 3852.365 ;
        RECT 87.120 3850.700 99.500 3852.300 ;
        RECT 95.280 3850.620 99.490 3850.700 ;
        RECT 89.285 3843.850 93.495 3843.890 ;
        RECT 87.120 3842.250 93.495 3843.850 ;
        RECT 89.285 3842.145 93.495 3842.250 ;
        RECT 95.265 3835.400 99.475 3835.475 ;
        RECT 87.120 3833.800 99.500 3835.400 ;
        RECT 3377.040 3834.240 3382.450 3839.730 ;
        RECT 95.265 3833.730 99.475 3833.800 ;
        RECT 89.265 3826.950 93.475 3827.025 ;
        RECT 87.120 3825.350 93.510 3826.950 ;
        RECT 3358.510 3826.150 3363.920 3831.640 ;
        RECT 89.265 3825.280 93.475 3825.350 ;
        RECT 3495.790 3819.780 3499.920 3819.840 ;
        RECT 95.310 3818.500 99.520 3818.575 ;
        RECT 87.120 3816.900 99.520 3818.500 ;
        RECT 3495.790 3818.180 3517.630 3819.780 ;
        RECT 3495.790 3818.125 3499.920 3818.180 ;
        RECT 95.310 3816.830 99.520 3816.900 ;
        RECT 3489.735 3816.280 3493.865 3816.355 ;
        RECT 3489.570 3814.680 3517.630 3816.280 ;
        RECT 3489.735 3814.640 3493.865 3814.680 ;
        RECT 3548.580 3800.990 3552.765 3801.075 ;
        RECT 3546.270 3799.390 3552.880 3800.990 ;
        RECT 3548.580 3799.300 3552.765 3799.390 ;
        RECT 3495.630 3795.750 3499.955 3795.850 ;
        RECT 3495.630 3794.150 3502.060 3795.750 ;
        RECT 3495.630 3794.080 3499.955 3794.150 ;
        RECT 3554.585 3792.540 3558.770 3792.620 ;
        RECT 3546.270 3790.940 3558.940 3792.540 ;
        RECT 3554.585 3790.845 3558.770 3790.940 ;
        RECT 3489.645 3787.300 3493.970 3787.360 ;
        RECT 3489.645 3785.700 3502.060 3787.300 ;
        RECT 3489.645 3785.590 3493.970 3785.700 ;
        RECT 3548.555 3784.090 3552.740 3784.205 ;
        RECT 3546.270 3782.490 3552.850 3784.090 ;
        RECT 3548.555 3782.430 3552.740 3782.490 ;
        RECT 3495.745 3778.850 3500.070 3778.935 ;
        RECT 3495.745 3777.250 3502.060 3778.850 ;
        RECT 3495.745 3777.165 3500.070 3777.250 ;
        RECT 3554.530 3775.640 3558.940 3775.750 ;
        RECT 3546.270 3774.140 3558.940 3775.640 ;
        RECT 3546.270 3774.060 3558.935 3774.140 ;
        RECT 3546.270 3774.040 3558.930 3774.060 ;
        RECT 3489.650 3770.400 3493.975 3770.460 ;
        RECT 3489.650 3768.800 3502.060 3770.400 ;
        RECT 3489.650 3768.690 3493.975 3768.800 ;
        RECT 3548.560 3767.190 3552.740 3767.280 ;
        RECT 3546.110 3765.590 3552.740 3767.190 ;
        RECT 3548.560 3765.480 3552.740 3765.590 ;
        RECT 3495.650 3761.950 3499.975 3762.055 ;
        RECT 3495.650 3760.350 3502.060 3761.950 ;
        RECT 3495.650 3760.285 3499.975 3760.350 ;
        RECT 3554.525 3758.740 3558.710 3758.820 ;
        RECT 3546.110 3757.140 3558.710 3758.740 ;
        RECT 3554.525 3757.045 3558.710 3757.140 ;
        RECT 3489.680 3753.500 3494.005 3753.600 ;
        RECT 3489.680 3751.900 3502.060 3753.500 ;
        RECT 3489.680 3751.830 3494.005 3751.900 ;
        RECT 221.390 3698.880 233.670 3704.150 ;
        RECT 205.340 3690.970 217.620 3696.240 ;
        RECT 89.230 3668.780 93.425 3668.895 ;
        RECT 71.550 3667.180 93.425 3668.780 ;
        RECT 89.230 3667.090 93.425 3667.180 ;
        RECT 95.260 3665.280 99.455 3665.350 ;
        RECT 71.550 3663.680 99.610 3665.280 ;
        RECT 95.260 3663.545 99.455 3663.680 ;
        RECT 89.245 3644.750 93.455 3644.840 ;
        RECT 87.120 3643.150 93.540 3644.750 ;
        RECT 89.245 3643.040 93.455 3643.150 ;
        RECT 95.280 3636.300 99.490 3636.365 ;
        RECT 87.120 3634.700 99.500 3636.300 ;
        RECT 95.280 3634.620 99.490 3634.700 ;
        RECT 89.285 3627.850 93.495 3627.890 ;
        RECT 87.120 3626.250 93.495 3627.850 ;
        RECT 89.285 3626.145 93.495 3626.250 ;
        RECT 95.265 3619.400 99.475 3619.475 ;
        RECT 87.120 3617.800 99.500 3619.400 ;
        RECT 95.265 3617.730 99.475 3617.800 ;
        RECT 89.265 3610.950 93.475 3611.025 ;
        RECT 87.120 3609.350 93.510 3610.950 ;
        RECT 89.265 3609.280 93.475 3609.350 ;
        RECT 3377.040 3609.240 3382.450 3614.730 ;
        RECT 95.310 3602.500 99.520 3602.575 ;
        RECT 87.120 3600.900 99.520 3602.500 ;
        RECT 3358.510 3601.150 3363.920 3606.640 ;
        RECT 95.310 3600.830 99.520 3600.900 ;
        RECT 3495.790 3594.780 3499.920 3594.840 ;
        RECT 3495.790 3593.180 3517.630 3594.780 ;
        RECT 3495.790 3593.125 3499.920 3593.180 ;
        RECT 3489.735 3591.280 3493.865 3591.355 ;
        RECT 3489.570 3589.680 3517.630 3591.280 ;
        RECT 3489.735 3589.640 3493.865 3589.680 ;
        RECT 3548.580 3575.990 3552.765 3576.075 ;
        RECT 3546.270 3574.390 3552.880 3575.990 ;
        RECT 3548.580 3574.300 3552.765 3574.390 ;
        RECT 3495.630 3570.750 3499.955 3570.850 ;
        RECT 3495.630 3569.150 3502.060 3570.750 ;
        RECT 3495.630 3569.080 3499.955 3569.150 ;
        RECT 3554.585 3567.540 3558.770 3567.620 ;
        RECT 3546.270 3565.940 3558.940 3567.540 ;
        RECT 3554.585 3565.845 3558.770 3565.940 ;
        RECT 3489.645 3562.300 3493.970 3562.360 ;
        RECT 3489.645 3560.700 3502.060 3562.300 ;
        RECT 3489.645 3560.590 3493.970 3560.700 ;
        RECT 3548.555 3559.090 3552.740 3559.205 ;
        RECT 3546.270 3557.490 3552.850 3559.090 ;
        RECT 3548.555 3557.430 3552.740 3557.490 ;
        RECT 3495.745 3553.850 3500.070 3553.935 ;
        RECT 3495.745 3552.250 3502.060 3553.850 ;
        RECT 3495.745 3552.165 3500.070 3552.250 ;
        RECT 3554.530 3550.640 3558.940 3550.750 ;
        RECT 3546.270 3549.140 3558.940 3550.640 ;
        RECT 3546.270 3549.060 3558.935 3549.140 ;
        RECT 3546.270 3549.040 3558.930 3549.060 ;
        RECT 3489.650 3545.400 3493.975 3545.460 ;
        RECT 3489.650 3543.800 3502.060 3545.400 ;
        RECT 3489.650 3543.690 3493.975 3543.800 ;
        RECT 3548.560 3542.190 3552.740 3542.280 ;
        RECT 3546.110 3540.590 3552.740 3542.190 ;
        RECT 3548.560 3540.480 3552.740 3540.590 ;
        RECT 3495.650 3536.950 3499.975 3537.055 ;
        RECT 3495.650 3535.350 3502.060 3536.950 ;
        RECT 3495.650 3535.285 3499.975 3535.350 ;
        RECT 3554.525 3533.740 3558.710 3533.820 ;
        RECT 3546.110 3532.140 3558.710 3533.740 ;
        RECT 3554.525 3532.045 3558.710 3532.140 ;
        RECT 3489.680 3528.500 3494.005 3528.600 ;
        RECT 3489.680 3526.900 3502.060 3528.500 ;
        RECT 3489.680 3526.830 3494.005 3526.900 ;
        RECT 221.390 3482.880 233.670 3488.150 ;
        RECT 205.340 3474.970 217.620 3480.240 ;
        RECT 89.230 3452.780 93.425 3452.895 ;
        RECT 71.550 3451.180 93.425 3452.780 ;
        RECT 89.230 3451.090 93.425 3451.180 ;
        RECT 95.260 3449.280 99.455 3449.350 ;
        RECT 71.550 3447.680 99.610 3449.280 ;
        RECT 95.260 3447.545 99.455 3447.680 ;
        RECT 89.245 3428.750 93.455 3428.840 ;
        RECT 87.120 3427.150 93.540 3428.750 ;
        RECT 89.245 3427.040 93.455 3427.150 ;
        RECT 95.280 3420.300 99.490 3420.365 ;
        RECT 87.120 3418.700 99.500 3420.300 ;
        RECT 95.280 3418.620 99.490 3418.700 ;
        RECT 89.285 3411.850 93.495 3411.890 ;
        RECT 87.120 3410.250 93.495 3411.850 ;
        RECT 89.285 3410.145 93.495 3410.250 ;
        RECT 95.265 3403.400 99.475 3403.475 ;
        RECT 87.120 3401.800 99.500 3403.400 ;
        RECT 95.265 3401.730 99.475 3401.800 ;
        RECT 89.265 3394.950 93.475 3395.025 ;
        RECT 87.120 3393.350 93.510 3394.950 ;
        RECT 89.265 3393.280 93.475 3393.350 ;
        RECT 95.310 3386.500 99.520 3386.575 ;
        RECT 87.120 3384.900 99.520 3386.500 ;
        RECT 95.310 3384.830 99.520 3384.900 ;
        RECT 3377.040 3383.240 3382.450 3388.730 ;
        RECT 3358.510 3375.150 3363.920 3380.640 ;
        RECT 3495.790 3368.780 3499.920 3368.840 ;
        RECT 3495.790 3367.180 3517.630 3368.780 ;
        RECT 3495.790 3367.125 3499.920 3367.180 ;
        RECT 3489.735 3365.280 3493.865 3365.355 ;
        RECT 3489.570 3363.680 3517.630 3365.280 ;
        RECT 3489.735 3363.640 3493.865 3363.680 ;
        RECT 3548.580 3349.990 3552.765 3350.075 ;
        RECT 3546.270 3348.390 3552.880 3349.990 ;
        RECT 3548.580 3348.300 3552.765 3348.390 ;
        RECT 3495.630 3344.750 3499.955 3344.850 ;
        RECT 3495.630 3343.150 3502.060 3344.750 ;
        RECT 3495.630 3343.080 3499.955 3343.150 ;
        RECT 3554.585 3341.540 3558.770 3341.620 ;
        RECT 3546.270 3339.940 3558.940 3341.540 ;
        RECT 3554.585 3339.845 3558.770 3339.940 ;
        RECT 3489.645 3336.300 3493.970 3336.360 ;
        RECT 3489.645 3334.700 3502.060 3336.300 ;
        RECT 3489.645 3334.590 3493.970 3334.700 ;
        RECT 3548.555 3333.090 3552.740 3333.205 ;
        RECT 3546.270 3331.490 3552.850 3333.090 ;
        RECT 3548.555 3331.430 3552.740 3331.490 ;
        RECT 3495.745 3327.850 3500.070 3327.935 ;
        RECT 3495.745 3326.250 3502.060 3327.850 ;
        RECT 3495.745 3326.165 3500.070 3326.250 ;
        RECT 3554.530 3324.640 3558.940 3324.750 ;
        RECT 3546.270 3323.140 3558.940 3324.640 ;
        RECT 3546.270 3323.060 3558.935 3323.140 ;
        RECT 3546.270 3323.040 3558.930 3323.060 ;
        RECT 3489.650 3319.400 3493.975 3319.460 ;
        RECT 3489.650 3317.800 3502.060 3319.400 ;
        RECT 3489.650 3317.690 3493.975 3317.800 ;
        RECT 3548.560 3316.190 3552.740 3316.280 ;
        RECT 3546.110 3314.590 3552.740 3316.190 ;
        RECT 3548.560 3314.480 3552.740 3314.590 ;
        RECT 3495.650 3310.950 3499.975 3311.055 ;
        RECT 3495.650 3309.350 3502.060 3310.950 ;
        RECT 3495.650 3309.285 3499.975 3309.350 ;
        RECT 3554.525 3307.740 3558.710 3307.820 ;
        RECT 3546.110 3306.140 3558.710 3307.740 ;
        RECT 3554.525 3306.045 3558.710 3306.140 ;
        RECT 3489.680 3302.500 3494.005 3302.600 ;
        RECT 3489.680 3300.900 3502.060 3302.500 ;
        RECT 3489.680 3300.830 3494.005 3300.900 ;
        RECT 221.390 3266.880 233.670 3272.150 ;
        RECT 205.340 3258.970 217.620 3264.240 ;
        RECT 89.230 3236.780 93.425 3236.895 ;
        RECT 71.550 3235.180 93.425 3236.780 ;
        RECT 89.230 3235.090 93.425 3235.180 ;
        RECT 95.260 3233.280 99.455 3233.350 ;
        RECT 71.550 3231.680 99.610 3233.280 ;
        RECT 95.260 3231.545 99.455 3231.680 ;
        RECT 89.245 3212.750 93.455 3212.840 ;
        RECT 87.120 3211.150 93.540 3212.750 ;
        RECT 89.245 3211.040 93.455 3211.150 ;
        RECT 95.280 3204.300 99.490 3204.365 ;
        RECT 87.120 3202.700 99.500 3204.300 ;
        RECT 95.280 3202.620 99.490 3202.700 ;
        RECT 89.285 3195.850 93.495 3195.890 ;
        RECT 87.120 3194.250 93.495 3195.850 ;
        RECT 89.285 3194.145 93.495 3194.250 ;
        RECT 95.265 3187.400 99.475 3187.475 ;
        RECT 87.120 3185.800 99.500 3187.400 ;
        RECT 95.265 3185.730 99.475 3185.800 ;
        RECT 89.265 3178.950 93.475 3179.025 ;
        RECT 87.120 3177.350 93.510 3178.950 ;
        RECT 89.265 3177.280 93.475 3177.350 ;
        RECT 95.310 3170.500 99.520 3170.575 ;
        RECT 87.120 3168.900 99.520 3170.500 ;
        RECT 95.310 3168.830 99.520 3168.900 ;
        RECT 3377.040 3158.240 3382.450 3163.730 ;
        RECT 3358.510 3150.150 3363.920 3155.640 ;
        RECT 3495.790 3143.780 3499.920 3143.840 ;
        RECT 3495.790 3142.180 3517.630 3143.780 ;
        RECT 3495.790 3142.125 3499.920 3142.180 ;
        RECT 3489.735 3140.280 3493.865 3140.355 ;
        RECT 3489.570 3138.680 3517.630 3140.280 ;
        RECT 3489.735 3138.640 3493.865 3138.680 ;
        RECT 3548.580 3124.990 3552.765 3125.075 ;
        RECT 3546.270 3123.390 3552.880 3124.990 ;
        RECT 3548.580 3123.300 3552.765 3123.390 ;
        RECT 3495.630 3119.750 3499.955 3119.850 ;
        RECT 3495.630 3118.150 3502.060 3119.750 ;
        RECT 3495.630 3118.080 3499.955 3118.150 ;
        RECT 3554.585 3116.540 3558.770 3116.620 ;
        RECT 3546.270 3114.940 3558.940 3116.540 ;
        RECT 3554.585 3114.845 3558.770 3114.940 ;
        RECT 3489.645 3111.300 3493.970 3111.360 ;
        RECT 3489.645 3109.700 3502.060 3111.300 ;
        RECT 3489.645 3109.590 3493.970 3109.700 ;
        RECT 3548.555 3108.090 3552.740 3108.205 ;
        RECT 3546.270 3106.490 3552.850 3108.090 ;
        RECT 3548.555 3106.430 3552.740 3106.490 ;
        RECT 3495.745 3102.850 3500.070 3102.935 ;
        RECT 3495.745 3101.250 3502.060 3102.850 ;
        RECT 3495.745 3101.165 3500.070 3101.250 ;
        RECT 3554.530 3099.640 3558.940 3099.750 ;
        RECT 3546.270 3098.140 3558.940 3099.640 ;
        RECT 3546.270 3098.060 3558.935 3098.140 ;
        RECT 3546.270 3098.040 3558.930 3098.060 ;
        RECT 3489.650 3094.400 3493.975 3094.460 ;
        RECT 3489.650 3092.800 3502.060 3094.400 ;
        RECT 3489.650 3092.690 3493.975 3092.800 ;
        RECT 3548.560 3091.190 3552.740 3091.280 ;
        RECT 3546.110 3089.590 3552.740 3091.190 ;
        RECT 3548.560 3089.480 3552.740 3089.590 ;
        RECT 3495.650 3085.950 3499.975 3086.055 ;
        RECT 3495.650 3084.350 3502.060 3085.950 ;
        RECT 3495.650 3084.285 3499.975 3084.350 ;
        RECT 3554.525 3082.740 3558.710 3082.820 ;
        RECT 3546.110 3081.140 3558.710 3082.740 ;
        RECT 3554.525 3081.045 3558.710 3081.140 ;
        RECT 3489.680 3077.500 3494.005 3077.600 ;
        RECT 3489.680 3075.900 3502.060 3077.500 ;
        RECT 3489.680 3075.830 3494.005 3075.900 ;
        RECT 221.390 3056.180 233.670 3061.450 ;
        RECT 205.340 3048.270 217.620 3053.540 ;
        RECT 89.230 3020.780 93.425 3020.895 ;
        RECT 71.550 3019.180 93.425 3020.780 ;
        RECT 89.230 3019.090 93.425 3019.180 ;
        RECT 95.260 3017.280 99.455 3017.350 ;
        RECT 71.550 3015.680 99.610 3017.280 ;
        RECT 95.260 3015.545 99.455 3015.680 ;
        RECT 89.245 2996.750 93.455 2996.840 ;
        RECT 87.120 2995.150 93.540 2996.750 ;
        RECT 89.245 2995.040 93.455 2995.150 ;
        RECT 95.280 2988.300 99.490 2988.365 ;
        RECT 87.120 2986.700 99.500 2988.300 ;
        RECT 95.280 2986.620 99.490 2986.700 ;
        RECT 89.285 2979.850 93.495 2979.890 ;
        RECT 87.120 2978.250 93.495 2979.850 ;
        RECT 89.285 2978.145 93.495 2978.250 ;
        RECT 95.265 2971.400 99.475 2971.475 ;
        RECT 87.120 2969.800 99.500 2971.400 ;
        RECT 95.265 2969.730 99.475 2969.800 ;
        RECT 89.265 2962.950 93.475 2963.025 ;
        RECT 87.120 2961.350 93.510 2962.950 ;
        RECT 89.265 2961.280 93.475 2961.350 ;
        RECT 95.310 2954.500 99.520 2954.575 ;
        RECT 87.120 2952.900 99.520 2954.500 ;
        RECT 95.310 2952.830 99.520 2952.900 ;
        RECT 3377.040 2932.240 3382.450 2937.730 ;
        RECT 3358.510 2924.150 3363.920 2929.640 ;
        RECT 3495.790 2917.780 3499.920 2917.840 ;
        RECT 3495.790 2916.180 3517.630 2917.780 ;
        RECT 3495.790 2916.125 3499.920 2916.180 ;
        RECT 3489.735 2914.280 3493.865 2914.355 ;
        RECT 3489.570 2912.680 3517.630 2914.280 ;
        RECT 3489.735 2912.640 3493.865 2912.680 ;
        RECT 3548.580 2898.990 3552.765 2899.075 ;
        RECT 3546.270 2897.390 3552.880 2898.990 ;
        RECT 3548.580 2897.300 3552.765 2897.390 ;
        RECT 3495.630 2893.750 3499.955 2893.850 ;
        RECT 3495.630 2892.150 3502.060 2893.750 ;
        RECT 3495.630 2892.080 3499.955 2892.150 ;
        RECT 3554.585 2890.540 3558.770 2890.620 ;
        RECT 3546.270 2888.940 3558.940 2890.540 ;
        RECT 3554.585 2888.845 3558.770 2888.940 ;
        RECT 3489.645 2885.300 3493.970 2885.360 ;
        RECT 3489.645 2883.700 3502.060 2885.300 ;
        RECT 3489.645 2883.590 3493.970 2883.700 ;
        RECT 3548.555 2882.090 3552.740 2882.205 ;
        RECT 3546.270 2880.490 3552.850 2882.090 ;
        RECT 3548.555 2880.430 3552.740 2880.490 ;
        RECT 3495.745 2876.850 3500.070 2876.935 ;
        RECT 3495.745 2875.250 3502.060 2876.850 ;
        RECT 3495.745 2875.165 3500.070 2875.250 ;
        RECT 3554.530 2873.640 3558.940 2873.750 ;
        RECT 3546.270 2872.140 3558.940 2873.640 ;
        RECT 3546.270 2872.060 3558.935 2872.140 ;
        RECT 3546.270 2872.040 3558.930 2872.060 ;
        RECT 3489.650 2868.400 3493.975 2868.460 ;
        RECT 3489.650 2866.800 3502.060 2868.400 ;
        RECT 3489.650 2866.690 3493.975 2866.800 ;
        RECT 3548.560 2865.190 3552.740 2865.280 ;
        RECT 3546.110 2863.590 3552.740 2865.190 ;
        RECT 3548.560 2863.480 3552.740 2863.590 ;
        RECT 3495.650 2859.950 3499.975 2860.055 ;
        RECT 3495.650 2858.350 3502.060 2859.950 ;
        RECT 3495.650 2858.285 3499.975 2858.350 ;
        RECT 3554.525 2856.740 3558.710 2856.820 ;
        RECT 3546.110 2855.140 3558.710 2856.740 ;
        RECT 3554.525 2855.045 3558.710 2855.140 ;
        RECT 3489.680 2851.500 3494.005 2851.600 ;
        RECT 3489.680 2849.900 3502.060 2851.500 ;
        RECT 3489.680 2849.830 3494.005 2849.900 ;
        RECT 221.390 2834.880 233.670 2840.150 ;
        RECT 205.340 2826.970 217.620 2832.240 ;
        RECT 89.230 2804.780 93.425 2804.895 ;
        RECT 71.550 2803.180 93.425 2804.780 ;
        RECT 89.230 2803.090 93.425 2803.180 ;
        RECT 95.260 2801.280 99.455 2801.350 ;
        RECT 71.550 2799.680 99.610 2801.280 ;
        RECT 95.260 2799.545 99.455 2799.680 ;
        RECT 89.245 2780.750 93.455 2780.840 ;
        RECT 87.120 2779.150 93.540 2780.750 ;
        RECT 89.245 2779.040 93.455 2779.150 ;
        RECT 95.280 2772.300 99.490 2772.365 ;
        RECT 87.120 2770.700 99.500 2772.300 ;
        RECT 95.280 2770.620 99.490 2770.700 ;
        RECT 89.285 2763.850 93.495 2763.890 ;
        RECT 87.120 2762.250 93.495 2763.850 ;
        RECT 89.285 2762.145 93.495 2762.250 ;
        RECT 95.265 2755.400 99.475 2755.475 ;
        RECT 87.120 2753.800 99.500 2755.400 ;
        RECT 95.265 2753.730 99.475 2753.800 ;
        RECT 89.265 2746.950 93.475 2747.025 ;
        RECT 87.120 2745.350 93.510 2746.950 ;
        RECT 89.265 2745.280 93.475 2745.350 ;
        RECT 95.310 2738.500 99.520 2738.575 ;
        RECT 87.120 2736.900 99.520 2738.500 ;
        RECT 95.310 2736.830 99.520 2736.900 ;
        RECT 3377.040 2707.240 3382.450 2712.730 ;
        RECT 3358.510 2699.150 3363.920 2704.640 ;
        RECT 3495.790 2692.780 3499.920 2692.840 ;
        RECT 3495.790 2691.180 3517.630 2692.780 ;
        RECT 3495.790 2691.125 3499.920 2691.180 ;
        RECT 3489.735 2689.280 3493.865 2689.355 ;
        RECT 3489.570 2687.680 3517.630 2689.280 ;
        RECT 3489.735 2687.640 3493.865 2687.680 ;
        RECT 3548.580 2673.990 3552.765 2674.075 ;
        RECT 3546.270 2672.390 3552.880 2673.990 ;
        RECT 3548.580 2672.300 3552.765 2672.390 ;
        RECT 3495.630 2668.750 3499.955 2668.850 ;
        RECT 3495.630 2667.150 3502.060 2668.750 ;
        RECT 3495.630 2667.080 3499.955 2667.150 ;
        RECT 3554.585 2665.540 3558.770 2665.620 ;
        RECT 3546.270 2663.940 3558.940 2665.540 ;
        RECT 3554.585 2663.845 3558.770 2663.940 ;
        RECT 3489.645 2660.300 3493.970 2660.360 ;
        RECT 3489.645 2658.700 3502.060 2660.300 ;
        RECT 3489.645 2658.590 3493.970 2658.700 ;
        RECT 3548.555 2657.090 3552.740 2657.205 ;
        RECT 3546.270 2655.490 3552.850 2657.090 ;
        RECT 3548.555 2655.430 3552.740 2655.490 ;
        RECT 3495.745 2651.850 3500.070 2651.935 ;
        RECT 3495.745 2650.250 3502.060 2651.850 ;
        RECT 3495.745 2650.165 3500.070 2650.250 ;
        RECT 3554.530 2648.640 3558.940 2648.750 ;
        RECT 3546.270 2647.140 3558.940 2648.640 ;
        RECT 3546.270 2647.060 3558.935 2647.140 ;
        RECT 3546.270 2647.040 3558.930 2647.060 ;
        RECT 3489.650 2643.400 3493.975 2643.460 ;
        RECT 3489.650 2641.800 3502.060 2643.400 ;
        RECT 3489.650 2641.690 3493.975 2641.800 ;
        RECT 3548.560 2640.190 3552.740 2640.280 ;
        RECT 3546.110 2638.590 3552.740 2640.190 ;
        RECT 3548.560 2638.480 3552.740 2638.590 ;
        RECT 3495.650 2634.950 3499.975 2635.055 ;
        RECT 3495.650 2633.350 3502.060 2634.950 ;
        RECT 3495.650 2633.285 3499.975 2633.350 ;
        RECT 3554.525 2631.740 3558.710 2631.820 ;
        RECT 3546.110 2630.140 3558.710 2631.740 ;
        RECT 3554.525 2630.045 3558.710 2630.140 ;
        RECT 3489.680 2626.500 3494.005 2626.600 ;
        RECT 3489.680 2624.900 3502.060 2626.500 ;
        RECT 3489.680 2624.830 3494.005 2624.900 ;
        RECT 3377.040 2487.240 3382.450 2492.730 ;
        RECT 3358.510 2479.150 3363.920 2484.640 ;
        RECT 3495.790 2472.780 3499.920 2472.840 ;
        RECT 3495.790 2471.180 3517.630 2472.780 ;
        RECT 3495.790 2471.125 3499.920 2471.180 ;
        RECT 3489.735 2469.280 3493.865 2469.355 ;
        RECT 3489.570 2467.680 3517.630 2469.280 ;
        RECT 3489.735 2467.640 3493.865 2467.680 ;
        RECT 3548.580 2453.990 3552.765 2454.075 ;
        RECT 3546.270 2452.390 3552.880 2453.990 ;
        RECT 3548.580 2452.300 3552.765 2452.390 ;
        RECT 3495.630 2448.750 3499.955 2448.850 ;
        RECT 3495.630 2447.150 3502.060 2448.750 ;
        RECT 3495.630 2447.080 3499.955 2447.150 ;
        RECT 3554.585 2445.540 3558.770 2445.620 ;
        RECT 3546.270 2443.940 3558.940 2445.540 ;
        RECT 3554.585 2443.845 3558.770 2443.940 ;
        RECT 3489.645 2440.300 3493.970 2440.360 ;
        RECT 3489.645 2438.700 3502.060 2440.300 ;
        RECT 3489.645 2438.590 3493.970 2438.700 ;
        RECT 3548.555 2437.090 3552.740 2437.205 ;
        RECT 3546.270 2435.490 3552.850 2437.090 ;
        RECT 3548.555 2435.430 3552.740 2435.490 ;
        RECT 3495.745 2431.850 3500.070 2431.935 ;
        RECT 3495.745 2430.250 3502.060 2431.850 ;
        RECT 3495.745 2430.165 3500.070 2430.250 ;
        RECT 3554.530 2428.640 3558.940 2428.750 ;
        RECT 3546.270 2427.140 3558.940 2428.640 ;
        RECT 3546.270 2427.060 3558.935 2427.140 ;
        RECT 3546.270 2427.040 3558.930 2427.060 ;
        RECT 3489.650 2423.400 3493.975 2423.460 ;
        RECT 3489.650 2421.800 3502.060 2423.400 ;
        RECT 3489.650 2421.690 3493.975 2421.800 ;
        RECT 3548.560 2420.190 3552.740 2420.280 ;
        RECT 3546.110 2418.590 3552.740 2420.190 ;
        RECT 3548.560 2418.480 3552.740 2418.590 ;
        RECT 3495.650 2414.950 3499.975 2415.055 ;
        RECT 3495.650 2413.350 3502.060 2414.950 ;
        RECT 3495.650 2413.285 3499.975 2413.350 ;
        RECT 3554.525 2411.740 3558.710 2411.820 ;
        RECT 3546.110 2410.140 3558.710 2411.740 ;
        RECT 3554.525 2410.045 3558.710 2410.140 ;
        RECT 3489.680 2406.500 3494.005 2406.600 ;
        RECT 3489.680 2404.900 3502.060 2406.500 ;
        RECT 3489.680 2404.830 3494.005 2404.900 ;
        RECT 221.390 2196.880 233.670 2202.150 ;
        RECT 205.340 2188.970 217.620 2194.240 ;
        RECT 89.230 2166.780 93.425 2166.895 ;
        RECT 71.550 2165.180 93.425 2166.780 ;
        RECT 89.230 2165.090 93.425 2165.180 ;
        RECT 95.260 2163.280 99.455 2163.350 ;
        RECT 71.550 2161.680 99.610 2163.280 ;
        RECT 95.260 2161.545 99.455 2161.680 ;
        RECT 89.245 2142.750 93.455 2142.840 ;
        RECT 87.120 2141.150 93.540 2142.750 ;
        RECT 89.245 2141.040 93.455 2141.150 ;
        RECT 95.280 2134.300 99.490 2134.365 ;
        RECT 87.120 2132.700 99.500 2134.300 ;
        RECT 95.280 2132.620 99.490 2132.700 ;
        RECT 89.285 2125.850 93.495 2125.890 ;
        RECT 87.120 2124.250 93.495 2125.850 ;
        RECT 89.285 2124.145 93.495 2124.250 ;
        RECT 95.265 2117.400 99.475 2117.475 ;
        RECT 87.120 2115.800 99.500 2117.400 ;
        RECT 95.265 2115.730 99.475 2115.800 ;
        RECT 89.265 2108.950 93.475 2109.025 ;
        RECT 87.120 2107.350 93.510 2108.950 ;
        RECT 89.265 2107.280 93.475 2107.350 ;
        RECT 95.310 2100.500 99.520 2100.575 ;
        RECT 87.120 2098.900 99.520 2100.500 ;
        RECT 95.310 2098.830 99.520 2098.900 ;
        RECT 3377.040 2046.240 3382.450 2051.730 ;
        RECT 3358.510 2038.150 3363.920 2043.640 ;
        RECT 3495.790 2031.780 3499.920 2031.840 ;
        RECT 3495.790 2030.180 3517.630 2031.780 ;
        RECT 3495.790 2030.125 3499.920 2030.180 ;
        RECT 3489.735 2028.280 3493.865 2028.355 ;
        RECT 3489.570 2026.680 3517.630 2028.280 ;
        RECT 3489.735 2026.640 3493.865 2026.680 ;
        RECT 3548.580 2012.990 3552.765 2013.075 ;
        RECT 3546.270 2011.390 3552.880 2012.990 ;
        RECT 3548.580 2011.300 3552.765 2011.390 ;
        RECT 3495.630 2007.750 3499.955 2007.850 ;
        RECT 3495.630 2006.150 3502.060 2007.750 ;
        RECT 3495.630 2006.080 3499.955 2006.150 ;
        RECT 3554.585 2004.540 3558.770 2004.620 ;
        RECT 3546.270 2002.940 3558.940 2004.540 ;
        RECT 3554.585 2002.845 3558.770 2002.940 ;
        RECT 3489.645 1999.300 3493.970 1999.360 ;
        RECT 3489.645 1997.700 3502.060 1999.300 ;
        RECT 3489.645 1997.590 3493.970 1997.700 ;
        RECT 3548.555 1996.090 3552.740 1996.205 ;
        RECT 3546.270 1994.490 3552.850 1996.090 ;
        RECT 3548.555 1994.430 3552.740 1994.490 ;
        RECT 3495.745 1990.850 3500.070 1990.935 ;
        RECT 3495.745 1989.250 3502.060 1990.850 ;
        RECT 3495.745 1989.165 3500.070 1989.250 ;
        RECT 3554.530 1987.640 3558.940 1987.750 ;
        RECT 221.390 1980.880 233.670 1986.150 ;
        RECT 3546.270 1986.140 3558.940 1987.640 ;
        RECT 3546.270 1986.060 3558.935 1986.140 ;
        RECT 3546.270 1986.040 3558.930 1986.060 ;
        RECT 3489.650 1982.400 3493.975 1982.460 ;
        RECT 3489.650 1980.800 3502.060 1982.400 ;
        RECT 3489.650 1980.690 3493.975 1980.800 ;
        RECT 3548.560 1979.190 3552.740 1979.280 ;
        RECT 205.340 1972.970 217.620 1978.240 ;
        RECT 3546.110 1977.590 3552.740 1979.190 ;
        RECT 3548.560 1977.480 3552.740 1977.590 ;
        RECT 3495.650 1973.950 3499.975 1974.055 ;
        RECT 3495.650 1972.350 3502.060 1973.950 ;
        RECT 3495.650 1972.285 3499.975 1972.350 ;
        RECT 3554.525 1970.740 3558.710 1970.820 ;
        RECT 3546.110 1969.140 3558.710 1970.740 ;
        RECT 3554.525 1969.045 3558.710 1969.140 ;
        RECT 3489.680 1965.500 3494.005 1965.600 ;
        RECT 3489.680 1963.900 3502.060 1965.500 ;
        RECT 3489.680 1963.830 3494.005 1963.900 ;
        RECT 89.230 1950.780 93.425 1950.895 ;
        RECT 71.550 1949.180 93.425 1950.780 ;
        RECT 89.230 1949.090 93.425 1949.180 ;
        RECT 95.260 1947.280 99.455 1947.350 ;
        RECT 71.550 1945.680 99.610 1947.280 ;
        RECT 95.260 1945.545 99.455 1945.680 ;
        RECT 89.245 1926.750 93.455 1926.840 ;
        RECT 87.120 1925.150 93.540 1926.750 ;
        RECT 89.245 1925.040 93.455 1925.150 ;
        RECT 95.280 1918.300 99.490 1918.365 ;
        RECT 87.120 1916.700 99.500 1918.300 ;
        RECT 95.280 1916.620 99.490 1916.700 ;
        RECT 89.285 1909.850 93.495 1909.890 ;
        RECT 87.120 1908.250 93.495 1909.850 ;
        RECT 89.285 1908.145 93.495 1908.250 ;
        RECT 95.265 1901.400 99.475 1901.475 ;
        RECT 87.120 1899.800 99.500 1901.400 ;
        RECT 95.265 1899.730 99.475 1899.800 ;
        RECT 89.265 1892.950 93.475 1893.025 ;
        RECT 87.120 1891.350 93.510 1892.950 ;
        RECT 89.265 1891.280 93.475 1891.350 ;
        RECT 95.310 1884.500 99.520 1884.575 ;
        RECT 87.120 1882.900 99.520 1884.500 ;
        RECT 95.310 1882.830 99.520 1882.900 ;
        RECT 3377.040 1820.240 3382.450 1825.730 ;
        RECT 3358.510 1812.150 3363.920 1817.640 ;
        RECT 3495.790 1805.780 3499.920 1805.840 ;
        RECT 3495.790 1804.180 3517.630 1805.780 ;
        RECT 3495.790 1804.125 3499.920 1804.180 ;
        RECT 3489.735 1802.280 3493.865 1802.355 ;
        RECT 3489.570 1800.680 3517.630 1802.280 ;
        RECT 3489.735 1800.640 3493.865 1800.680 ;
        RECT 3548.580 1786.990 3552.765 1787.075 ;
        RECT 3546.270 1785.390 3552.880 1786.990 ;
        RECT 3548.580 1785.300 3552.765 1785.390 ;
        RECT 3495.630 1781.750 3499.955 1781.850 ;
        RECT 3495.630 1780.150 3502.060 1781.750 ;
        RECT 3495.630 1780.080 3499.955 1780.150 ;
        RECT 3554.585 1778.540 3558.770 1778.620 ;
        RECT 3546.270 1776.940 3558.940 1778.540 ;
        RECT 3554.585 1776.845 3558.770 1776.940 ;
        RECT 221.390 1769.880 233.670 1775.150 ;
        RECT 3489.645 1773.300 3493.970 1773.360 ;
        RECT 3489.645 1771.700 3502.060 1773.300 ;
        RECT 3489.645 1771.590 3493.970 1771.700 ;
        RECT 3548.555 1770.090 3552.740 1770.205 ;
        RECT 3546.270 1768.490 3552.850 1770.090 ;
        RECT 3548.555 1768.430 3552.740 1768.490 ;
        RECT 205.340 1761.970 217.620 1767.240 ;
        RECT 3495.745 1764.850 3500.070 1764.935 ;
        RECT 3495.745 1763.250 3502.060 1764.850 ;
        RECT 3495.745 1763.165 3500.070 1763.250 ;
        RECT 3554.530 1761.640 3558.940 1761.750 ;
        RECT 3546.270 1760.140 3558.940 1761.640 ;
        RECT 3546.270 1760.060 3558.935 1760.140 ;
        RECT 3546.270 1760.040 3558.930 1760.060 ;
        RECT 3489.650 1756.400 3493.975 1756.460 ;
        RECT 3489.650 1754.800 3502.060 1756.400 ;
        RECT 3489.650 1754.690 3493.975 1754.800 ;
        RECT 3548.560 1753.190 3552.740 1753.280 ;
        RECT 3546.110 1751.590 3552.740 1753.190 ;
        RECT 3548.560 1751.480 3552.740 1751.590 ;
        RECT 3495.650 1747.950 3499.975 1748.055 ;
        RECT 3495.650 1746.350 3502.060 1747.950 ;
        RECT 3495.650 1746.285 3499.975 1746.350 ;
        RECT 3554.525 1744.740 3558.710 1744.820 ;
        RECT 3546.110 1743.140 3558.710 1744.740 ;
        RECT 3554.525 1743.045 3558.710 1743.140 ;
        RECT 3489.680 1739.500 3494.005 1739.600 ;
        RECT 3489.680 1737.900 3502.060 1739.500 ;
        RECT 3489.680 1737.830 3494.005 1737.900 ;
        RECT 89.230 1734.780 93.425 1734.895 ;
        RECT 71.550 1733.180 93.425 1734.780 ;
        RECT 89.230 1733.090 93.425 1733.180 ;
        RECT 95.260 1731.280 99.455 1731.350 ;
        RECT 71.550 1729.680 99.610 1731.280 ;
        RECT 95.260 1729.545 99.455 1729.680 ;
        RECT 89.245 1710.750 93.455 1710.840 ;
        RECT 87.120 1709.150 93.540 1710.750 ;
        RECT 89.245 1709.040 93.455 1709.150 ;
        RECT 95.280 1702.300 99.490 1702.365 ;
        RECT 87.120 1700.700 99.500 1702.300 ;
        RECT 95.280 1700.620 99.490 1700.700 ;
        RECT 89.285 1693.850 93.495 1693.890 ;
        RECT 87.120 1692.250 93.495 1693.850 ;
        RECT 89.285 1692.145 93.495 1692.250 ;
        RECT 95.265 1685.400 99.475 1685.475 ;
        RECT 87.120 1683.800 99.500 1685.400 ;
        RECT 95.265 1683.730 99.475 1683.800 ;
        RECT 89.265 1676.950 93.475 1677.025 ;
        RECT 87.120 1675.350 93.510 1676.950 ;
        RECT 89.265 1675.280 93.475 1675.350 ;
        RECT 95.310 1668.500 99.520 1668.575 ;
        RECT 87.120 1666.900 99.520 1668.500 ;
        RECT 95.310 1666.830 99.520 1666.900 ;
        RECT 3377.040 1595.240 3382.450 1600.730 ;
        RECT 3358.510 1587.150 3363.920 1592.640 ;
        RECT 3495.790 1580.780 3499.920 1580.840 ;
        RECT 3495.790 1579.180 3517.630 1580.780 ;
        RECT 3495.790 1579.125 3499.920 1579.180 ;
        RECT 3489.735 1577.280 3493.865 1577.355 ;
        RECT 3489.570 1575.680 3517.630 1577.280 ;
        RECT 3489.735 1575.640 3493.865 1575.680 ;
        RECT 3548.580 1561.990 3552.765 1562.075 ;
        RECT 3546.270 1560.390 3552.880 1561.990 ;
        RECT 3548.580 1560.300 3552.765 1560.390 ;
        RECT 3495.630 1556.750 3499.955 1556.850 ;
        RECT 3495.630 1555.150 3502.060 1556.750 ;
        RECT 3495.630 1555.080 3499.955 1555.150 ;
        RECT 221.390 1548.880 233.670 1554.150 ;
        RECT 3554.585 1553.540 3558.770 1553.620 ;
        RECT 3546.270 1551.940 3558.940 1553.540 ;
        RECT 3554.585 1551.845 3558.770 1551.940 ;
        RECT 3489.645 1548.300 3493.970 1548.360 ;
        RECT 3489.645 1546.700 3502.060 1548.300 ;
        RECT 3489.645 1546.590 3493.970 1546.700 ;
        RECT 205.340 1540.970 217.620 1546.240 ;
        RECT 3548.555 1545.090 3552.740 1545.205 ;
        RECT 3546.270 1543.490 3552.850 1545.090 ;
        RECT 3548.555 1543.430 3552.740 1543.490 ;
        RECT 3495.745 1539.850 3500.070 1539.935 ;
        RECT 3495.745 1538.250 3502.060 1539.850 ;
        RECT 3495.745 1538.165 3500.070 1538.250 ;
        RECT 3554.530 1536.640 3558.940 1536.750 ;
        RECT 3546.270 1535.140 3558.940 1536.640 ;
        RECT 3546.270 1535.060 3558.935 1535.140 ;
        RECT 3546.270 1535.040 3558.930 1535.060 ;
        RECT 3489.650 1531.400 3493.975 1531.460 ;
        RECT 3489.650 1529.800 3502.060 1531.400 ;
        RECT 3489.650 1529.690 3493.975 1529.800 ;
        RECT 3548.560 1528.190 3552.740 1528.280 ;
        RECT 3546.110 1526.590 3552.740 1528.190 ;
        RECT 3548.560 1526.480 3552.740 1526.590 ;
        RECT 3495.650 1522.950 3499.975 1523.055 ;
        RECT 3495.650 1521.350 3502.060 1522.950 ;
        RECT 3495.650 1521.285 3499.975 1521.350 ;
        RECT 3554.525 1519.740 3558.710 1519.820 ;
        RECT 89.230 1518.780 93.425 1518.895 ;
        RECT 71.550 1517.180 93.425 1518.780 ;
        RECT 3546.110 1518.140 3558.710 1519.740 ;
        RECT 3554.525 1518.045 3558.710 1518.140 ;
        RECT 89.230 1517.090 93.425 1517.180 ;
        RECT 95.260 1515.280 99.455 1515.350 ;
        RECT 71.550 1513.680 99.610 1515.280 ;
        RECT 3489.680 1514.500 3494.005 1514.600 ;
        RECT 95.260 1513.545 99.455 1513.680 ;
        RECT 3489.680 1512.900 3502.060 1514.500 ;
        RECT 3489.680 1512.830 3494.005 1512.900 ;
        RECT 89.245 1494.750 93.455 1494.840 ;
        RECT 87.120 1493.150 93.540 1494.750 ;
        RECT 89.245 1493.040 93.455 1493.150 ;
        RECT 95.280 1486.300 99.490 1486.365 ;
        RECT 87.120 1484.700 99.500 1486.300 ;
        RECT 95.280 1484.620 99.490 1484.700 ;
        RECT 89.285 1477.850 93.495 1477.890 ;
        RECT 87.120 1476.250 93.495 1477.850 ;
        RECT 89.285 1476.145 93.495 1476.250 ;
        RECT 95.265 1469.400 99.475 1469.475 ;
        RECT 87.120 1467.800 99.500 1469.400 ;
        RECT 95.265 1467.730 99.475 1467.800 ;
        RECT 89.265 1460.950 93.475 1461.025 ;
        RECT 87.120 1459.350 93.510 1460.950 ;
        RECT 89.265 1459.280 93.475 1459.350 ;
        RECT 95.310 1452.500 99.520 1452.575 ;
        RECT 87.120 1450.900 99.520 1452.500 ;
        RECT 95.310 1450.830 99.520 1450.900 ;
        RECT 3256.130 1388.920 3315.790 1392.020 ;
        RECT 221.140 1379.440 233.810 1386.310 ;
        RECT 3260.940 1384.120 3315.790 1387.220 ;
        RECT 278.770 1379.320 306.940 1382.420 ;
        RECT 3354.420 1380.370 3366.820 1387.050 ;
        RECT 3370.420 1384.100 3382.820 1391.780 ;
        RECT 214.150 1346.890 217.640 1377.290 ;
        RECT 278.770 1374.520 302.140 1377.620 ;
        RECT 3377.040 1370.240 3382.450 1375.730 ;
        RECT 3358.510 1362.150 3363.920 1367.640 ;
        RECT 3495.790 1355.780 3499.920 1355.840 ;
        RECT 3495.790 1354.180 3517.630 1355.780 ;
        RECT 3495.790 1354.125 3499.920 1354.180 ;
        RECT 3489.735 1352.280 3493.865 1352.355 ;
        RECT 3489.570 1350.680 3517.630 1352.280 ;
        RECT 3489.735 1350.640 3493.865 1350.680 ;
        RECT 3548.580 1336.990 3552.765 1337.075 ;
        RECT 3546.270 1335.390 3552.880 1336.990 ;
        RECT 3548.580 1335.300 3552.765 1335.390 ;
        RECT 3495.630 1331.750 3499.955 1331.850 ;
        RECT 3495.630 1330.150 3502.060 1331.750 ;
        RECT 3495.630 1330.080 3499.955 1330.150 ;
        RECT 3554.585 1328.540 3558.770 1328.620 ;
        RECT 3546.270 1326.940 3558.940 1328.540 ;
        RECT 3554.585 1326.845 3558.770 1326.940 ;
        RECT 3489.645 1323.300 3493.970 1323.360 ;
        RECT 3489.645 1321.700 3502.060 1323.300 ;
        RECT 3489.645 1321.590 3493.970 1321.700 ;
        RECT 3548.555 1320.090 3552.740 1320.205 ;
        RECT 3546.270 1318.490 3552.850 1320.090 ;
        RECT 3548.555 1318.430 3552.740 1318.490 ;
        RECT 3495.745 1314.850 3500.070 1314.935 ;
        RECT 3495.745 1313.250 3502.060 1314.850 ;
        RECT 3495.745 1313.165 3500.070 1313.250 ;
        RECT 3554.530 1311.640 3558.940 1311.750 ;
        RECT 3546.270 1310.140 3558.940 1311.640 ;
        RECT 3546.270 1310.060 3558.935 1310.140 ;
        RECT 3546.270 1310.040 3558.930 1310.060 ;
        RECT 3489.650 1306.400 3493.975 1306.460 ;
        RECT 3489.650 1304.800 3502.060 1306.400 ;
        RECT 3489.650 1304.690 3493.975 1304.800 ;
        RECT 3548.560 1303.190 3552.740 1303.280 ;
        RECT 89.230 1302.780 93.425 1302.895 ;
        RECT 71.550 1301.180 93.425 1302.780 ;
        RECT 3546.110 1301.590 3552.740 1303.190 ;
        RECT 3548.560 1301.480 3552.740 1301.590 ;
        RECT 89.230 1301.090 93.425 1301.180 ;
        RECT 95.260 1299.280 99.455 1299.350 ;
        RECT 71.550 1297.680 99.610 1299.280 ;
        RECT 3495.650 1297.950 3499.975 1298.055 ;
        RECT 95.260 1297.545 99.455 1297.680 ;
        RECT 3495.650 1296.350 3502.060 1297.950 ;
        RECT 3495.650 1296.285 3499.975 1296.350 ;
        RECT 3554.525 1294.740 3558.710 1294.820 ;
        RECT 3546.110 1293.140 3558.710 1294.740 ;
        RECT 3554.525 1293.045 3558.710 1293.140 ;
        RECT 3489.680 1289.500 3494.005 1289.600 ;
        RECT 3489.680 1287.900 3502.060 1289.500 ;
        RECT 3489.680 1287.830 3494.005 1287.900 ;
        RECT 89.245 1278.750 93.455 1278.840 ;
        RECT 87.120 1277.150 93.540 1278.750 ;
        RECT 89.245 1277.040 93.455 1277.150 ;
        RECT 95.280 1270.300 99.490 1270.365 ;
        RECT 87.120 1268.700 99.500 1270.300 ;
        RECT 95.280 1268.620 99.490 1268.700 ;
        RECT 89.285 1261.850 93.495 1261.890 ;
        RECT 87.120 1260.250 93.495 1261.850 ;
        RECT 89.285 1260.145 93.495 1260.250 ;
        RECT 95.265 1253.400 99.475 1253.475 ;
        RECT 87.120 1251.800 99.500 1253.400 ;
        RECT 95.265 1251.730 99.475 1251.800 ;
        RECT 89.265 1244.950 93.475 1245.025 ;
        RECT 87.120 1243.350 93.510 1244.950 ;
        RECT 89.265 1243.280 93.475 1243.350 ;
        RECT 95.310 1236.500 99.520 1236.575 ;
        RECT 87.120 1234.900 99.520 1236.500 ;
        RECT 95.310 1234.830 99.520 1234.900 ;
        RECT 3377.040 1144.240 3382.450 1149.730 ;
        RECT 3358.510 1136.150 3363.920 1141.640 ;
        RECT 3495.790 1129.780 3499.920 1129.840 ;
        RECT 3495.790 1128.180 3517.630 1129.780 ;
        RECT 3495.790 1128.125 3499.920 1128.180 ;
        RECT 3489.735 1126.280 3493.865 1126.355 ;
        RECT 3489.570 1124.680 3517.630 1126.280 ;
        RECT 3489.735 1124.640 3493.865 1124.680 ;
        RECT 3548.580 1110.990 3552.765 1111.075 ;
        RECT 3546.270 1109.390 3552.880 1110.990 ;
        RECT 3548.580 1109.300 3552.765 1109.390 ;
        RECT 3495.630 1105.750 3499.955 1105.850 ;
        RECT 3495.630 1104.150 3502.060 1105.750 ;
        RECT 3495.630 1104.080 3499.955 1104.150 ;
        RECT 3554.585 1102.540 3558.770 1102.620 ;
        RECT 3546.270 1100.940 3558.940 1102.540 ;
        RECT 3554.585 1100.845 3558.770 1100.940 ;
        RECT 3489.645 1097.300 3493.970 1097.360 ;
        RECT 3489.645 1095.700 3502.060 1097.300 ;
        RECT 3489.645 1095.590 3493.970 1095.700 ;
        RECT 3548.555 1094.090 3552.740 1094.205 ;
        RECT 3546.270 1092.490 3552.850 1094.090 ;
        RECT 3548.555 1092.430 3552.740 1092.490 ;
        RECT 3495.745 1088.850 3500.070 1088.935 ;
        RECT 3495.745 1087.250 3502.060 1088.850 ;
        RECT 3495.745 1087.165 3500.070 1087.250 ;
        RECT 89.230 1086.780 93.425 1086.895 ;
        RECT 71.550 1085.180 93.425 1086.780 ;
        RECT 3554.530 1085.640 3558.940 1085.750 ;
        RECT 89.230 1085.090 93.425 1085.180 ;
        RECT 3546.270 1084.140 3558.940 1085.640 ;
        RECT 3546.270 1084.060 3558.935 1084.140 ;
        RECT 3546.270 1084.040 3558.930 1084.060 ;
        RECT 95.260 1083.280 99.455 1083.350 ;
        RECT 71.550 1081.680 99.610 1083.280 ;
        RECT 95.260 1081.545 99.455 1081.680 ;
        RECT 3489.650 1080.400 3493.975 1080.460 ;
        RECT 3489.650 1078.800 3502.060 1080.400 ;
        RECT 3489.650 1078.690 3493.975 1078.800 ;
        RECT 3548.560 1077.190 3552.740 1077.280 ;
        RECT 3546.110 1075.590 3552.740 1077.190 ;
        RECT 3548.560 1075.480 3552.740 1075.590 ;
        RECT 3495.650 1071.950 3499.975 1072.055 ;
        RECT 3495.650 1070.350 3502.060 1071.950 ;
        RECT 3495.650 1070.285 3499.975 1070.350 ;
        RECT 3554.525 1068.740 3558.710 1068.820 ;
        RECT 3546.110 1067.140 3558.710 1068.740 ;
        RECT 3554.525 1067.045 3558.710 1067.140 ;
        RECT 3489.680 1063.500 3494.005 1063.600 ;
        RECT 89.245 1062.750 93.455 1062.840 ;
        RECT 87.120 1061.150 93.540 1062.750 ;
        RECT 3489.680 1061.900 3502.060 1063.500 ;
        RECT 3489.680 1061.830 3494.005 1061.900 ;
        RECT 89.245 1061.040 93.455 1061.150 ;
        RECT 95.280 1054.300 99.490 1054.365 ;
        RECT 87.120 1052.700 99.500 1054.300 ;
        RECT 95.280 1052.620 99.490 1052.700 ;
        RECT 89.285 1045.850 93.495 1045.890 ;
        RECT 87.120 1044.250 93.495 1045.850 ;
        RECT 89.285 1044.145 93.495 1044.250 ;
        RECT 95.265 1037.400 99.475 1037.475 ;
        RECT 87.120 1035.800 99.500 1037.400 ;
        RECT 95.265 1035.730 99.475 1035.800 ;
        RECT 89.265 1028.950 93.475 1029.025 ;
        RECT 87.120 1027.350 93.510 1028.950 ;
        RECT 89.265 1027.280 93.475 1027.350 ;
        RECT 95.310 1020.500 99.520 1020.575 ;
        RECT 87.120 1018.900 99.520 1020.500 ;
        RECT 95.310 1018.830 99.520 1018.900 ;
        RECT 3377.040 919.240 3382.450 924.730 ;
        RECT 3358.510 911.150 3363.920 916.640 ;
        RECT 3495.790 904.780 3499.920 904.840 ;
        RECT 3495.790 903.180 3517.630 904.780 ;
        RECT 3495.790 903.125 3499.920 903.180 ;
        RECT 3489.735 901.280 3493.865 901.355 ;
        RECT 3489.570 899.680 3517.630 901.280 ;
        RECT 3489.735 899.640 3493.865 899.680 ;
        RECT 3548.580 885.990 3552.765 886.075 ;
        RECT 3546.270 884.390 3552.880 885.990 ;
        RECT 3548.580 884.300 3552.765 884.390 ;
        RECT 3495.630 880.750 3499.955 880.850 ;
        RECT 3495.630 879.150 3502.060 880.750 ;
        RECT 3495.630 879.080 3499.955 879.150 ;
        RECT 3554.585 877.540 3558.770 877.620 ;
        RECT 3546.270 875.940 3558.940 877.540 ;
        RECT 3554.585 875.845 3558.770 875.940 ;
        RECT 3489.645 872.300 3493.970 872.360 ;
        RECT 3489.645 870.700 3502.060 872.300 ;
        RECT 3489.645 870.590 3493.970 870.700 ;
        RECT 3548.555 869.090 3552.740 869.205 ;
        RECT 3546.270 867.490 3552.850 869.090 ;
        RECT 3548.555 867.430 3552.740 867.490 ;
        RECT 3495.745 863.850 3500.070 863.935 ;
        RECT 3495.745 862.250 3502.060 863.850 ;
        RECT 3495.745 862.165 3500.070 862.250 ;
        RECT 3554.530 860.640 3558.940 860.750 ;
        RECT 3546.270 859.140 3558.940 860.640 ;
        RECT 3546.270 859.060 3558.935 859.140 ;
        RECT 3546.270 859.040 3558.930 859.060 ;
        RECT 3489.650 855.400 3493.975 855.460 ;
        RECT 3489.650 853.800 3502.060 855.400 ;
        RECT 3489.650 853.690 3493.975 853.800 ;
        RECT 3548.560 852.190 3552.740 852.280 ;
        RECT 3546.110 850.590 3552.740 852.190 ;
        RECT 3548.560 850.480 3552.740 850.590 ;
        RECT 3495.650 846.950 3499.975 847.055 ;
        RECT 3495.650 845.350 3502.060 846.950 ;
        RECT 3495.650 845.285 3499.975 845.350 ;
        RECT 3554.525 843.740 3558.710 843.820 ;
        RECT 3546.110 842.140 3558.710 843.740 ;
        RECT 3554.525 842.045 3558.710 842.140 ;
        RECT 3489.680 838.500 3494.005 838.600 ;
        RECT 3489.680 836.900 3502.060 838.500 ;
        RECT 3489.680 836.830 3494.005 836.900 ;
        RECT 3377.040 693.240 3382.450 698.730 ;
        RECT 3358.510 685.150 3363.920 690.640 ;
        RECT 3495.790 678.780 3499.920 678.840 ;
        RECT 3495.790 677.180 3517.630 678.780 ;
        RECT 3495.790 677.125 3499.920 677.180 ;
        RECT 3489.735 675.280 3493.865 675.355 ;
        RECT 3489.570 673.680 3517.630 675.280 ;
        RECT 3489.735 673.640 3493.865 673.680 ;
        RECT 3548.580 659.990 3552.765 660.075 ;
        RECT 3546.270 658.390 3552.880 659.990 ;
        RECT 3548.580 658.300 3552.765 658.390 ;
        RECT 3495.630 654.750 3499.955 654.850 ;
        RECT 3495.630 653.150 3502.060 654.750 ;
        RECT 3495.630 653.080 3499.955 653.150 ;
        RECT 3554.585 651.540 3558.770 651.620 ;
        RECT 3546.270 649.940 3558.940 651.540 ;
        RECT 3554.585 649.845 3558.770 649.940 ;
        RECT 3489.645 646.300 3493.970 646.360 ;
        RECT 3489.645 644.700 3502.060 646.300 ;
        RECT 3489.645 644.590 3493.970 644.700 ;
        RECT 3548.555 643.090 3552.740 643.205 ;
        RECT 3546.270 641.490 3552.850 643.090 ;
        RECT 3548.555 641.430 3552.740 641.490 ;
        RECT 3495.745 637.850 3500.070 637.935 ;
        RECT 3495.745 636.250 3502.060 637.850 ;
        RECT 3495.745 636.165 3500.070 636.250 ;
        RECT 3554.530 634.640 3558.940 634.750 ;
        RECT 3546.270 633.140 3558.940 634.640 ;
        RECT 3546.270 633.060 3558.935 633.140 ;
        RECT 3546.270 633.040 3558.930 633.060 ;
        RECT 3489.650 629.400 3493.975 629.460 ;
        RECT 3489.650 627.800 3502.060 629.400 ;
        RECT 3489.650 627.690 3493.975 627.800 ;
        RECT 3548.560 626.190 3552.740 626.280 ;
        RECT 3546.110 624.590 3552.740 626.190 ;
        RECT 3548.560 624.480 3552.740 624.590 ;
        RECT 3495.650 620.950 3499.975 621.055 ;
        RECT 3495.650 619.350 3502.060 620.950 ;
        RECT 3495.650 619.285 3499.975 619.350 ;
        RECT 3554.525 617.740 3558.710 617.820 ;
        RECT 3546.110 616.140 3558.710 617.740 ;
        RECT 3554.525 616.045 3558.710 616.140 ;
        RECT 3489.680 612.500 3494.005 612.600 ;
        RECT 3489.680 610.900 3502.060 612.500 ;
        RECT 3489.680 610.830 3494.005 610.900 ;
        RECT 3209.530 465.770 3232.720 467.370 ;
        RECT 643.050 206.310 718.230 208.000 ;
        RECT 650.710 202.910 724.725 204.610 ;
  END
END ./mag/caravel_power_routing
END LIBRARY

