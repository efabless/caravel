magic
tech sky130A
magscale 1 2
timestamp 1607107372
<< obsli1 >>
rect 1104 1071 5980 6001
<< obsm1 >>
rect 566 1040 6518 6032
<< metal2 >>
rect 1122 6277 1178 7077
rect 1674 6277 1730 7077
rect 2226 6277 2282 7077
rect 2962 6277 3018 7077
rect 3514 6277 3570 7077
rect 4066 6277 4122 7077
rect 4802 6277 4858 7077
rect 5354 6277 5410 7077
rect 5906 6277 5962 7077
rect 6458 6277 6514 7077
rect 570 0 626 800
rect 1122 0 1178 800
rect 1674 0 1730 800
rect 2226 0 2282 800
rect 2962 0 3018 800
rect 3514 0 3570 800
rect 4066 0 4122 800
rect 4802 0 4858 800
rect 5354 0 5410 800
rect 5906 0 5962 800
<< obsm2 >>
rect 572 6221 1066 6277
rect 1234 6221 1618 6277
rect 1786 6221 2170 6277
rect 2338 6221 2906 6277
rect 3074 6221 3458 6277
rect 3626 6221 4010 6277
rect 4178 6221 4746 6277
rect 4914 6221 5298 6277
rect 5466 6221 5850 6277
rect 6018 6221 6402 6277
rect 572 856 6512 6221
rect 682 800 1066 856
rect 1234 800 1618 856
rect 1786 800 2170 856
rect 2338 800 2906 856
rect 3074 800 3458 856
rect 3626 800 4010 856
rect 4178 800 4746 856
rect 4914 800 5298 856
rect 5466 800 5850 856
rect 6018 800 6512 856
<< metal3 >>
rect 0 5992 800 6112
rect 0 5176 800 5296
rect 6309 5176 7109 5296
rect 0 4360 800 4480
rect 6309 4360 7109 4480
rect 6309 3544 7109 3664
rect 0 3272 800 3392
rect 0 2456 800 2576
rect 6309 2456 7109 2576
rect 0 1640 800 1760
rect 6309 1640 7109 1760
rect 6309 824 7109 944
<< obsm3 >>
rect 880 5912 6309 6082
rect 800 5376 6309 5912
rect 880 5096 6229 5376
rect 800 4560 6309 5096
rect 880 4280 6229 4560
rect 800 3744 6309 4280
rect 800 3472 6229 3744
rect 880 3464 6229 3472
rect 880 3192 6309 3464
rect 800 2656 6309 3192
rect 880 2376 6229 2656
rect 800 1840 6309 2376
rect 880 1560 6229 1840
rect 800 1024 6309 1560
rect 800 851 6229 1024
<< obsm4 >>
rect 1756 1040 5327 6032
<< metal5 >>
rect 1104 2512 5980 2832
rect 1104 1696 5980 2016
<< obsm5 >>
rect 1104 3328 5980 5280
<< labels >>
rlabel metal2 s 4066 6277 4122 7077 6 mask_rev[0]
port 1 nsew
rlabel metal2 s 4066 0 4122 800 6 mask_rev[10]
port 2 nsew
rlabel metal2 s 1122 0 1178 800 6 mask_rev[11]
port 3 nsew
rlabel metal2 s 570 0 626 800 6 mask_rev[12]
port 4 nsew
rlabel metal2 s 5354 6277 5410 7077 6 mask_rev[13]
port 5 nsew
rlabel metal2 s 5906 0 5962 800 6 mask_rev[14]
port 6 nsew
rlabel metal3 s 6309 1640 7109 1760 6 mask_rev[15]
port 7 nsew
rlabel metal2 s 2226 0 2282 800 6 mask_rev[16]
port 8 nsew
rlabel metal2 s 1674 6277 1730 7077 6 mask_rev[17]
port 9 nsew
rlabel metal3 s 0 5176 800 5296 6 mask_rev[18]
port 10 nsew
rlabel metal2 s 2962 6277 3018 7077 6 mask_rev[19]
port 11 nsew
rlabel metal3 s 0 3272 800 3392 6 mask_rev[1]
port 12 nsew
rlabel metal3 s 6309 2456 7109 2576 6 mask_rev[20]
port 13 nsew
rlabel metal3 s 6309 824 7109 944 6 mask_rev[21]
port 14 nsew
rlabel metal3 s 0 5992 800 6112 6 mask_rev[22]
port 15 nsew
rlabel metal2 s 1674 0 1730 800 6 mask_rev[23]
port 16 nsew
rlabel metal2 s 5906 6277 5962 7077 6 mask_rev[24]
port 17 nsew
rlabel metal3 s 0 1640 800 1760 6 mask_rev[25]
port 18 nsew
rlabel metal2 s 4802 6277 4858 7077 6 mask_rev[26]
port 19 nsew
rlabel metal2 s 1122 6277 1178 7077 6 mask_rev[27]
port 20 nsew
rlabel metal2 s 6458 6277 6514 7077 6 mask_rev[28]
port 21 nsew
rlabel metal2 s 5354 0 5410 800 6 mask_rev[29]
port 22 nsew
rlabel metal3 s 0 2456 800 2576 6 mask_rev[2]
port 23 nsew
rlabel metal3 s 6309 5176 7109 5296 6 mask_rev[30]
port 24 nsew
rlabel metal2 s 2962 0 3018 800 6 mask_rev[31]
port 25 nsew
rlabel metal2 s 3514 0 3570 800 6 mask_rev[3]
port 26 nsew
rlabel metal3 s 6309 3544 7109 3664 6 mask_rev[4]
port 27 nsew
rlabel metal3 s 6309 4360 7109 4480 6 mask_rev[5]
port 28 nsew
rlabel metal3 s 0 4360 800 4480 6 mask_rev[6]
port 29 nsew
rlabel metal2 s 3514 6277 3570 7077 6 mask_rev[7]
port 30 nsew
rlabel metal2 s 4802 0 4858 800 6 mask_rev[8]
port 31 nsew
rlabel metal2 s 2226 6277 2282 7077 6 mask_rev[9]
port 32 nsew
rlabel metal5 s 1104 1696 5980 2016 6 VPWR
port 33 nsew power default
rlabel metal5 s 1104 2512 5980 2832 6 VGND
port 34 nsew ground default
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 7109 7077
string LEFview TRUE
string GDS_FILE ../gds/user_id_programming.gds
string GDS_START 0
<< end >>

