magic
tech sky130A
magscale 1 2
timestamp 1677507609
<< obsli1 >>
rect 92 527 4232 3825
<< obsm1 >>
rect 92 496 4232 3856
<< metal2 >>
rect 132 496 452 3944
rect 852 496 1172 3856
rect 1652 496 1972 3944
rect 2372 496 2692 3856
rect 3172 496 3492 3944
rect 3892 496 4212 3856
rect 2134 0 2190 400
<< obsm2 >>
rect 2136 456 2188 3534
<< metal3 >>
rect 44 3624 4280 3944
rect 44 2824 4280 3144
rect 44 2104 4280 2424
rect 44 1304 4280 1624
rect 44 584 4280 904
<< labels >>
rlabel metal2 s 2134 0 2190 400 6 gpio_logic1
port 1 nsew signal output
rlabel metal2 s 132 496 452 3944 6 vccd1
port 2 nsew power bidirectional
rlabel metal2 s 1652 496 1972 3944 6 vccd1
port 2 nsew power bidirectional
rlabel metal2 s 3172 496 3492 3944 6 vccd1
port 2 nsew power bidirectional
rlabel metal3 s 44 584 4280 904 6 vccd1
port 2 nsew power bidirectional
rlabel metal3 s 44 2104 4280 2424 6 vccd1
port 2 nsew power bidirectional
rlabel metal3 s 44 3624 4280 3944 6 vccd1
port 2 nsew power bidirectional
rlabel metal2 s 852 496 1172 3856 6 vssd1
port 3 nsew ground bidirectional
rlabel metal2 s 2372 496 2692 3856 6 vssd1
port 3 nsew ground bidirectional
rlabel metal2 s 3892 496 4212 3856 6 vssd1
port 3 nsew ground bidirectional
rlabel metal3 s 44 1304 4280 1624 6 vssd1
port 3 nsew ground bidirectional
rlabel metal3 s 44 2824 4280 3144 6 vssd1
port 3 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 4400 4400
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 51880
string GDS_FILE /home/hosni/caravel_sky130/caravel_redesign-2/caravel/openlane/gpio_logic_high/runs/23_02_27_06_19/results/signoff/gpio_logic_high.magic.gds
string GDS_START 20238
<< end >>

