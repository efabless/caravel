magic
tech sky130A
timestamp 0
<< properties >>
string FIXED_BBOX 0 0 0 0
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 257538366
string GDS_FILE /home/hosni/caravan/caravan-mpw9-PnR/caravel/openlane/caravan_core/runs/23_05_24_09_10/results/signoff/caravan_core.magic.gds
string GDS_START 62452332
<< end >>

